module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 ;
  assign n129 = x0 &  x64 ;
  assign n130 = ( x2 & ~n129 ) | ( x2 & 1'b0 ) | ( ~n129 & 1'b0 ) ;
  assign n131 = ~x1 |  x0 ;
  assign n132 = ( x64 & ~n131 ) | ( x64 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n133 = ~x1 & x2 ;
  assign n134 = ( x1 & ~x2 ) | ( x1 & 1'b0 ) | ( ~x2 & 1'b0 ) ;
  assign n135 = n133 | n134 ;
  assign n136 = x0 &  ~n135 ;
  assign n137 = x65 &  n136 ;
  assign n138 = n132 | n137 ;
  assign n139 = ~x0 | ~n135 ;
  assign n140 = ( x64 & ~x65 ) | ( x64 & 1'b0 ) | ( ~x65 & 1'b0 ) ;
  assign n141 = ~x64 & x65 ;
  assign n142 = n140 | n141 ;
  assign n143 = n139 &  n142 ;
  assign n144 = ( n138 & ~n143 ) | ( n138 & n142 ) | ( ~n143 & n142 ) ;
  assign n146 = ( x2 & n130 ) | ( x2 & n144 ) | ( n130 & n144 ) ;
  assign n145 = ( x2 & ~n130 ) | ( x2 & n144 ) | ( ~n130 & n144 ) ;
  assign n147 = ( n130 & ~n146 ) | ( n130 & n145 ) | ( ~n146 & n145 ) ;
  assign n148 = x66 &  n136 ;
  assign n149 = ( x0 & ~x1 ) | ( x0 & x2 ) | ( ~x1 & x2 ) ;
  assign n150 = ~n149 |  x0 ;
  assign n151 = ( x64 & ~n150 ) | ( x64 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n152 = ( x65 & ~n131 ) | ( x65 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n153 = n151 | n152 ;
  assign n154 = n148 | n153 ;
  assign n155 = ~x66 & n141 ;
  assign n156 = ( x66 & ~n141 ) | ( x66 & 1'b0 ) | ( ~n141 & 1'b0 ) ;
  assign n157 = n155 | n156 ;
  assign n158 = n139 | n157 ;
  assign n159 = ( n154 & ~n139 ) | ( n154 & n158 ) | ( ~n139 & n158 ) ;
  assign n160 = ( x2 & ~n144 ) | ( x2 & 1'b0 ) | ( ~n144 & 1'b0 ) ;
  assign n162 = ( n146 & n159 ) | ( n146 & n160 ) | ( n159 & n160 ) ;
  assign n161 = ( n159 & ~n146 ) | ( n159 & n160 ) | ( ~n146 & n160 ) ;
  assign n163 = ( n146 & ~n162 ) | ( n146 & n161 ) | ( ~n162 & n161 ) ;
  assign n167 = ~n136 & x67 ;
  assign n164 = ( x65 & ~n150 ) | ( x65 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n165 = ( x66 & ~n131 ) | ( x66 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n166 = n164 | n165 ;
  assign n168 = ( x67 & ~n167 ) | ( x67 & n166 ) | ( ~n167 & n166 ) ;
  assign n169 = ~x64 & x66 ;
  assign n170 = ( x64 & n169 ) | ( x64 & x65 ) | ( n169 & x65 ) ;
  assign n171 = ( x66 & ~x67 ) | ( x66 & n170 ) | ( ~x67 & n170 ) ;
  assign n172 = ( x66 & x67 ) | ( x66 & n170 ) | ( x67 & n170 ) ;
  assign n173 = ( ~x67 & ~n171 ) | ( ~x67 & n172 ) | ( ~n171 & n172 ) ;
  assign n174 = ( n173 & ~n139 ) | ( n173 & n168 ) | ( ~n139 & n168 ) ;
  assign n175 = n174 | n139 ;
  assign n176 = ( x2 & ~n168 ) | ( x2 & n175 ) | ( ~n168 & n175 ) ;
  assign n177 = ( n168 & ~x2 ) | ( n168 & n175 ) | ( ~x2 & n175 ) ;
  assign n178 = ( n176 & ~n175 ) | ( n176 & n177 ) | ( ~n175 & n177 ) ;
  assign n179 = ( n129 & ~n144 ) | ( n129 & n159 ) | ( ~n144 & n159 ) ;
  assign n180 = ( x2 & n144 ) | ( x2 & n179 ) | ( n144 & n179 ) ;
  assign n181 = ( x2 & ~n180 ) | ( x2 & 1'b0 ) | ( ~n180 & 1'b0 ) ;
  assign n182 = ( x2 & ~x3 ) | ( x2 & 1'b0 ) | ( ~x3 & 1'b0 ) ;
  assign n183 = ~x2 & x3 ;
  assign n184 = n182 | n183 ;
  assign n185 = x64 &  n184 ;
  assign n186 = ( n178 & ~n181 ) | ( n178 & n185 ) | ( ~n181 & n185 ) ;
  assign n187 = ( n178 & ~n185 ) | ( n178 & n181 ) | ( ~n185 & n181 ) ;
  assign n188 = ( n186 & ~n178 ) | ( n186 & n187 ) | ( ~n178 & n187 ) ;
  assign n189 = ( x5 & ~n185 ) | ( x5 & 1'b0 ) | ( ~n185 & 1'b0 ) ;
  assign n190 = ( x3 & x4 ) | ( x3 & n182 ) | ( x4 & n182 ) ;
  assign n191 = ( x3 & ~n183 ) | ( x3 & x4 ) | ( ~n183 & x4 ) ;
  assign n192 = ~n190 &  n191 ;
  assign n193 = x64 &  n192 ;
  assign n194 = ~x4 & x5 ;
  assign n195 = ( x4 & ~x5 ) | ( x4 & 1'b0 ) | ( ~x5 & 1'b0 ) ;
  assign n196 = n194 | n195 ;
  assign n197 = ~n184 |  n196 ;
  assign n198 = ( x65 & ~n197 ) | ( x65 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n199 = n193 | n198 ;
  assign n200 = ~n184 | ~n196 ;
  assign n201 = ( n142 & ~n200 ) | ( n142 & 1'b0 ) | ( ~n200 & 1'b0 ) ;
  assign n202 = n199 | n201 ;
  assign n204 = ( x5 & n189 ) | ( x5 & n202 ) | ( n189 & n202 ) ;
  assign n203 = ( x5 & ~n189 ) | ( x5 & n202 ) | ( ~n189 & n202 ) ;
  assign n205 = ( n189 & ~n204 ) | ( n189 & n203 ) | ( ~n204 & n203 ) ;
  assign n219 = ( n181 & ~n178 ) | ( n181 & n185 ) | ( ~n178 & n185 ) ;
  assign n209 = ~n136 & x68 ;
  assign n206 = ( x66 & ~n150 ) | ( x66 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n207 = ( x67 & ~n131 ) | ( x67 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n208 = n206 | n207 ;
  assign n210 = ( x68 & ~n209 ) | ( x68 & n208 ) | ( ~n209 & n208 ) ;
  assign n212 = ( x67 & x68 ) | ( x67 & n172 ) | ( x68 & n172 ) ;
  assign n211 = ( x67 & ~x68 ) | ( x67 & n172 ) | ( ~x68 & n172 ) ;
  assign n213 = ( x68 & ~n212 ) | ( x68 & n211 ) | ( ~n212 & n211 ) ;
  assign n214 = ( n139 & ~n210 ) | ( n139 & n213 ) | ( ~n210 & n213 ) ;
  assign n215 = ~n139 & n214 ;
  assign n216 = ( x2 & n210 ) | ( x2 & n215 ) | ( n210 & n215 ) ;
  assign n217 = ( x2 & ~n215 ) | ( x2 & n210 ) | ( ~n215 & n210 ) ;
  assign n218 = ( n215 & ~n216 ) | ( n215 & n217 ) | ( ~n216 & n217 ) ;
  assign n220 = ( n205 & ~n219 ) | ( n205 & n218 ) | ( ~n219 & n218 ) ;
  assign n221 = ( n205 & ~n218 ) | ( n205 & n219 ) | ( ~n218 & n219 ) ;
  assign n222 = ( n220 & ~n205 ) | ( n220 & n221 ) | ( ~n205 & n221 ) ;
  assign n233 = ( x5 & ~n185 ) | ( x5 & n202 ) | ( ~n185 & n202 ) ;
  assign n234 = ~n202 & n233 ;
  assign n231 = n200 &  n157 ;
  assign n224 = ( x3 & ~x4 ) | ( x3 & n196 ) | ( ~x4 & n196 ) ;
  assign n223 = ( x3 & ~x4 ) | ( x3 & n184 ) | ( ~x4 & n184 ) ;
  assign n225 = ~n224 |  n223 ;
  assign n229 = x64 &  n225 ;
  assign n226 = ( x66 & ~n197 ) | ( x66 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n227 = x65 &  n192 ;
  assign n228 = n226 | n227 ;
  assign n230 = ( x64 & ~n229 ) | ( x64 & n228 ) | ( ~n229 & n228 ) ;
  assign n232 = ( n157 & ~n231 ) | ( n157 & n230 ) | ( ~n231 & n230 ) ;
  assign n236 = ( x5 & n232 ) | ( x5 & n234 ) | ( n232 & n234 ) ;
  assign n235 = ( x5 & ~n234 ) | ( x5 & n232 ) | ( ~n234 & n232 ) ;
  assign n237 = ( n234 & ~n236 ) | ( n234 & n235 ) | ( ~n236 & n235 ) ;
  assign n238 = ( n205 & n218 ) | ( n205 & n219 ) | ( n218 & n219 ) ;
  assign n242 = ~n136 & x69 ;
  assign n239 = ( x67 & ~n150 ) | ( x67 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n240 = ( x68 & ~n131 ) | ( x68 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n241 = n239 | n240 ;
  assign n243 = ( x69 & ~n242 ) | ( x69 & n241 ) | ( ~n242 & n241 ) ;
  assign n245 = ( x68 & x69 ) | ( x68 & n212 ) | ( x69 & n212 ) ;
  assign n244 = ( x68 & ~x69 ) | ( x68 & n212 ) | ( ~x69 & n212 ) ;
  assign n246 = ( x69 & ~n245 ) | ( x69 & n244 ) | ( ~n245 & n244 ) ;
  assign n247 = ( n139 & ~n243 ) | ( n139 & n246 ) | ( ~n243 & n246 ) ;
  assign n248 = ~n139 & n247 ;
  assign n249 = ( n243 & ~x2 ) | ( n243 & n248 ) | ( ~x2 & n248 ) ;
  assign n250 = ( x2 & ~n243 ) | ( x2 & n248 ) | ( ~n243 & n248 ) ;
  assign n251 = ( n249 & ~n248 ) | ( n249 & n250 ) | ( ~n248 & n250 ) ;
  assign n252 = ( n237 & n238 ) | ( n237 & n251 ) | ( n238 & n251 ) ;
  assign n253 = ( n238 & ~n237 ) | ( n238 & n251 ) | ( ~n237 & n251 ) ;
  assign n254 = ( n237 & ~n252 ) | ( n237 & n253 ) | ( ~n252 & n253 ) ;
  assign n278 = ~n136 & x70 ;
  assign n275 = ( x68 & ~n150 ) | ( x68 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n276 = ( x69 & ~n131 ) | ( x69 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n277 = n275 | n276 ;
  assign n279 = ( x70 & ~n278 ) | ( x70 & n277 ) | ( ~n278 & n277 ) ;
  assign n281 = ( x69 & x70 ) | ( x69 & n245 ) | ( x70 & n245 ) ;
  assign n280 = ( x69 & ~x70 ) | ( x69 & n245 ) | ( ~x70 & n245 ) ;
  assign n282 = ( x70 & ~n281 ) | ( x70 & n280 ) | ( ~n281 & n280 ) ;
  assign n283 = ( n139 & ~n279 ) | ( n139 & n282 ) | ( ~n279 & n282 ) ;
  assign n284 = ~n139 & n283 ;
  assign n285 = ( x2 & n279 ) | ( x2 & n284 ) | ( n279 & n284 ) ;
  assign n286 = ( x2 & ~n284 ) | ( x2 & n279 ) | ( ~n284 & n279 ) ;
  assign n287 = ( n284 & ~n285 ) | ( n284 & n286 ) | ( ~n285 & n286 ) ;
  assign n265 = x65 &  n225 ;
  assign n262 = ( x67 & ~n197 ) | ( x67 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n263 = x66 &  n192 ;
  assign n264 = n262 | n263 ;
  assign n266 = ( x65 & ~n265 ) | ( x65 & n264 ) | ( ~n265 & n264 ) ;
  assign n267 = n173 | n200 ;
  assign n268 = ~n266 & n267 ;
  assign n269 = x5 &  n268 ;
  assign n270 = x5 | n268 ;
  assign n271 = ~n269 & n270 ;
  assign n255 = ( n185 & ~n202 ) | ( n185 & n232 ) | ( ~n202 & n232 ) ;
  assign n256 = ( x5 & n202 ) | ( x5 & n255 ) | ( n202 & n255 ) ;
  assign n257 = ( x5 & ~n256 ) | ( x5 & 1'b0 ) | ( ~n256 & 1'b0 ) ;
  assign n258 = ( x5 & ~x6 ) | ( x5 & 1'b0 ) | ( ~x6 & 1'b0 ) ;
  assign n259 = ~x5 & x6 ;
  assign n260 = n258 | n259 ;
  assign n261 = x64 &  n260 ;
  assign n272 = ( n257 & n261 ) | ( n257 & n271 ) | ( n261 & n271 ) ;
  assign n273 = ( n257 & ~n271 ) | ( n257 & n261 ) | ( ~n271 & n261 ) ;
  assign n274 = ( n271 & ~n272 ) | ( n271 & n273 ) | ( ~n272 & n273 ) ;
  assign n288 = ( n252 & ~n287 ) | ( n252 & n274 ) | ( ~n287 & n274 ) ;
  assign n289 = ( n274 & ~n252 ) | ( n274 & n287 ) | ( ~n252 & n287 ) ;
  assign n290 = ( n288 & ~n274 ) | ( n288 & n289 ) | ( ~n274 & n289 ) ;
  assign n305 = ( x8 & ~n261 ) | ( x8 & 1'b0 ) | ( ~n261 & 1'b0 ) ;
  assign n306 = ( x6 & x7 ) | ( x6 & n258 ) | ( x7 & n258 ) ;
  assign n307 = ( x6 & ~n259 ) | ( x6 & x7 ) | ( ~n259 & x7 ) ;
  assign n308 = ~n306 &  n307 ;
  assign n309 = x64 &  n308 ;
  assign n310 = ~x7 & x8 ;
  assign n311 = ( x7 & ~x8 ) | ( x7 & 1'b0 ) | ( ~x8 & 1'b0 ) ;
  assign n312 = n310 | n311 ;
  assign n313 = ~n260 |  n312 ;
  assign n314 = ( x65 & ~n313 ) | ( x65 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n315 = n309 | n314 ;
  assign n316 = ~n260 | ~n312 ;
  assign n317 = ( n142 & ~n316 ) | ( n142 & 1'b0 ) | ( ~n316 & 1'b0 ) ;
  assign n318 = n315 | n317 ;
  assign n320 = ( x8 & n305 ) | ( x8 & n318 ) | ( n305 & n318 ) ;
  assign n319 = ( x8 & ~n305 ) | ( x8 & n318 ) | ( ~n305 & n318 ) ;
  assign n321 = ( n305 & ~n320 ) | ( n305 & n319 ) | ( ~n320 & n319 ) ;
  assign n325 = x66 &  n225 ;
  assign n322 = ( x68 & ~n197 ) | ( x68 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n323 = x67 &  n192 ;
  assign n324 = n322 | n323 ;
  assign n326 = ( x66 & ~n325 ) | ( x66 & n324 ) | ( ~n325 & n324 ) ;
  assign n327 = ~n200 & n213 ;
  assign n328 = n326 | n327 ;
  assign n329 = ( x5 & ~n328 ) | ( x5 & 1'b0 ) | ( ~n328 & 1'b0 ) ;
  assign n330 = ~x5 & n328 ;
  assign n331 = n329 | n330 ;
  assign n332 = ( n273 & n321 ) | ( n273 & n331 ) | ( n321 & n331 ) ;
  assign n333 = ( n273 & ~n321 ) | ( n273 & n331 ) | ( ~n321 & n331 ) ;
  assign n334 = ( n321 & ~n332 ) | ( n321 & n333 ) | ( ~n332 & n333 ) ;
  assign n294 = ~n136 & x71 ;
  assign n291 = ( x69 & ~n150 ) | ( x69 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n292 = ( x70 & ~n131 ) | ( x70 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n293 = n291 | n292 ;
  assign n295 = ( x71 & ~n294 ) | ( x71 & n293 ) | ( ~n294 & n293 ) ;
  assign n297 = ( x70 & x71 ) | ( x70 & n281 ) | ( x71 & n281 ) ;
  assign n296 = ( x70 & ~x71 ) | ( x70 & n281 ) | ( ~x71 & n281 ) ;
  assign n298 = ( x71 & ~n297 ) | ( x71 & n296 ) | ( ~n297 & n296 ) ;
  assign n299 = ( n139 & ~n295 ) | ( n139 & n298 ) | ( ~n295 & n298 ) ;
  assign n300 = ~n139 & n299 ;
  assign n301 = ( n295 & ~x2 ) | ( n295 & n300 ) | ( ~x2 & n300 ) ;
  assign n302 = ( x2 & ~n295 ) | ( x2 & n300 ) | ( ~n295 & n300 ) ;
  assign n303 = ( n301 & ~n300 ) | ( n301 & n302 ) | ( ~n300 & n302 ) ;
  assign n304 = ( n252 & ~n274 ) | ( n252 & n287 ) | ( ~n274 & n287 ) ;
  assign n335 = ( n303 & n304 ) | ( n303 & n334 ) | ( n304 & n334 ) ;
  assign n336 = ( n303 & ~n334 ) | ( n303 & n304 ) | ( ~n334 & n304 ) ;
  assign n337 = ( n334 & ~n335 ) | ( n334 & n336 ) | ( ~n335 & n336 ) ;
  assign n341 = ~n136 & x72 ;
  assign n338 = ( x70 & ~n150 ) | ( x70 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n339 = ( x71 & ~n131 ) | ( x71 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n340 = n338 | n339 ;
  assign n342 = ( x72 & ~n341 ) | ( x72 & n340 ) | ( ~n341 & n340 ) ;
  assign n344 = ( x71 & x72 ) | ( x71 & n297 ) | ( x72 & n297 ) ;
  assign n343 = ( x71 & ~x72 ) | ( x71 & n297 ) | ( ~x72 & n297 ) ;
  assign n345 = ( x72 & ~n344 ) | ( x72 & n343 ) | ( ~n344 & n343 ) ;
  assign n346 = ( n139 & ~n342 ) | ( n139 & n345 ) | ( ~n342 & n345 ) ;
  assign n347 = ~n139 & n346 ;
  assign n348 = ( x2 & n342 ) | ( x2 & n347 ) | ( n342 & n347 ) ;
  assign n349 = ( x2 & ~n347 ) | ( x2 & n342 ) | ( ~n347 & n342 ) ;
  assign n350 = ( n347 & ~n348 ) | ( n347 & n349 ) | ( ~n348 & n349 ) ;
  assign n352 = ( x6 & ~x7 ) | ( x6 & n312 ) | ( ~x7 & n312 ) ;
  assign n351 = ( x6 & ~x7 ) | ( x6 & n260 ) | ( ~x7 & n260 ) ;
  assign n353 = ~n352 |  n351 ;
  assign n357 = x64 &  n353 ;
  assign n354 = ( x66 & ~n313 ) | ( x66 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n355 = x65 &  n308 ;
  assign n356 = n354 | n355 ;
  assign n358 = ( x64 & ~n357 ) | ( x64 & n356 ) | ( ~n357 & n356 ) ;
  assign n359 = ( n157 & ~n316 ) | ( n157 & 1'b0 ) | ( ~n316 & 1'b0 ) ;
  assign n360 = n358 | n359 ;
  assign n361 = ( x8 & ~n261 ) | ( x8 & n318 ) | ( ~n261 & n318 ) ;
  assign n362 = ~n318 & n361 ;
  assign n363 = ( n360 & ~x8 ) | ( n360 & n362 ) | ( ~x8 & n362 ) ;
  assign n364 = ( x8 & ~n360 ) | ( x8 & n362 ) | ( ~n360 & n362 ) ;
  assign n365 = ( n363 & ~n362 ) | ( n363 & n364 ) | ( ~n362 & n364 ) ;
  assign n369 = x67 &  n225 ;
  assign n366 = ( x69 & ~n197 ) | ( x69 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n367 = x68 &  n192 ;
  assign n368 = n366 | n367 ;
  assign n370 = ( x67 & ~n369 ) | ( x67 & n368 ) | ( ~n369 & n368 ) ;
  assign n371 = ~n200 & n246 ;
  assign n372 = n370 | n371 ;
  assign n373 = ( x5 & ~n372 ) | ( x5 & 1'b0 ) | ( ~n372 & 1'b0 ) ;
  assign n374 = ~x5 & n372 ;
  assign n375 = n373 | n374 ;
  assign n376 = ( n332 & ~n365 ) | ( n332 & n375 ) | ( ~n365 & n375 ) ;
  assign n377 = ( n332 & ~n375 ) | ( n332 & n365 ) | ( ~n375 & n365 ) ;
  assign n378 = ( n376 & ~n332 ) | ( n376 & n377 ) | ( ~n332 & n377 ) ;
  assign n379 = ( n335 & n350 ) | ( n335 & n378 ) | ( n350 & n378 ) ;
  assign n380 = ( n335 & ~n350 ) | ( n335 & n378 ) | ( ~n350 & n378 ) ;
  assign n381 = ( n350 & ~n379 ) | ( n350 & n380 ) | ( ~n379 & n380 ) ;
  assign n395 = ( x8 & ~x9 ) | ( x8 & 1'b0 ) | ( ~x9 & 1'b0 ) ;
  assign n396 = ~x8 & x9 ;
  assign n397 = n395 | n396 ;
  assign n398 = x64 &  n397 ;
  assign n399 = ( n261 & ~n318 ) | ( n261 & n360 ) | ( ~n318 & n360 ) ;
  assign n400 = ( x8 & n318 ) | ( x8 & n399 ) | ( n318 & n399 ) ;
  assign n401 = ( x8 & ~n400 ) | ( x8 & 1'b0 ) | ( ~n400 & 1'b0 ) ;
  assign n405 = x65 &  n353 ;
  assign n402 = ( x67 & ~n313 ) | ( x67 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n403 = x66 &  n308 ;
  assign n404 = n402 | n403 ;
  assign n406 = ( x65 & ~n405 ) | ( x65 & n404 ) | ( ~n405 & n404 ) ;
  assign n407 = n173 | n316 ;
  assign n408 = ~n406 & n407 ;
  assign n409 = x8 &  n408 ;
  assign n410 = x8 | n408 ;
  assign n411 = ~n409 & n410 ;
  assign n412 = ( n398 & ~n401 ) | ( n398 & n411 ) | ( ~n401 & n411 ) ;
  assign n413 = ( n398 & ~n411 ) | ( n398 & n401 ) | ( ~n411 & n401 ) ;
  assign n414 = ( n412 & ~n398 ) | ( n412 & n413 ) | ( ~n398 & n413 ) ;
  assign n415 = ( n332 & n365 ) | ( n332 & n375 ) | ( n365 & n375 ) ;
  assign n419 = x68 &  n225 ;
  assign n416 = ( x70 & ~n197 ) | ( x70 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n417 = x69 &  n192 ;
  assign n418 = n416 | n417 ;
  assign n420 = ( x68 & ~n419 ) | ( x68 & n418 ) | ( ~n419 & n418 ) ;
  assign n421 = ~n200 & n282 ;
  assign n422 = n420 | n421 ;
  assign n423 = ( x5 & ~n422 ) | ( x5 & 1'b0 ) | ( ~n422 & 1'b0 ) ;
  assign n424 = ~x5 & n422 ;
  assign n425 = n423 | n424 ;
  assign n427 = ( n414 & n415 ) | ( n414 & n425 ) | ( n415 & n425 ) ;
  assign n426 = ( n415 & ~n414 ) | ( n415 & n425 ) | ( ~n414 & n425 ) ;
  assign n428 = ( n414 & ~n427 ) | ( n414 & n426 ) | ( ~n427 & n426 ) ;
  assign n385 = ~n136 & x73 ;
  assign n382 = ( x71 & ~n150 ) | ( x71 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n383 = ( x72 & ~n131 ) | ( x72 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n384 = n382 | n383 ;
  assign n386 = ( x73 & ~n385 ) | ( x73 & n384 ) | ( ~n385 & n384 ) ;
  assign n388 = ( x72 & x73 ) | ( x72 & n344 ) | ( x73 & n344 ) ;
  assign n387 = ( x72 & ~x73 ) | ( x72 & n344 ) | ( ~x73 & n344 ) ;
  assign n389 = ( x73 & ~n388 ) | ( x73 & n387 ) | ( ~n388 & n387 ) ;
  assign n390 = ( n139 & ~n386 ) | ( n139 & n389 ) | ( ~n386 & n389 ) ;
  assign n391 = ~n139 & n390 ;
  assign n392 = ( x2 & n386 ) | ( x2 & n391 ) | ( n386 & n391 ) ;
  assign n393 = ( x2 & ~n391 ) | ( x2 & n386 ) | ( ~n391 & n386 ) ;
  assign n394 = ( n391 & ~n392 ) | ( n391 & n393 ) | ( ~n392 & n393 ) ;
  assign n429 = ( n379 & ~n428 ) | ( n379 & n394 ) | ( ~n428 & n394 ) ;
  assign n430 = ( n394 & ~n379 ) | ( n394 & n428 ) | ( ~n379 & n428 ) ;
  assign n431 = ( n429 & ~n394 ) | ( n429 & n430 ) | ( ~n394 & n430 ) ;
  assign n478 = ~n136 & x74 ;
  assign n475 = ( x72 & ~n150 ) | ( x72 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n476 = ( x73 & ~n131 ) | ( x73 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n477 = n475 | n476 ;
  assign n479 = ( x74 & ~n478 ) | ( x74 & n477 ) | ( ~n478 & n477 ) ;
  assign n481 = ( x73 & x74 ) | ( x73 & n388 ) | ( x74 & n388 ) ;
  assign n480 = ( x73 & ~x74 ) | ( x73 & n388 ) | ( ~x74 & n388 ) ;
  assign n482 = ( x74 & ~n481 ) | ( x74 & n480 ) | ( ~n481 & n480 ) ;
  assign n483 = ( n139 & ~n479 ) | ( n139 & n482 ) | ( ~n479 & n482 ) ;
  assign n484 = ~n139 & n483 ;
  assign n485 = ( x2 & n479 ) | ( x2 & n484 ) | ( n479 & n484 ) ;
  assign n486 = ( x2 & ~n484 ) | ( x2 & n479 ) | ( ~n484 & n479 ) ;
  assign n487 = ( n484 & ~n485 ) | ( n484 & n486 ) | ( ~n485 & n486 ) ;
  assign n435 = x66 &  n353 ;
  assign n432 = ( x68 & ~n313 ) | ( x68 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n433 = x67 &  n308 ;
  assign n434 = n432 | n433 ;
  assign n436 = ( x66 & ~n435 ) | ( x66 & n434 ) | ( ~n435 & n434 ) ;
  assign n437 = ( n213 & ~n316 ) | ( n213 & 1'b0 ) | ( ~n316 & 1'b0 ) ;
  assign n438 = n436 | n437 ;
  assign n439 = ( x8 & ~n438 ) | ( x8 & 1'b0 ) | ( ~n438 & 1'b0 ) ;
  assign n440 = ~x8 & n438 ;
  assign n441 = n439 | n440 ;
  assign n442 = ( x11 & ~n398 ) | ( x11 & 1'b0 ) | ( ~n398 & 1'b0 ) ;
  assign n443 = ( x9 & x10 ) | ( x9 & n395 ) | ( x10 & n395 ) ;
  assign n444 = ( x9 & ~n396 ) | ( x9 & x10 ) | ( ~n396 & x10 ) ;
  assign n445 = ~n443 &  n444 ;
  assign n446 = x64 &  n445 ;
  assign n447 = ~x10 & x11 ;
  assign n448 = ( x10 & ~x11 ) | ( x10 & 1'b0 ) | ( ~x11 & 1'b0 ) ;
  assign n449 = n447 | n448 ;
  assign n450 = ~n397 |  n449 ;
  assign n451 = ( x65 & ~n450 ) | ( x65 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n452 = n446 | n451 ;
  assign n453 = ~n397 | ~n449 ;
  assign n454 = ( n142 & ~n453 ) | ( n142 & 1'b0 ) | ( ~n453 & 1'b0 ) ;
  assign n455 = n452 | n454 ;
  assign n457 = ( x11 & n442 ) | ( x11 & n455 ) | ( n442 & n455 ) ;
  assign n456 = ( x11 & ~n442 ) | ( x11 & n455 ) | ( ~n442 & n455 ) ;
  assign n458 = ( n442 & ~n457 ) | ( n442 & n456 ) | ( ~n457 & n456 ) ;
  assign n460 = ( n413 & n441 ) | ( n413 & n458 ) | ( n441 & n458 ) ;
  assign n459 = ( n413 & ~n441 ) | ( n413 & n458 ) | ( ~n441 & n458 ) ;
  assign n461 = ( n441 & ~n460 ) | ( n441 & n459 ) | ( ~n460 & n459 ) ;
  assign n465 = x69 &  n225 ;
  assign n462 = ( x71 & ~n197 ) | ( x71 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n463 = x70 &  n192 ;
  assign n464 = n462 | n463 ;
  assign n466 = ( x69 & ~n465 ) | ( x69 & n464 ) | ( ~n465 & n464 ) ;
  assign n467 = ~n200 & n298 ;
  assign n468 = n466 | n467 ;
  assign n469 = ( x5 & ~n468 ) | ( x5 & 1'b0 ) | ( ~n468 & 1'b0 ) ;
  assign n470 = ~x5 & n468 ;
  assign n471 = n469 | n470 ;
  assign n472 = ( n426 & n461 ) | ( n426 & n471 ) | ( n461 & n471 ) ;
  assign n473 = ( n426 & ~n461 ) | ( n426 & n471 ) | ( ~n461 & n471 ) ;
  assign n474 = ( n461 & ~n472 ) | ( n461 & n473 ) | ( ~n472 & n473 ) ;
  assign n488 = ( n429 & ~n487 ) | ( n429 & n474 ) | ( ~n487 & n474 ) ;
  assign n489 = ( n474 & ~n429 ) | ( n474 & n487 ) | ( ~n429 & n487 ) ;
  assign n490 = ( n488 & ~n474 ) | ( n488 & n489 ) | ( ~n474 & n489 ) ;
  assign n519 = x67 &  n353 ;
  assign n516 = ( x69 & ~n313 ) | ( x69 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n517 = x68 &  n308 ;
  assign n518 = n516 | n517 ;
  assign n520 = ( x67 & ~n519 ) | ( x67 & n518 ) | ( ~n519 & n518 ) ;
  assign n521 = ( n246 & ~n316 ) | ( n246 & 1'b0 ) | ( ~n316 & 1'b0 ) ;
  assign n522 = n520 | n521 ;
  assign n523 = ( x8 & ~n522 ) | ( x8 & 1'b0 ) | ( ~n522 & 1'b0 ) ;
  assign n524 = ~x8 & n522 ;
  assign n525 = n523 | n524 ;
  assign n502 = ( x9 & ~x10 ) | ( x9 & n449 ) | ( ~x10 & n449 ) ;
  assign n501 = ( x9 & ~x10 ) | ( x9 & n397 ) | ( ~x10 & n397 ) ;
  assign n503 = ~n502 |  n501 ;
  assign n507 = x64 &  n503 ;
  assign n504 = ( x66 & ~n450 ) | ( x66 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n505 = x65 &  n445 ;
  assign n506 = n504 | n505 ;
  assign n508 = ( x64 & ~n507 ) | ( x64 & n506 ) | ( ~n507 & n506 ) ;
  assign n509 = ( n157 & ~n453 ) | ( n157 & 1'b0 ) | ( ~n453 & 1'b0 ) ;
  assign n510 = n508 | n509 ;
  assign n511 = ( x11 & n398 ) | ( x11 & n455 ) | ( n398 & n455 ) ;
  assign n512 = ( x11 & ~n511 ) | ( x11 & 1'b0 ) | ( ~n511 & 1'b0 ) ;
  assign n514 = ( x11 & n510 ) | ( x11 & n512 ) | ( n510 & n512 ) ;
  assign n513 = ( n510 & ~x11 ) | ( n510 & n512 ) | ( ~x11 & n512 ) ;
  assign n515 = ( x11 & ~n514 ) | ( x11 & n513 ) | ( ~n514 & n513 ) ;
  assign n526 = ( n460 & ~n525 ) | ( n460 & n515 ) | ( ~n525 & n515 ) ;
  assign n527 = ( n515 & ~n460 ) | ( n515 & n525 ) | ( ~n460 & n525 ) ;
  assign n528 = ( n526 & ~n515 ) | ( n526 & n527 ) | ( ~n515 & n527 ) ;
  assign n494 = x70 &  n225 ;
  assign n491 = ( x72 & ~n197 ) | ( x72 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n492 = x71 &  n192 ;
  assign n493 = n491 | n492 ;
  assign n495 = ( x70 & ~n494 ) | ( x70 & n493 ) | ( ~n494 & n493 ) ;
  assign n496 = ~n200 & n345 ;
  assign n497 = n495 | n496 ;
  assign n498 = ( x5 & ~n497 ) | ( x5 & 1'b0 ) | ( ~n497 & 1'b0 ) ;
  assign n499 = ~x5 & n497 ;
  assign n500 = n498 | n499 ;
  assign n529 = ( n472 & n500 ) | ( n472 & n528 ) | ( n500 & n528 ) ;
  assign n530 = ( n472 & ~n528 ) | ( n472 & n500 ) | ( ~n528 & n500 ) ;
  assign n531 = ( n528 & ~n529 ) | ( n528 & n530 ) | ( ~n529 & n530 ) ;
  assign n532 = ( n429 & n474 ) | ( n429 & n487 ) | ( n474 & n487 ) ;
  assign n536 = ~n136 & x75 ;
  assign n533 = ( x73 & ~n150 ) | ( x73 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n534 = ( x74 & ~n131 ) | ( x74 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n535 = n533 | n534 ;
  assign n537 = ( x75 & ~n536 ) | ( x75 & n535 ) | ( ~n536 & n535 ) ;
  assign n539 = ( x74 & x75 ) | ( x74 & n481 ) | ( x75 & n481 ) ;
  assign n538 = ( x74 & ~x75 ) | ( x74 & n481 ) | ( ~x75 & n481 ) ;
  assign n540 = ( x75 & ~n539 ) | ( x75 & n538 ) | ( ~n539 & n538 ) ;
  assign n541 = ( n139 & ~n537 ) | ( n139 & n540 ) | ( ~n537 & n540 ) ;
  assign n542 = ~n139 & n541 ;
  assign n543 = ( x2 & n537 ) | ( x2 & n542 ) | ( n537 & n542 ) ;
  assign n544 = ( x2 & ~n542 ) | ( x2 & n537 ) | ( ~n542 & n537 ) ;
  assign n545 = ( n542 & ~n543 ) | ( n542 & n544 ) | ( ~n543 & n544 ) ;
  assign n546 = ( n531 & ~n532 ) | ( n531 & n545 ) | ( ~n532 & n545 ) ;
  assign n547 = ( n531 & ~n545 ) | ( n531 & n532 ) | ( ~n545 & n532 ) ;
  assign n548 = ( n546 & ~n531 ) | ( n546 & n547 ) | ( ~n531 & n547 ) ;
  assign n549 = ( x11 & ~x12 ) | ( x11 & 1'b0 ) | ( ~x12 & 1'b0 ) ;
  assign n550 = ~x11 & x12 ;
  assign n551 = n549 | n550 ;
  assign n552 = x64 &  n551 ;
  assign n553 = ( x11 & n510 ) | ( x11 & n511 ) | ( n510 & n511 ) ;
  assign n554 = ( x11 & ~n553 ) | ( x11 & 1'b0 ) | ( ~n553 & 1'b0 ) ;
  assign n558 = x65 &  n503 ;
  assign n555 = ( x67 & ~n450 ) | ( x67 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n556 = x66 &  n445 ;
  assign n557 = n555 | n556 ;
  assign n559 = ( x65 & ~n558 ) | ( x65 & n557 ) | ( ~n558 & n557 ) ;
  assign n560 = n173 | n453 ;
  assign n561 = ~n559 & n560 ;
  assign n562 = x11 &  n561 ;
  assign n563 = x11 | n561 ;
  assign n564 = ~n562 & n563 ;
  assign n565 = ( n552 & ~n554 ) | ( n552 & n564 ) | ( ~n554 & n564 ) ;
  assign n566 = ( n552 & ~n564 ) | ( n552 & n554 ) | ( ~n564 & n554 ) ;
  assign n567 = ( n565 & ~n552 ) | ( n565 & n566 ) | ( ~n552 & n566 ) ;
  assign n571 = x68 &  n353 ;
  assign n568 = ( x70 & ~n313 ) | ( x70 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n569 = x69 &  n308 ;
  assign n570 = n568 | n569 ;
  assign n572 = ( x68 & ~n571 ) | ( x68 & n570 ) | ( ~n571 & n570 ) ;
  assign n573 = ( n282 & ~n316 ) | ( n282 & 1'b0 ) | ( ~n316 & 1'b0 ) ;
  assign n574 = n572 | n573 ;
  assign n575 = ( x8 & ~n574 ) | ( x8 & 1'b0 ) | ( ~n574 & 1'b0 ) ;
  assign n576 = ~x8 & n574 ;
  assign n577 = n575 | n576 ;
  assign n578 = ( n460 & n515 ) | ( n460 & n525 ) | ( n515 & n525 ) ;
  assign n579 = ( n567 & ~n577 ) | ( n567 & n578 ) | ( ~n577 & n578 ) ;
  assign n580 = ( n567 & ~n578 ) | ( n567 & n577 ) | ( ~n578 & n577 ) ;
  assign n581 = ( n579 & ~n567 ) | ( n579 & n580 ) | ( ~n567 & n580 ) ;
  assign n585 = x71 &  n225 ;
  assign n582 = ( x73 & ~n197 ) | ( x73 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n583 = x72 &  n192 ;
  assign n584 = n582 | n583 ;
  assign n586 = ( x71 & ~n585 ) | ( x71 & n584 ) | ( ~n585 & n584 ) ;
  assign n587 = ~n200 & n389 ;
  assign n588 = n586 | n587 ;
  assign n589 = ( x5 & ~n588 ) | ( x5 & 1'b0 ) | ( ~n588 & 1'b0 ) ;
  assign n590 = ~x5 & n588 ;
  assign n591 = n589 | n590 ;
  assign n592 = ( n529 & n581 ) | ( n529 & n591 ) | ( n581 & n591 ) ;
  assign n593 = ( n581 & ~n529 ) | ( n581 & n591 ) | ( ~n529 & n591 ) ;
  assign n594 = ( n529 & ~n592 ) | ( n529 & n593 ) | ( ~n592 & n593 ) ;
  assign n595 = ( n531 & n532 ) | ( n531 & n545 ) | ( n532 & n545 ) ;
  assign n599 = ~n136 & x76 ;
  assign n596 = ( x74 & ~n150 ) | ( x74 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n597 = ( x75 & ~n131 ) | ( x75 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n598 = n596 | n597 ;
  assign n600 = ( x76 & ~n599 ) | ( x76 & n598 ) | ( ~n599 & n598 ) ;
  assign n602 = ( x75 & x76 ) | ( x75 & n539 ) | ( x76 & n539 ) ;
  assign n601 = ( x75 & ~x76 ) | ( x75 & n539 ) | ( ~x76 & n539 ) ;
  assign n603 = ( x76 & ~n602 ) | ( x76 & n601 ) | ( ~n602 & n601 ) ;
  assign n604 = ( n139 & ~n600 ) | ( n139 & n603 ) | ( ~n600 & n603 ) ;
  assign n605 = ~n139 & n604 ;
  assign n606 = ( n600 & ~x2 ) | ( n600 & n605 ) | ( ~x2 & n605 ) ;
  assign n607 = ( x2 & ~n600 ) | ( x2 & n605 ) | ( ~n600 & n605 ) ;
  assign n608 = ( n606 & ~n605 ) | ( n606 & n607 ) | ( ~n605 & n607 ) ;
  assign n610 = ( n594 & n595 ) | ( n594 & n608 ) | ( n595 & n608 ) ;
  assign n609 = ( n595 & ~n594 ) | ( n595 & n608 ) | ( ~n594 & n608 ) ;
  assign n611 = ( n594 & ~n610 ) | ( n594 & n609 ) | ( ~n610 & n609 ) ;
  assign n612 = ( n529 & ~n581 ) | ( n529 & n591 ) | ( ~n581 & n591 ) ;
  assign n626 = x66 &  n503 ;
  assign n623 = ( x68 & ~n450 ) | ( x68 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n624 = x67 &  n445 ;
  assign n625 = n623 | n624 ;
  assign n627 = ( x66 & ~n626 ) | ( x66 & n625 ) | ( ~n626 & n625 ) ;
  assign n628 = ( n213 & ~n453 ) | ( n213 & 1'b0 ) | ( ~n453 & 1'b0 ) ;
  assign n629 = n627 | n628 ;
  assign n630 = ( x11 & ~n629 ) | ( x11 & 1'b0 ) | ( ~n629 & 1'b0 ) ;
  assign n631 = ~x11 & n629 ;
  assign n632 = n630 | n631 ;
  assign n633 = ( x14 & ~n552 ) | ( x14 & 1'b0 ) | ( ~n552 & 1'b0 ) ;
  assign n634 = ( x12 & x13 ) | ( x12 & n549 ) | ( x13 & n549 ) ;
  assign n635 = ( x12 & ~n550 ) | ( x12 & x13 ) | ( ~n550 & x13 ) ;
  assign n636 = ~n634 &  n635 ;
  assign n637 = x64 &  n636 ;
  assign n638 = ~x13 & x14 ;
  assign n639 = ( x13 & ~x14 ) | ( x13 & 1'b0 ) | ( ~x14 & 1'b0 ) ;
  assign n640 = n638 | n639 ;
  assign n641 = ~n551 |  n640 ;
  assign n642 = ( x65 & ~n641 ) | ( x65 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n643 = n637 | n642 ;
  assign n644 = ~n551 | ~n640 ;
  assign n645 = ( n142 & ~n644 ) | ( n142 & 1'b0 ) | ( ~n644 & 1'b0 ) ;
  assign n646 = n643 | n645 ;
  assign n648 = ( x14 & n633 ) | ( x14 & n646 ) | ( n633 & n646 ) ;
  assign n647 = ( x14 & ~n633 ) | ( x14 & n646 ) | ( ~n633 & n646 ) ;
  assign n649 = ( n633 & ~n648 ) | ( n633 & n647 ) | ( ~n648 & n647 ) ;
  assign n651 = ( n566 & n632 ) | ( n566 & n649 ) | ( n632 & n649 ) ;
  assign n650 = ( n566 & ~n632 ) | ( n566 & n649 ) | ( ~n632 & n649 ) ;
  assign n652 = ( n632 & ~n651 ) | ( n632 & n650 ) | ( ~n651 & n650 ) ;
  assign n663 = ( n577 & ~n567 ) | ( n577 & n578 ) | ( ~n567 & n578 ) ;
  assign n656 = x69 &  n353 ;
  assign n653 = ( x71 & ~n313 ) | ( x71 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n654 = x70 &  n308 ;
  assign n655 = n653 | n654 ;
  assign n657 = ( x69 & ~n656 ) | ( x69 & n655 ) | ( ~n656 & n655 ) ;
  assign n658 = ( n298 & ~n316 ) | ( n298 & 1'b0 ) | ( ~n316 & 1'b0 ) ;
  assign n659 = n657 | n658 ;
  assign n660 = ( x8 & ~n659 ) | ( x8 & 1'b0 ) | ( ~n659 & 1'b0 ) ;
  assign n661 = ~x8 & n659 ;
  assign n662 = n660 | n661 ;
  assign n664 = ( n652 & ~n663 ) | ( n652 & n662 ) | ( ~n663 & n662 ) ;
  assign n665 = ( n652 & ~n662 ) | ( n652 & n663 ) | ( ~n662 & n663 ) ;
  assign n666 = ( n664 & ~n652 ) | ( n664 & n665 ) | ( ~n652 & n665 ) ;
  assign n616 = x72 &  n225 ;
  assign n613 = ( x74 & ~n197 ) | ( x74 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n614 = x73 &  n192 ;
  assign n615 = n613 | n614 ;
  assign n617 = ( x72 & ~n616 ) | ( x72 & n615 ) | ( ~n616 & n615 ) ;
  assign n618 = ~n200 & n482 ;
  assign n619 = n617 | n618 ;
  assign n620 = ( x5 & ~n619 ) | ( x5 & 1'b0 ) | ( ~n619 & 1'b0 ) ;
  assign n621 = ~x5 & n619 ;
  assign n622 = n620 | n621 ;
  assign n667 = ( n612 & ~n666 ) | ( n612 & n622 ) | ( ~n666 & n622 ) ;
  assign n668 = ( n612 & ~n622 ) | ( n612 & n666 ) | ( ~n622 & n666 ) ;
  assign n669 = ( n667 & ~n612 ) | ( n667 & n668 ) | ( ~n612 & n668 ) ;
  assign n673 = ~n136 & x77 ;
  assign n670 = ( x75 & ~n150 ) | ( x75 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n671 = ( x76 & ~n131 ) | ( x76 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n672 = n670 | n671 ;
  assign n674 = ( x77 & ~n673 ) | ( x77 & n672 ) | ( ~n673 & n672 ) ;
  assign n676 = ( x76 & x77 ) | ( x76 & n602 ) | ( x77 & n602 ) ;
  assign n675 = ( x76 & ~x77 ) | ( x76 & n602 ) | ( ~x77 & n602 ) ;
  assign n677 = ( x77 & ~n676 ) | ( x77 & n675 ) | ( ~n676 & n675 ) ;
  assign n678 = ( n139 & ~n674 ) | ( n139 & n677 ) | ( ~n674 & n677 ) ;
  assign n679 = ~n139 & n678 ;
  assign n680 = ( x2 & n674 ) | ( x2 & n679 ) | ( n674 & n679 ) ;
  assign n681 = ( x2 & ~n679 ) | ( x2 & n674 ) | ( ~n679 & n674 ) ;
  assign n682 = ( n679 & ~n680 ) | ( n679 & n681 ) | ( ~n680 & n681 ) ;
  assign n683 = ( n669 & ~n609 ) | ( n669 & n682 ) | ( ~n609 & n682 ) ;
  assign n684 = ( n609 & ~n682 ) | ( n609 & n669 ) | ( ~n682 & n669 ) ;
  assign n685 = ( n683 & ~n669 ) | ( n683 & n684 ) | ( ~n669 & n684 ) ;
  assign n689 = ~n136 & x78 ;
  assign n686 = ( x76 & ~n150 ) | ( x76 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n687 = ( x77 & ~n131 ) | ( x77 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n688 = n686 | n687 ;
  assign n690 = ( x78 & ~n689 ) | ( x78 & n688 ) | ( ~n689 & n688 ) ;
  assign n692 = ( x77 & x78 ) | ( x77 & n676 ) | ( x78 & n676 ) ;
  assign n691 = ( x77 & ~x78 ) | ( x77 & n676 ) | ( ~x78 & n676 ) ;
  assign n693 = ( x78 & ~n692 ) | ( x78 & n691 ) | ( ~n692 & n691 ) ;
  assign n694 = ( n139 & ~n690 ) | ( n139 & n693 ) | ( ~n690 & n693 ) ;
  assign n695 = ~n139 & n694 ;
  assign n696 = ( x2 & n690 ) | ( x2 & n695 ) | ( n690 & n695 ) ;
  assign n697 = ( x2 & ~n695 ) | ( x2 & n690 ) | ( ~n695 & n690 ) ;
  assign n698 = ( n695 & ~n696 ) | ( n695 & n697 ) | ( ~n696 & n697 ) ;
  assign n699 = ( n609 & n669 ) | ( n609 & n682 ) | ( n669 & n682 ) ;
  assign n729 = x67 &  n503 ;
  assign n726 = ( x69 & ~n450 ) | ( x69 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n727 = x68 &  n445 ;
  assign n728 = n726 | n727 ;
  assign n730 = ( x67 & ~n729 ) | ( x67 & n728 ) | ( ~n729 & n728 ) ;
  assign n731 = ( n246 & ~n453 ) | ( n246 & 1'b0 ) | ( ~n453 & 1'b0 ) ;
  assign n732 = n730 | n731 ;
  assign n733 = ( x11 & ~n732 ) | ( x11 & 1'b0 ) | ( ~n732 & 1'b0 ) ;
  assign n734 = ~x11 & n732 ;
  assign n735 = n733 | n734 ;
  assign n712 = ( x12 & ~x13 ) | ( x12 & n640 ) | ( ~x13 & n640 ) ;
  assign n711 = ( x12 & ~x13 ) | ( x12 & n551 ) | ( ~x13 & n551 ) ;
  assign n713 = ~n712 |  n711 ;
  assign n717 = x64 &  n713 ;
  assign n714 = ( x66 & ~n641 ) | ( x66 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n715 = x65 &  n636 ;
  assign n716 = n714 | n715 ;
  assign n718 = ( x64 & ~n717 ) | ( x64 & n716 ) | ( ~n717 & n716 ) ;
  assign n719 = ( n157 & ~n644 ) | ( n157 & 1'b0 ) | ( ~n644 & 1'b0 ) ;
  assign n720 = n718 | n719 ;
  assign n721 = ( x14 & n552 ) | ( x14 & n646 ) | ( n552 & n646 ) ;
  assign n722 = ( x14 & ~n721 ) | ( x14 & 1'b0 ) | ( ~n721 & 1'b0 ) ;
  assign n724 = ( x14 & n720 ) | ( x14 & n722 ) | ( n720 & n722 ) ;
  assign n723 = ( n720 & ~x14 ) | ( n720 & n722 ) | ( ~x14 & n722 ) ;
  assign n725 = ( x14 & ~n724 ) | ( x14 & n723 ) | ( ~n724 & n723 ) ;
  assign n736 = ( n651 & ~n735 ) | ( n651 & n725 ) | ( ~n735 & n725 ) ;
  assign n737 = ( n725 & ~n651 ) | ( n725 & n735 ) | ( ~n651 & n735 ) ;
  assign n738 = ( n736 & ~n725 ) | ( n736 & n737 ) | ( ~n725 & n737 ) ;
  assign n739 = ( n652 & n662 ) | ( n652 & n663 ) | ( n662 & n663 ) ;
  assign n743 = x70 &  n353 ;
  assign n740 = ( x72 & ~n313 ) | ( x72 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n741 = x71 &  n308 ;
  assign n742 = n740 | n741 ;
  assign n744 = ( x70 & ~n743 ) | ( x70 & n742 ) | ( ~n743 & n742 ) ;
  assign n745 = ~n316 & n345 ;
  assign n746 = n744 | n745 ;
  assign n747 = ( x8 & ~n746 ) | ( x8 & 1'b0 ) | ( ~n746 & 1'b0 ) ;
  assign n748 = ~x8 & n746 ;
  assign n749 = n747 | n748 ;
  assign n750 = ( n738 & ~n739 ) | ( n738 & n749 ) | ( ~n739 & n749 ) ;
  assign n751 = ( n738 & ~n749 ) | ( n738 & n739 ) | ( ~n749 & n739 ) ;
  assign n752 = ( n750 & ~n738 ) | ( n750 & n751 ) | ( ~n738 & n751 ) ;
  assign n703 = x73 &  n225 ;
  assign n700 = ( x75 & ~n197 ) | ( x75 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n701 = x74 &  n192 ;
  assign n702 = n700 | n701 ;
  assign n704 = ( x73 & ~n703 ) | ( x73 & n702 ) | ( ~n703 & n702 ) ;
  assign n705 = ~n200 & n540 ;
  assign n706 = n704 | n705 ;
  assign n707 = ( x5 & ~n706 ) | ( x5 & 1'b0 ) | ( ~n706 & 1'b0 ) ;
  assign n708 = ~x5 & n706 ;
  assign n709 = n707 | n708 ;
  assign n710 = ( n612 & n622 ) | ( n612 & n666 ) | ( n622 & n666 ) ;
  assign n753 = ( n709 & n710 ) | ( n709 & n752 ) | ( n710 & n752 ) ;
  assign n754 = ( n709 & ~n752 ) | ( n709 & n710 ) | ( ~n752 & n710 ) ;
  assign n755 = ( n752 & ~n753 ) | ( n752 & n754 ) | ( ~n753 & n754 ) ;
  assign n757 = ( n698 & n699 ) | ( n698 & n755 ) | ( n699 & n755 ) ;
  assign n756 = ( n699 & ~n698 ) | ( n699 & n755 ) | ( ~n698 & n755 ) ;
  assign n758 = ( n698 & ~n757 ) | ( n698 & n756 ) | ( ~n757 & n756 ) ;
  assign n762 = ~n136 & x79 ;
  assign n759 = ( x77 & ~n150 ) | ( x77 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n760 = ( x78 & ~n131 ) | ( x78 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n761 = n759 | n760 ;
  assign n763 = ( x79 & ~n762 ) | ( x79 & n761 ) | ( ~n762 & n761 ) ;
  assign n765 = ( x78 & x79 ) | ( x78 & n692 ) | ( x79 & n692 ) ;
  assign n764 = ( x78 & ~x79 ) | ( x78 & n692 ) | ( ~x79 & n692 ) ;
  assign n766 = ( x79 & ~n765 ) | ( x79 & n764 ) | ( ~n765 & n764 ) ;
  assign n767 = ( n139 & ~n763 ) | ( n139 & n766 ) | ( ~n763 & n766 ) ;
  assign n768 = ~n139 & n767 ;
  assign n769 = ( x2 & n763 ) | ( x2 & n768 ) | ( n763 & n768 ) ;
  assign n770 = ( x2 & ~n768 ) | ( x2 & n763 ) | ( ~n768 & n763 ) ;
  assign n771 = ( n768 & ~n769 ) | ( n768 & n770 ) | ( ~n769 & n770 ) ;
  assign n785 = x71 &  n353 ;
  assign n782 = ( x73 & ~n313 ) | ( x73 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n783 = x72 &  n308 ;
  assign n784 = n782 | n783 ;
  assign n786 = ( x71 & ~n785 ) | ( x71 & n784 ) | ( ~n785 & n784 ) ;
  assign n787 = ~n316 & n389 ;
  assign n788 = n786 | n787 ;
  assign n789 = ( x8 & ~n788 ) | ( x8 & 1'b0 ) | ( ~n788 & 1'b0 ) ;
  assign n790 = ~x8 & n788 ;
  assign n791 = n789 | n790 ;
  assign n792 = ( n738 & n739 ) | ( n738 & n749 ) | ( n739 & n749 ) ;
  assign n793 = ( x14 & ~x15 ) | ( x14 & 1'b0 ) | ( ~x15 & 1'b0 ) ;
  assign n794 = ~x14 & x15 ;
  assign n795 = n793 | n794 ;
  assign n796 = x64 &  n795 ;
  assign n797 = ( x14 & n720 ) | ( x14 & n721 ) | ( n720 & n721 ) ;
  assign n798 = ( x14 & ~n797 ) | ( x14 & 1'b0 ) | ( ~n797 & 1'b0 ) ;
  assign n802 = x65 &  n713 ;
  assign n799 = ( x67 & ~n641 ) | ( x67 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n800 = x66 &  n636 ;
  assign n801 = n799 | n800 ;
  assign n803 = ( x65 & ~n802 ) | ( x65 & n801 ) | ( ~n802 & n801 ) ;
  assign n804 = n173 | n644 ;
  assign n805 = ~n803 & n804 ;
  assign n806 = x14 &  n805 ;
  assign n807 = x14 | n805 ;
  assign n808 = ~n806 & n807 ;
  assign n809 = ( n796 & ~n798 ) | ( n796 & n808 ) | ( ~n798 & n808 ) ;
  assign n810 = ( n796 & ~n808 ) | ( n796 & n798 ) | ( ~n808 & n798 ) ;
  assign n811 = ( n809 & ~n796 ) | ( n809 & n810 ) | ( ~n796 & n810 ) ;
  assign n812 = ( n651 & n725 ) | ( n651 & n735 ) | ( n725 & n735 ) ;
  assign n816 = x68 &  n503 ;
  assign n813 = ( x70 & ~n450 ) | ( x70 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n814 = x69 &  n445 ;
  assign n815 = n813 | n814 ;
  assign n817 = ( x68 & ~n816 ) | ( x68 & n815 ) | ( ~n816 & n815 ) ;
  assign n818 = ( n282 & ~n453 ) | ( n282 & 1'b0 ) | ( ~n453 & 1'b0 ) ;
  assign n819 = n817 | n818 ;
  assign n820 = ( x11 & ~n819 ) | ( x11 & 1'b0 ) | ( ~n819 & 1'b0 ) ;
  assign n821 = ~x11 & n819 ;
  assign n822 = n820 | n821 ;
  assign n823 = ( n811 & ~n812 ) | ( n811 & n822 ) | ( ~n812 & n822 ) ;
  assign n824 = ( n812 & ~n811 ) | ( n812 & n822 ) | ( ~n811 & n822 ) ;
  assign n825 = ( n823 & ~n822 ) | ( n823 & n824 ) | ( ~n822 & n824 ) ;
  assign n826 = ( n791 & ~n792 ) | ( n791 & n825 ) | ( ~n792 & n825 ) ;
  assign n827 = ( n791 & ~n825 ) | ( n791 & n792 ) | ( ~n825 & n792 ) ;
  assign n828 = ( n826 & ~n791 ) | ( n826 & n827 ) | ( ~n791 & n827 ) ;
  assign n775 = x74 &  n225 ;
  assign n772 = ( x76 & ~n197 ) | ( x76 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n773 = x75 &  n192 ;
  assign n774 = n772 | n773 ;
  assign n776 = ( x74 & ~n775 ) | ( x74 & n774 ) | ( ~n775 & n774 ) ;
  assign n777 = ~n200 & n603 ;
  assign n778 = n776 | n777 ;
  assign n779 = ( x5 & ~n778 ) | ( x5 & 1'b0 ) | ( ~n778 & 1'b0 ) ;
  assign n780 = ~x5 & n778 ;
  assign n781 = n779 | n780 ;
  assign n830 = ( n753 & n781 ) | ( n753 & n828 ) | ( n781 & n828 ) ;
  assign n829 = ( n753 & ~n828 ) | ( n753 & n781 ) | ( ~n828 & n781 ) ;
  assign n831 = ( n828 & ~n830 ) | ( n828 & n829 ) | ( ~n830 & n829 ) ;
  assign n832 = ( n771 & ~n757 ) | ( n771 & n831 ) | ( ~n757 & n831 ) ;
  assign n833 = ( n757 & ~n831 ) | ( n757 & n771 ) | ( ~n831 & n771 ) ;
  assign n834 = ( n832 & ~n771 ) | ( n832 & n833 ) | ( ~n771 & n833 ) ;
  assign n838 = ~n136 & x80 ;
  assign n835 = ( x78 & ~n150 ) | ( x78 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n836 = ( x79 & ~n131 ) | ( x79 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n837 = n835 | n836 ;
  assign n839 = ( x80 & ~n838 ) | ( x80 & n837 ) | ( ~n838 & n837 ) ;
  assign n841 = ( x79 & x80 ) | ( x79 & n765 ) | ( x80 & n765 ) ;
  assign n840 = ( x79 & ~x80 ) | ( x79 & n765 ) | ( ~x80 & n765 ) ;
  assign n842 = ( x80 & ~n841 ) | ( x80 & n840 ) | ( ~n841 & n840 ) ;
  assign n843 = ( n139 & ~n839 ) | ( n139 & n842 ) | ( ~n839 & n842 ) ;
  assign n844 = ~n139 & n843 ;
  assign n845 = ( x2 & n839 ) | ( x2 & n844 ) | ( n839 & n844 ) ;
  assign n846 = ( x2 & ~n844 ) | ( x2 & n839 ) | ( ~n844 & n839 ) ;
  assign n847 = ( n844 & ~n845 ) | ( n844 & n846 ) | ( ~n845 & n846 ) ;
  assign n861 = x72 &  n353 ;
  assign n858 = ( x74 & ~n313 ) | ( x74 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n859 = x73 &  n308 ;
  assign n860 = n858 | n859 ;
  assign n862 = ( x72 & ~n861 ) | ( x72 & n860 ) | ( ~n861 & n860 ) ;
  assign n863 = ~n316 & n482 ;
  assign n864 = n862 | n863 ;
  assign n865 = ( x8 & ~n864 ) | ( x8 & 1'b0 ) | ( ~n864 & 1'b0 ) ;
  assign n866 = ~x8 & n864 ;
  assign n867 = n865 | n866 ;
  assign n871 = x69 &  n503 ;
  assign n868 = ( x71 & ~n450 ) | ( x71 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n869 = x70 &  n445 ;
  assign n870 = n868 | n869 ;
  assign n872 = ( x69 & ~n871 ) | ( x69 & n870 ) | ( ~n871 & n870 ) ;
  assign n873 = ( n298 & ~n453 ) | ( n298 & 1'b0 ) | ( ~n453 & 1'b0 ) ;
  assign n874 = n872 | n873 ;
  assign n875 = ( x11 & ~n874 ) | ( x11 & 1'b0 ) | ( ~n874 & 1'b0 ) ;
  assign n876 = ~x11 & n874 ;
  assign n877 = n875 | n876 ;
  assign n881 = x66 &  n713 ;
  assign n878 = ( x68 & ~n641 ) | ( x68 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n879 = x67 &  n636 ;
  assign n880 = n878 | n879 ;
  assign n882 = ( x66 & ~n881 ) | ( x66 & n880 ) | ( ~n881 & n880 ) ;
  assign n883 = ( n644 & ~n882 ) | ( n644 & n213 ) | ( ~n882 & n213 ) ;
  assign n884 = ~n644 & n883 ;
  assign n885 = ( n882 & ~x14 ) | ( n882 & n884 ) | ( ~x14 & n884 ) ;
  assign n886 = ( x14 & ~n882 ) | ( x14 & n884 ) | ( ~n882 & n884 ) ;
  assign n887 = ( n885 & ~n884 ) | ( n885 & n886 ) | ( ~n884 & n886 ) ;
  assign n888 = ( x17 & ~n796 ) | ( x17 & 1'b0 ) | ( ~n796 & 1'b0 ) ;
  assign n889 = ( x15 & x16 ) | ( x15 & n793 ) | ( x16 & n793 ) ;
  assign n890 = ( x15 & ~n794 ) | ( x15 & x16 ) | ( ~n794 & x16 ) ;
  assign n891 = ~n889 &  n890 ;
  assign n892 = x64 &  n891 ;
  assign n893 = ~x16 & x17 ;
  assign n894 = ( x16 & ~x17 ) | ( x16 & 1'b0 ) | ( ~x17 & 1'b0 ) ;
  assign n895 = n893 | n894 ;
  assign n896 = ~n795 |  n895 ;
  assign n897 = ( x65 & ~n896 ) | ( x65 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n898 = n892 | n897 ;
  assign n899 = ~n795 | ~n895 ;
  assign n900 = ( n142 & ~n899 ) | ( n142 & 1'b0 ) | ( ~n899 & 1'b0 ) ;
  assign n901 = n898 | n900 ;
  assign n903 = ( x17 & n888 ) | ( x17 & n901 ) | ( n888 & n901 ) ;
  assign n902 = ( x17 & ~n888 ) | ( x17 & n901 ) | ( ~n888 & n901 ) ;
  assign n904 = ( n888 & ~n903 ) | ( n888 & n902 ) | ( ~n903 & n902 ) ;
  assign n906 = ( n810 & n887 ) | ( n810 & n904 ) | ( n887 & n904 ) ;
  assign n905 = ( n810 & ~n887 ) | ( n810 & n904 ) | ( ~n887 & n904 ) ;
  assign n907 = ( n887 & ~n906 ) | ( n887 & n905 ) | ( ~n906 & n905 ) ;
  assign n909 = ( n824 & n877 ) | ( n824 & n907 ) | ( n877 & n907 ) ;
  assign n908 = ( n824 & ~n877 ) | ( n824 & n907 ) | ( ~n877 & n907 ) ;
  assign n910 = ( n877 & ~n909 ) | ( n877 & n908 ) | ( ~n909 & n908 ) ;
  assign n912 = ( n827 & n867 ) | ( n827 & n910 ) | ( n867 & n910 ) ;
  assign n911 = ( n827 & ~n867 ) | ( n827 & n910 ) | ( ~n867 & n910 ) ;
  assign n913 = ( n867 & ~n912 ) | ( n867 & n911 ) | ( ~n912 & n911 ) ;
  assign n851 = x75 &  n225 ;
  assign n848 = ( x77 & ~n197 ) | ( x77 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n849 = x76 &  n192 ;
  assign n850 = n848 | n849 ;
  assign n852 = ( x75 & ~n851 ) | ( x75 & n850 ) | ( ~n851 & n850 ) ;
  assign n853 = ~n200 & n677 ;
  assign n854 = n852 | n853 ;
  assign n855 = ( x5 & ~n854 ) | ( x5 & 1'b0 ) | ( ~n854 & 1'b0 ) ;
  assign n856 = ~x5 & n854 ;
  assign n857 = n855 | n856 ;
  assign n914 = ( n829 & n857 ) | ( n829 & n913 ) | ( n857 & n913 ) ;
  assign n915 = ( n829 & ~n913 ) | ( n829 & n857 ) | ( ~n913 & n857 ) ;
  assign n916 = ( n913 & ~n914 ) | ( n913 & n915 ) | ( ~n914 & n915 ) ;
  assign n918 = ( n833 & n847 ) | ( n833 & n916 ) | ( n847 & n916 ) ;
  assign n917 = ( n833 & ~n847 ) | ( n833 & n916 ) | ( ~n847 & n916 ) ;
  assign n919 = ( n847 & ~n918 ) | ( n847 & n917 ) | ( ~n918 & n917 ) ;
  assign n933 = x73 &  n353 ;
  assign n930 = ( x75 & ~n313 ) | ( x75 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n931 = x74 &  n308 ;
  assign n932 = n930 | n931 ;
  assign n934 = ( x73 & ~n933 ) | ( x73 & n932 ) | ( ~n933 & n932 ) ;
  assign n935 = ~n316 & n540 ;
  assign n936 = n934 | n935 ;
  assign n937 = ( x8 & ~n936 ) | ( x8 & 1'b0 ) | ( ~n936 & 1'b0 ) ;
  assign n938 = ~x8 & n936 ;
  assign n939 = n937 | n938 ;
  assign n958 = x67 &  n713 ;
  assign n955 = ( x69 & ~n641 ) | ( x69 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n956 = x68 &  n636 ;
  assign n957 = n955 | n956 ;
  assign n959 = ( x67 & ~n958 ) | ( x67 & n957 ) | ( ~n958 & n957 ) ;
  assign n960 = ( n246 & ~n644 ) | ( n246 & 1'b0 ) | ( ~n644 & 1'b0 ) ;
  assign n961 = n959 | n960 ;
  assign n962 = ( x14 & ~n961 ) | ( x14 & 1'b0 ) | ( ~n961 & 1'b0 ) ;
  assign n963 = ~x14 & n961 ;
  assign n964 = n962 | n963 ;
  assign n941 = ( x15 & ~x16 ) | ( x15 & n895 ) | ( ~x16 & n895 ) ;
  assign n940 = ( x15 & ~x16 ) | ( x15 & n795 ) | ( ~x16 & n795 ) ;
  assign n942 = ~n941 |  n940 ;
  assign n946 = x64 &  n942 ;
  assign n943 = ( x66 & ~n896 ) | ( x66 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n944 = x65 &  n891 ;
  assign n945 = n943 | n944 ;
  assign n947 = ( x64 & ~n946 ) | ( x64 & n945 ) | ( ~n946 & n945 ) ;
  assign n948 = ( n157 & ~n899 ) | ( n157 & 1'b0 ) | ( ~n899 & 1'b0 ) ;
  assign n949 = n947 | n948 ;
  assign n950 = ( x17 & ~n796 ) | ( x17 & n901 ) | ( ~n796 & n901 ) ;
  assign n951 = ~n901 & n950 ;
  assign n952 = ( n949 & ~x17 ) | ( n949 & n951 ) | ( ~x17 & n951 ) ;
  assign n953 = ( x17 & ~n949 ) | ( x17 & n951 ) | ( ~n949 & n951 ) ;
  assign n954 = ( n952 & ~n951 ) | ( n952 & n953 ) | ( ~n951 & n953 ) ;
  assign n965 = ( n906 & ~n964 ) | ( n906 & n954 ) | ( ~n964 & n954 ) ;
  assign n966 = ( n954 & ~n906 ) | ( n954 & n964 ) | ( ~n906 & n964 ) ;
  assign n967 = ( n965 & ~n954 ) | ( n965 & n966 ) | ( ~n954 & n966 ) ;
  assign n971 = x70 &  n503 ;
  assign n968 = ( x72 & ~n450 ) | ( x72 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n969 = x71 &  n445 ;
  assign n970 = n968 | n969 ;
  assign n972 = ( x70 & ~n971 ) | ( x70 & n970 ) | ( ~n971 & n970 ) ;
  assign n973 = ( n345 & ~n453 ) | ( n345 & 1'b0 ) | ( ~n453 & 1'b0 ) ;
  assign n974 = n972 | n973 ;
  assign n975 = ( x11 & ~n974 ) | ( x11 & 1'b0 ) | ( ~n974 & 1'b0 ) ;
  assign n976 = ~x11 & n974 ;
  assign n977 = n975 | n976 ;
  assign n978 = ( n967 & ~n909 ) | ( n967 & n977 ) | ( ~n909 & n977 ) ;
  assign n979 = ( n909 & ~n977 ) | ( n909 & n967 ) | ( ~n977 & n967 ) ;
  assign n980 = ( n978 & ~n967 ) | ( n978 & n979 ) | ( ~n967 & n979 ) ;
  assign n982 = ( n912 & n939 ) | ( n912 & n980 ) | ( n939 & n980 ) ;
  assign n981 = ( n912 & ~n939 ) | ( n912 & n980 ) | ( ~n939 & n980 ) ;
  assign n983 = ( n939 & ~n982 ) | ( n939 & n981 ) | ( ~n982 & n981 ) ;
  assign n923 = x76 &  n225 ;
  assign n920 = ( x78 & ~n197 ) | ( x78 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n921 = x77 &  n192 ;
  assign n922 = n920 | n921 ;
  assign n924 = ( x76 & ~n923 ) | ( x76 & n922 ) | ( ~n923 & n922 ) ;
  assign n925 = ~n200 & n693 ;
  assign n926 = n924 | n925 ;
  assign n927 = ( x5 & ~n926 ) | ( x5 & 1'b0 ) | ( ~n926 & 1'b0 ) ;
  assign n928 = ~x5 & n926 ;
  assign n929 = n927 | n928 ;
  assign n984 = ( n914 & n929 ) | ( n914 & n983 ) | ( n929 & n983 ) ;
  assign n985 = ( n914 & ~n983 ) | ( n914 & n929 ) | ( ~n983 & n929 ) ;
  assign n986 = ( n983 & ~n984 ) | ( n983 & n985 ) | ( ~n984 & n985 ) ;
  assign n990 = ~n136 & x81 ;
  assign n987 = ( x79 & ~n150 ) | ( x79 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n988 = ( x80 & ~n131 ) | ( x80 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n989 = n987 | n988 ;
  assign n991 = ( x81 & ~n990 ) | ( x81 & n989 ) | ( ~n990 & n989 ) ;
  assign n993 = ( x80 & x81 ) | ( x80 & n841 ) | ( x81 & n841 ) ;
  assign n992 = ( x80 & ~x81 ) | ( x80 & n841 ) | ( ~x81 & n841 ) ;
  assign n994 = ( x81 & ~n993 ) | ( x81 & n992 ) | ( ~n993 & n992 ) ;
  assign n995 = ( n139 & ~n991 ) | ( n139 & n994 ) | ( ~n991 & n994 ) ;
  assign n996 = ~n139 & n995 ;
  assign n997 = ( n991 & ~x2 ) | ( n991 & n996 ) | ( ~x2 & n996 ) ;
  assign n998 = ( x2 & ~n991 ) | ( x2 & n996 ) | ( ~n991 & n996 ) ;
  assign n999 = ( n997 & ~n996 ) | ( n997 & n998 ) | ( ~n996 & n998 ) ;
  assign n1000 = ( n918 & n986 ) | ( n918 & n999 ) | ( n986 & n999 ) ;
  assign n1001 = ( n918 & ~n986 ) | ( n918 & n999 ) | ( ~n986 & n999 ) ;
  assign n1002 = ( n986 & ~n1000 ) | ( n986 & n1001 ) | ( ~n1000 & n1001 ) ;
  assign n1016 = x74 &  n353 ;
  assign n1013 = ( x76 & ~n313 ) | ( x76 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n1014 = x75 &  n308 ;
  assign n1015 = n1013 | n1014 ;
  assign n1017 = ( x74 & ~n1016 ) | ( x74 & n1015 ) | ( ~n1016 & n1015 ) ;
  assign n1018 = ~n316 & n603 ;
  assign n1019 = n1017 | n1018 ;
  assign n1020 = ( x8 & ~n1019 ) | ( x8 & 1'b0 ) | ( ~n1019 & 1'b0 ) ;
  assign n1021 = ~x8 & n1019 ;
  assign n1022 = n1020 | n1021 ;
  assign n1023 = ( x17 & ~x18 ) | ( x17 & 1'b0 ) | ( ~x18 & 1'b0 ) ;
  assign n1024 = ~x17 & x18 ;
  assign n1025 = n1023 | n1024 ;
  assign n1026 = x64 &  n1025 ;
  assign n1027 = ( n796 & ~n901 ) | ( n796 & n949 ) | ( ~n901 & n949 ) ;
  assign n1028 = ( x17 & n901 ) | ( x17 & n1027 ) | ( n901 & n1027 ) ;
  assign n1029 = ( x17 & ~n1028 ) | ( x17 & 1'b0 ) | ( ~n1028 & 1'b0 ) ;
  assign n1033 = x65 &  n942 ;
  assign n1030 = ( x67 & ~n896 ) | ( x67 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n1031 = x66 &  n891 ;
  assign n1032 = n1030 | n1031 ;
  assign n1034 = ( x65 & ~n1033 ) | ( x65 & n1032 ) | ( ~n1033 & n1032 ) ;
  assign n1035 = n173 | n899 ;
  assign n1036 = ~n1034 & n1035 ;
  assign n1037 = x17 &  n1036 ;
  assign n1038 = x17 | n1036 ;
  assign n1039 = ~n1037 & n1038 ;
  assign n1040 = ( n1026 & ~n1029 ) | ( n1026 & n1039 ) | ( ~n1029 & n1039 ) ;
  assign n1041 = ( n1026 & ~n1039 ) | ( n1026 & n1029 ) | ( ~n1039 & n1029 ) ;
  assign n1042 = ( n1040 & ~n1026 ) | ( n1040 & n1041 ) | ( ~n1026 & n1041 ) ;
  assign n1043 = ( n906 & n954 ) | ( n906 & n964 ) | ( n954 & n964 ) ;
  assign n1047 = x68 &  n713 ;
  assign n1044 = ( x70 & ~n641 ) | ( x70 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n1045 = x69 &  n636 ;
  assign n1046 = n1044 | n1045 ;
  assign n1048 = ( x68 & ~n1047 ) | ( x68 & n1046 ) | ( ~n1047 & n1046 ) ;
  assign n1049 = ( n282 & ~n644 ) | ( n282 & 1'b0 ) | ( ~n644 & 1'b0 ) ;
  assign n1050 = n1048 | n1049 ;
  assign n1051 = ( x14 & ~n1050 ) | ( x14 & 1'b0 ) | ( ~n1050 & 1'b0 ) ;
  assign n1052 = ~x14 & n1050 ;
  assign n1053 = n1051 | n1052 ;
  assign n1054 = ( n1042 & ~n1043 ) | ( n1042 & n1053 ) | ( ~n1043 & n1053 ) ;
  assign n1055 = ( n1043 & ~n1042 ) | ( n1043 & n1053 ) | ( ~n1042 & n1053 ) ;
  assign n1056 = ( n1054 & ~n1053 ) | ( n1054 & n1055 ) | ( ~n1053 & n1055 ) ;
  assign n1061 = x71 &  n503 ;
  assign n1058 = ( x73 & ~n450 ) | ( x73 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n1059 = x72 &  n445 ;
  assign n1060 = n1058 | n1059 ;
  assign n1062 = ( x71 & ~n1061 ) | ( x71 & n1060 ) | ( ~n1061 & n1060 ) ;
  assign n1063 = ( n389 & ~n453 ) | ( n389 & 1'b0 ) | ( ~n453 & 1'b0 ) ;
  assign n1064 = n1062 | n1063 ;
  assign n1065 = ( x11 & ~n1064 ) | ( x11 & 1'b0 ) | ( ~n1064 & 1'b0 ) ;
  assign n1066 = ~x11 & n1064 ;
  assign n1067 = n1065 | n1066 ;
  assign n1057 = ( n909 & n967 ) | ( n909 & n977 ) | ( n967 & n977 ) ;
  assign n1068 = ( n1056 & ~n1067 ) | ( n1056 & n1057 ) | ( ~n1067 & n1057 ) ;
  assign n1069 = ( n1056 & ~n1057 ) | ( n1056 & n1067 ) | ( ~n1057 & n1067 ) ;
  assign n1070 = ( n1068 & ~n1056 ) | ( n1068 & n1069 ) | ( ~n1056 & n1069 ) ;
  assign n1071 = ( n1022 & ~n982 ) | ( n1022 & n1070 ) | ( ~n982 & n1070 ) ;
  assign n1072 = ( n982 & ~n1070 ) | ( n982 & n1022 ) | ( ~n1070 & n1022 ) ;
  assign n1073 = ( n1071 & ~n1022 ) | ( n1071 & n1072 ) | ( ~n1022 & n1072 ) ;
  assign n1006 = x77 &  n225 ;
  assign n1003 = ( x79 & ~n197 ) | ( x79 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n1004 = x78 &  n192 ;
  assign n1005 = n1003 | n1004 ;
  assign n1007 = ( x77 & ~n1006 ) | ( x77 & n1005 ) | ( ~n1006 & n1005 ) ;
  assign n1008 = ~n200 & n766 ;
  assign n1009 = n1007 | n1008 ;
  assign n1010 = ( x5 & ~n1009 ) | ( x5 & 1'b0 ) | ( ~n1009 & 1'b0 ) ;
  assign n1011 = ~x5 & n1009 ;
  assign n1012 = n1010 | n1011 ;
  assign n1075 = ( n984 & n1012 ) | ( n984 & n1073 ) | ( n1012 & n1073 ) ;
  assign n1074 = ( n984 & ~n1073 ) | ( n984 & n1012 ) | ( ~n1073 & n1012 ) ;
  assign n1076 = ( n1073 & ~n1075 ) | ( n1073 & n1074 ) | ( ~n1075 & n1074 ) ;
  assign n1080 = ~n136 & x82 ;
  assign n1077 = ( x80 & ~n150 ) | ( x80 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n1078 = ( x81 & ~n131 ) | ( x81 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n1079 = n1077 | n1078 ;
  assign n1081 = ( x82 & ~n1080 ) | ( x82 & n1079 ) | ( ~n1080 & n1079 ) ;
  assign n1083 = ( x81 & x82 ) | ( x81 & n993 ) | ( x82 & n993 ) ;
  assign n1082 = ( x81 & ~x82 ) | ( x81 & n993 ) | ( ~x82 & n993 ) ;
  assign n1084 = ( x82 & ~n1083 ) | ( x82 & n1082 ) | ( ~n1083 & n1082 ) ;
  assign n1085 = ( n139 & ~n1081 ) | ( n139 & n1084 ) | ( ~n1081 & n1084 ) ;
  assign n1086 = ~n139 & n1085 ;
  assign n1087 = ( x2 & n1081 ) | ( x2 & n1086 ) | ( n1081 & n1086 ) ;
  assign n1088 = ( x2 & ~n1086 ) | ( x2 & n1081 ) | ( ~n1086 & n1081 ) ;
  assign n1089 = ( n1086 & ~n1087 ) | ( n1086 & n1088 ) | ( ~n1087 & n1088 ) ;
  assign n1090 = ( n1000 & ~n1076 ) | ( n1000 & n1089 ) | ( ~n1076 & n1089 ) ;
  assign n1091 = ( n1076 & ~n1000 ) | ( n1076 & n1089 ) | ( ~n1000 & n1089 ) ;
  assign n1092 = ( n1090 & ~n1089 ) | ( n1090 & n1091 ) | ( ~n1089 & n1091 ) ;
  assign n1096 = ~n136 & x83 ;
  assign n1093 = ( x81 & ~n150 ) | ( x81 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n1094 = ( x82 & ~n131 ) | ( x82 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n1095 = n1093 | n1094 ;
  assign n1097 = ( x83 & ~n1096 ) | ( x83 & n1095 ) | ( ~n1096 & n1095 ) ;
  assign n1099 = ( x82 & x83 ) | ( x82 & n1083 ) | ( x83 & n1083 ) ;
  assign n1098 = ( x82 & ~x83 ) | ( x82 & n1083 ) | ( ~x83 & n1083 ) ;
  assign n1100 = ( x83 & ~n1099 ) | ( x83 & n1098 ) | ( ~n1099 & n1098 ) ;
  assign n1101 = ( n139 & ~n1097 ) | ( n139 & n1100 ) | ( ~n1097 & n1100 ) ;
  assign n1102 = ~n139 & n1101 ;
  assign n1103 = ( x2 & n1097 ) | ( x2 & n1102 ) | ( n1097 & n1102 ) ;
  assign n1104 = ( x2 & ~n1102 ) | ( x2 & n1097 ) | ( ~n1102 & n1097 ) ;
  assign n1105 = ( n1102 & ~n1103 ) | ( n1102 & n1104 ) | ( ~n1103 & n1104 ) ;
  assign n1109 = x75 &  n353 ;
  assign n1106 = ( x77 & ~n313 ) | ( x77 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n1107 = x76 &  n308 ;
  assign n1108 = n1106 | n1107 ;
  assign n1110 = ( x75 & ~n1109 ) | ( x75 & n1108 ) | ( ~n1109 & n1108 ) ;
  assign n1111 = ~n316 & n677 ;
  assign n1112 = n1110 | n1111 ;
  assign n1113 = ( x8 & ~n1112 ) | ( x8 & 1'b0 ) | ( ~n1112 & 1'b0 ) ;
  assign n1114 = ~x8 & n1112 ;
  assign n1115 = n1113 | n1114 ;
  assign n1119 = x72 &  n503 ;
  assign n1116 = ( x74 & ~n450 ) | ( x74 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n1117 = x73 &  n445 ;
  assign n1118 = n1116 | n1117 ;
  assign n1120 = ( x72 & ~n1119 ) | ( x72 & n1118 ) | ( ~n1119 & n1118 ) ;
  assign n1121 = ~n453 & n482 ;
  assign n1122 = n1120 | n1121 ;
  assign n1123 = ( x11 & ~n1122 ) | ( x11 & 1'b0 ) | ( ~n1122 & 1'b0 ) ;
  assign n1124 = ~x11 & n1122 ;
  assign n1125 = n1123 | n1124 ;
  assign n1129 = x69 &  n713 ;
  assign n1126 = ( x71 & ~n641 ) | ( x71 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n1127 = x70 &  n636 ;
  assign n1128 = n1126 | n1127 ;
  assign n1130 = ( x69 & ~n1129 ) | ( x69 & n1128 ) | ( ~n1129 & n1128 ) ;
  assign n1131 = ( n298 & ~n644 ) | ( n298 & 1'b0 ) | ( ~n644 & 1'b0 ) ;
  assign n1132 = n1130 | n1131 ;
  assign n1133 = ( x14 & ~n1132 ) | ( x14 & 1'b0 ) | ( ~n1132 & 1'b0 ) ;
  assign n1134 = ~x14 & n1132 ;
  assign n1135 = n1133 | n1134 ;
  assign n1139 = x66 &  n942 ;
  assign n1136 = ( x68 & ~n896 ) | ( x68 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n1137 = x67 &  n891 ;
  assign n1138 = n1136 | n1137 ;
  assign n1140 = ( x66 & ~n1139 ) | ( x66 & n1138 ) | ( ~n1139 & n1138 ) ;
  assign n1141 = ( n899 & ~n1140 ) | ( n899 & n213 ) | ( ~n1140 & n213 ) ;
  assign n1142 = ~n899 & n1141 ;
  assign n1143 = ( n1140 & ~x17 ) | ( n1140 & n1142 ) | ( ~x17 & n1142 ) ;
  assign n1144 = ( x17 & ~n1140 ) | ( x17 & n1142 ) | ( ~n1140 & n1142 ) ;
  assign n1145 = ( n1143 & ~n1142 ) | ( n1143 & n1144 ) | ( ~n1142 & n1144 ) ;
  assign n1146 = ( x20 & ~n1026 ) | ( x20 & 1'b0 ) | ( ~n1026 & 1'b0 ) ;
  assign n1147 = ( x18 & x19 ) | ( x18 & n1023 ) | ( x19 & n1023 ) ;
  assign n1148 = ( x18 & ~n1024 ) | ( x18 & x19 ) | ( ~n1024 & x19 ) ;
  assign n1149 = ~n1147 &  n1148 ;
  assign n1150 = x64 &  n1149 ;
  assign n1151 = ~x19 & x20 ;
  assign n1152 = ( x19 & ~x20 ) | ( x19 & 1'b0 ) | ( ~x20 & 1'b0 ) ;
  assign n1153 = n1151 | n1152 ;
  assign n1154 = ~n1025 |  n1153 ;
  assign n1155 = ( x65 & ~n1154 ) | ( x65 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n1156 = n1150 | n1155 ;
  assign n1157 = ~n1025 | ~n1153 ;
  assign n1158 = ( n142 & ~n1157 ) | ( n142 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n1159 = n1156 | n1158 ;
  assign n1161 = ( x20 & n1146 ) | ( x20 & n1159 ) | ( n1146 & n1159 ) ;
  assign n1160 = ( x20 & ~n1146 ) | ( x20 & n1159 ) | ( ~n1146 & n1159 ) ;
  assign n1162 = ( n1146 & ~n1161 ) | ( n1146 & n1160 ) | ( ~n1161 & n1160 ) ;
  assign n1164 = ( n1041 & n1145 ) | ( n1041 & n1162 ) | ( n1145 & n1162 ) ;
  assign n1163 = ( n1041 & ~n1145 ) | ( n1041 & n1162 ) | ( ~n1145 & n1162 ) ;
  assign n1165 = ( n1145 & ~n1164 ) | ( n1145 & n1163 ) | ( ~n1164 & n1163 ) ;
  assign n1167 = ( n1055 & n1135 ) | ( n1055 & n1165 ) | ( n1135 & n1165 ) ;
  assign n1166 = ( n1055 & ~n1135 ) | ( n1055 & n1165 ) | ( ~n1135 & n1165 ) ;
  assign n1168 = ( n1135 & ~n1167 ) | ( n1135 & n1166 ) | ( ~n1167 & n1166 ) ;
  assign n1169 = ( n1057 & ~n1056 ) | ( n1057 & n1067 ) | ( ~n1056 & n1067 ) ;
  assign n1170 = ( n1125 & n1168 ) | ( n1125 & n1169 ) | ( n1168 & n1169 ) ;
  assign n1171 = ( n1168 & ~n1125 ) | ( n1168 & n1169 ) | ( ~n1125 & n1169 ) ;
  assign n1172 = ( n1125 & ~n1170 ) | ( n1125 & n1171 ) | ( ~n1170 & n1171 ) ;
  assign n1173 = ( n1072 & n1115 ) | ( n1072 & n1172 ) | ( n1115 & n1172 ) ;
  assign n1174 = ( n1072 & ~n1115 ) | ( n1072 & n1172 ) | ( ~n1115 & n1172 ) ;
  assign n1175 = ( n1115 & ~n1173 ) | ( n1115 & n1174 ) | ( ~n1173 & n1174 ) ;
  assign n1179 = x78 &  n225 ;
  assign n1176 = ( x80 & ~n197 ) | ( x80 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n1177 = x79 &  n192 ;
  assign n1178 = n1176 | n1177 ;
  assign n1180 = ( x78 & ~n1179 ) | ( x78 & n1178 ) | ( ~n1179 & n1178 ) ;
  assign n1181 = ~n200 & n842 ;
  assign n1182 = n1180 | n1181 ;
  assign n1183 = ( x5 & ~n1182 ) | ( x5 & 1'b0 ) | ( ~n1182 & 1'b0 ) ;
  assign n1184 = ~x5 & n1182 ;
  assign n1185 = n1183 | n1184 ;
  assign n1186 = ( n1074 & n1175 ) | ( n1074 & n1185 ) | ( n1175 & n1185 ) ;
  assign n1187 = ( n1074 & ~n1175 ) | ( n1074 & n1185 ) | ( ~n1175 & n1185 ) ;
  assign n1188 = ( n1175 & ~n1186 ) | ( n1175 & n1187 ) | ( ~n1186 & n1187 ) ;
  assign n1189 = ( n1090 & n1105 ) | ( n1090 & n1188 ) | ( n1105 & n1188 ) ;
  assign n1190 = ( n1090 & ~n1105 ) | ( n1090 & n1188 ) | ( ~n1105 & n1188 ) ;
  assign n1191 = ( n1105 & ~n1189 ) | ( n1105 & n1190 ) | ( ~n1189 & n1190 ) ;
  assign n1218 = x73 &  n503 ;
  assign n1215 = ( x75 & ~n450 ) | ( x75 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n1216 = x74 &  n445 ;
  assign n1217 = n1215 | n1216 ;
  assign n1219 = ( x73 & ~n1218 ) | ( x73 & n1217 ) | ( ~n1218 & n1217 ) ;
  assign n1220 = ~n453 & n540 ;
  assign n1221 = n1219 | n1220 ;
  assign n1222 = ( x11 & ~n1221 ) | ( x11 & 1'b0 ) | ( ~n1221 & 1'b0 ) ;
  assign n1223 = ~x11 & n1221 ;
  assign n1224 = n1222 | n1223 ;
  assign n1243 = x67 &  n942 ;
  assign n1240 = ( x69 & ~n896 ) | ( x69 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n1241 = x68 &  n891 ;
  assign n1242 = n1240 | n1241 ;
  assign n1244 = ( x67 & ~n1243 ) | ( x67 & n1242 ) | ( ~n1243 & n1242 ) ;
  assign n1245 = ( n246 & ~n899 ) | ( n246 & 1'b0 ) | ( ~n899 & 1'b0 ) ;
  assign n1246 = n1244 | n1245 ;
  assign n1247 = ( x17 & ~n1246 ) | ( x17 & 1'b0 ) | ( ~n1246 & 1'b0 ) ;
  assign n1248 = ~x17 & n1246 ;
  assign n1249 = n1247 | n1248 ;
  assign n1226 = ( x18 & ~x19 ) | ( x18 & n1153 ) | ( ~x19 & n1153 ) ;
  assign n1225 = ( x18 & ~x19 ) | ( x18 & n1025 ) | ( ~x19 & n1025 ) ;
  assign n1227 = ~n1226 |  n1225 ;
  assign n1231 = x64 &  n1227 ;
  assign n1228 = ( x66 & ~n1154 ) | ( x66 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n1229 = x65 &  n1149 ;
  assign n1230 = n1228 | n1229 ;
  assign n1232 = ( x64 & ~n1231 ) | ( x64 & n1230 ) | ( ~n1231 & n1230 ) ;
  assign n1233 = ( n157 & ~n1157 ) | ( n157 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n1234 = n1232 | n1233 ;
  assign n1235 = ( x20 & n1026 ) | ( x20 & n1159 ) | ( n1026 & n1159 ) ;
  assign n1236 = ( x20 & ~n1235 ) | ( x20 & 1'b0 ) | ( ~n1235 & 1'b0 ) ;
  assign n1238 = ( x20 & n1234 ) | ( x20 & n1236 ) | ( n1234 & n1236 ) ;
  assign n1237 = ( n1234 & ~x20 ) | ( n1234 & n1236 ) | ( ~x20 & n1236 ) ;
  assign n1239 = ( x20 & ~n1238 ) | ( x20 & n1237 ) | ( ~n1238 & n1237 ) ;
  assign n1250 = ( n1164 & ~n1249 ) | ( n1164 & n1239 ) | ( ~n1249 & n1239 ) ;
  assign n1251 = ( n1239 & ~n1164 ) | ( n1239 & n1249 ) | ( ~n1164 & n1249 ) ;
  assign n1252 = ( n1250 & ~n1239 ) | ( n1250 & n1251 ) | ( ~n1239 & n1251 ) ;
  assign n1256 = x70 &  n713 ;
  assign n1253 = ( x72 & ~n641 ) | ( x72 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n1254 = x71 &  n636 ;
  assign n1255 = n1253 | n1254 ;
  assign n1257 = ( x70 & ~n1256 ) | ( x70 & n1255 ) | ( ~n1256 & n1255 ) ;
  assign n1258 = ( n345 & ~n644 ) | ( n345 & 1'b0 ) | ( ~n644 & 1'b0 ) ;
  assign n1259 = n1257 | n1258 ;
  assign n1260 = ( x14 & ~n1259 ) | ( x14 & 1'b0 ) | ( ~n1259 & 1'b0 ) ;
  assign n1261 = ~x14 & n1259 ;
  assign n1262 = n1260 | n1261 ;
  assign n1263 = ( n1252 & ~n1167 ) | ( n1252 & n1262 ) | ( ~n1167 & n1262 ) ;
  assign n1264 = ( n1167 & ~n1262 ) | ( n1167 & n1252 ) | ( ~n1262 & n1252 ) ;
  assign n1265 = ( n1263 & ~n1252 ) | ( n1263 & n1264 ) | ( ~n1252 & n1264 ) ;
  assign n1267 = ( n1170 & n1224 ) | ( n1170 & n1265 ) | ( n1224 & n1265 ) ;
  assign n1266 = ( n1170 & ~n1224 ) | ( n1170 & n1265 ) | ( ~n1224 & n1265 ) ;
  assign n1268 = ( n1224 & ~n1267 ) | ( n1224 & n1266 ) | ( ~n1267 & n1266 ) ;
  assign n1272 = x76 &  n353 ;
  assign n1269 = ( x78 & ~n313 ) | ( x78 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n1270 = x77 &  n308 ;
  assign n1271 = n1269 | n1270 ;
  assign n1273 = ( x76 & ~n1272 ) | ( x76 & n1271 ) | ( ~n1272 & n1271 ) ;
  assign n1274 = ~n316 & n693 ;
  assign n1275 = n1273 | n1274 ;
  assign n1276 = ( x8 & ~n1275 ) | ( x8 & 1'b0 ) | ( ~n1275 & 1'b0 ) ;
  assign n1277 = ~x8 & n1275 ;
  assign n1278 = n1276 | n1277 ;
  assign n1279 = ( n1268 & ~n1173 ) | ( n1268 & n1278 ) | ( ~n1173 & n1278 ) ;
  assign n1280 = ( n1173 & ~n1278 ) | ( n1173 & n1268 ) | ( ~n1278 & n1268 ) ;
  assign n1281 = ( n1279 & ~n1268 ) | ( n1279 & n1280 ) | ( ~n1268 & n1280 ) ;
  assign n1208 = x79 &  n225 ;
  assign n1205 = ( x81 & ~n197 ) | ( x81 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n1206 = x80 &  n192 ;
  assign n1207 = n1205 | n1206 ;
  assign n1209 = ( x79 & ~n1208 ) | ( x79 & n1207 ) | ( ~n1208 & n1207 ) ;
  assign n1210 = ~n200 & n994 ;
  assign n1211 = n1209 | n1210 ;
  assign n1212 = ( x5 & ~n1211 ) | ( x5 & 1'b0 ) | ( ~n1211 & 1'b0 ) ;
  assign n1213 = ~x5 & n1211 ;
  assign n1214 = n1212 | n1213 ;
  assign n1282 = ( n1186 & n1214 ) | ( n1186 & n1281 ) | ( n1214 & n1281 ) ;
  assign n1283 = ( n1186 & ~n1281 ) | ( n1186 & n1214 ) | ( ~n1281 & n1214 ) ;
  assign n1284 = ( n1281 & ~n1282 ) | ( n1281 & n1283 ) | ( ~n1282 & n1283 ) ;
  assign n1195 = ~n136 & x84 ;
  assign n1192 = ( x82 & ~n150 ) | ( x82 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n1193 = ( x83 & ~n131 ) | ( x83 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n1194 = n1192 | n1193 ;
  assign n1196 = ( x84 & ~n1195 ) | ( x84 & n1194 ) | ( ~n1195 & n1194 ) ;
  assign n1198 = ( x83 & x84 ) | ( x83 & n1099 ) | ( x84 & n1099 ) ;
  assign n1197 = ( x83 & ~x84 ) | ( x83 & n1099 ) | ( ~x84 & n1099 ) ;
  assign n1199 = ( x84 & ~n1198 ) | ( x84 & n1197 ) | ( ~n1198 & n1197 ) ;
  assign n1200 = ( n139 & ~n1196 ) | ( n139 & n1199 ) | ( ~n1196 & n1199 ) ;
  assign n1201 = ~n139 & n1200 ;
  assign n1202 = ( x2 & n1196 ) | ( x2 & n1201 ) | ( n1196 & n1201 ) ;
  assign n1203 = ( x2 & ~n1201 ) | ( x2 & n1196 ) | ( ~n1201 & n1196 ) ;
  assign n1204 = ( n1201 & ~n1202 ) | ( n1201 & n1203 ) | ( ~n1202 & n1203 ) ;
  assign n1285 = ( n1189 & ~n1284 ) | ( n1189 & n1204 ) | ( ~n1284 & n1204 ) ;
  assign n1286 = ( n1204 & ~n1189 ) | ( n1204 & n1284 ) | ( ~n1189 & n1284 ) ;
  assign n1287 = ( n1285 & ~n1204 ) | ( n1285 & n1286 ) | ( ~n1204 & n1286 ) ;
  assign n1291 = ~n136 & x85 ;
  assign n1288 = ( x83 & ~n150 ) | ( x83 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n1289 = ( x84 & ~n131 ) | ( x84 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n1290 = n1288 | n1289 ;
  assign n1292 = ( x85 & ~n1291 ) | ( x85 & n1290 ) | ( ~n1291 & n1290 ) ;
  assign n1294 = ( x84 & x85 ) | ( x84 & n1198 ) | ( x85 & n1198 ) ;
  assign n1293 = ( x84 & ~x85 ) | ( x84 & n1198 ) | ( ~x85 & n1198 ) ;
  assign n1295 = ( x85 & ~n1294 ) | ( x85 & n1293 ) | ( ~n1294 & n1293 ) ;
  assign n1296 = ( n139 & ~n1292 ) | ( n139 & n1295 ) | ( ~n1292 & n1295 ) ;
  assign n1297 = ~n139 & n1296 ;
  assign n1298 = ( x2 & n1292 ) | ( x2 & n1297 ) | ( n1292 & n1297 ) ;
  assign n1299 = ( x2 & ~n1297 ) | ( x2 & n1292 ) | ( ~n1297 & n1292 ) ;
  assign n1300 = ( n1297 & ~n1298 ) | ( n1297 & n1299 ) | ( ~n1298 & n1299 ) ;
  assign n1304 = x77 &  n353 ;
  assign n1301 = ( x79 & ~n313 ) | ( x79 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n1302 = x78 &  n308 ;
  assign n1303 = n1301 | n1302 ;
  assign n1305 = ( x77 & ~n1304 ) | ( x77 & n1303 ) | ( ~n1304 & n1303 ) ;
  assign n1306 = ~n316 & n766 ;
  assign n1307 = n1305 | n1306 ;
  assign n1308 = ( x8 & ~n1307 ) | ( x8 & 1'b0 ) | ( ~n1307 & 1'b0 ) ;
  assign n1309 = ~x8 & n1307 ;
  assign n1310 = n1308 | n1309 ;
  assign n1311 = ( n1173 & n1268 ) | ( n1173 & n1278 ) | ( n1268 & n1278 ) ;
  assign n1315 = x74 &  n503 ;
  assign n1312 = ( x76 & ~n450 ) | ( x76 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n1313 = x75 &  n445 ;
  assign n1314 = n1312 | n1313 ;
  assign n1316 = ( x74 & ~n1315 ) | ( x74 & n1314 ) | ( ~n1315 & n1314 ) ;
  assign n1317 = ~n453 & n603 ;
  assign n1318 = n1316 | n1317 ;
  assign n1319 = ( x11 & ~n1318 ) | ( x11 & 1'b0 ) | ( ~n1318 & 1'b0 ) ;
  assign n1320 = ~x11 & n1318 ;
  assign n1321 = n1319 | n1320 ;
  assign n1322 = ( x20 & ~x21 ) | ( x20 & 1'b0 ) | ( ~x21 & 1'b0 ) ;
  assign n1323 = ~x20 & x21 ;
  assign n1324 = n1322 | n1323 ;
  assign n1325 = x64 &  n1324 ;
  assign n1326 = ( x20 & n1234 ) | ( x20 & n1235 ) | ( n1234 & n1235 ) ;
  assign n1327 = ( x20 & ~n1326 ) | ( x20 & 1'b0 ) | ( ~n1326 & 1'b0 ) ;
  assign n1331 = x65 &  n1227 ;
  assign n1328 = ( x67 & ~n1154 ) | ( x67 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n1329 = x66 &  n1149 ;
  assign n1330 = n1328 | n1329 ;
  assign n1332 = ( x65 & ~n1331 ) | ( x65 & n1330 ) | ( ~n1331 & n1330 ) ;
  assign n1333 = n173 | n1157 ;
  assign n1334 = ~n1332 & n1333 ;
  assign n1335 = x20 &  n1334 ;
  assign n1336 = x20 | n1334 ;
  assign n1337 = ~n1335 & n1336 ;
  assign n1338 = ( n1325 & ~n1327 ) | ( n1325 & n1337 ) | ( ~n1327 & n1337 ) ;
  assign n1339 = ( n1325 & ~n1337 ) | ( n1325 & n1327 ) | ( ~n1337 & n1327 ) ;
  assign n1340 = ( n1338 & ~n1325 ) | ( n1338 & n1339 ) | ( ~n1325 & n1339 ) ;
  assign n1341 = ( n1164 & n1239 ) | ( n1164 & n1249 ) | ( n1239 & n1249 ) ;
  assign n1345 = x68 &  n942 ;
  assign n1342 = ( x70 & ~n896 ) | ( x70 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n1343 = x69 &  n891 ;
  assign n1344 = n1342 | n1343 ;
  assign n1346 = ( x68 & ~n1345 ) | ( x68 & n1344 ) | ( ~n1345 & n1344 ) ;
  assign n1347 = ( n282 & ~n899 ) | ( n282 & 1'b0 ) | ( ~n899 & 1'b0 ) ;
  assign n1348 = n1346 | n1347 ;
  assign n1349 = ( x17 & ~n1348 ) | ( x17 & 1'b0 ) | ( ~n1348 & 1'b0 ) ;
  assign n1350 = ~x17 & n1348 ;
  assign n1351 = n1349 | n1350 ;
  assign n1352 = ( n1340 & ~n1341 ) | ( n1340 & n1351 ) | ( ~n1341 & n1351 ) ;
  assign n1353 = ( n1341 & ~n1340 ) | ( n1341 & n1351 ) | ( ~n1340 & n1351 ) ;
  assign n1354 = ( n1352 & ~n1351 ) | ( n1352 & n1353 ) | ( ~n1351 & n1353 ) ;
  assign n1359 = x71 &  n713 ;
  assign n1356 = ( x73 & ~n641 ) | ( x73 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n1357 = x72 &  n636 ;
  assign n1358 = n1356 | n1357 ;
  assign n1360 = ( x71 & ~n1359 ) | ( x71 & n1358 ) | ( ~n1359 & n1358 ) ;
  assign n1361 = ( n389 & ~n644 ) | ( n389 & 1'b0 ) | ( ~n644 & 1'b0 ) ;
  assign n1362 = n1360 | n1361 ;
  assign n1363 = ( x14 & ~n1362 ) | ( x14 & 1'b0 ) | ( ~n1362 & 1'b0 ) ;
  assign n1364 = ~x14 & n1362 ;
  assign n1365 = n1363 | n1364 ;
  assign n1355 = ( n1167 & n1252 ) | ( n1167 & n1262 ) | ( n1252 & n1262 ) ;
  assign n1366 = ( n1354 & ~n1365 ) | ( n1354 & n1355 ) | ( ~n1365 & n1355 ) ;
  assign n1367 = ( n1354 & ~n1355 ) | ( n1354 & n1365 ) | ( ~n1355 & n1365 ) ;
  assign n1368 = ( n1366 & ~n1354 ) | ( n1366 & n1367 ) | ( ~n1354 & n1367 ) ;
  assign n1369 = ( n1321 & ~n1267 ) | ( n1321 & n1368 ) | ( ~n1267 & n1368 ) ;
  assign n1370 = ( n1267 & ~n1368 ) | ( n1267 & n1321 ) | ( ~n1368 & n1321 ) ;
  assign n1371 = ( n1369 & ~n1321 ) | ( n1369 & n1370 ) | ( ~n1321 & n1370 ) ;
  assign n1372 = ( n1310 & ~n1311 ) | ( n1310 & n1371 ) | ( ~n1311 & n1371 ) ;
  assign n1373 = ( n1310 & ~n1371 ) | ( n1310 & n1311 ) | ( ~n1371 & n1311 ) ;
  assign n1374 = ( n1372 & ~n1310 ) | ( n1372 & n1373 ) | ( ~n1310 & n1373 ) ;
  assign n1378 = x80 &  n225 ;
  assign n1375 = ( x82 & ~n197 ) | ( x82 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n1376 = x81 &  n192 ;
  assign n1377 = n1375 | n1376 ;
  assign n1379 = ( x80 & ~n1378 ) | ( x80 & n1377 ) | ( ~n1378 & n1377 ) ;
  assign n1380 = ~n200 & n1084 ;
  assign n1381 = n1379 | n1380 ;
  assign n1382 = ( x5 & ~n1381 ) | ( x5 & 1'b0 ) | ( ~n1381 & 1'b0 ) ;
  assign n1383 = ~x5 & n1381 ;
  assign n1384 = n1382 | n1383 ;
  assign n1385 = ( n1282 & n1374 ) | ( n1282 & n1384 ) | ( n1374 & n1384 ) ;
  assign n1386 = ( n1374 & ~n1282 ) | ( n1374 & n1384 ) | ( ~n1282 & n1384 ) ;
  assign n1387 = ( n1282 & ~n1385 ) | ( n1282 & n1386 ) | ( ~n1385 & n1386 ) ;
  assign n1388 = ( n1189 & n1204 ) | ( n1189 & n1284 ) | ( n1204 & n1284 ) ;
  assign n1389 = ( n1300 & ~n1387 ) | ( n1300 & n1388 ) | ( ~n1387 & n1388 ) ;
  assign n1390 = ( n1300 & ~n1388 ) | ( n1300 & n1387 ) | ( ~n1388 & n1387 ) ;
  assign n1391 = ( n1389 & ~n1300 ) | ( n1389 & n1390 ) | ( ~n1300 & n1390 ) ;
  assign n1492 = ~n136 & x86 ;
  assign n1489 = ( x84 & ~n150 ) | ( x84 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n1490 = ( x85 & ~n131 ) | ( x85 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n1491 = n1489 | n1490 ;
  assign n1493 = ( x86 & ~n1492 ) | ( x86 & n1491 ) | ( ~n1492 & n1491 ) ;
  assign n1495 = ( x85 & x86 ) | ( x85 & n1294 ) | ( x86 & n1294 ) ;
  assign n1494 = ( x85 & ~x86 ) | ( x85 & n1294 ) | ( ~x86 & n1294 ) ;
  assign n1496 = ( x86 & ~n1495 ) | ( x86 & n1494 ) | ( ~n1495 & n1494 ) ;
  assign n1497 = ( n139 & ~n1493 ) | ( n139 & n1496 ) | ( ~n1493 & n1496 ) ;
  assign n1498 = ~n139 & n1497 ;
  assign n1499 = ( x2 & n1493 ) | ( x2 & n1498 ) | ( n1493 & n1498 ) ;
  assign n1500 = ( x2 & ~n1498 ) | ( x2 & n1493 ) | ( ~n1498 & n1493 ) ;
  assign n1501 = ( n1498 & ~n1499 ) | ( n1498 & n1500 ) | ( ~n1499 & n1500 ) ;
  assign n1392 = ( n1282 & ~n1374 ) | ( n1282 & n1384 ) | ( ~n1374 & n1384 ) ;
  assign n1406 = x78 &  n353 ;
  assign n1403 = ( x80 & ~n313 ) | ( x80 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n1404 = x79 &  n308 ;
  assign n1405 = n1403 | n1404 ;
  assign n1407 = ( x78 & ~n1406 ) | ( x78 & n1405 ) | ( ~n1406 & n1405 ) ;
  assign n1408 = ~n316 & n842 ;
  assign n1409 = n1407 | n1408 ;
  assign n1410 = ( x8 & ~n1409 ) | ( x8 & 1'b0 ) | ( ~n1409 & 1'b0 ) ;
  assign n1411 = ~x8 & n1409 ;
  assign n1412 = n1410 | n1411 ;
  assign n1473 = x75 &  n503 ;
  assign n1470 = ( x77 & ~n450 ) | ( x77 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n1471 = x76 &  n445 ;
  assign n1472 = n1470 | n1471 ;
  assign n1474 = ( x75 & ~n1473 ) | ( x75 & n1472 ) | ( ~n1473 & n1472 ) ;
  assign n1475 = ~n453 & n677 ;
  assign n1476 = n1474 | n1475 ;
  assign n1477 = ( x11 & ~n1476 ) | ( x11 & 1'b0 ) | ( ~n1476 & 1'b0 ) ;
  assign n1478 = ~x11 & n1476 ;
  assign n1479 = n1477 | n1478 ;
  assign n1416 = x72 &  n713 ;
  assign n1413 = ( x74 & ~n641 ) | ( x74 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n1414 = x73 &  n636 ;
  assign n1415 = n1413 | n1414 ;
  assign n1417 = ( x72 & ~n1416 ) | ( x72 & n1415 ) | ( ~n1416 & n1415 ) ;
  assign n1418 = ( n482 & ~n644 ) | ( n482 & 1'b0 ) | ( ~n644 & 1'b0 ) ;
  assign n1419 = n1417 | n1418 ;
  assign n1420 = ( x14 & ~n1419 ) | ( x14 & 1'b0 ) | ( ~n1419 & 1'b0 ) ;
  assign n1421 = ~x14 & n1419 ;
  assign n1422 = n1420 | n1421 ;
  assign n1426 = x69 &  n942 ;
  assign n1423 = ( x71 & ~n896 ) | ( x71 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n1424 = x70 &  n891 ;
  assign n1425 = n1423 | n1424 ;
  assign n1427 = ( x69 & ~n1426 ) | ( x69 & n1425 ) | ( ~n1426 & n1425 ) ;
  assign n1428 = ( n298 & ~n899 ) | ( n298 & 1'b0 ) | ( ~n899 & 1'b0 ) ;
  assign n1429 = n1427 | n1428 ;
  assign n1430 = ( x17 & ~n1429 ) | ( x17 & 1'b0 ) | ( ~n1429 & 1'b0 ) ;
  assign n1431 = ~x17 & n1429 ;
  assign n1432 = n1430 | n1431 ;
  assign n1436 = x66 &  n1227 ;
  assign n1433 = ( x68 & ~n1154 ) | ( x68 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n1434 = x67 &  n1149 ;
  assign n1435 = n1433 | n1434 ;
  assign n1437 = ( x66 & ~n1436 ) | ( x66 & n1435 ) | ( ~n1436 & n1435 ) ;
  assign n1438 = ( n1157 & ~n1437 ) | ( n1157 & n213 ) | ( ~n1437 & n213 ) ;
  assign n1439 = ~n1157 & n1438 ;
  assign n1440 = ( n1437 & ~x20 ) | ( n1437 & n1439 ) | ( ~x20 & n1439 ) ;
  assign n1441 = ( x20 & ~n1437 ) | ( x20 & n1439 ) | ( ~n1437 & n1439 ) ;
  assign n1442 = ( n1440 & ~n1439 ) | ( n1440 & n1441 ) | ( ~n1439 & n1441 ) ;
  assign n1443 = ( x23 & ~n1325 ) | ( x23 & 1'b0 ) | ( ~n1325 & 1'b0 ) ;
  assign n1444 = ( x21 & x22 ) | ( x21 & n1322 ) | ( x22 & n1322 ) ;
  assign n1445 = ( x21 & ~n1323 ) | ( x21 & x22 ) | ( ~n1323 & x22 ) ;
  assign n1446 = ~n1444 &  n1445 ;
  assign n1447 = x64 &  n1446 ;
  assign n1448 = ~x22 & x23 ;
  assign n1449 = ( x22 & ~x23 ) | ( x22 & 1'b0 ) | ( ~x23 & 1'b0 ) ;
  assign n1450 = n1448 | n1449 ;
  assign n1451 = ~n1324 |  n1450 ;
  assign n1452 = ( x65 & ~n1451 ) | ( x65 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n1453 = n1447 | n1452 ;
  assign n1454 = ~n1324 | ~n1450 ;
  assign n1455 = ( n142 & ~n1454 ) | ( n142 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n1456 = n1453 | n1455 ;
  assign n1458 = ( x23 & n1443 ) | ( x23 & n1456 ) | ( n1443 & n1456 ) ;
  assign n1457 = ( x23 & ~n1443 ) | ( x23 & n1456 ) | ( ~n1443 & n1456 ) ;
  assign n1459 = ( n1443 & ~n1458 ) | ( n1443 & n1457 ) | ( ~n1458 & n1457 ) ;
  assign n1461 = ( n1339 & n1442 ) | ( n1339 & n1459 ) | ( n1442 & n1459 ) ;
  assign n1460 = ( n1339 & ~n1442 ) | ( n1339 & n1459 ) | ( ~n1442 & n1459 ) ;
  assign n1462 = ( n1442 & ~n1461 ) | ( n1442 & n1460 ) | ( ~n1461 & n1460 ) ;
  assign n1464 = ( n1353 & n1432 ) | ( n1353 & n1462 ) | ( n1432 & n1462 ) ;
  assign n1463 = ( n1353 & ~n1432 ) | ( n1353 & n1462 ) | ( ~n1432 & n1462 ) ;
  assign n1465 = ( n1432 & ~n1464 ) | ( n1432 & n1463 ) | ( ~n1464 & n1463 ) ;
  assign n1466 = ( n1355 & ~n1354 ) | ( n1355 & n1365 ) | ( ~n1354 & n1365 ) ;
  assign n1467 = ( n1422 & n1465 ) | ( n1422 & n1466 ) | ( n1465 & n1466 ) ;
  assign n1468 = ( n1465 & ~n1422 ) | ( n1465 & n1466 ) | ( ~n1422 & n1466 ) ;
  assign n1469 = ( n1422 & ~n1467 ) | ( n1422 & n1468 ) | ( ~n1467 & n1468 ) ;
  assign n1480 = ( n1370 & ~n1479 ) | ( n1370 & n1469 ) | ( ~n1479 & n1469 ) ;
  assign n1481 = ( n1469 & ~n1370 ) | ( n1469 & n1479 ) | ( ~n1370 & n1479 ) ;
  assign n1482 = ( n1480 & ~n1469 ) | ( n1480 & n1481 ) | ( ~n1469 & n1481 ) ;
  assign n1484 = ( n1373 & n1412 ) | ( n1373 & n1482 ) | ( n1412 & n1482 ) ;
  assign n1483 = ( n1373 & ~n1412 ) | ( n1373 & n1482 ) | ( ~n1412 & n1482 ) ;
  assign n1485 = ( n1412 & ~n1484 ) | ( n1412 & n1483 ) | ( ~n1484 & n1483 ) ;
  assign n1396 = x81 &  n225 ;
  assign n1393 = ( x83 & ~n197 ) | ( x83 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n1394 = x82 &  n192 ;
  assign n1395 = n1393 | n1394 ;
  assign n1397 = ( x81 & ~n1396 ) | ( x81 & n1395 ) | ( ~n1396 & n1395 ) ;
  assign n1398 = ~n200 & n1100 ;
  assign n1399 = n1397 | n1398 ;
  assign n1400 = ( x5 & ~n1399 ) | ( x5 & 1'b0 ) | ( ~n1399 & 1'b0 ) ;
  assign n1401 = ~x5 & n1399 ;
  assign n1402 = n1400 | n1401 ;
  assign n1486 = ( n1392 & ~n1485 ) | ( n1392 & n1402 ) | ( ~n1485 & n1402 ) ;
  assign n1487 = ( n1392 & ~n1402 ) | ( n1392 & n1485 ) | ( ~n1402 & n1485 ) ;
  assign n1488 = ( n1486 & ~n1392 ) | ( n1486 & n1487 ) | ( ~n1392 & n1487 ) ;
  assign n1502 = ( n1389 & ~n1501 ) | ( n1389 & n1488 ) | ( ~n1501 & n1488 ) ;
  assign n1503 = ( n1488 & ~n1389 ) | ( n1488 & n1501 ) | ( ~n1389 & n1501 ) ;
  assign n1504 = ( n1502 & ~n1488 ) | ( n1502 & n1503 ) | ( ~n1488 & n1503 ) ;
  assign n1508 = ~n136 & x87 ;
  assign n1505 = ( x85 & ~n150 ) | ( x85 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n1506 = ( x86 & ~n131 ) | ( x86 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n1507 = n1505 | n1506 ;
  assign n1509 = ( x87 & ~n1508 ) | ( x87 & n1507 ) | ( ~n1508 & n1507 ) ;
  assign n1511 = ( x86 & x87 ) | ( x86 & n1495 ) | ( x87 & n1495 ) ;
  assign n1510 = ( x86 & ~x87 ) | ( x86 & n1495 ) | ( ~x87 & n1495 ) ;
  assign n1512 = ( x87 & ~n1511 ) | ( x87 & n1510 ) | ( ~n1511 & n1510 ) ;
  assign n1513 = ( n139 & ~n1509 ) | ( n139 & n1512 ) | ( ~n1509 & n1512 ) ;
  assign n1514 = ~n139 & n1513 ;
  assign n1515 = ( x2 & n1509 ) | ( x2 & n1514 ) | ( n1509 & n1514 ) ;
  assign n1516 = ( x2 & ~n1514 ) | ( x2 & n1509 ) | ( ~n1514 & n1509 ) ;
  assign n1517 = ( n1514 & ~n1515 ) | ( n1514 & n1516 ) | ( ~n1515 & n1516 ) ;
  assign n1518 = ( n1392 & n1402 ) | ( n1392 & n1485 ) | ( n1402 & n1485 ) ;
  assign n1522 = x82 &  n225 ;
  assign n1519 = ( x84 & ~n197 ) | ( x84 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n1520 = x83 &  n192 ;
  assign n1521 = n1519 | n1520 ;
  assign n1523 = ( x82 & ~n1522 ) | ( x82 & n1521 ) | ( ~n1522 & n1521 ) ;
  assign n1524 = ~n200 & n1199 ;
  assign n1525 = n1523 | n1524 ;
  assign n1526 = ( x5 & ~n1525 ) | ( x5 & 1'b0 ) | ( ~n1525 & 1'b0 ) ;
  assign n1527 = ~x5 & n1525 ;
  assign n1528 = n1526 | n1527 ;
  assign n1532 = x79 &  n353 ;
  assign n1529 = ( x81 & ~n313 ) | ( x81 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n1530 = x80 &  n308 ;
  assign n1531 = n1529 | n1530 ;
  assign n1533 = ( x79 & ~n1532 ) | ( x79 & n1531 ) | ( ~n1532 & n1531 ) ;
  assign n1534 = ~n316 & n994 ;
  assign n1535 = n1533 | n1534 ;
  assign n1536 = ( x8 & ~n1535 ) | ( x8 & 1'b0 ) | ( ~n1535 & 1'b0 ) ;
  assign n1537 = ~x8 & n1535 ;
  assign n1538 = n1536 | n1537 ;
  assign n1542 = x73 &  n713 ;
  assign n1539 = ( x75 & ~n641 ) | ( x75 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n1540 = x74 &  n636 ;
  assign n1541 = n1539 | n1540 ;
  assign n1543 = ( x73 & ~n1542 ) | ( x73 & n1541 ) | ( ~n1542 & n1541 ) ;
  assign n1544 = ( n540 & ~n644 ) | ( n540 & 1'b0 ) | ( ~n644 & 1'b0 ) ;
  assign n1545 = n1543 | n1544 ;
  assign n1546 = ( x14 & ~n1545 ) | ( x14 & 1'b0 ) | ( ~n1545 & 1'b0 ) ;
  assign n1547 = ~x14 & n1545 ;
  assign n1548 = n1546 | n1547 ;
  assign n1567 = x67 &  n1227 ;
  assign n1564 = ( x69 & ~n1154 ) | ( x69 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n1565 = x68 &  n1149 ;
  assign n1566 = n1564 | n1565 ;
  assign n1568 = ( x67 & ~n1567 ) | ( x67 & n1566 ) | ( ~n1567 & n1566 ) ;
  assign n1569 = ( n246 & ~n1157 ) | ( n246 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n1570 = n1568 | n1569 ;
  assign n1571 = ( x20 & ~n1570 ) | ( x20 & 1'b0 ) | ( ~n1570 & 1'b0 ) ;
  assign n1572 = ~x20 & n1570 ;
  assign n1573 = n1571 | n1572 ;
  assign n1550 = ( x21 & ~x22 ) | ( x21 & n1450 ) | ( ~x22 & n1450 ) ;
  assign n1549 = ( x21 & ~x22 ) | ( x21 & n1324 ) | ( ~x22 & n1324 ) ;
  assign n1551 = ~n1550 |  n1549 ;
  assign n1555 = x64 &  n1551 ;
  assign n1552 = ( x66 & ~n1451 ) | ( x66 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n1553 = x65 &  n1446 ;
  assign n1554 = n1552 | n1553 ;
  assign n1556 = ( x64 & ~n1555 ) | ( x64 & n1554 ) | ( ~n1555 & n1554 ) ;
  assign n1557 = ( n157 & ~n1454 ) | ( n157 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n1558 = n1556 | n1557 ;
  assign n1559 = ( x23 & ~n1325 ) | ( x23 & n1456 ) | ( ~n1325 & n1456 ) ;
  assign n1560 = ~n1456 & n1559 ;
  assign n1561 = ( n1558 & ~x23 ) | ( n1558 & n1560 ) | ( ~x23 & n1560 ) ;
  assign n1562 = ( x23 & ~n1558 ) | ( x23 & n1560 ) | ( ~n1558 & n1560 ) ;
  assign n1563 = ( n1561 & ~n1560 ) | ( n1561 & n1562 ) | ( ~n1560 & n1562 ) ;
  assign n1574 = ( n1461 & ~n1573 ) | ( n1461 & n1563 ) | ( ~n1573 & n1563 ) ;
  assign n1575 = ( n1563 & ~n1461 ) | ( n1563 & n1573 ) | ( ~n1461 & n1573 ) ;
  assign n1576 = ( n1574 & ~n1563 ) | ( n1574 & n1575 ) | ( ~n1563 & n1575 ) ;
  assign n1580 = x70 &  n942 ;
  assign n1577 = ( x72 & ~n896 ) | ( x72 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n1578 = x71 &  n891 ;
  assign n1579 = n1577 | n1578 ;
  assign n1581 = ( x70 & ~n1580 ) | ( x70 & n1579 ) | ( ~n1580 & n1579 ) ;
  assign n1582 = ( n345 & ~n899 ) | ( n345 & 1'b0 ) | ( ~n899 & 1'b0 ) ;
  assign n1583 = n1581 | n1582 ;
  assign n1584 = ( x17 & ~n1583 ) | ( x17 & 1'b0 ) | ( ~n1583 & 1'b0 ) ;
  assign n1585 = ~x17 & n1583 ;
  assign n1586 = n1584 | n1585 ;
  assign n1587 = ( n1576 & ~n1464 ) | ( n1576 & n1586 ) | ( ~n1464 & n1586 ) ;
  assign n1588 = ( n1464 & ~n1586 ) | ( n1464 & n1576 ) | ( ~n1586 & n1576 ) ;
  assign n1589 = ( n1587 & ~n1576 ) | ( n1587 & n1588 ) | ( ~n1576 & n1588 ) ;
  assign n1591 = ( n1467 & n1548 ) | ( n1467 & n1589 ) | ( n1548 & n1589 ) ;
  assign n1590 = ( n1467 & ~n1548 ) | ( n1467 & n1589 ) | ( ~n1548 & n1589 ) ;
  assign n1592 = ( n1548 & ~n1591 ) | ( n1548 & n1590 ) | ( ~n1591 & n1590 ) ;
  assign n1603 = ( n1370 & n1469 ) | ( n1370 & n1479 ) | ( n1469 & n1479 ) ;
  assign n1596 = x76 &  n503 ;
  assign n1593 = ( x78 & ~n450 ) | ( x78 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n1594 = x77 &  n445 ;
  assign n1595 = n1593 | n1594 ;
  assign n1597 = ( x76 & ~n1596 ) | ( x76 & n1595 ) | ( ~n1596 & n1595 ) ;
  assign n1598 = ~n453 & n693 ;
  assign n1599 = n1597 | n1598 ;
  assign n1600 = ( x11 & ~n1599 ) | ( x11 & 1'b0 ) | ( ~n1599 & 1'b0 ) ;
  assign n1601 = ~x11 & n1599 ;
  assign n1602 = n1600 | n1601 ;
  assign n1604 = ( n1592 & ~n1603 ) | ( n1592 & n1602 ) | ( ~n1603 & n1602 ) ;
  assign n1605 = ( n1592 & ~n1602 ) | ( n1592 & n1603 ) | ( ~n1602 & n1603 ) ;
  assign n1606 = ( n1604 & ~n1592 ) | ( n1604 & n1605 ) | ( ~n1592 & n1605 ) ;
  assign n1608 = ( n1484 & n1538 ) | ( n1484 & n1606 ) | ( n1538 & n1606 ) ;
  assign n1607 = ( n1484 & ~n1538 ) | ( n1484 & n1606 ) | ( ~n1538 & n1606 ) ;
  assign n1609 = ( n1538 & ~n1608 ) | ( n1538 & n1607 ) | ( ~n1608 & n1607 ) ;
  assign n1610 = ( n1518 & n1528 ) | ( n1518 & n1609 ) | ( n1528 & n1609 ) ;
  assign n1611 = ( n1528 & ~n1518 ) | ( n1528 & n1609 ) | ( ~n1518 & n1609 ) ;
  assign n1612 = ( n1518 & ~n1610 ) | ( n1518 & n1611 ) | ( ~n1610 & n1611 ) ;
  assign n1613 = ( n1389 & n1488 ) | ( n1389 & n1501 ) | ( n1488 & n1501 ) ;
  assign n1614 = ( n1517 & n1612 ) | ( n1517 & n1613 ) | ( n1612 & n1613 ) ;
  assign n1615 = ( n1612 & ~n1517 ) | ( n1612 & n1613 ) | ( ~n1517 & n1613 ) ;
  assign n1616 = ( n1517 & ~n1614 ) | ( n1517 & n1615 ) | ( ~n1614 & n1615 ) ;
  assign n1620 = ~n136 & x88 ;
  assign n1617 = ( x86 & ~n150 ) | ( x86 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n1618 = ( x87 & ~n131 ) | ( x87 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n1619 = n1617 | n1618 ;
  assign n1621 = ( x88 & ~n1620 ) | ( x88 & n1619 ) | ( ~n1620 & n1619 ) ;
  assign n1623 = ( x87 & x88 ) | ( x87 & n1511 ) | ( x88 & n1511 ) ;
  assign n1622 = ( x87 & ~x88 ) | ( x87 & n1511 ) | ( ~x88 & n1511 ) ;
  assign n1624 = ( x88 & ~n1623 ) | ( x88 & n1622 ) | ( ~n1623 & n1622 ) ;
  assign n1625 = ( n139 & ~n1621 ) | ( n139 & n1624 ) | ( ~n1621 & n1624 ) ;
  assign n1626 = ~n139 & n1625 ;
  assign n1627 = ( x2 & n1621 ) | ( x2 & n1626 ) | ( n1621 & n1626 ) ;
  assign n1628 = ( x2 & ~n1626 ) | ( x2 & n1621 ) | ( ~n1626 & n1621 ) ;
  assign n1629 = ( n1626 & ~n1627 ) | ( n1626 & n1628 ) | ( ~n1627 & n1628 ) ;
  assign n1643 = x74 &  n713 ;
  assign n1640 = ( x76 & ~n641 ) | ( x76 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n1641 = x75 &  n636 ;
  assign n1642 = n1640 | n1641 ;
  assign n1644 = ( x74 & ~n1643 ) | ( x74 & n1642 ) | ( ~n1643 & n1642 ) ;
  assign n1645 = ( n603 & ~n644 ) | ( n603 & 1'b0 ) | ( ~n644 & 1'b0 ) ;
  assign n1646 = n1644 | n1645 ;
  assign n1647 = ( x14 & ~n1646 ) | ( x14 & 1'b0 ) | ( ~n1646 & 1'b0 ) ;
  assign n1648 = ~x14 & n1646 ;
  assign n1649 = n1647 | n1648 ;
  assign n1650 = ( x23 & ~x24 ) | ( x23 & 1'b0 ) | ( ~x24 & 1'b0 ) ;
  assign n1651 = ~x23 & x24 ;
  assign n1652 = n1650 | n1651 ;
  assign n1653 = x64 &  n1652 ;
  assign n1654 = ( n1325 & ~n1456 ) | ( n1325 & n1558 ) | ( ~n1456 & n1558 ) ;
  assign n1655 = ( x23 & n1456 ) | ( x23 & n1654 ) | ( n1456 & n1654 ) ;
  assign n1656 = ( x23 & ~n1655 ) | ( x23 & 1'b0 ) | ( ~n1655 & 1'b0 ) ;
  assign n1660 = x65 &  n1551 ;
  assign n1657 = ( x67 & ~n1451 ) | ( x67 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n1658 = x66 &  n1446 ;
  assign n1659 = n1657 | n1658 ;
  assign n1661 = ( x65 & ~n1660 ) | ( x65 & n1659 ) | ( ~n1660 & n1659 ) ;
  assign n1662 = n173 | n1454 ;
  assign n1663 = ~n1661 & n1662 ;
  assign n1664 = x23 &  n1663 ;
  assign n1665 = x23 | n1663 ;
  assign n1666 = ~n1664 & n1665 ;
  assign n1667 = ( n1653 & ~n1656 ) | ( n1653 & n1666 ) | ( ~n1656 & n1666 ) ;
  assign n1668 = ( n1653 & ~n1666 ) | ( n1653 & n1656 ) | ( ~n1666 & n1656 ) ;
  assign n1669 = ( n1667 & ~n1653 ) | ( n1667 & n1668 ) | ( ~n1653 & n1668 ) ;
  assign n1670 = ( n1461 & n1563 ) | ( n1461 & n1573 ) | ( n1563 & n1573 ) ;
  assign n1674 = x68 &  n1227 ;
  assign n1671 = ( x70 & ~n1154 ) | ( x70 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n1672 = x69 &  n1149 ;
  assign n1673 = n1671 | n1672 ;
  assign n1675 = ( x68 & ~n1674 ) | ( x68 & n1673 ) | ( ~n1674 & n1673 ) ;
  assign n1676 = ( n282 & ~n1157 ) | ( n282 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n1677 = n1675 | n1676 ;
  assign n1678 = ( x20 & ~n1677 ) | ( x20 & 1'b0 ) | ( ~n1677 & 1'b0 ) ;
  assign n1679 = ~x20 & n1677 ;
  assign n1680 = n1678 | n1679 ;
  assign n1681 = ( n1669 & ~n1670 ) | ( n1669 & n1680 ) | ( ~n1670 & n1680 ) ;
  assign n1682 = ( n1670 & ~n1669 ) | ( n1670 & n1680 ) | ( ~n1669 & n1680 ) ;
  assign n1683 = ( n1681 & ~n1680 ) | ( n1681 & n1682 ) | ( ~n1680 & n1682 ) ;
  assign n1688 = x71 &  n942 ;
  assign n1685 = ( x73 & ~n896 ) | ( x73 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n1686 = x72 &  n891 ;
  assign n1687 = n1685 | n1686 ;
  assign n1689 = ( x71 & ~n1688 ) | ( x71 & n1687 ) | ( ~n1688 & n1687 ) ;
  assign n1690 = ( n389 & ~n899 ) | ( n389 & 1'b0 ) | ( ~n899 & 1'b0 ) ;
  assign n1691 = n1689 | n1690 ;
  assign n1692 = ( x17 & ~n1691 ) | ( x17 & 1'b0 ) | ( ~n1691 & 1'b0 ) ;
  assign n1693 = ~x17 & n1691 ;
  assign n1694 = n1692 | n1693 ;
  assign n1684 = ( n1464 & n1576 ) | ( n1464 & n1586 ) | ( n1576 & n1586 ) ;
  assign n1695 = ( n1683 & ~n1694 ) | ( n1683 & n1684 ) | ( ~n1694 & n1684 ) ;
  assign n1696 = ( n1683 & ~n1684 ) | ( n1683 & n1694 ) | ( ~n1684 & n1694 ) ;
  assign n1697 = ( n1695 & ~n1683 ) | ( n1695 & n1696 ) | ( ~n1683 & n1696 ) ;
  assign n1698 = ( n1649 & ~n1591 ) | ( n1649 & n1697 ) | ( ~n1591 & n1697 ) ;
  assign n1699 = ( n1591 & ~n1697 ) | ( n1591 & n1649 ) | ( ~n1697 & n1649 ) ;
  assign n1700 = ( n1698 & ~n1649 ) | ( n1698 & n1699 ) | ( ~n1649 & n1699 ) ;
  assign n1704 = x77 &  n503 ;
  assign n1701 = ( x79 & ~n450 ) | ( x79 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n1702 = x78 &  n445 ;
  assign n1703 = n1701 | n1702 ;
  assign n1705 = ( x77 & ~n1704 ) | ( x77 & n1703 ) | ( ~n1704 & n1703 ) ;
  assign n1706 = ~n453 & n766 ;
  assign n1707 = n1705 | n1706 ;
  assign n1708 = ( x11 & ~n1707 ) | ( x11 & 1'b0 ) | ( ~n1707 & 1'b0 ) ;
  assign n1709 = ~x11 & n1707 ;
  assign n1710 = n1708 | n1709 ;
  assign n1711 = ( n1592 & n1602 ) | ( n1592 & n1603 ) | ( n1602 & n1603 ) ;
  assign n1712 = ( n1700 & ~n1710 ) | ( n1700 & n1711 ) | ( ~n1710 & n1711 ) ;
  assign n1713 = ( n1700 & ~n1711 ) | ( n1700 & n1710 ) | ( ~n1711 & n1710 ) ;
  assign n1714 = ( n1712 & ~n1700 ) | ( n1712 & n1713 ) | ( ~n1700 & n1713 ) ;
  assign n1718 = x80 &  n353 ;
  assign n1715 = ( x82 & ~n313 ) | ( x82 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n1716 = x81 &  n308 ;
  assign n1717 = n1715 | n1716 ;
  assign n1719 = ( x80 & ~n1718 ) | ( x80 & n1717 ) | ( ~n1718 & n1717 ) ;
  assign n1720 = ~n316 & n1084 ;
  assign n1721 = n1719 | n1720 ;
  assign n1722 = ( x8 & ~n1721 ) | ( x8 & 1'b0 ) | ( ~n1721 & 1'b0 ) ;
  assign n1723 = ~x8 & n1721 ;
  assign n1724 = n1722 | n1723 ;
  assign n1725 = ( n1714 & ~n1608 ) | ( n1714 & n1724 ) | ( ~n1608 & n1724 ) ;
  assign n1726 = ( n1608 & ~n1724 ) | ( n1608 & n1714 ) | ( ~n1724 & n1714 ) ;
  assign n1727 = ( n1725 & ~n1714 ) | ( n1725 & n1726 ) | ( ~n1714 & n1726 ) ;
  assign n1633 = x83 &  n225 ;
  assign n1630 = ( x85 & ~n197 ) | ( x85 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n1631 = x84 &  n192 ;
  assign n1632 = n1630 | n1631 ;
  assign n1634 = ( x83 & ~n1633 ) | ( x83 & n1632 ) | ( ~n1633 & n1632 ) ;
  assign n1635 = ~n200 & n1295 ;
  assign n1636 = n1634 | n1635 ;
  assign n1637 = ( x5 & ~n1636 ) | ( x5 & 1'b0 ) | ( ~n1636 & 1'b0 ) ;
  assign n1638 = ~x5 & n1636 ;
  assign n1639 = n1637 | n1638 ;
  assign n1729 = ( n1610 & n1639 ) | ( n1610 & n1727 ) | ( n1639 & n1727 ) ;
  assign n1728 = ( n1610 & ~n1727 ) | ( n1610 & n1639 ) | ( ~n1727 & n1639 ) ;
  assign n1730 = ( n1727 & ~n1729 ) | ( n1727 & n1728 ) | ( ~n1729 & n1728 ) ;
  assign n1731 = ( n1614 & n1629 ) | ( n1614 & n1730 ) | ( n1629 & n1730 ) ;
  assign n1732 = ( n1614 & ~n1629 ) | ( n1614 & n1730 ) | ( ~n1629 & n1730 ) ;
  assign n1733 = ( n1629 & ~n1731 ) | ( n1629 & n1732 ) | ( ~n1731 & n1732 ) ;
  assign n1737 = ~n136 & x89 ;
  assign n1734 = ( x87 & ~n150 ) | ( x87 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n1735 = ( x88 & ~n131 ) | ( x88 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n1736 = n1734 | n1735 ;
  assign n1738 = ( x89 & ~n1737 ) | ( x89 & n1736 ) | ( ~n1737 & n1736 ) ;
  assign n1740 = ( x88 & x89 ) | ( x88 & n1623 ) | ( x89 & n1623 ) ;
  assign n1739 = ( x88 & ~x89 ) | ( x88 & n1623 ) | ( ~x89 & n1623 ) ;
  assign n1741 = ( x89 & ~n1740 ) | ( x89 & n1739 ) | ( ~n1740 & n1739 ) ;
  assign n1742 = ( n139 & ~n1738 ) | ( n139 & n1741 ) | ( ~n1738 & n1741 ) ;
  assign n1743 = ~n139 & n1742 ;
  assign n1744 = ( x2 & n1738 ) | ( x2 & n1743 ) | ( n1738 & n1743 ) ;
  assign n1745 = ( x2 & ~n1743 ) | ( x2 & n1738 ) | ( ~n1743 & n1738 ) ;
  assign n1746 = ( n1743 & ~n1744 ) | ( n1743 & n1745 ) | ( ~n1744 & n1745 ) ;
  assign n1747 = ( n1614 & ~n1730 ) | ( n1614 & n1629 ) | ( ~n1730 & n1629 ) ;
  assign n1751 = x84 &  n225 ;
  assign n1748 = ( x86 & ~n197 ) | ( x86 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n1749 = x85 &  n192 ;
  assign n1750 = n1748 | n1749 ;
  assign n1752 = ( x84 & ~n1751 ) | ( x84 & n1750 ) | ( ~n1751 & n1750 ) ;
  assign n1753 = ~n200 & n1496 ;
  assign n1754 = n1752 | n1753 ;
  assign n1755 = ( x5 & ~n1754 ) | ( x5 & 1'b0 ) | ( ~n1754 & 1'b0 ) ;
  assign n1756 = ~x5 & n1754 ;
  assign n1757 = n1755 | n1756 ;
  assign n1761 = x81 &  n353 ;
  assign n1758 = ( x83 & ~n313 ) | ( x83 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n1759 = x82 &  n308 ;
  assign n1760 = n1758 | n1759 ;
  assign n1762 = ( x81 & ~n1761 ) | ( x81 & n1760 ) | ( ~n1761 & n1760 ) ;
  assign n1763 = ~n316 & n1100 ;
  assign n1764 = n1762 | n1763 ;
  assign n1765 = ( x8 & ~n1764 ) | ( x8 & 1'b0 ) | ( ~n1764 & 1'b0 ) ;
  assign n1766 = ~x8 & n1764 ;
  assign n1767 = n1765 | n1766 ;
  assign n1771 = x75 &  n713 ;
  assign n1768 = ( x77 & ~n641 ) | ( x77 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n1769 = x76 &  n636 ;
  assign n1770 = n1768 | n1769 ;
  assign n1772 = ( x75 & ~n1771 ) | ( x75 & n1770 ) | ( ~n1771 & n1770 ) ;
  assign n1773 = ~n644 & n677 ;
  assign n1774 = n1772 | n1773 ;
  assign n1775 = ( x14 & ~n1774 ) | ( x14 & 1'b0 ) | ( ~n1774 & 1'b0 ) ;
  assign n1776 = ~x14 & n1774 ;
  assign n1777 = n1775 | n1776 ;
  assign n1781 = x72 &  n942 ;
  assign n1778 = ( x74 & ~n896 ) | ( x74 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n1779 = x73 &  n891 ;
  assign n1780 = n1778 | n1779 ;
  assign n1782 = ( x72 & ~n1781 ) | ( x72 & n1780 ) | ( ~n1781 & n1780 ) ;
  assign n1783 = ( n482 & ~n899 ) | ( n482 & 1'b0 ) | ( ~n899 & 1'b0 ) ;
  assign n1784 = n1782 | n1783 ;
  assign n1785 = ( x17 & ~n1784 ) | ( x17 & 1'b0 ) | ( ~n1784 & 1'b0 ) ;
  assign n1786 = ~x17 & n1784 ;
  assign n1787 = n1785 | n1786 ;
  assign n1791 = x69 &  n1227 ;
  assign n1788 = ( x71 & ~n1154 ) | ( x71 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n1789 = x70 &  n1149 ;
  assign n1790 = n1788 | n1789 ;
  assign n1792 = ( x69 & ~n1791 ) | ( x69 & n1790 ) | ( ~n1791 & n1790 ) ;
  assign n1793 = ( n298 & ~n1157 ) | ( n298 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n1794 = n1792 | n1793 ;
  assign n1795 = ( x20 & ~n1794 ) | ( x20 & 1'b0 ) | ( ~n1794 & 1'b0 ) ;
  assign n1796 = ~x20 & n1794 ;
  assign n1797 = n1795 | n1796 ;
  assign n1801 = x66 &  n1551 ;
  assign n1798 = ( x68 & ~n1451 ) | ( x68 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n1799 = x67 &  n1446 ;
  assign n1800 = n1798 | n1799 ;
  assign n1802 = ( x66 & ~n1801 ) | ( x66 & n1800 ) | ( ~n1801 & n1800 ) ;
  assign n1803 = ( n1454 & ~n1802 ) | ( n1454 & n213 ) | ( ~n1802 & n213 ) ;
  assign n1804 = ~n1454 & n1803 ;
  assign n1805 = ( n1802 & ~x23 ) | ( n1802 & n1804 ) | ( ~x23 & n1804 ) ;
  assign n1806 = ( x23 & ~n1802 ) | ( x23 & n1804 ) | ( ~n1802 & n1804 ) ;
  assign n1807 = ( n1805 & ~n1804 ) | ( n1805 & n1806 ) | ( ~n1804 & n1806 ) ;
  assign n1808 = ( x26 & ~n1653 ) | ( x26 & 1'b0 ) | ( ~n1653 & 1'b0 ) ;
  assign n1809 = ( x24 & x25 ) | ( x24 & n1650 ) | ( x25 & n1650 ) ;
  assign n1810 = ( x24 & ~n1651 ) | ( x24 & x25 ) | ( ~n1651 & x25 ) ;
  assign n1811 = ~n1809 &  n1810 ;
  assign n1812 = x64 &  n1811 ;
  assign n1813 = ~x25 & x26 ;
  assign n1814 = ( x25 & ~x26 ) | ( x25 & 1'b0 ) | ( ~x26 & 1'b0 ) ;
  assign n1815 = n1813 | n1814 ;
  assign n1816 = ~n1652 |  n1815 ;
  assign n1817 = ( x65 & ~n1816 ) | ( x65 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n1818 = n1812 | n1817 ;
  assign n1819 = ~n1652 | ~n1815 ;
  assign n1820 = ( n142 & ~n1819 ) | ( n142 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n1821 = n1818 | n1820 ;
  assign n1823 = ( x26 & n1808 ) | ( x26 & n1821 ) | ( n1808 & n1821 ) ;
  assign n1822 = ( x26 & ~n1808 ) | ( x26 & n1821 ) | ( ~n1808 & n1821 ) ;
  assign n1824 = ( n1808 & ~n1823 ) | ( n1808 & n1822 ) | ( ~n1823 & n1822 ) ;
  assign n1826 = ( n1668 & n1807 ) | ( n1668 & n1824 ) | ( n1807 & n1824 ) ;
  assign n1825 = ( n1668 & ~n1807 ) | ( n1668 & n1824 ) | ( ~n1807 & n1824 ) ;
  assign n1827 = ( n1807 & ~n1826 ) | ( n1807 & n1825 ) | ( ~n1826 & n1825 ) ;
  assign n1829 = ( n1682 & n1797 ) | ( n1682 & n1827 ) | ( n1797 & n1827 ) ;
  assign n1828 = ( n1682 & ~n1797 ) | ( n1682 & n1827 ) | ( ~n1797 & n1827 ) ;
  assign n1830 = ( n1797 & ~n1829 ) | ( n1797 & n1828 ) | ( ~n1829 & n1828 ) ;
  assign n1831 = ( n1684 & ~n1683 ) | ( n1684 & n1694 ) | ( ~n1683 & n1694 ) ;
  assign n1832 = ( n1787 & n1830 ) | ( n1787 & n1831 ) | ( n1830 & n1831 ) ;
  assign n1833 = ( n1830 & ~n1787 ) | ( n1830 & n1831 ) | ( ~n1787 & n1831 ) ;
  assign n1834 = ( n1787 & ~n1832 ) | ( n1787 & n1833 ) | ( ~n1832 & n1833 ) ;
  assign n1835 = ( n1699 & n1777 ) | ( n1699 & n1834 ) | ( n1777 & n1834 ) ;
  assign n1836 = ( n1699 & ~n1777 ) | ( n1699 & n1834 ) | ( ~n1777 & n1834 ) ;
  assign n1837 = ( n1777 & ~n1835 ) | ( n1777 & n1836 ) | ( ~n1835 & n1836 ) ;
  assign n1848 = ( n1710 & ~n1700 ) | ( n1710 & n1711 ) | ( ~n1700 & n1711 ) ;
  assign n1841 = x78 &  n503 ;
  assign n1838 = ( x80 & ~n450 ) | ( x80 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n1839 = x79 &  n445 ;
  assign n1840 = n1838 | n1839 ;
  assign n1842 = ( x78 & ~n1841 ) | ( x78 & n1840 ) | ( ~n1841 & n1840 ) ;
  assign n1843 = ~n453 & n842 ;
  assign n1844 = n1842 | n1843 ;
  assign n1845 = ( x11 & ~n1844 ) | ( x11 & 1'b0 ) | ( ~n1844 & 1'b0 ) ;
  assign n1846 = ~x11 & n1844 ;
  assign n1847 = n1845 | n1846 ;
  assign n1849 = ( n1837 & ~n1848 ) | ( n1837 & n1847 ) | ( ~n1848 & n1847 ) ;
  assign n1850 = ( n1837 & ~n1847 ) | ( n1837 & n1848 ) | ( ~n1847 & n1848 ) ;
  assign n1851 = ( n1849 & ~n1837 ) | ( n1849 & n1850 ) | ( ~n1837 & n1850 ) ;
  assign n1852 = ( n1608 & ~n1714 ) | ( n1608 & n1724 ) | ( ~n1714 & n1724 ) ;
  assign n1853 = ( n1767 & n1851 ) | ( n1767 & n1852 ) | ( n1851 & n1852 ) ;
  assign n1854 = ( n1851 & ~n1767 ) | ( n1851 & n1852 ) | ( ~n1767 & n1852 ) ;
  assign n1855 = ( n1767 & ~n1853 ) | ( n1767 & n1854 ) | ( ~n1853 & n1854 ) ;
  assign n1856 = ( n1728 & n1757 ) | ( n1728 & n1855 ) | ( n1757 & n1855 ) ;
  assign n1857 = ( n1757 & ~n1728 ) | ( n1757 & n1855 ) | ( ~n1728 & n1855 ) ;
  assign n1858 = ( n1728 & ~n1856 ) | ( n1728 & n1857 ) | ( ~n1856 & n1857 ) ;
  assign n1860 = ( n1746 & n1747 ) | ( n1746 & n1858 ) | ( n1747 & n1858 ) ;
  assign n1859 = ( n1747 & ~n1746 ) | ( n1747 & n1858 ) | ( ~n1746 & n1858 ) ;
  assign n1861 = ( n1746 & ~n1860 ) | ( n1746 & n1859 ) | ( ~n1860 & n1859 ) ;
  assign n1875 = x82 &  n353 ;
  assign n1872 = ( x84 & ~n313 ) | ( x84 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n1873 = x83 &  n308 ;
  assign n1874 = n1872 | n1873 ;
  assign n1876 = ( x82 & ~n1875 ) | ( x82 & n1874 ) | ( ~n1875 & n1874 ) ;
  assign n1877 = ~n316 & n1199 ;
  assign n1878 = n1876 | n1877 ;
  assign n1879 = ( x8 & ~n1878 ) | ( x8 & 1'b0 ) | ( ~n1878 & 1'b0 ) ;
  assign n1880 = ~x8 & n1878 ;
  assign n1881 = n1879 | n1880 ;
  assign n1939 = x76 &  n713 ;
  assign n1936 = ( x78 & ~n641 ) | ( x78 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n1937 = x77 &  n636 ;
  assign n1938 = n1936 | n1937 ;
  assign n1940 = ( x76 & ~n1939 ) | ( x76 & n1938 ) | ( ~n1939 & n1938 ) ;
  assign n1941 = ~n644 & n693 ;
  assign n1942 = n1940 | n1941 ;
  assign n1943 = ( x14 & ~n1942 ) | ( x14 & 1'b0 ) | ( ~n1942 & 1'b0 ) ;
  assign n1944 = ~x14 & n1942 ;
  assign n1945 = n1943 | n1944 ;
  assign n1885 = x73 &  n942 ;
  assign n1882 = ( x75 & ~n896 ) | ( x75 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n1883 = x74 &  n891 ;
  assign n1884 = n1882 | n1883 ;
  assign n1886 = ( x73 & ~n1885 ) | ( x73 & n1884 ) | ( ~n1885 & n1884 ) ;
  assign n1887 = ( n540 & ~n899 ) | ( n540 & 1'b0 ) | ( ~n899 & 1'b0 ) ;
  assign n1888 = n1886 | n1887 ;
  assign n1889 = ( x17 & ~n1888 ) | ( x17 & 1'b0 ) | ( ~n1888 & 1'b0 ) ;
  assign n1890 = ~x17 & n1888 ;
  assign n1891 = n1889 | n1890 ;
  assign n1910 = x67 &  n1551 ;
  assign n1907 = ( x69 & ~n1451 ) | ( x69 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n1908 = x68 &  n1446 ;
  assign n1909 = n1907 | n1908 ;
  assign n1911 = ( x67 & ~n1910 ) | ( x67 & n1909 ) | ( ~n1910 & n1909 ) ;
  assign n1912 = ( n246 & ~n1454 ) | ( n246 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n1913 = n1911 | n1912 ;
  assign n1914 = ( x23 & ~n1913 ) | ( x23 & 1'b0 ) | ( ~n1913 & 1'b0 ) ;
  assign n1915 = ~x23 & n1913 ;
  assign n1916 = n1914 | n1915 ;
  assign n1893 = ( x24 & ~x25 ) | ( x24 & n1815 ) | ( ~x25 & n1815 ) ;
  assign n1892 = ( x24 & ~x25 ) | ( x24 & n1652 ) | ( ~x25 & n1652 ) ;
  assign n1894 = ~n1893 |  n1892 ;
  assign n1898 = x64 &  n1894 ;
  assign n1895 = ( x66 & ~n1816 ) | ( x66 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n1896 = x65 &  n1811 ;
  assign n1897 = n1895 | n1896 ;
  assign n1899 = ( x64 & ~n1898 ) | ( x64 & n1897 ) | ( ~n1898 & n1897 ) ;
  assign n1900 = ( n157 & ~n1819 ) | ( n157 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n1901 = n1899 | n1900 ;
  assign n1902 = ( x26 & ~n1653 ) | ( x26 & n1821 ) | ( ~n1653 & n1821 ) ;
  assign n1903 = ~n1821 & n1902 ;
  assign n1904 = ( n1901 & ~x26 ) | ( n1901 & n1903 ) | ( ~x26 & n1903 ) ;
  assign n1905 = ( x26 & ~n1901 ) | ( x26 & n1903 ) | ( ~n1901 & n1903 ) ;
  assign n1906 = ( n1904 & ~n1903 ) | ( n1904 & n1905 ) | ( ~n1903 & n1905 ) ;
  assign n1917 = ( n1826 & ~n1916 ) | ( n1826 & n1906 ) | ( ~n1916 & n1906 ) ;
  assign n1918 = ( n1906 & ~n1826 ) | ( n1906 & n1916 ) | ( ~n1826 & n1916 ) ;
  assign n1919 = ( n1917 & ~n1906 ) | ( n1917 & n1918 ) | ( ~n1906 & n1918 ) ;
  assign n1923 = x70 &  n1227 ;
  assign n1920 = ( x72 & ~n1154 ) | ( x72 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n1921 = x71 &  n1149 ;
  assign n1922 = n1920 | n1921 ;
  assign n1924 = ( x70 & ~n1923 ) | ( x70 & n1922 ) | ( ~n1923 & n1922 ) ;
  assign n1925 = ( n345 & ~n1157 ) | ( n345 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n1926 = n1924 | n1925 ;
  assign n1927 = ( x20 & ~n1926 ) | ( x20 & 1'b0 ) | ( ~n1926 & 1'b0 ) ;
  assign n1928 = ~x20 & n1926 ;
  assign n1929 = n1927 | n1928 ;
  assign n1930 = ( n1919 & ~n1829 ) | ( n1919 & n1929 ) | ( ~n1829 & n1929 ) ;
  assign n1931 = ( n1829 & ~n1929 ) | ( n1829 & n1919 ) | ( ~n1929 & n1919 ) ;
  assign n1932 = ( n1930 & ~n1919 ) | ( n1930 & n1931 ) | ( ~n1919 & n1931 ) ;
  assign n1934 = ( n1832 & n1891 ) | ( n1832 & n1932 ) | ( n1891 & n1932 ) ;
  assign n1933 = ( n1832 & ~n1891 ) | ( n1832 & n1932 ) | ( ~n1891 & n1932 ) ;
  assign n1935 = ( n1891 & ~n1934 ) | ( n1891 & n1933 ) | ( ~n1934 & n1933 ) ;
  assign n1947 = ( n1835 & n1935 ) | ( n1835 & n1945 ) | ( n1935 & n1945 ) ;
  assign n1946 = ( n1835 & ~n1945 ) | ( n1835 & n1935 ) | ( ~n1945 & n1935 ) ;
  assign n1948 = ( n1945 & ~n1947 ) | ( n1945 & n1946 ) | ( ~n1947 & n1946 ) ;
  assign n1949 = ( n1837 & n1847 ) | ( n1837 & n1848 ) | ( n1847 & n1848 ) ;
  assign n1953 = x79 &  n503 ;
  assign n1950 = ( x81 & ~n450 ) | ( x81 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n1951 = x80 &  n445 ;
  assign n1952 = n1950 | n1951 ;
  assign n1954 = ( x79 & ~n1953 ) | ( x79 & n1952 ) | ( ~n1953 & n1952 ) ;
  assign n1955 = ~n453 & n994 ;
  assign n1956 = n1954 | n1955 ;
  assign n1957 = ( x11 & ~n1956 ) | ( x11 & 1'b0 ) | ( ~n1956 & 1'b0 ) ;
  assign n1958 = ~x11 & n1956 ;
  assign n1959 = n1957 | n1958 ;
  assign n1960 = ( n1948 & ~n1949 ) | ( n1948 & n1959 ) | ( ~n1949 & n1959 ) ;
  assign n1961 = ( n1948 & ~n1959 ) | ( n1948 & n1949 ) | ( ~n1959 & n1949 ) ;
  assign n1962 = ( n1960 & ~n1948 ) | ( n1960 & n1961 ) | ( ~n1948 & n1961 ) ;
  assign n1963 = ( n1853 & n1881 ) | ( n1853 & n1962 ) | ( n1881 & n1962 ) ;
  assign n1964 = ( n1853 & ~n1881 ) | ( n1853 & n1962 ) | ( ~n1881 & n1962 ) ;
  assign n1965 = ( n1881 & ~n1963 ) | ( n1881 & n1964 ) | ( ~n1963 & n1964 ) ;
  assign n1865 = x85 &  n225 ;
  assign n1862 = ( x87 & ~n197 ) | ( x87 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n1863 = x86 &  n192 ;
  assign n1864 = n1862 | n1863 ;
  assign n1866 = ( x85 & ~n1865 ) | ( x85 & n1864 ) | ( ~n1865 & n1864 ) ;
  assign n1867 = ~n200 & n1512 ;
  assign n1868 = n1866 | n1867 ;
  assign n1869 = ( x5 & ~n1868 ) | ( x5 & 1'b0 ) | ( ~n1868 & 1'b0 ) ;
  assign n1870 = ~x5 & n1868 ;
  assign n1871 = n1869 | n1870 ;
  assign n1966 = ( n1856 & ~n1965 ) | ( n1856 & n1871 ) | ( ~n1965 & n1871 ) ;
  assign n1967 = ( n1856 & ~n1871 ) | ( n1856 & n1965 ) | ( ~n1871 & n1965 ) ;
  assign n1968 = ( n1966 & ~n1856 ) | ( n1966 & n1967 ) | ( ~n1856 & n1967 ) ;
  assign n1972 = ~n136 & x90 ;
  assign n1969 = ( x88 & ~n150 ) | ( x88 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n1970 = ( x89 & ~n131 ) | ( x89 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n1971 = n1969 | n1970 ;
  assign n1973 = ( x90 & ~n1972 ) | ( x90 & n1971 ) | ( ~n1972 & n1971 ) ;
  assign n1975 = ( x89 & x90 ) | ( x89 & n1740 ) | ( x90 & n1740 ) ;
  assign n1974 = ( x89 & ~x90 ) | ( x89 & n1740 ) | ( ~x90 & n1740 ) ;
  assign n1976 = ( x90 & ~n1975 ) | ( x90 & n1974 ) | ( ~n1975 & n1974 ) ;
  assign n1977 = ( n139 & ~n1973 ) | ( n139 & n1976 ) | ( ~n1973 & n1976 ) ;
  assign n1978 = ~n139 & n1977 ;
  assign n1979 = ( x2 & n1973 ) | ( x2 & n1978 ) | ( n1973 & n1978 ) ;
  assign n1980 = ( x2 & ~n1978 ) | ( x2 & n1973 ) | ( ~n1978 & n1973 ) ;
  assign n1981 = ( n1978 & ~n1979 ) | ( n1978 & n1980 ) | ( ~n1979 & n1980 ) ;
  assign n1982 = ( n1968 & ~n1860 ) | ( n1968 & n1981 ) | ( ~n1860 & n1981 ) ;
  assign n1983 = ( n1860 & ~n1981 ) | ( n1860 & n1968 ) | ( ~n1981 & n1968 ) ;
  assign n1984 = ( n1982 & ~n1968 ) | ( n1982 & n1983 ) | ( ~n1968 & n1983 ) ;
  assign n1998 = x80 &  n503 ;
  assign n1995 = ( x82 & ~n450 ) | ( x82 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n1996 = x81 &  n445 ;
  assign n1997 = n1995 | n1996 ;
  assign n1999 = ( x80 & ~n1998 ) | ( x80 & n1997 ) | ( ~n1998 & n1997 ) ;
  assign n2000 = ~n453 & n1084 ;
  assign n2001 = n1999 | n2000 ;
  assign n2002 = ( x11 & ~n2001 ) | ( x11 & 1'b0 ) | ( ~n2001 & 1'b0 ) ;
  assign n2003 = ~x11 & n2001 ;
  assign n2004 = n2002 | n2003 ;
  assign n2069 = x77 &  n713 ;
  assign n2066 = ( x79 & ~n641 ) | ( x79 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n2067 = x78 &  n636 ;
  assign n2068 = n2066 | n2067 ;
  assign n2070 = ( x77 & ~n2069 ) | ( x77 & n2068 ) | ( ~n2069 & n2068 ) ;
  assign n2071 = ~n644 & n766 ;
  assign n2072 = n2070 | n2071 ;
  assign n2073 = ( x14 & ~n2072 ) | ( x14 & 1'b0 ) | ( ~n2072 & 1'b0 ) ;
  assign n2074 = ~x14 & n2072 ;
  assign n2075 = n2073 | n2074 ;
  assign n2008 = x74 &  n942 ;
  assign n2005 = ( x76 & ~n896 ) | ( x76 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n2006 = x75 &  n891 ;
  assign n2007 = n2005 | n2006 ;
  assign n2009 = ( x74 & ~n2008 ) | ( x74 & n2007 ) | ( ~n2008 & n2007 ) ;
  assign n2010 = ( n603 & ~n899 ) | ( n603 & 1'b0 ) | ( ~n899 & 1'b0 ) ;
  assign n2011 = n2009 | n2010 ;
  assign n2012 = ( x17 & ~n2011 ) | ( x17 & 1'b0 ) | ( ~n2011 & 1'b0 ) ;
  assign n2013 = ~x17 & n2011 ;
  assign n2014 = n2012 | n2013 ;
  assign n2015 = ( x26 & ~x27 ) | ( x26 & 1'b0 ) | ( ~x27 & 1'b0 ) ;
  assign n2016 = ~x26 & x27 ;
  assign n2017 = n2015 | n2016 ;
  assign n2018 = x64 &  n2017 ;
  assign n2019 = ( n1653 & ~n1821 ) | ( n1653 & n1901 ) | ( ~n1821 & n1901 ) ;
  assign n2020 = ( x26 & n1821 ) | ( x26 & n2019 ) | ( n1821 & n2019 ) ;
  assign n2021 = ( x26 & ~n2020 ) | ( x26 & 1'b0 ) | ( ~n2020 & 1'b0 ) ;
  assign n2025 = x65 &  n1894 ;
  assign n2022 = ( x67 & ~n1816 ) | ( x67 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n2023 = x66 &  n1811 ;
  assign n2024 = n2022 | n2023 ;
  assign n2026 = ( x65 & ~n2025 ) | ( x65 & n2024 ) | ( ~n2025 & n2024 ) ;
  assign n2027 = n173 | n1819 ;
  assign n2028 = ~n2026 & n2027 ;
  assign n2029 = x26 &  n2028 ;
  assign n2030 = x26 | n2028 ;
  assign n2031 = ~n2029 & n2030 ;
  assign n2032 = ( n2018 & ~n2021 ) | ( n2018 & n2031 ) | ( ~n2021 & n2031 ) ;
  assign n2033 = ( n2018 & ~n2031 ) | ( n2018 & n2021 ) | ( ~n2031 & n2021 ) ;
  assign n2034 = ( n2032 & ~n2018 ) | ( n2032 & n2033 ) | ( ~n2018 & n2033 ) ;
  assign n2035 = ( n1826 & n1906 ) | ( n1826 & n1916 ) | ( n1906 & n1916 ) ;
  assign n2039 = x68 &  n1551 ;
  assign n2036 = ( x70 & ~n1451 ) | ( x70 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n2037 = x69 &  n1446 ;
  assign n2038 = n2036 | n2037 ;
  assign n2040 = ( x68 & ~n2039 ) | ( x68 & n2038 ) | ( ~n2039 & n2038 ) ;
  assign n2041 = ( n282 & ~n1454 ) | ( n282 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n2042 = n2040 | n2041 ;
  assign n2043 = ( x23 & ~n2042 ) | ( x23 & 1'b0 ) | ( ~n2042 & 1'b0 ) ;
  assign n2044 = ~x23 & n2042 ;
  assign n2045 = n2043 | n2044 ;
  assign n2046 = ( n2034 & ~n2035 ) | ( n2034 & n2045 ) | ( ~n2035 & n2045 ) ;
  assign n2047 = ( n2035 & ~n2034 ) | ( n2035 & n2045 ) | ( ~n2034 & n2045 ) ;
  assign n2048 = ( n2046 & ~n2045 ) | ( n2046 & n2047 ) | ( ~n2045 & n2047 ) ;
  assign n2053 = x71 &  n1227 ;
  assign n2050 = ( x73 & ~n1154 ) | ( x73 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n2051 = x72 &  n1149 ;
  assign n2052 = n2050 | n2051 ;
  assign n2054 = ( x71 & ~n2053 ) | ( x71 & n2052 ) | ( ~n2053 & n2052 ) ;
  assign n2055 = ( n389 & ~n1157 ) | ( n389 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n2056 = n2054 | n2055 ;
  assign n2057 = ( x20 & ~n2056 ) | ( x20 & 1'b0 ) | ( ~n2056 & 1'b0 ) ;
  assign n2058 = ~x20 & n2056 ;
  assign n2059 = n2057 | n2058 ;
  assign n2049 = ( n1829 & n1919 ) | ( n1829 & n1929 ) | ( n1919 & n1929 ) ;
  assign n2060 = ( n2048 & ~n2059 ) | ( n2048 & n2049 ) | ( ~n2059 & n2049 ) ;
  assign n2061 = ( n2048 & ~n2049 ) | ( n2048 & n2059 ) | ( ~n2049 & n2059 ) ;
  assign n2062 = ( n2060 & ~n2048 ) | ( n2060 & n2061 ) | ( ~n2048 & n2061 ) ;
  assign n2063 = ( n2014 & ~n1934 ) | ( n2014 & n2062 ) | ( ~n1934 & n2062 ) ;
  assign n2064 = ( n1934 & ~n2062 ) | ( n1934 & n2014 ) | ( ~n2062 & n2014 ) ;
  assign n2065 = ( n2063 & ~n2014 ) | ( n2063 & n2064 ) | ( ~n2014 & n2064 ) ;
  assign n2076 = ( n1947 & ~n2075 ) | ( n1947 & n2065 ) | ( ~n2075 & n2065 ) ;
  assign n2077 = ( n2065 & ~n1947 ) | ( n2065 & n2075 ) | ( ~n1947 & n2075 ) ;
  assign n2078 = ( n2076 & ~n2065 ) | ( n2076 & n2077 ) | ( ~n2065 & n2077 ) ;
  assign n2079 = ( n1948 & n1949 ) | ( n1948 & n1959 ) | ( n1949 & n1959 ) ;
  assign n2080 = ( n2004 & ~n2078 ) | ( n2004 & n2079 ) | ( ~n2078 & n2079 ) ;
  assign n2081 = ( n2004 & ~n2079 ) | ( n2004 & n2078 ) | ( ~n2079 & n2078 ) ;
  assign n2082 = ( n2080 & ~n2004 ) | ( n2080 & n2081 ) | ( ~n2004 & n2081 ) ;
  assign n1988 = x83 &  n353 ;
  assign n1985 = ( x85 & ~n313 ) | ( x85 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n1986 = x84 &  n308 ;
  assign n1987 = n1985 | n1986 ;
  assign n1989 = ( x83 & ~n1988 ) | ( x83 & n1987 ) | ( ~n1988 & n1987 ) ;
  assign n1990 = ~n316 & n1295 ;
  assign n1991 = n1989 | n1990 ;
  assign n1992 = ( x8 & ~n1991 ) | ( x8 & 1'b0 ) | ( ~n1991 & 1'b0 ) ;
  assign n1993 = ~x8 & n1991 ;
  assign n1994 = n1992 | n1993 ;
  assign n2083 = ( n1963 & ~n2082 ) | ( n1963 & n1994 ) | ( ~n2082 & n1994 ) ;
  assign n2084 = ( n1994 & ~n1963 ) | ( n1994 & n2082 ) | ( ~n1963 & n2082 ) ;
  assign n2085 = ( n2083 & ~n1994 ) | ( n2083 & n2084 ) | ( ~n1994 & n2084 ) ;
  assign n2086 = ( n1856 & n1871 ) | ( n1856 & n1965 ) | ( n1871 & n1965 ) ;
  assign n2090 = x86 &  n225 ;
  assign n2087 = ( x88 & ~n197 ) | ( x88 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n2088 = x87 &  n192 ;
  assign n2089 = n2087 | n2088 ;
  assign n2091 = ( x86 & ~n2090 ) | ( x86 & n2089 ) | ( ~n2090 & n2089 ) ;
  assign n2092 = ~n200 & n1624 ;
  assign n2093 = n2091 | n2092 ;
  assign n2094 = ( x5 & ~n2093 ) | ( x5 & 1'b0 ) | ( ~n2093 & 1'b0 ) ;
  assign n2095 = ~x5 & n2093 ;
  assign n2096 = n2094 | n2095 ;
  assign n2098 = ( n2085 & n2086 ) | ( n2085 & n2096 ) | ( n2086 & n2096 ) ;
  assign n2097 = ( n2086 & ~n2085 ) | ( n2086 & n2096 ) | ( ~n2085 & n2096 ) ;
  assign n2099 = ( n2085 & ~n2098 ) | ( n2085 & n2097 ) | ( ~n2098 & n2097 ) ;
  assign n2100 = ( n1860 & n1968 ) | ( n1860 & n1981 ) | ( n1968 & n1981 ) ;
  assign n2104 = ~n136 & x91 ;
  assign n2101 = ( x89 & ~n150 ) | ( x89 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n2102 = ( x90 & ~n131 ) | ( x90 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n2103 = n2101 | n2102 ;
  assign n2105 = ( x91 & ~n2104 ) | ( x91 & n2103 ) | ( ~n2104 & n2103 ) ;
  assign n2107 = ( x90 & x91 ) | ( x90 & n1975 ) | ( x91 & n1975 ) ;
  assign n2106 = ( x90 & ~x91 ) | ( x90 & n1975 ) | ( ~x91 & n1975 ) ;
  assign n2108 = ( x91 & ~n2107 ) | ( x91 & n2106 ) | ( ~n2107 & n2106 ) ;
  assign n2109 = ( n139 & ~n2105 ) | ( n139 & n2108 ) | ( ~n2105 & n2108 ) ;
  assign n2110 = ~n139 & n2109 ;
  assign n2111 = ( x2 & n2105 ) | ( x2 & n2110 ) | ( n2105 & n2110 ) ;
  assign n2112 = ( x2 & ~n2110 ) | ( x2 & n2105 ) | ( ~n2110 & n2105 ) ;
  assign n2113 = ( n2110 & ~n2111 ) | ( n2110 & n2112 ) | ( ~n2111 & n2112 ) ;
  assign n2114 = ( n2099 & ~n2100 ) | ( n2099 & n2113 ) | ( ~n2100 & n2113 ) ;
  assign n2115 = ( n2099 & ~n2113 ) | ( n2099 & n2100 ) | ( ~n2113 & n2100 ) ;
  assign n2116 = ( n2114 & ~n2099 ) | ( n2114 & n2115 ) | ( ~n2099 & n2115 ) ;
  assign n2120 = x84 &  n353 ;
  assign n2117 = ( x86 & ~n313 ) | ( x86 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n2118 = x85 &  n308 ;
  assign n2119 = n2117 | n2118 ;
  assign n2121 = ( x84 & ~n2120 ) | ( x84 & n2119 ) | ( ~n2120 & n2119 ) ;
  assign n2122 = ~n316 & n1496 ;
  assign n2123 = n2121 | n2122 ;
  assign n2124 = ( x8 & ~n2123 ) | ( x8 & 1'b0 ) | ( ~n2123 & 1'b0 ) ;
  assign n2125 = ~x8 & n2123 ;
  assign n2126 = n2124 | n2125 ;
  assign n2130 = x81 &  n503 ;
  assign n2127 = ( x83 & ~n450 ) | ( x83 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n2128 = x82 &  n445 ;
  assign n2129 = n2127 | n2128 ;
  assign n2131 = ( x81 & ~n2130 ) | ( x81 & n2129 ) | ( ~n2130 & n2129 ) ;
  assign n2132 = ~n453 & n1100 ;
  assign n2133 = n2131 | n2132 ;
  assign n2134 = ( x11 & ~n2133 ) | ( x11 & 1'b0 ) | ( ~n2133 & 1'b0 ) ;
  assign n2135 = ~x11 & n2133 ;
  assign n2136 = n2134 | n2135 ;
  assign n2140 = x78 &  n713 ;
  assign n2137 = ( x80 & ~n641 ) | ( x80 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n2138 = x79 &  n636 ;
  assign n2139 = n2137 | n2138 ;
  assign n2141 = ( x78 & ~n2140 ) | ( x78 & n2139 ) | ( ~n2140 & n2139 ) ;
  assign n2142 = ~n644 & n842 ;
  assign n2143 = n2141 | n2142 ;
  assign n2144 = ( x14 & ~n2143 ) | ( x14 & 1'b0 ) | ( ~n2143 & 1'b0 ) ;
  assign n2145 = ~x14 & n2143 ;
  assign n2146 = n2144 | n2145 ;
  assign n2150 = x75 &  n942 ;
  assign n2147 = ( x77 & ~n896 ) | ( x77 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n2148 = x76 &  n891 ;
  assign n2149 = n2147 | n2148 ;
  assign n2151 = ( x75 & ~n2150 ) | ( x75 & n2149 ) | ( ~n2150 & n2149 ) ;
  assign n2152 = ( n677 & ~n899 ) | ( n677 & 1'b0 ) | ( ~n899 & 1'b0 ) ;
  assign n2153 = n2151 | n2152 ;
  assign n2154 = ( x17 & ~n2153 ) | ( x17 & 1'b0 ) | ( ~n2153 & 1'b0 ) ;
  assign n2155 = ~x17 & n2153 ;
  assign n2156 = n2154 | n2155 ;
  assign n2160 = x72 &  n1227 ;
  assign n2157 = ( x74 & ~n1154 ) | ( x74 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n2158 = x73 &  n1149 ;
  assign n2159 = n2157 | n2158 ;
  assign n2161 = ( x72 & ~n2160 ) | ( x72 & n2159 ) | ( ~n2160 & n2159 ) ;
  assign n2162 = ( n482 & ~n1157 ) | ( n482 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n2163 = n2161 | n2162 ;
  assign n2164 = ( x20 & ~n2163 ) | ( x20 & 1'b0 ) | ( ~n2163 & 1'b0 ) ;
  assign n2165 = ~x20 & n2163 ;
  assign n2166 = n2164 | n2165 ;
  assign n2170 = x69 &  n1551 ;
  assign n2167 = ( x71 & ~n1451 ) | ( x71 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n2168 = x70 &  n1446 ;
  assign n2169 = n2167 | n2168 ;
  assign n2171 = ( x69 & ~n2170 ) | ( x69 & n2169 ) | ( ~n2170 & n2169 ) ;
  assign n2172 = ( n298 & ~n1454 ) | ( n298 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n2173 = n2171 | n2172 ;
  assign n2174 = ( x23 & ~n2173 ) | ( x23 & 1'b0 ) | ( ~n2173 & 1'b0 ) ;
  assign n2175 = ~x23 & n2173 ;
  assign n2176 = n2174 | n2175 ;
  assign n2180 = x66 &  n1894 ;
  assign n2177 = ( x68 & ~n1816 ) | ( x68 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n2178 = x67 &  n1811 ;
  assign n2179 = n2177 | n2178 ;
  assign n2181 = ( x66 & ~n2180 ) | ( x66 & n2179 ) | ( ~n2180 & n2179 ) ;
  assign n2182 = ( n1819 & ~n2181 ) | ( n1819 & n213 ) | ( ~n2181 & n213 ) ;
  assign n2183 = ~n1819 & n2182 ;
  assign n2184 = ( n2181 & ~x26 ) | ( n2181 & n2183 ) | ( ~x26 & n2183 ) ;
  assign n2185 = ( x26 & ~n2181 ) | ( x26 & n2183 ) | ( ~n2181 & n2183 ) ;
  assign n2186 = ( n2184 & ~n2183 ) | ( n2184 & n2185 ) | ( ~n2183 & n2185 ) ;
  assign n2187 = ( x29 & ~n2018 ) | ( x29 & 1'b0 ) | ( ~n2018 & 1'b0 ) ;
  assign n2188 = ( x27 & x28 ) | ( x27 & n2015 ) | ( x28 & n2015 ) ;
  assign n2189 = ( x27 & ~n2016 ) | ( x27 & x28 ) | ( ~n2016 & x28 ) ;
  assign n2190 = ~n2188 &  n2189 ;
  assign n2191 = x64 &  n2190 ;
  assign n2192 = ~x28 & x29 ;
  assign n2193 = ( x28 & ~x29 ) | ( x28 & 1'b0 ) | ( ~x29 & 1'b0 ) ;
  assign n2194 = n2192 | n2193 ;
  assign n2195 = ~n2017 |  n2194 ;
  assign n2196 = ( x65 & ~n2195 ) | ( x65 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n2197 = n2191 | n2196 ;
  assign n2198 = ~n2017 | ~n2194 ;
  assign n2199 = ( n142 & ~n2198 ) | ( n142 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n2200 = n2197 | n2199 ;
  assign n2202 = ( x29 & n2187 ) | ( x29 & n2200 ) | ( n2187 & n2200 ) ;
  assign n2201 = ( x29 & ~n2187 ) | ( x29 & n2200 ) | ( ~n2187 & n2200 ) ;
  assign n2203 = ( n2187 & ~n2202 ) | ( n2187 & n2201 ) | ( ~n2202 & n2201 ) ;
  assign n2205 = ( n2033 & n2186 ) | ( n2033 & n2203 ) | ( n2186 & n2203 ) ;
  assign n2204 = ( n2033 & ~n2186 ) | ( n2033 & n2203 ) | ( ~n2186 & n2203 ) ;
  assign n2206 = ( n2186 & ~n2205 ) | ( n2186 & n2204 ) | ( ~n2205 & n2204 ) ;
  assign n2208 = ( n2047 & n2176 ) | ( n2047 & n2206 ) | ( n2176 & n2206 ) ;
  assign n2207 = ( n2047 & ~n2176 ) | ( n2047 & n2206 ) | ( ~n2176 & n2206 ) ;
  assign n2209 = ( n2176 & ~n2208 ) | ( n2176 & n2207 ) | ( ~n2208 & n2207 ) ;
  assign n2210 = ( n2049 & ~n2048 ) | ( n2049 & n2059 ) | ( ~n2048 & n2059 ) ;
  assign n2211 = ( n2166 & n2209 ) | ( n2166 & n2210 ) | ( n2209 & n2210 ) ;
  assign n2212 = ( n2209 & ~n2166 ) | ( n2209 & n2210 ) | ( ~n2166 & n2210 ) ;
  assign n2213 = ( n2166 & ~n2211 ) | ( n2166 & n2212 ) | ( ~n2211 & n2212 ) ;
  assign n2214 = ( n2064 & n2156 ) | ( n2064 & n2213 ) | ( n2156 & n2213 ) ;
  assign n2215 = ( n2064 & ~n2156 ) | ( n2064 & n2213 ) | ( ~n2156 & n2213 ) ;
  assign n2216 = ( n2156 & ~n2214 ) | ( n2156 & n2215 ) | ( ~n2214 & n2215 ) ;
  assign n2217 = ( n1947 & ~n2065 ) | ( n1947 & n2075 ) | ( ~n2065 & n2075 ) ;
  assign n2218 = ( n2146 & ~n2216 ) | ( n2146 & n2217 ) | ( ~n2216 & n2217 ) ;
  assign n2219 = ( n2146 & ~n2217 ) | ( n2146 & n2216 ) | ( ~n2217 & n2216 ) ;
  assign n2220 = ( n2218 & ~n2146 ) | ( n2218 & n2219 ) | ( ~n2146 & n2219 ) ;
  assign n2221 = ( n2080 & n2136 ) | ( n2080 & n2220 ) | ( n2136 & n2220 ) ;
  assign n2222 = ( n2080 & ~n2136 ) | ( n2080 & n2220 ) | ( ~n2136 & n2220 ) ;
  assign n2223 = ( n2136 & ~n2221 ) | ( n2136 & n2222 ) | ( ~n2221 & n2222 ) ;
  assign n2224 = ( n2083 & n2126 ) | ( n2083 & n2223 ) | ( n2126 & n2223 ) ;
  assign n2225 = ( n2083 & ~n2126 ) | ( n2083 & n2223 ) | ( ~n2126 & n2223 ) ;
  assign n2226 = ( n2126 & ~n2224 ) | ( n2126 & n2225 ) | ( ~n2224 & n2225 ) ;
  assign n2230 = x87 &  n225 ;
  assign n2227 = ( x89 & ~n197 ) | ( x89 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n2228 = x88 &  n192 ;
  assign n2229 = n2227 | n2228 ;
  assign n2231 = ( x87 & ~n2230 ) | ( x87 & n2229 ) | ( ~n2230 & n2229 ) ;
  assign n2232 = ~n200 & n1741 ;
  assign n2233 = n2231 | n2232 ;
  assign n2234 = ( x5 & ~n2233 ) | ( x5 & 1'b0 ) | ( ~n2233 & 1'b0 ) ;
  assign n2235 = ~x5 & n2233 ;
  assign n2236 = n2234 | n2235 ;
  assign n2237 = ( n2097 & n2226 ) | ( n2097 & n2236 ) | ( n2226 & n2236 ) ;
  assign n2238 = ( n2097 & ~n2226 ) | ( n2097 & n2236 ) | ( ~n2226 & n2236 ) ;
  assign n2239 = ( n2226 & ~n2237 ) | ( n2226 & n2238 ) | ( ~n2237 & n2238 ) ;
  assign n2244 = ~n136 & x92 ;
  assign n2241 = ( x90 & ~n150 ) | ( x90 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n2242 = ( x91 & ~n131 ) | ( x91 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n2243 = n2241 | n2242 ;
  assign n2245 = ( x92 & ~n2244 ) | ( x92 & n2243 ) | ( ~n2244 & n2243 ) ;
  assign n2247 = ( x91 & x92 ) | ( x91 & n2107 ) | ( x92 & n2107 ) ;
  assign n2246 = ( x91 & ~x92 ) | ( x91 & n2107 ) | ( ~x92 & n2107 ) ;
  assign n2248 = ( x92 & ~n2247 ) | ( x92 & n2246 ) | ( ~n2247 & n2246 ) ;
  assign n2249 = ( n139 & ~n2245 ) | ( n139 & n2248 ) | ( ~n2245 & n2248 ) ;
  assign n2250 = ~n139 & n2249 ;
  assign n2251 = ( x2 & n2245 ) | ( x2 & n2250 ) | ( n2245 & n2250 ) ;
  assign n2252 = ( x2 & ~n2250 ) | ( x2 & n2245 ) | ( ~n2250 & n2245 ) ;
  assign n2253 = ( n2250 & ~n2251 ) | ( n2250 & n2252 ) | ( ~n2251 & n2252 ) ;
  assign n2240 = ( n2100 & ~n2099 ) | ( n2100 & n2113 ) | ( ~n2099 & n2113 ) ;
  assign n2254 = ( n2239 & ~n2253 ) | ( n2239 & n2240 ) | ( ~n2253 & n2240 ) ;
  assign n2255 = ( n2239 & ~n2240 ) | ( n2239 & n2253 ) | ( ~n2240 & n2253 ) ;
  assign n2256 = ( n2254 & ~n2239 ) | ( n2254 & n2255 ) | ( ~n2239 & n2255 ) ;
  assign n2260 = ~n136 & x93 ;
  assign n2257 = ( x91 & ~n150 ) | ( x91 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n2258 = ( x92 & ~n131 ) | ( x92 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n2259 = n2257 | n2258 ;
  assign n2261 = ( x93 & ~n2260 ) | ( x93 & n2259 ) | ( ~n2260 & n2259 ) ;
  assign n2262 = ( x92 & ~x93 ) | ( x92 & n2247 ) | ( ~x93 & n2247 ) ;
  assign n2263 = ( x92 & x93 ) | ( x92 & n2247 ) | ( x93 & n2247 ) ;
  assign n2264 = ( ~x93 & ~n2262 ) | ( ~x93 & n2263 ) | ( ~n2262 & n2263 ) ;
  assign n2265 = ( n2261 & ~n139 ) | ( n2261 & n2264 ) | ( ~n139 & n2264 ) ;
  assign n2266 = n139 | n2265 ;
  assign n2268 = ( x2 & n2261 ) | ( x2 & n2266 ) | ( n2261 & n2266 ) ;
  assign n2267 = ( x2 & ~n2266 ) | ( x2 & n2261 ) | ( ~n2266 & n2261 ) ;
  assign n2269 = ( n2266 & ~n2268 ) | ( n2266 & n2267 ) | ( ~n2268 & n2267 ) ;
  assign n2390 = ( n2239 & n2240 ) | ( n2239 & n2253 ) | ( n2240 & n2253 ) ;
  assign n2374 = x82 &  n503 ;
  assign n2371 = ( x84 & ~n450 ) | ( x84 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n2372 = x83 &  n445 ;
  assign n2373 = n2371 | n2372 ;
  assign n2375 = ( x82 & ~n2374 ) | ( x82 & n2373 ) | ( ~n2374 & n2373 ) ;
  assign n2376 = ~n453 & n1199 ;
  assign n2377 = n2375 | n2376 ;
  assign n2378 = ( x11 & ~n2377 ) | ( x11 & 1'b0 ) | ( ~n2377 & 1'b0 ) ;
  assign n2379 = ~x11 & n2377 ;
  assign n2380 = n2378 | n2379 ;
  assign n2293 = x79 &  n713 ;
  assign n2290 = ( x81 & ~n641 ) | ( x81 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n2291 = x80 &  n636 ;
  assign n2292 = n2290 | n2291 ;
  assign n2294 = ( x79 & ~n2293 ) | ( x79 & n2292 ) | ( ~n2293 & n2292 ) ;
  assign n2295 = ~n644 & n994 ;
  assign n2296 = n2294 | n2295 ;
  assign n2297 = ( x14 & ~n2296 ) | ( x14 & 1'b0 ) | ( ~n2296 & 1'b0 ) ;
  assign n2298 = ~x14 & n2296 ;
  assign n2299 = n2297 | n2298 ;
  assign n2303 = x73 &  n1227 ;
  assign n2300 = ( x75 & ~n1154 ) | ( x75 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n2301 = x74 &  n1149 ;
  assign n2302 = n2300 | n2301 ;
  assign n2304 = ( x73 & ~n2303 ) | ( x73 & n2302 ) | ( ~n2303 & n2302 ) ;
  assign n2305 = ( n540 & ~n1157 ) | ( n540 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n2306 = n2304 | n2305 ;
  assign n2307 = ( x20 & ~n2306 ) | ( x20 & 1'b0 ) | ( ~n2306 & 1'b0 ) ;
  assign n2308 = ~x20 & n2306 ;
  assign n2309 = n2307 | n2308 ;
  assign n2328 = x67 &  n1894 ;
  assign n2325 = ( x69 & ~n1816 ) | ( x69 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n2326 = x68 &  n1811 ;
  assign n2327 = n2325 | n2326 ;
  assign n2329 = ( x67 & ~n2328 ) | ( x67 & n2327 ) | ( ~n2328 & n2327 ) ;
  assign n2330 = ( n246 & ~n1819 ) | ( n246 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n2331 = n2329 | n2330 ;
  assign n2332 = ( x26 & ~n2331 ) | ( x26 & 1'b0 ) | ( ~n2331 & 1'b0 ) ;
  assign n2333 = ~x26 & n2331 ;
  assign n2334 = n2332 | n2333 ;
  assign n2311 = ( x27 & ~x28 ) | ( x27 & n2194 ) | ( ~x28 & n2194 ) ;
  assign n2310 = ( x27 & ~x28 ) | ( x27 & n2017 ) | ( ~x28 & n2017 ) ;
  assign n2312 = ~n2311 |  n2310 ;
  assign n2316 = x64 &  n2312 ;
  assign n2313 = ( x66 & ~n2195 ) | ( x66 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n2314 = x65 &  n2190 ;
  assign n2315 = n2313 | n2314 ;
  assign n2317 = ( x64 & ~n2316 ) | ( x64 & n2315 ) | ( ~n2316 & n2315 ) ;
  assign n2318 = ( n157 & ~n2198 ) | ( n157 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n2319 = n2317 | n2318 ;
  assign n2320 = ( x29 & ~n2018 ) | ( x29 & n2200 ) | ( ~n2018 & n2200 ) ;
  assign n2321 = ~n2200 & n2320 ;
  assign n2322 = ( n2319 & ~x29 ) | ( n2319 & n2321 ) | ( ~x29 & n2321 ) ;
  assign n2323 = ( x29 & ~n2319 ) | ( x29 & n2321 ) | ( ~n2319 & n2321 ) ;
  assign n2324 = ( n2322 & ~n2321 ) | ( n2322 & n2323 ) | ( ~n2321 & n2323 ) ;
  assign n2335 = ( n2205 & ~n2334 ) | ( n2205 & n2324 ) | ( ~n2334 & n2324 ) ;
  assign n2336 = ( n2324 & ~n2205 ) | ( n2324 & n2334 ) | ( ~n2205 & n2334 ) ;
  assign n2337 = ( n2335 & ~n2324 ) | ( n2335 & n2336 ) | ( ~n2324 & n2336 ) ;
  assign n2341 = x70 &  n1551 ;
  assign n2338 = ( x72 & ~n1451 ) | ( x72 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n2339 = x71 &  n1446 ;
  assign n2340 = n2338 | n2339 ;
  assign n2342 = ( x70 & ~n2341 ) | ( x70 & n2340 ) | ( ~n2341 & n2340 ) ;
  assign n2343 = ( n345 & ~n1454 ) | ( n345 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n2344 = n2342 | n2343 ;
  assign n2345 = ( x23 & ~n2344 ) | ( x23 & 1'b0 ) | ( ~n2344 & 1'b0 ) ;
  assign n2346 = ~x23 & n2344 ;
  assign n2347 = n2345 | n2346 ;
  assign n2348 = ( n2337 & ~n2208 ) | ( n2337 & n2347 ) | ( ~n2208 & n2347 ) ;
  assign n2349 = ( n2208 & ~n2347 ) | ( n2208 & n2337 ) | ( ~n2347 & n2337 ) ;
  assign n2350 = ( n2348 & ~n2337 ) | ( n2348 & n2349 ) | ( ~n2337 & n2349 ) ;
  assign n2352 = ( n2211 & n2309 ) | ( n2211 & n2350 ) | ( n2309 & n2350 ) ;
  assign n2351 = ( n2211 & ~n2309 ) | ( n2211 & n2350 ) | ( ~n2309 & n2350 ) ;
  assign n2353 = ( n2309 & ~n2352 ) | ( n2309 & n2351 ) | ( ~n2352 & n2351 ) ;
  assign n2357 = x76 &  n942 ;
  assign n2354 = ( x78 & ~n896 ) | ( x78 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n2355 = x77 &  n891 ;
  assign n2356 = n2354 | n2355 ;
  assign n2358 = ( x76 & ~n2357 ) | ( x76 & n2356 ) | ( ~n2357 & n2356 ) ;
  assign n2359 = ( n693 & ~n899 ) | ( n693 & 1'b0 ) | ( ~n899 & 1'b0 ) ;
  assign n2360 = n2358 | n2359 ;
  assign n2361 = ( x17 & ~n2360 ) | ( x17 & 1'b0 ) | ( ~n2360 & 1'b0 ) ;
  assign n2362 = ~x17 & n2360 ;
  assign n2363 = n2361 | n2362 ;
  assign n2364 = ( n2353 & ~n2214 ) | ( n2353 & n2363 ) | ( ~n2214 & n2363 ) ;
  assign n2365 = ( n2214 & ~n2363 ) | ( n2214 & n2353 ) | ( ~n2363 & n2353 ) ;
  assign n2366 = ( n2364 & ~n2353 ) | ( n2364 & n2365 ) | ( ~n2353 & n2365 ) ;
  assign n2367 = ( n2146 & n2216 ) | ( n2146 & n2217 ) | ( n2216 & n2217 ) ;
  assign n2368 = ( n2299 & n2366 ) | ( n2299 & n2367 ) | ( n2366 & n2367 ) ;
  assign n2369 = ( n2366 & ~n2299 ) | ( n2366 & n2367 ) | ( ~n2299 & n2367 ) ;
  assign n2370 = ( n2299 & ~n2368 ) | ( n2299 & n2369 ) | ( ~n2368 & n2369 ) ;
  assign n2381 = ( n2221 & ~n2380 ) | ( n2221 & n2370 ) | ( ~n2380 & n2370 ) ;
  assign n2382 = ( n2370 & ~n2221 ) | ( n2370 & n2380 ) | ( ~n2221 & n2380 ) ;
  assign n2383 = ( n2381 & ~n2370 ) | ( n2381 & n2382 ) | ( ~n2370 & n2382 ) ;
  assign n2283 = x85 &  n353 ;
  assign n2280 = ( x87 & ~n313 ) | ( x87 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n2281 = x86 &  n308 ;
  assign n2282 = n2280 | n2281 ;
  assign n2284 = ( x85 & ~n2283 ) | ( x85 & n2282 ) | ( ~n2283 & n2282 ) ;
  assign n2285 = ~n316 & n1512 ;
  assign n2286 = n2284 | n2285 ;
  assign n2287 = ( x8 & ~n2286 ) | ( x8 & 1'b0 ) | ( ~n2286 & 1'b0 ) ;
  assign n2288 = ~x8 & n2286 ;
  assign n2289 = n2287 | n2288 ;
  assign n2384 = ( n2224 & ~n2383 ) | ( n2224 & n2289 ) | ( ~n2383 & n2289 ) ;
  assign n2385 = ( n2289 & ~n2224 ) | ( n2289 & n2383 ) | ( ~n2224 & n2383 ) ;
  assign n2386 = ( n2384 & ~n2289 ) | ( n2384 & n2385 ) | ( ~n2289 & n2385 ) ;
  assign n2273 = x88 &  n225 ;
  assign n2270 = ( x90 & ~n197 ) | ( x90 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n2271 = x89 &  n192 ;
  assign n2272 = n2270 | n2271 ;
  assign n2274 = ( x88 & ~n2273 ) | ( x88 & n2272 ) | ( ~n2273 & n2272 ) ;
  assign n2275 = ~n200 & n1976 ;
  assign n2276 = n2274 | n2275 ;
  assign n2277 = ( x5 & ~n2276 ) | ( x5 & 1'b0 ) | ( ~n2276 & 1'b0 ) ;
  assign n2278 = ~x5 & n2276 ;
  assign n2279 = n2277 | n2278 ;
  assign n2387 = ( n2237 & n2279 ) | ( n2237 & n2386 ) | ( n2279 & n2386 ) ;
  assign n2388 = ( n2237 & ~n2386 ) | ( n2237 & n2279 ) | ( ~n2386 & n2279 ) ;
  assign n2389 = ( n2386 & ~n2387 ) | ( n2386 & n2388 ) | ( ~n2387 & n2388 ) ;
  assign n2391 = ( n2269 & ~n2390 ) | ( n2269 & n2389 ) | ( ~n2390 & n2389 ) ;
  assign n2392 = ( n2269 & ~n2389 ) | ( n2269 & n2390 ) | ( ~n2389 & n2390 ) ;
  assign n2393 = ( n2391 & ~n2269 ) | ( n2391 & n2392 ) | ( ~n2269 & n2392 ) ;
  assign n2397 = ~n136 & x94 ;
  assign n2394 = ( x92 & ~n150 ) | ( x92 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n2395 = ( x93 & ~n131 ) | ( x93 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n2396 = n2394 | n2395 ;
  assign n2398 = ( x94 & ~n2397 ) | ( x94 & n2396 ) | ( ~n2397 & n2396 ) ;
  assign n2400 = ( x93 & x94 ) | ( x93 & n2263 ) | ( x94 & n2263 ) ;
  assign n2399 = ( x93 & ~x94 ) | ( x93 & n2263 ) | ( ~x94 & n2263 ) ;
  assign n2401 = ( x94 & ~n2400 ) | ( x94 & n2399 ) | ( ~n2400 & n2399 ) ;
  assign n2402 = ( n139 & ~n2398 ) | ( n139 & n2401 ) | ( ~n2398 & n2401 ) ;
  assign n2403 = ~n139 & n2402 ;
  assign n2404 = ( x2 & n2398 ) | ( x2 & n2403 ) | ( n2398 & n2403 ) ;
  assign n2405 = ( x2 & ~n2403 ) | ( x2 & n2398 ) | ( ~n2403 & n2398 ) ;
  assign n2406 = ( n2403 & ~n2404 ) | ( n2403 & n2405 ) | ( ~n2404 & n2405 ) ;
  assign n2420 = x74 &  n1227 ;
  assign n2417 = ( x76 & ~n1154 ) | ( x76 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n2418 = x75 &  n1149 ;
  assign n2419 = n2417 | n2418 ;
  assign n2421 = ( x74 & ~n2420 ) | ( x74 & n2419 ) | ( ~n2420 & n2419 ) ;
  assign n2422 = ( n603 & ~n1157 ) | ( n603 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n2423 = n2421 | n2422 ;
  assign n2424 = ( x20 & ~n2423 ) | ( x20 & 1'b0 ) | ( ~n2423 & 1'b0 ) ;
  assign n2425 = ~x20 & n2423 ;
  assign n2426 = n2424 | n2425 ;
  assign n2427 = ( x29 & ~x30 ) | ( x29 & 1'b0 ) | ( ~x30 & 1'b0 ) ;
  assign n2428 = ~x29 & x30 ;
  assign n2429 = n2427 | n2428 ;
  assign n2430 = x64 &  n2429 ;
  assign n2431 = ( n2018 & ~n2200 ) | ( n2018 & n2319 ) | ( ~n2200 & n2319 ) ;
  assign n2432 = ( x29 & n2200 ) | ( x29 & n2431 ) | ( n2200 & n2431 ) ;
  assign n2433 = ( x29 & ~n2432 ) | ( x29 & 1'b0 ) | ( ~n2432 & 1'b0 ) ;
  assign n2437 = x65 &  n2312 ;
  assign n2434 = ( x67 & ~n2195 ) | ( x67 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n2435 = x66 &  n2190 ;
  assign n2436 = n2434 | n2435 ;
  assign n2438 = ( x65 & ~n2437 ) | ( x65 & n2436 ) | ( ~n2437 & n2436 ) ;
  assign n2439 = n173 | n2198 ;
  assign n2440 = ~n2438 & n2439 ;
  assign n2441 = x29 &  n2440 ;
  assign n2442 = x29 | n2440 ;
  assign n2443 = ~n2441 & n2442 ;
  assign n2444 = ( n2430 & ~n2433 ) | ( n2430 & n2443 ) | ( ~n2433 & n2443 ) ;
  assign n2445 = ( n2430 & ~n2443 ) | ( n2430 & n2433 ) | ( ~n2443 & n2433 ) ;
  assign n2446 = ( n2444 & ~n2430 ) | ( n2444 & n2445 ) | ( ~n2430 & n2445 ) ;
  assign n2447 = ( n2205 & n2324 ) | ( n2205 & n2334 ) | ( n2324 & n2334 ) ;
  assign n2451 = x68 &  n1894 ;
  assign n2448 = ( x70 & ~n1816 ) | ( x70 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n2449 = x69 &  n1811 ;
  assign n2450 = n2448 | n2449 ;
  assign n2452 = ( x68 & ~n2451 ) | ( x68 & n2450 ) | ( ~n2451 & n2450 ) ;
  assign n2453 = ( n282 & ~n1819 ) | ( n282 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n2454 = n2452 | n2453 ;
  assign n2455 = ( x26 & ~n2454 ) | ( x26 & 1'b0 ) | ( ~n2454 & 1'b0 ) ;
  assign n2456 = ~x26 & n2454 ;
  assign n2457 = n2455 | n2456 ;
  assign n2458 = ( n2446 & ~n2447 ) | ( n2446 & n2457 ) | ( ~n2447 & n2457 ) ;
  assign n2459 = ( n2447 & ~n2446 ) | ( n2447 & n2457 ) | ( ~n2446 & n2457 ) ;
  assign n2460 = ( n2458 & ~n2457 ) | ( n2458 & n2459 ) | ( ~n2457 & n2459 ) ;
  assign n2465 = x71 &  n1551 ;
  assign n2462 = ( x73 & ~n1451 ) | ( x73 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n2463 = x72 &  n1446 ;
  assign n2464 = n2462 | n2463 ;
  assign n2466 = ( x71 & ~n2465 ) | ( x71 & n2464 ) | ( ~n2465 & n2464 ) ;
  assign n2467 = ( n389 & ~n1454 ) | ( n389 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n2468 = n2466 | n2467 ;
  assign n2469 = ( x23 & ~n2468 ) | ( x23 & 1'b0 ) | ( ~n2468 & 1'b0 ) ;
  assign n2470 = ~x23 & n2468 ;
  assign n2471 = n2469 | n2470 ;
  assign n2461 = ( n2208 & n2337 ) | ( n2208 & n2347 ) | ( n2337 & n2347 ) ;
  assign n2472 = ( n2460 & ~n2471 ) | ( n2460 & n2461 ) | ( ~n2471 & n2461 ) ;
  assign n2473 = ( n2460 & ~n2461 ) | ( n2460 & n2471 ) | ( ~n2461 & n2471 ) ;
  assign n2474 = ( n2472 & ~n2460 ) | ( n2472 & n2473 ) | ( ~n2460 & n2473 ) ;
  assign n2475 = ( n2426 & ~n2352 ) | ( n2426 & n2474 ) | ( ~n2352 & n2474 ) ;
  assign n2476 = ( n2352 & ~n2474 ) | ( n2352 & n2426 ) | ( ~n2474 & n2426 ) ;
  assign n2477 = ( n2475 & ~n2426 ) | ( n2475 & n2476 ) | ( ~n2426 & n2476 ) ;
  assign n2481 = x77 &  n942 ;
  assign n2478 = ( x79 & ~n896 ) | ( x79 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n2479 = x78 &  n891 ;
  assign n2480 = n2478 | n2479 ;
  assign n2482 = ( x77 & ~n2481 ) | ( x77 & n2480 ) | ( ~n2481 & n2480 ) ;
  assign n2483 = ( n766 & ~n899 ) | ( n766 & 1'b0 ) | ( ~n899 & 1'b0 ) ;
  assign n2484 = n2482 | n2483 ;
  assign n2485 = ( x17 & ~n2484 ) | ( x17 & 1'b0 ) | ( ~n2484 & 1'b0 ) ;
  assign n2486 = ~x17 & n2484 ;
  assign n2487 = n2485 | n2486 ;
  assign n2488 = ( n2214 & n2353 ) | ( n2214 & n2363 ) | ( n2353 & n2363 ) ;
  assign n2489 = ( n2477 & ~n2487 ) | ( n2477 & n2488 ) | ( ~n2487 & n2488 ) ;
  assign n2490 = ( n2477 & ~n2488 ) | ( n2477 & n2487 ) | ( ~n2488 & n2487 ) ;
  assign n2491 = ( n2489 & ~n2477 ) | ( n2489 & n2490 ) | ( ~n2477 & n2490 ) ;
  assign n2410 = x80 &  n713 ;
  assign n2407 = ( x82 & ~n641 ) | ( x82 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n2408 = x81 &  n636 ;
  assign n2409 = n2407 | n2408 ;
  assign n2411 = ( x80 & ~n2410 ) | ( x80 & n2409 ) | ( ~n2410 & n2409 ) ;
  assign n2412 = ~n644 & n1084 ;
  assign n2413 = n2411 | n2412 ;
  assign n2414 = ( x14 & ~n2413 ) | ( x14 & 1'b0 ) | ( ~n2413 & 1'b0 ) ;
  assign n2415 = ~x14 & n2413 ;
  assign n2416 = n2414 | n2415 ;
  assign n2492 = ( n2368 & ~n2491 ) | ( n2368 & n2416 ) | ( ~n2491 & n2416 ) ;
  assign n2493 = ( n2416 & ~n2368 ) | ( n2416 & n2491 ) | ( ~n2368 & n2491 ) ;
  assign n2494 = ( n2492 & ~n2416 ) | ( n2492 & n2493 ) | ( ~n2416 & n2493 ) ;
  assign n2495 = ( n2221 & n2370 ) | ( n2221 & n2380 ) | ( n2370 & n2380 ) ;
  assign n2499 = x83 &  n503 ;
  assign n2496 = ( x85 & ~n450 ) | ( x85 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n2497 = x84 &  n445 ;
  assign n2498 = n2496 | n2497 ;
  assign n2500 = ( x83 & ~n2499 ) | ( x83 & n2498 ) | ( ~n2499 & n2498 ) ;
  assign n2501 = ~n453 & n1295 ;
  assign n2502 = n2500 | n2501 ;
  assign n2503 = ( x11 & ~n2502 ) | ( x11 & 1'b0 ) | ( ~n2502 & 1'b0 ) ;
  assign n2504 = ~x11 & n2502 ;
  assign n2505 = n2503 | n2504 ;
  assign n2506 = ( n2494 & ~n2495 ) | ( n2494 & n2505 ) | ( ~n2495 & n2505 ) ;
  assign n2507 = ( n2494 & ~n2505 ) | ( n2494 & n2495 ) | ( ~n2505 & n2495 ) ;
  assign n2508 = ( n2506 & ~n2494 ) | ( n2506 & n2507 ) | ( ~n2494 & n2507 ) ;
  assign n2513 = x86 &  n353 ;
  assign n2510 = ( x88 & ~n313 ) | ( x88 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n2511 = x87 &  n308 ;
  assign n2512 = n2510 | n2511 ;
  assign n2514 = ( x86 & ~n2513 ) | ( x86 & n2512 ) | ( ~n2513 & n2512 ) ;
  assign n2515 = ~n316 & n1624 ;
  assign n2516 = n2514 | n2515 ;
  assign n2517 = ( x8 & ~n2516 ) | ( x8 & 1'b0 ) | ( ~n2516 & 1'b0 ) ;
  assign n2518 = ~x8 & n2516 ;
  assign n2519 = n2517 | n2518 ;
  assign n2509 = ( n2224 & n2289 ) | ( n2224 & n2383 ) | ( n2289 & n2383 ) ;
  assign n2520 = ( n2508 & ~n2519 ) | ( n2508 & n2509 ) | ( ~n2519 & n2509 ) ;
  assign n2521 = ( n2508 & ~n2509 ) | ( n2508 & n2519 ) | ( ~n2509 & n2519 ) ;
  assign n2522 = ( n2520 & ~n2508 ) | ( n2520 & n2521 ) | ( ~n2508 & n2521 ) ;
  assign n2526 = x89 &  n225 ;
  assign n2523 = ( x91 & ~n197 ) | ( x91 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n2524 = x90 &  n192 ;
  assign n2525 = n2523 | n2524 ;
  assign n2527 = ( x89 & ~n2526 ) | ( x89 & n2525 ) | ( ~n2526 & n2525 ) ;
  assign n2528 = ~n200 & n2108 ;
  assign n2529 = n2527 | n2528 ;
  assign n2530 = ( x5 & ~n2529 ) | ( x5 & 1'b0 ) | ( ~n2529 & 1'b0 ) ;
  assign n2531 = ~x5 & n2529 ;
  assign n2532 = n2530 | n2531 ;
  assign n2533 = ( n2387 & n2522 ) | ( n2387 & n2532 ) | ( n2522 & n2532 ) ;
  assign n2534 = ( n2522 & ~n2387 ) | ( n2522 & n2532 ) | ( ~n2387 & n2532 ) ;
  assign n2535 = ( n2387 & ~n2533 ) | ( n2387 & n2534 ) | ( ~n2533 & n2534 ) ;
  assign n2536 = ( n2389 & ~n2269 ) | ( n2389 & n2390 ) | ( ~n2269 & n2390 ) ;
  assign n2537 = ( n2406 & ~n2535 ) | ( n2406 & n2536 ) | ( ~n2535 & n2536 ) ;
  assign n2538 = ( n2406 & ~n2536 ) | ( n2406 & n2535 ) | ( ~n2536 & n2535 ) ;
  assign n2539 = ( n2537 & ~n2406 ) | ( n2537 & n2538 ) | ( ~n2406 & n2538 ) ;
  assign n2543 = ~n136 & x95 ;
  assign n2540 = ( x93 & ~n150 ) | ( x93 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n2541 = ( x94 & ~n131 ) | ( x94 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n2542 = n2540 | n2541 ;
  assign n2544 = ( x95 & ~n2543 ) | ( x95 & n2542 ) | ( ~n2543 & n2542 ) ;
  assign n2546 = ( x94 & x95 ) | ( x94 & n2400 ) | ( x95 & n2400 ) ;
  assign n2545 = ( x94 & ~x95 ) | ( x94 & n2400 ) | ( ~x95 & n2400 ) ;
  assign n2547 = ( x95 & ~n2546 ) | ( x95 & n2545 ) | ( ~n2546 & n2545 ) ;
  assign n2548 = ( n139 & ~n2544 ) | ( n139 & n2547 ) | ( ~n2544 & n2547 ) ;
  assign n2549 = ~n139 & n2548 ;
  assign n2550 = ( x2 & n2544 ) | ( x2 & n2549 ) | ( n2544 & n2549 ) ;
  assign n2551 = ( x2 & ~n2549 ) | ( x2 & n2544 ) | ( ~n2549 & n2544 ) ;
  assign n2552 = ( n2549 & ~n2550 ) | ( n2549 & n2551 ) | ( ~n2550 & n2551 ) ;
  assign n2553 = ( n2387 & ~n2522 ) | ( n2387 & n2532 ) | ( ~n2522 & n2532 ) ;
  assign n2567 = x87 &  n353 ;
  assign n2564 = ( x89 & ~n313 ) | ( x89 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n2565 = x88 &  n308 ;
  assign n2566 = n2564 | n2565 ;
  assign n2568 = ( x87 & ~n2567 ) | ( x87 & n2566 ) | ( ~n2567 & n2566 ) ;
  assign n2569 = ~n316 & n1741 ;
  assign n2570 = n2568 | n2569 ;
  assign n2571 = ( x8 & ~n2570 ) | ( x8 & 1'b0 ) | ( ~n2570 & 1'b0 ) ;
  assign n2572 = ~x8 & n2570 ;
  assign n2573 = n2571 | n2572 ;
  assign n2577 = x84 &  n503 ;
  assign n2574 = ( x86 & ~n450 ) | ( x86 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n2575 = x85 &  n445 ;
  assign n2576 = n2574 | n2575 ;
  assign n2578 = ( x84 & ~n2577 ) | ( x84 & n2576 ) | ( ~n2577 & n2576 ) ;
  assign n2579 = ~n453 & n1496 ;
  assign n2580 = n2578 | n2579 ;
  assign n2581 = ( x11 & ~n2580 ) | ( x11 & 1'b0 ) | ( ~n2580 & 1'b0 ) ;
  assign n2582 = ~x11 & n2580 ;
  assign n2583 = n2581 | n2582 ;
  assign n2587 = x81 &  n713 ;
  assign n2584 = ( x83 & ~n641 ) | ( x83 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n2585 = x82 &  n636 ;
  assign n2586 = n2584 | n2585 ;
  assign n2588 = ( x81 & ~n2587 ) | ( x81 & n2586 ) | ( ~n2587 & n2586 ) ;
  assign n2589 = ~n644 & n1100 ;
  assign n2590 = n2588 | n2589 ;
  assign n2591 = ( x14 & ~n2590 ) | ( x14 & 1'b0 ) | ( ~n2590 & 1'b0 ) ;
  assign n2592 = ~x14 & n2590 ;
  assign n2593 = n2591 | n2592 ;
  assign n2597 = x75 &  n1227 ;
  assign n2594 = ( x77 & ~n1154 ) | ( x77 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n2595 = x76 &  n1149 ;
  assign n2596 = n2594 | n2595 ;
  assign n2598 = ( x75 & ~n2597 ) | ( x75 & n2596 ) | ( ~n2597 & n2596 ) ;
  assign n2599 = ( n677 & ~n1157 ) | ( n677 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n2600 = n2598 | n2599 ;
  assign n2601 = ( x20 & ~n2600 ) | ( x20 & 1'b0 ) | ( ~n2600 & 1'b0 ) ;
  assign n2602 = ~x20 & n2600 ;
  assign n2603 = n2601 | n2602 ;
  assign n2607 = x72 &  n1551 ;
  assign n2604 = ( x74 & ~n1451 ) | ( x74 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n2605 = x73 &  n1446 ;
  assign n2606 = n2604 | n2605 ;
  assign n2608 = ( x72 & ~n2607 ) | ( x72 & n2606 ) | ( ~n2607 & n2606 ) ;
  assign n2609 = ( n482 & ~n1454 ) | ( n482 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n2610 = n2608 | n2609 ;
  assign n2611 = ( x23 & ~n2610 ) | ( x23 & 1'b0 ) | ( ~n2610 & 1'b0 ) ;
  assign n2612 = ~x23 & n2610 ;
  assign n2613 = n2611 | n2612 ;
  assign n2617 = x69 &  n1894 ;
  assign n2614 = ( x71 & ~n1816 ) | ( x71 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n2615 = x70 &  n1811 ;
  assign n2616 = n2614 | n2615 ;
  assign n2618 = ( x69 & ~n2617 ) | ( x69 & n2616 ) | ( ~n2617 & n2616 ) ;
  assign n2619 = ( n298 & ~n1819 ) | ( n298 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n2620 = n2618 | n2619 ;
  assign n2621 = ( x26 & ~n2620 ) | ( x26 & 1'b0 ) | ( ~n2620 & 1'b0 ) ;
  assign n2622 = ~x26 & n2620 ;
  assign n2623 = n2621 | n2622 ;
  assign n2627 = x66 &  n2312 ;
  assign n2624 = ( x68 & ~n2195 ) | ( x68 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n2625 = x67 &  n2190 ;
  assign n2626 = n2624 | n2625 ;
  assign n2628 = ( x66 & ~n2627 ) | ( x66 & n2626 ) | ( ~n2627 & n2626 ) ;
  assign n2629 = ( n2198 & ~n2628 ) | ( n2198 & n213 ) | ( ~n2628 & n213 ) ;
  assign n2630 = ~n2198 & n2629 ;
  assign n2631 = ( n2628 & ~x29 ) | ( n2628 & n2630 ) | ( ~x29 & n2630 ) ;
  assign n2632 = ( x29 & ~n2628 ) | ( x29 & n2630 ) | ( ~n2628 & n2630 ) ;
  assign n2633 = ( n2631 & ~n2630 ) | ( n2631 & n2632 ) | ( ~n2630 & n2632 ) ;
  assign n2634 = ( x32 & ~n2430 ) | ( x32 & 1'b0 ) | ( ~n2430 & 1'b0 ) ;
  assign n2635 = ( x30 & x31 ) | ( x30 & n2427 ) | ( x31 & n2427 ) ;
  assign n2636 = ( x30 & ~n2428 ) | ( x30 & x31 ) | ( ~n2428 & x31 ) ;
  assign n2637 = ~n2635 &  n2636 ;
  assign n2638 = x64 &  n2637 ;
  assign n2639 = ~x31 & x32 ;
  assign n2640 = ( x31 & ~x32 ) | ( x31 & 1'b0 ) | ( ~x32 & 1'b0 ) ;
  assign n2641 = n2639 | n2640 ;
  assign n2642 = ~n2429 |  n2641 ;
  assign n2643 = ( x65 & ~n2642 ) | ( x65 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n2644 = n2638 | n2643 ;
  assign n2645 = ~n2429 | ~n2641 ;
  assign n2646 = ( n142 & ~n2645 ) | ( n142 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n2647 = n2644 | n2646 ;
  assign n2649 = ( x32 & n2634 ) | ( x32 & n2647 ) | ( n2634 & n2647 ) ;
  assign n2648 = ( x32 & ~n2634 ) | ( x32 & n2647 ) | ( ~n2634 & n2647 ) ;
  assign n2650 = ( n2634 & ~n2649 ) | ( n2634 & n2648 ) | ( ~n2649 & n2648 ) ;
  assign n2652 = ( n2445 & n2633 ) | ( n2445 & n2650 ) | ( n2633 & n2650 ) ;
  assign n2651 = ( n2445 & ~n2633 ) | ( n2445 & n2650 ) | ( ~n2633 & n2650 ) ;
  assign n2653 = ( n2633 & ~n2652 ) | ( n2633 & n2651 ) | ( ~n2652 & n2651 ) ;
  assign n2655 = ( n2459 & n2623 ) | ( n2459 & n2653 ) | ( n2623 & n2653 ) ;
  assign n2654 = ( n2459 & ~n2623 ) | ( n2459 & n2653 ) | ( ~n2623 & n2653 ) ;
  assign n2656 = ( n2623 & ~n2655 ) | ( n2623 & n2654 ) | ( ~n2655 & n2654 ) ;
  assign n2657 = ( n2461 & ~n2460 ) | ( n2461 & n2471 ) | ( ~n2460 & n2471 ) ;
  assign n2658 = ( n2613 & n2656 ) | ( n2613 & n2657 ) | ( n2656 & n2657 ) ;
  assign n2659 = ( n2656 & ~n2613 ) | ( n2656 & n2657 ) | ( ~n2613 & n2657 ) ;
  assign n2660 = ( n2613 & ~n2658 ) | ( n2613 & n2659 ) | ( ~n2658 & n2659 ) ;
  assign n2661 = ( n2476 & n2603 ) | ( n2476 & n2660 ) | ( n2603 & n2660 ) ;
  assign n2662 = ( n2476 & ~n2603 ) | ( n2476 & n2660 ) | ( ~n2603 & n2660 ) ;
  assign n2663 = ( n2603 & ~n2661 ) | ( n2603 & n2662 ) | ( ~n2661 & n2662 ) ;
  assign n2674 = ( n2487 & ~n2477 ) | ( n2487 & n2488 ) | ( ~n2477 & n2488 ) ;
  assign n2667 = x78 &  n942 ;
  assign n2664 = ( x80 & ~n896 ) | ( x80 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n2665 = x79 &  n891 ;
  assign n2666 = n2664 | n2665 ;
  assign n2668 = ( x78 & ~n2667 ) | ( x78 & n2666 ) | ( ~n2667 & n2666 ) ;
  assign n2669 = ( n842 & ~n899 ) | ( n842 & 1'b0 ) | ( ~n899 & 1'b0 ) ;
  assign n2670 = n2668 | n2669 ;
  assign n2671 = ( x17 & ~n2670 ) | ( x17 & 1'b0 ) | ( ~n2670 & 1'b0 ) ;
  assign n2672 = ~x17 & n2670 ;
  assign n2673 = n2671 | n2672 ;
  assign n2675 = ( n2663 & ~n2674 ) | ( n2663 & n2673 ) | ( ~n2674 & n2673 ) ;
  assign n2676 = ( n2663 & ~n2673 ) | ( n2663 & n2674 ) | ( ~n2673 & n2674 ) ;
  assign n2677 = ( n2675 & ~n2663 ) | ( n2675 & n2676 ) | ( ~n2663 & n2676 ) ;
  assign n2678 = ( n2492 & n2593 ) | ( n2492 & n2677 ) | ( n2593 & n2677 ) ;
  assign n2679 = ( n2492 & ~n2593 ) | ( n2492 & n2677 ) | ( ~n2593 & n2677 ) ;
  assign n2680 = ( n2593 & ~n2678 ) | ( n2593 & n2679 ) | ( ~n2678 & n2679 ) ;
  assign n2681 = ( n2495 & ~n2494 ) | ( n2495 & n2505 ) | ( ~n2494 & n2505 ) ;
  assign n2682 = ( n2583 & n2680 ) | ( n2583 & n2681 ) | ( n2680 & n2681 ) ;
  assign n2683 = ( n2680 & ~n2583 ) | ( n2680 & n2681 ) | ( ~n2583 & n2681 ) ;
  assign n2684 = ( n2583 & ~n2682 ) | ( n2583 & n2683 ) | ( ~n2682 & n2683 ) ;
  assign n2685 = ( n2509 & ~n2508 ) | ( n2509 & n2519 ) | ( ~n2508 & n2519 ) ;
  assign n2686 = ( n2573 & n2684 ) | ( n2573 & n2685 ) | ( n2684 & n2685 ) ;
  assign n2687 = ( n2684 & ~n2573 ) | ( n2684 & n2685 ) | ( ~n2573 & n2685 ) ;
  assign n2688 = ( n2573 & ~n2686 ) | ( n2573 & n2687 ) | ( ~n2686 & n2687 ) ;
  assign n2557 = x90 &  n225 ;
  assign n2554 = ( x92 & ~n197 ) | ( x92 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n2555 = x91 &  n192 ;
  assign n2556 = n2554 | n2555 ;
  assign n2558 = ( x90 & ~n2557 ) | ( x90 & n2556 ) | ( ~n2557 & n2556 ) ;
  assign n2559 = ~n200 & n2248 ;
  assign n2560 = n2558 | n2559 ;
  assign n2561 = ( x5 & ~n2560 ) | ( x5 & 1'b0 ) | ( ~n2560 & 1'b0 ) ;
  assign n2562 = ~x5 & n2560 ;
  assign n2563 = n2561 | n2562 ;
  assign n2689 = ( n2553 & ~n2688 ) | ( n2553 & n2563 ) | ( ~n2688 & n2563 ) ;
  assign n2690 = ( n2553 & ~n2563 ) | ( n2553 & n2688 ) | ( ~n2563 & n2688 ) ;
  assign n2691 = ( n2689 & ~n2553 ) | ( n2689 & n2690 ) | ( ~n2553 & n2690 ) ;
  assign n2692 = ( n2537 & n2552 ) | ( n2537 & n2691 ) | ( n2552 & n2691 ) ;
  assign n2693 = ( n2537 & ~n2552 ) | ( n2537 & n2691 ) | ( ~n2552 & n2691 ) ;
  assign n2694 = ( n2552 & ~n2692 ) | ( n2552 & n2693 ) | ( ~n2692 & n2693 ) ;
  assign n2832 = ~n136 & x96 ;
  assign n2829 = ( x94 & ~n150 ) | ( x94 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n2830 = ( x95 & ~n131 ) | ( x95 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n2831 = n2829 | n2830 ;
  assign n2833 = ( x96 & ~n2832 ) | ( x96 & n2831 ) | ( ~n2832 & n2831 ) ;
  assign n2835 = ( x95 & x96 ) | ( x95 & n2546 ) | ( x96 & n2546 ) ;
  assign n2834 = ( x95 & ~x96 ) | ( x95 & n2546 ) | ( ~x96 & n2546 ) ;
  assign n2836 = ( x96 & ~n2835 ) | ( x96 & n2834 ) | ( ~n2835 & n2834 ) ;
  assign n2837 = ( n139 & ~n2833 ) | ( n139 & n2836 ) | ( ~n2833 & n2836 ) ;
  assign n2838 = ~n139 & n2837 ;
  assign n2839 = ( x2 & n2833 ) | ( x2 & n2838 ) | ( n2833 & n2838 ) ;
  assign n2840 = ( x2 & ~n2838 ) | ( x2 & n2833 ) | ( ~n2838 & n2833 ) ;
  assign n2841 = ( n2838 & ~n2839 ) | ( n2838 & n2840 ) | ( ~n2839 & n2840 ) ;
  assign n2695 = ( n2553 & n2563 ) | ( n2553 & n2688 ) | ( n2563 & n2688 ) ;
  assign n2699 = x91 &  n225 ;
  assign n2696 = ( x93 & ~n197 ) | ( x93 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n2697 = x92 &  n192 ;
  assign n2698 = n2696 | n2697 ;
  assign n2700 = ( x91 & ~n2699 ) | ( x91 & n2698 ) | ( ~n2699 & n2698 ) ;
  assign n2701 = n200 | n2264 ;
  assign n2702 = ~n2700 & n2701 ;
  assign n2703 = x5 &  n2702 ;
  assign n2704 = x5 | n2702 ;
  assign n2705 = ~n2703 & n2704 ;
  assign n2790 = x82 &  n713 ;
  assign n2787 = ( x84 & ~n641 ) | ( x84 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n2788 = x83 &  n636 ;
  assign n2789 = n2787 | n2788 ;
  assign n2791 = ( x82 & ~n2790 ) | ( x82 & n2789 ) | ( ~n2790 & n2789 ) ;
  assign n2792 = ~n644 & n1199 ;
  assign n2793 = n2791 | n2792 ;
  assign n2794 = ( x14 & ~n2793 ) | ( x14 & 1'b0 ) | ( ~n2793 & 1'b0 ) ;
  assign n2795 = ~x14 & n2793 ;
  assign n2796 = n2794 | n2795 ;
  assign n2750 = x73 &  n1551 ;
  assign n2747 = ( x75 & ~n1451 ) | ( x75 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n2748 = x74 &  n1446 ;
  assign n2749 = n2747 | n2748 ;
  assign n2751 = ( x73 & ~n2750 ) | ( x73 & n2749 ) | ( ~n2750 & n2749 ) ;
  assign n2752 = ( n540 & ~n1454 ) | ( n540 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n2753 = n2751 | n2752 ;
  assign n2754 = ( x23 & ~n2753 ) | ( x23 & 1'b0 ) | ( ~n2753 & 1'b0 ) ;
  assign n2755 = ~x23 & n2753 ;
  assign n2756 = n2754 | n2755 ;
  assign n2734 = x67 &  n2312 ;
  assign n2731 = ( x69 & ~n2195 ) | ( x69 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n2732 = x68 &  n2190 ;
  assign n2733 = n2731 | n2732 ;
  assign n2735 = ( x67 & ~n2734 ) | ( x67 & n2733 ) | ( ~n2734 & n2733 ) ;
  assign n2736 = ( n246 & ~n2198 ) | ( n246 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n2737 = n2735 | n2736 ;
  assign n2738 = ( x29 & ~n2737 ) | ( x29 & 1'b0 ) | ( ~n2737 & 1'b0 ) ;
  assign n2739 = ~x29 & n2737 ;
  assign n2740 = n2738 | n2739 ;
  assign n2717 = ( x30 & ~x31 ) | ( x30 & n2641 ) | ( ~x31 & n2641 ) ;
  assign n2716 = ( x30 & ~x31 ) | ( x30 & n2429 ) | ( ~x31 & n2429 ) ;
  assign n2718 = ~n2717 |  n2716 ;
  assign n2722 = x64 &  n2718 ;
  assign n2719 = ( x66 & ~n2642 ) | ( x66 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n2720 = x65 &  n2637 ;
  assign n2721 = n2719 | n2720 ;
  assign n2723 = ( x64 & ~n2722 ) | ( x64 & n2721 ) | ( ~n2722 & n2721 ) ;
  assign n2724 = ( n157 & ~n2645 ) | ( n157 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n2725 = n2723 | n2724 ;
  assign n2726 = ( x32 & ~n2430 ) | ( x32 & n2647 ) | ( ~n2430 & n2647 ) ;
  assign n2727 = ~n2647 & n2726 ;
  assign n2728 = ( n2725 & ~x32 ) | ( n2725 & n2727 ) | ( ~x32 & n2727 ) ;
  assign n2729 = ( x32 & ~n2725 ) | ( x32 & n2727 ) | ( ~n2725 & n2727 ) ;
  assign n2730 = ( n2728 & ~n2727 ) | ( n2728 & n2729 ) | ( ~n2727 & n2729 ) ;
  assign n2741 = ( n2652 & ~n2740 ) | ( n2652 & n2730 ) | ( ~n2740 & n2730 ) ;
  assign n2742 = ( n2730 & ~n2652 ) | ( n2730 & n2740 ) | ( ~n2652 & n2740 ) ;
  assign n2743 = ( n2741 & ~n2730 ) | ( n2741 & n2742 ) | ( ~n2730 & n2742 ) ;
  assign n2709 = x70 &  n1894 ;
  assign n2706 = ( x72 & ~n1816 ) | ( x72 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n2707 = x71 &  n1811 ;
  assign n2708 = n2706 | n2707 ;
  assign n2710 = ( x70 & ~n2709 ) | ( x70 & n2708 ) | ( ~n2709 & n2708 ) ;
  assign n2711 = ( n345 & ~n1819 ) | ( n345 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n2712 = n2710 | n2711 ;
  assign n2713 = ( x26 & ~n2712 ) | ( x26 & 1'b0 ) | ( ~n2712 & 1'b0 ) ;
  assign n2714 = ~x26 & n2712 ;
  assign n2715 = n2713 | n2714 ;
  assign n2744 = ( n2655 & ~n2743 ) | ( n2655 & n2715 ) | ( ~n2743 & n2715 ) ;
  assign n2745 = ( n2715 & ~n2655 ) | ( n2715 & n2743 ) | ( ~n2655 & n2743 ) ;
  assign n2746 = ( n2744 & ~n2715 ) | ( n2744 & n2745 ) | ( ~n2715 & n2745 ) ;
  assign n2757 = ( n2658 & ~n2756 ) | ( n2658 & n2746 ) | ( ~n2756 & n2746 ) ;
  assign n2758 = ( n2746 & ~n2658 ) | ( n2746 & n2756 ) | ( ~n2658 & n2756 ) ;
  assign n2759 = ( n2757 & ~n2746 ) | ( n2757 & n2758 ) | ( ~n2746 & n2758 ) ;
  assign n2763 = x76 &  n1227 ;
  assign n2760 = ( x78 & ~n1154 ) | ( x78 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n2761 = x77 &  n1149 ;
  assign n2762 = n2760 | n2761 ;
  assign n2764 = ( x76 & ~n2763 ) | ( x76 & n2762 ) | ( ~n2763 & n2762 ) ;
  assign n2765 = ( n693 & ~n1157 ) | ( n693 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n2766 = n2764 | n2765 ;
  assign n2767 = ( x20 & ~n2766 ) | ( x20 & 1'b0 ) | ( ~n2766 & 1'b0 ) ;
  assign n2768 = ~x20 & n2766 ;
  assign n2769 = n2767 | n2768 ;
  assign n2770 = ( n2759 & ~n2661 ) | ( n2759 & n2769 ) | ( ~n2661 & n2769 ) ;
  assign n2771 = ( n2661 & ~n2769 ) | ( n2661 & n2759 ) | ( ~n2769 & n2759 ) ;
  assign n2772 = ( n2770 & ~n2759 ) | ( n2770 & n2771 ) | ( ~n2759 & n2771 ) ;
  assign n2783 = ( n2663 & n2673 ) | ( n2663 & n2674 ) | ( n2673 & n2674 ) ;
  assign n2776 = x79 &  n942 ;
  assign n2773 = ( x81 & ~n896 ) | ( x81 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n2774 = x80 &  n891 ;
  assign n2775 = n2773 | n2774 ;
  assign n2777 = ( x79 & ~n2776 ) | ( x79 & n2775 ) | ( ~n2776 & n2775 ) ;
  assign n2778 = ~n899 & n994 ;
  assign n2779 = n2777 | n2778 ;
  assign n2780 = ( x17 & ~n2779 ) | ( x17 & 1'b0 ) | ( ~n2779 & 1'b0 ) ;
  assign n2781 = ~x17 & n2779 ;
  assign n2782 = n2780 | n2781 ;
  assign n2784 = ( n2772 & ~n2783 ) | ( n2772 & n2782 ) | ( ~n2783 & n2782 ) ;
  assign n2785 = ( n2772 & ~n2782 ) | ( n2772 & n2783 ) | ( ~n2782 & n2783 ) ;
  assign n2786 = ( n2784 & ~n2772 ) | ( n2784 & n2785 ) | ( ~n2772 & n2785 ) ;
  assign n2797 = ( n2678 & ~n2796 ) | ( n2678 & n2786 ) | ( ~n2796 & n2786 ) ;
  assign n2798 = ( n2786 & ~n2678 ) | ( n2786 & n2796 ) | ( ~n2678 & n2796 ) ;
  assign n2799 = ( n2797 & ~n2786 ) | ( n2797 & n2798 ) | ( ~n2786 & n2798 ) ;
  assign n2803 = x85 &  n503 ;
  assign n2800 = ( x87 & ~n450 ) | ( x87 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n2801 = x86 &  n445 ;
  assign n2802 = n2800 | n2801 ;
  assign n2804 = ( x85 & ~n2803 ) | ( x85 & n2802 ) | ( ~n2803 & n2802 ) ;
  assign n2805 = ~n453 & n1512 ;
  assign n2806 = n2804 | n2805 ;
  assign n2807 = ( x11 & ~n2806 ) | ( x11 & 1'b0 ) | ( ~n2806 & 1'b0 ) ;
  assign n2808 = ~x11 & n2806 ;
  assign n2809 = n2807 | n2808 ;
  assign n2810 = ( n2799 & ~n2682 ) | ( n2799 & n2809 ) | ( ~n2682 & n2809 ) ;
  assign n2811 = ( n2682 & ~n2809 ) | ( n2682 & n2799 ) | ( ~n2809 & n2799 ) ;
  assign n2812 = ( n2810 & ~n2799 ) | ( n2810 & n2811 ) | ( ~n2799 & n2811 ) ;
  assign n2816 = x88 &  n353 ;
  assign n2813 = ( x90 & ~n313 ) | ( x90 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n2814 = x89 &  n308 ;
  assign n2815 = n2813 | n2814 ;
  assign n2817 = ( x88 & ~n2816 ) | ( x88 & n2815 ) | ( ~n2816 & n2815 ) ;
  assign n2818 = ~n316 & n1976 ;
  assign n2819 = n2817 | n2818 ;
  assign n2820 = ( x8 & ~n2819 ) | ( x8 & 1'b0 ) | ( ~n2819 & 1'b0 ) ;
  assign n2821 = ~x8 & n2819 ;
  assign n2822 = n2820 | n2821 ;
  assign n2823 = ( n2812 & ~n2686 ) | ( n2812 & n2822 ) | ( ~n2686 & n2822 ) ;
  assign n2824 = ( n2686 & ~n2822 ) | ( n2686 & n2812 ) | ( ~n2822 & n2812 ) ;
  assign n2825 = ( n2823 & ~n2812 ) | ( n2823 & n2824 ) | ( ~n2812 & n2824 ) ;
  assign n2827 = ( n2695 & n2705 ) | ( n2695 & n2825 ) | ( n2705 & n2825 ) ;
  assign n2826 = ( n2705 & ~n2695 ) | ( n2705 & n2825 ) | ( ~n2695 & n2825 ) ;
  assign n2828 = ( n2695 & ~n2827 ) | ( n2695 & n2826 ) | ( ~n2827 & n2826 ) ;
  assign n2842 = ( n2692 & ~n2841 ) | ( n2692 & n2828 ) | ( ~n2841 & n2828 ) ;
  assign n2843 = ( n2828 & ~n2692 ) | ( n2828 & n2841 ) | ( ~n2692 & n2841 ) ;
  assign n2844 = ( n2842 & ~n2828 ) | ( n2842 & n2843 ) | ( ~n2828 & n2843 ) ;
  assign n2845 = ( n2695 & ~n2705 ) | ( n2695 & n2825 ) | ( ~n2705 & n2825 ) ;
  assign n2849 = x92 &  n225 ;
  assign n2846 = ( x94 & ~n197 ) | ( x94 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n2847 = x93 &  n192 ;
  assign n2848 = n2846 | n2847 ;
  assign n2850 = ( x92 & ~n2849 ) | ( x92 & n2848 ) | ( ~n2849 & n2848 ) ;
  assign n2851 = ~n200 & n2401 ;
  assign n2852 = n2850 | n2851 ;
  assign n2853 = ( x5 & ~n2852 ) | ( x5 & 1'b0 ) | ( ~n2852 & 1'b0 ) ;
  assign n2854 = ~x5 & n2852 ;
  assign n2855 = n2853 | n2854 ;
  assign n2856 = ( x32 & ~x33 ) | ( x32 & 1'b0 ) | ( ~x33 & 1'b0 ) ;
  assign n2857 = ~x32 & x33 ;
  assign n2858 = n2856 | n2857 ;
  assign n2859 = x64 &  n2858 ;
  assign n2860 = ( n2430 & ~n2647 ) | ( n2430 & n2725 ) | ( ~n2647 & n2725 ) ;
  assign n2861 = ( x32 & n2647 ) | ( x32 & n2860 ) | ( n2647 & n2860 ) ;
  assign n2862 = ( x32 & ~n2861 ) | ( x32 & 1'b0 ) | ( ~n2861 & 1'b0 ) ;
  assign n2866 = x65 &  n2718 ;
  assign n2863 = ( x67 & ~n2642 ) | ( x67 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n2864 = x66 &  n2637 ;
  assign n2865 = n2863 | n2864 ;
  assign n2867 = ( x65 & ~n2866 ) | ( x65 & n2865 ) | ( ~n2866 & n2865 ) ;
  assign n2868 = n173 | n2645 ;
  assign n2869 = ~n2867 & n2868 ;
  assign n2870 = x32 &  n2869 ;
  assign n2871 = x32 | n2869 ;
  assign n2872 = ~n2870 & n2871 ;
  assign n2873 = ( n2859 & ~n2862 ) | ( n2859 & n2872 ) | ( ~n2862 & n2872 ) ;
  assign n2874 = ( n2859 & ~n2872 ) | ( n2859 & n2862 ) | ( ~n2872 & n2862 ) ;
  assign n2875 = ( n2873 & ~n2859 ) | ( n2873 & n2874 ) | ( ~n2859 & n2874 ) ;
  assign n2876 = ( n2652 & n2730 ) | ( n2652 & n2740 ) | ( n2730 & n2740 ) ;
  assign n2880 = x68 &  n2312 ;
  assign n2877 = ( x70 & ~n2195 ) | ( x70 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n2878 = x69 &  n2190 ;
  assign n2879 = n2877 | n2878 ;
  assign n2881 = ( x68 & ~n2880 ) | ( x68 & n2879 ) | ( ~n2880 & n2879 ) ;
  assign n2882 = ( n282 & ~n2198 ) | ( n282 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n2883 = n2881 | n2882 ;
  assign n2884 = ( x29 & ~n2883 ) | ( x29 & 1'b0 ) | ( ~n2883 & 1'b0 ) ;
  assign n2885 = ~x29 & n2883 ;
  assign n2886 = n2884 | n2885 ;
  assign n2887 = ( n2875 & ~n2876 ) | ( n2875 & n2886 ) | ( ~n2876 & n2886 ) ;
  assign n2888 = ( n2876 & ~n2875 ) | ( n2876 & n2886 ) | ( ~n2875 & n2886 ) ;
  assign n2889 = ( n2887 & ~n2886 ) | ( n2887 & n2888 ) | ( ~n2886 & n2888 ) ;
  assign n2894 = x71 &  n1894 ;
  assign n2891 = ( x73 & ~n1816 ) | ( x73 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n2892 = x72 &  n1811 ;
  assign n2893 = n2891 | n2892 ;
  assign n2895 = ( x71 & ~n2894 ) | ( x71 & n2893 ) | ( ~n2894 & n2893 ) ;
  assign n2896 = ( n389 & ~n1819 ) | ( n389 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n2897 = n2895 | n2896 ;
  assign n2898 = ( x26 & ~n2897 ) | ( x26 & 1'b0 ) | ( ~n2897 & 1'b0 ) ;
  assign n2899 = ~x26 & n2897 ;
  assign n2900 = n2898 | n2899 ;
  assign n2890 = ( n2655 & n2715 ) | ( n2655 & n2743 ) | ( n2715 & n2743 ) ;
  assign n2901 = ( n2889 & ~n2900 ) | ( n2889 & n2890 ) | ( ~n2900 & n2890 ) ;
  assign n2902 = ( n2889 & ~n2890 ) | ( n2889 & n2900 ) | ( ~n2890 & n2900 ) ;
  assign n2903 = ( n2901 & ~n2889 ) | ( n2901 & n2902 ) | ( ~n2889 & n2902 ) ;
  assign n2904 = ( n2658 & n2746 ) | ( n2658 & n2756 ) | ( n2746 & n2756 ) ;
  assign n2908 = x74 &  n1551 ;
  assign n2905 = ( x76 & ~n1451 ) | ( x76 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n2906 = x75 &  n1446 ;
  assign n2907 = n2905 | n2906 ;
  assign n2909 = ( x74 & ~n2908 ) | ( x74 & n2907 ) | ( ~n2908 & n2907 ) ;
  assign n2910 = ( n603 & ~n1454 ) | ( n603 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n2911 = n2909 | n2910 ;
  assign n2912 = ( x23 & ~n2911 ) | ( x23 & 1'b0 ) | ( ~n2911 & 1'b0 ) ;
  assign n2913 = ~x23 & n2911 ;
  assign n2914 = n2912 | n2913 ;
  assign n2915 = ( n2903 & ~n2904 ) | ( n2903 & n2914 ) | ( ~n2904 & n2914 ) ;
  assign n2916 = ( n2903 & ~n2914 ) | ( n2903 & n2904 ) | ( ~n2914 & n2904 ) ;
  assign n2917 = ( n2915 & ~n2903 ) | ( n2915 & n2916 ) | ( ~n2903 & n2916 ) ;
  assign n2918 = ( n2661 & n2759 ) | ( n2661 & n2769 ) | ( n2759 & n2769 ) ;
  assign n2922 = x77 &  n1227 ;
  assign n2919 = ( x79 & ~n1154 ) | ( x79 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n2920 = x78 &  n1149 ;
  assign n2921 = n2919 | n2920 ;
  assign n2923 = ( x77 & ~n2922 ) | ( x77 & n2921 ) | ( ~n2922 & n2921 ) ;
  assign n2924 = ( n766 & ~n1157 ) | ( n766 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n2925 = n2923 | n2924 ;
  assign n2926 = ( x20 & ~n2925 ) | ( x20 & 1'b0 ) | ( ~n2925 & 1'b0 ) ;
  assign n2927 = ~x20 & n2925 ;
  assign n2928 = n2926 | n2927 ;
  assign n2929 = ( n2917 & ~n2918 ) | ( n2917 & n2928 ) | ( ~n2918 & n2928 ) ;
  assign n2930 = ( n2918 & ~n2917 ) | ( n2918 & n2928 ) | ( ~n2917 & n2928 ) ;
  assign n2931 = ( n2929 & ~n2928 ) | ( n2929 & n2930 ) | ( ~n2928 & n2930 ) ;
  assign n2936 = x80 &  n942 ;
  assign n2933 = ( x82 & ~n896 ) | ( x82 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n2934 = x81 &  n891 ;
  assign n2935 = n2933 | n2934 ;
  assign n2937 = ( x80 & ~n2936 ) | ( x80 & n2935 ) | ( ~n2936 & n2935 ) ;
  assign n2938 = ~n899 & n1084 ;
  assign n2939 = n2937 | n2938 ;
  assign n2940 = ( x17 & ~n2939 ) | ( x17 & 1'b0 ) | ( ~n2939 & 1'b0 ) ;
  assign n2941 = ~x17 & n2939 ;
  assign n2942 = n2940 | n2941 ;
  assign n2932 = ( n2772 & n2782 ) | ( n2772 & n2783 ) | ( n2782 & n2783 ) ;
  assign n2943 = ( n2931 & ~n2942 ) | ( n2931 & n2932 ) | ( ~n2942 & n2932 ) ;
  assign n2944 = ( n2931 & ~n2932 ) | ( n2931 & n2942 ) | ( ~n2932 & n2942 ) ;
  assign n2945 = ( n2943 & ~n2931 ) | ( n2943 & n2944 ) | ( ~n2931 & n2944 ) ;
  assign n2946 = ( n2678 & n2786 ) | ( n2678 & n2796 ) | ( n2786 & n2796 ) ;
  assign n2950 = x83 &  n713 ;
  assign n2947 = ( x85 & ~n641 ) | ( x85 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n2948 = x84 &  n636 ;
  assign n2949 = n2947 | n2948 ;
  assign n2951 = ( x83 & ~n2950 ) | ( x83 & n2949 ) | ( ~n2950 & n2949 ) ;
  assign n2952 = ~n644 & n1295 ;
  assign n2953 = n2951 | n2952 ;
  assign n2954 = ( x14 & ~n2953 ) | ( x14 & 1'b0 ) | ( ~n2953 & 1'b0 ) ;
  assign n2955 = ~x14 & n2953 ;
  assign n2956 = n2954 | n2955 ;
  assign n2957 = ( n2945 & ~n2946 ) | ( n2945 & n2956 ) | ( ~n2946 & n2956 ) ;
  assign n2958 = ( n2945 & ~n2956 ) | ( n2945 & n2946 ) | ( ~n2956 & n2946 ) ;
  assign n2959 = ( n2957 & ~n2945 ) | ( n2957 & n2958 ) | ( ~n2945 & n2958 ) ;
  assign n2964 = x86 &  n503 ;
  assign n2961 = ( x88 & ~n450 ) | ( x88 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n2962 = x87 &  n445 ;
  assign n2963 = n2961 | n2962 ;
  assign n2965 = ( x86 & ~n2964 ) | ( x86 & n2963 ) | ( ~n2964 & n2963 ) ;
  assign n2966 = ~n453 & n1624 ;
  assign n2967 = n2965 | n2966 ;
  assign n2968 = ( x11 & ~n2967 ) | ( x11 & 1'b0 ) | ( ~n2967 & 1'b0 ) ;
  assign n2969 = ~x11 & n2967 ;
  assign n2970 = n2968 | n2969 ;
  assign n2960 = ( n2682 & n2799 ) | ( n2682 & n2809 ) | ( n2799 & n2809 ) ;
  assign n2971 = ( n2959 & ~n2970 ) | ( n2959 & n2960 ) | ( ~n2970 & n2960 ) ;
  assign n2972 = ( n2959 & ~n2960 ) | ( n2959 & n2970 ) | ( ~n2960 & n2970 ) ;
  assign n2973 = ( n2971 & ~n2959 ) | ( n2971 & n2972 ) | ( ~n2959 & n2972 ) ;
  assign n2977 = x89 &  n353 ;
  assign n2974 = ( x91 & ~n313 ) | ( x91 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n2975 = x90 &  n308 ;
  assign n2976 = n2974 | n2975 ;
  assign n2978 = ( x89 & ~n2977 ) | ( x89 & n2976 ) | ( ~n2977 & n2976 ) ;
  assign n2979 = ~n316 & n2108 ;
  assign n2980 = n2978 | n2979 ;
  assign n2981 = ( x8 & ~n2980 ) | ( x8 & 1'b0 ) | ( ~n2980 & 1'b0 ) ;
  assign n2982 = ~x8 & n2980 ;
  assign n2983 = n2981 | n2982 ;
  assign n2984 = ( n2686 & n2812 ) | ( n2686 & n2822 ) | ( n2812 & n2822 ) ;
  assign n2985 = ( n2973 & ~n2983 ) | ( n2973 & n2984 ) | ( ~n2983 & n2984 ) ;
  assign n2986 = ( n2973 & ~n2984 ) | ( n2973 & n2983 ) | ( ~n2984 & n2983 ) ;
  assign n2987 = ( n2985 & ~n2973 ) | ( n2985 & n2986 ) | ( ~n2973 & n2986 ) ;
  assign n2988 = ( n2845 & n2855 ) | ( n2845 & n2987 ) | ( n2855 & n2987 ) ;
  assign n2989 = ( n2855 & ~n2845 ) | ( n2855 & n2987 ) | ( ~n2845 & n2987 ) ;
  assign n2990 = ( n2845 & ~n2988 ) | ( n2845 & n2989 ) | ( ~n2988 & n2989 ) ;
  assign n2995 = ~n136 & x97 ;
  assign n2992 = ( x95 & ~n150 ) | ( x95 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n2993 = ( x96 & ~n131 ) | ( x96 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n2994 = n2992 | n2993 ;
  assign n2996 = ( x97 & ~n2995 ) | ( x97 & n2994 ) | ( ~n2995 & n2994 ) ;
  assign n2998 = ( x96 & x97 ) | ( x96 & n2835 ) | ( x97 & n2835 ) ;
  assign n2997 = ( x96 & ~x97 ) | ( x96 & n2835 ) | ( ~x97 & n2835 ) ;
  assign n2999 = ( x97 & ~n2998 ) | ( x97 & n2997 ) | ( ~n2998 & n2997 ) ;
  assign n3000 = ( n139 & ~n2996 ) | ( n139 & n2999 ) | ( ~n2996 & n2999 ) ;
  assign n3001 = ~n139 & n3000 ;
  assign n3002 = ( x2 & n2996 ) | ( x2 & n3001 ) | ( n2996 & n3001 ) ;
  assign n3003 = ( x2 & ~n3001 ) | ( x2 & n2996 ) | ( ~n3001 & n2996 ) ;
  assign n3004 = ( n3001 & ~n3002 ) | ( n3001 & n3003 ) | ( ~n3002 & n3003 ) ;
  assign n2991 = ( n2692 & ~n2828 ) | ( n2692 & n2841 ) | ( ~n2828 & n2841 ) ;
  assign n3005 = ( n2990 & ~n3004 ) | ( n2990 & n2991 ) | ( ~n3004 & n2991 ) ;
  assign n3006 = ( n2990 & ~n2991 ) | ( n2990 & n3004 ) | ( ~n2991 & n3004 ) ;
  assign n3007 = ( n3005 & ~n2990 ) | ( n3005 & n3006 ) | ( ~n2990 & n3006 ) ;
  assign n3008 = ( n2845 & ~n2987 ) | ( n2845 & n2855 ) | ( ~n2987 & n2855 ) ;
  assign n3022 = x90 &  n353 ;
  assign n3019 = ( x92 & ~n313 ) | ( x92 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n3020 = x91 &  n308 ;
  assign n3021 = n3019 | n3020 ;
  assign n3023 = ( x90 & ~n3022 ) | ( x90 & n3021 ) | ( ~n3022 & n3021 ) ;
  assign n3024 = ~n316 & n2248 ;
  assign n3025 = n3023 | n3024 ;
  assign n3026 = ( x8 & ~n3025 ) | ( x8 & 1'b0 ) | ( ~n3025 & 1'b0 ) ;
  assign n3027 = ~x8 & n3025 ;
  assign n3028 = n3026 | n3027 ;
  assign n3032 = x84 &  n713 ;
  assign n3029 = ( x86 & ~n641 ) | ( x86 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n3030 = x85 &  n636 ;
  assign n3031 = n3029 | n3030 ;
  assign n3033 = ( x84 & ~n3032 ) | ( x84 & n3031 ) | ( ~n3032 & n3031 ) ;
  assign n3034 = ~n644 & n1496 ;
  assign n3035 = n3033 | n3034 ;
  assign n3036 = ( x14 & ~n3035 ) | ( x14 & 1'b0 ) | ( ~n3035 & 1'b0 ) ;
  assign n3037 = ~x14 & n3035 ;
  assign n3038 = n3036 | n3037 ;
  assign n3042 = x81 &  n942 ;
  assign n3039 = ( x83 & ~n896 ) | ( x83 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n3040 = x82 &  n891 ;
  assign n3041 = n3039 | n3040 ;
  assign n3043 = ( x81 & ~n3042 ) | ( x81 & n3041 ) | ( ~n3042 & n3041 ) ;
  assign n3044 = ~n899 & n1100 ;
  assign n3045 = n3043 | n3044 ;
  assign n3046 = ( x17 & ~n3045 ) | ( x17 & 1'b0 ) | ( ~n3045 & 1'b0 ) ;
  assign n3047 = ~x17 & n3045 ;
  assign n3048 = n3046 | n3047 ;
  assign n3062 = x69 &  n2312 ;
  assign n3059 = ( x71 & ~n2195 ) | ( x71 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n3060 = x70 &  n2190 ;
  assign n3061 = n3059 | n3060 ;
  assign n3063 = ( x69 & ~n3062 ) | ( x69 & n3061 ) | ( ~n3062 & n3061 ) ;
  assign n3064 = ( n298 & ~n2198 ) | ( n298 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n3065 = n3063 | n3064 ;
  assign n3066 = ( x29 & ~n3065 ) | ( x29 & 1'b0 ) | ( ~n3065 & 1'b0 ) ;
  assign n3067 = ~x29 & n3065 ;
  assign n3068 = n3066 | n3067 ;
  assign n3072 = x66 &  n2718 ;
  assign n3069 = ( x68 & ~n2642 ) | ( x68 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n3070 = x67 &  n2637 ;
  assign n3071 = n3069 | n3070 ;
  assign n3073 = ( x66 & ~n3072 ) | ( x66 & n3071 ) | ( ~n3072 & n3071 ) ;
  assign n3074 = ( n213 & ~n2645 ) | ( n213 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n3075 = n3073 | n3074 ;
  assign n3076 = ( x32 & ~n3075 ) | ( x32 & 1'b0 ) | ( ~n3075 & 1'b0 ) ;
  assign n3077 = ~x32 & n3075 ;
  assign n3078 = n3076 | n3077 ;
  assign n3079 = ( x35 & ~n2859 ) | ( x35 & 1'b0 ) | ( ~n2859 & 1'b0 ) ;
  assign n3080 = ( x33 & x34 ) | ( x33 & n2856 ) | ( x34 & n2856 ) ;
  assign n3081 = ( x33 & ~n2857 ) | ( x33 & x34 ) | ( ~n2857 & x34 ) ;
  assign n3082 = ~n3080 &  n3081 ;
  assign n3083 = x64 &  n3082 ;
  assign n3084 = ~x34 & x35 ;
  assign n3085 = ( x34 & ~x35 ) | ( x34 & 1'b0 ) | ( ~x35 & 1'b0 ) ;
  assign n3086 = n3084 | n3085 ;
  assign n3087 = ~n2858 |  n3086 ;
  assign n3088 = ( x65 & ~n3087 ) | ( x65 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n3089 = n3083 | n3088 ;
  assign n3090 = ~n2858 | ~n3086 ;
  assign n3091 = ( n142 & ~n3090 ) | ( n142 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n3092 = n3089 | n3091 ;
  assign n3094 = ( x35 & n3079 ) | ( x35 & n3092 ) | ( n3079 & n3092 ) ;
  assign n3093 = ( x35 & ~n3079 ) | ( x35 & n3092 ) | ( ~n3079 & n3092 ) ;
  assign n3095 = ( n3079 & ~n3094 ) | ( n3079 & n3093 ) | ( ~n3094 & n3093 ) ;
  assign n3097 = ( n2874 & n3078 ) | ( n2874 & n3095 ) | ( n3078 & n3095 ) ;
  assign n3096 = ( n2874 & ~n3078 ) | ( n2874 & n3095 ) | ( ~n3078 & n3095 ) ;
  assign n3098 = ( n3078 & ~n3097 ) | ( n3078 & n3096 ) | ( ~n3097 & n3096 ) ;
  assign n3100 = ( n2888 & n3068 ) | ( n2888 & n3098 ) | ( n3068 & n3098 ) ;
  assign n3099 = ( n2888 & ~n3068 ) | ( n2888 & n3098 ) | ( ~n3068 & n3098 ) ;
  assign n3101 = ( n3068 & ~n3100 ) | ( n3068 & n3099 ) | ( ~n3100 & n3099 ) ;
  assign n3112 = ( n2890 & ~n2889 ) | ( n2890 & n2900 ) | ( ~n2889 & n2900 ) ;
  assign n3105 = x72 &  n1894 ;
  assign n3102 = ( x74 & ~n1816 ) | ( x74 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n3103 = x73 &  n1811 ;
  assign n3104 = n3102 | n3103 ;
  assign n3106 = ( x72 & ~n3105 ) | ( x72 & n3104 ) | ( ~n3105 & n3104 ) ;
  assign n3107 = ( n482 & ~n1819 ) | ( n482 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n3108 = n3106 | n3107 ;
  assign n3109 = ( x26 & ~n3108 ) | ( x26 & 1'b0 ) | ( ~n3108 & 1'b0 ) ;
  assign n3110 = ~x26 & n3108 ;
  assign n3111 = n3109 | n3110 ;
  assign n3113 = ( n3101 & ~n3112 ) | ( n3101 & n3111 ) | ( ~n3112 & n3111 ) ;
  assign n3114 = ( n3101 & ~n3111 ) | ( n3101 & n3112 ) | ( ~n3111 & n3112 ) ;
  assign n3115 = ( n3113 & ~n3101 ) | ( n3113 & n3114 ) | ( ~n3101 & n3114 ) ;
  assign n3120 = x75 &  n1551 ;
  assign n3117 = ( x77 & ~n1451 ) | ( x77 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n3118 = x76 &  n1446 ;
  assign n3119 = n3117 | n3118 ;
  assign n3121 = ( x75 & ~n3120 ) | ( x75 & n3119 ) | ( ~n3120 & n3119 ) ;
  assign n3122 = ( n677 & ~n1454 ) | ( n677 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n3123 = n3121 | n3122 ;
  assign n3124 = ( x23 & ~n3123 ) | ( x23 & 1'b0 ) | ( ~n3123 & 1'b0 ) ;
  assign n3125 = ~x23 & n3123 ;
  assign n3126 = n3124 | n3125 ;
  assign n3116 = ( n2904 & ~n2903 ) | ( n2904 & n2914 ) | ( ~n2903 & n2914 ) ;
  assign n3127 = ( n3115 & ~n3126 ) | ( n3115 & n3116 ) | ( ~n3126 & n3116 ) ;
  assign n3128 = ( n3115 & ~n3116 ) | ( n3115 & n3126 ) | ( ~n3116 & n3126 ) ;
  assign n3129 = ( n3127 & ~n3115 ) | ( n3127 & n3128 ) | ( ~n3115 & n3128 ) ;
  assign n3052 = x78 &  n1227 ;
  assign n3049 = ( x80 & ~n1154 ) | ( x80 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n3050 = x79 &  n1149 ;
  assign n3051 = n3049 | n3050 ;
  assign n3053 = ( x78 & ~n3052 ) | ( x78 & n3051 ) | ( ~n3052 & n3051 ) ;
  assign n3054 = ( n842 & ~n1157 ) | ( n842 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n3055 = n3053 | n3054 ;
  assign n3056 = ( x20 & ~n3055 ) | ( x20 & 1'b0 ) | ( ~n3055 & 1'b0 ) ;
  assign n3057 = ~x20 & n3055 ;
  assign n3058 = n3056 | n3057 ;
  assign n3130 = ( n2930 & ~n3129 ) | ( n2930 & n3058 ) | ( ~n3129 & n3058 ) ;
  assign n3131 = ( n3058 & ~n2930 ) | ( n3058 & n3129 ) | ( ~n2930 & n3129 ) ;
  assign n3132 = ( n3130 & ~n3058 ) | ( n3130 & n3131 ) | ( ~n3058 & n3131 ) ;
  assign n3133 = ( n2932 & ~n2931 ) | ( n2932 & n2942 ) | ( ~n2931 & n2942 ) ;
  assign n3134 = ( n3048 & n3132 ) | ( n3048 & n3133 ) | ( n3132 & n3133 ) ;
  assign n3135 = ( n3132 & ~n3048 ) | ( n3132 & n3133 ) | ( ~n3048 & n3133 ) ;
  assign n3136 = ( n3048 & ~n3134 ) | ( n3048 & n3135 ) | ( ~n3134 & n3135 ) ;
  assign n3137 = ( n2946 & ~n2945 ) | ( n2946 & n2956 ) | ( ~n2945 & n2956 ) ;
  assign n3138 = ( n3038 & n3136 ) | ( n3038 & n3137 ) | ( n3136 & n3137 ) ;
  assign n3139 = ( n3136 & ~n3038 ) | ( n3136 & n3137 ) | ( ~n3038 & n3137 ) ;
  assign n3140 = ( n3038 & ~n3138 ) | ( n3038 & n3139 ) | ( ~n3138 & n3139 ) ;
  assign n3145 = x87 &  n503 ;
  assign n3142 = ( x89 & ~n450 ) | ( x89 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n3143 = x88 &  n445 ;
  assign n3144 = n3142 | n3143 ;
  assign n3146 = ( x87 & ~n3145 ) | ( x87 & n3144 ) | ( ~n3145 & n3144 ) ;
  assign n3147 = ~n453 & n1741 ;
  assign n3148 = n3146 | n3147 ;
  assign n3149 = ( x11 & ~n3148 ) | ( x11 & 1'b0 ) | ( ~n3148 & 1'b0 ) ;
  assign n3150 = ~x11 & n3148 ;
  assign n3151 = n3149 | n3150 ;
  assign n3141 = ( n2960 & ~n2959 ) | ( n2960 & n2970 ) | ( ~n2959 & n2970 ) ;
  assign n3152 = ( n3140 & ~n3151 ) | ( n3140 & n3141 ) | ( ~n3151 & n3141 ) ;
  assign n3153 = ( n3140 & ~n3141 ) | ( n3140 & n3151 ) | ( ~n3141 & n3151 ) ;
  assign n3154 = ( n3152 & ~n3140 ) | ( n3152 & n3153 ) | ( ~n3140 & n3153 ) ;
  assign n3155 = ( n2983 & ~n2973 ) | ( n2983 & n2984 ) | ( ~n2973 & n2984 ) ;
  assign n3156 = ( n3028 & ~n3154 ) | ( n3028 & n3155 ) | ( ~n3154 & n3155 ) ;
  assign n3157 = ( n3028 & ~n3155 ) | ( n3028 & n3154 ) | ( ~n3155 & n3154 ) ;
  assign n3158 = ( n3156 & ~n3028 ) | ( n3156 & n3157 ) | ( ~n3028 & n3157 ) ;
  assign n3012 = x93 &  n225 ;
  assign n3009 = ( x95 & ~n197 ) | ( x95 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n3010 = x94 &  n192 ;
  assign n3011 = n3009 | n3010 ;
  assign n3013 = ( x93 & ~n3012 ) | ( x93 & n3011 ) | ( ~n3012 & n3011 ) ;
  assign n3014 = ~n200 & n2547 ;
  assign n3015 = n3013 | n3014 ;
  assign n3016 = ( x5 & ~n3015 ) | ( x5 & 1'b0 ) | ( ~n3015 & 1'b0 ) ;
  assign n3017 = ~x5 & n3015 ;
  assign n3018 = n3016 | n3017 ;
  assign n3159 = ( n3008 & ~n3158 ) | ( n3008 & n3018 ) | ( ~n3158 & n3018 ) ;
  assign n3160 = ( n3008 & ~n3018 ) | ( n3008 & n3158 ) | ( ~n3018 & n3158 ) ;
  assign n3161 = ( n3159 & ~n3008 ) | ( n3159 & n3160 ) | ( ~n3008 & n3160 ) ;
  assign n3162 = ( n2991 & ~n2990 ) | ( n2991 & n3004 ) | ( ~n2990 & n3004 ) ;
  assign n3166 = ~n136 & x98 ;
  assign n3163 = ( x96 & ~n150 ) | ( x96 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n3164 = ( x97 & ~n131 ) | ( x97 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n3165 = n3163 | n3164 ;
  assign n3167 = ( x98 & ~n3166 ) | ( x98 & n3165 ) | ( ~n3166 & n3165 ) ;
  assign n3169 = ( x97 & x98 ) | ( x97 & n2998 ) | ( x98 & n2998 ) ;
  assign n3168 = ( x97 & ~x98 ) | ( x97 & n2998 ) | ( ~x98 & n2998 ) ;
  assign n3170 = ( x98 & ~n3169 ) | ( x98 & n3168 ) | ( ~n3169 & n3168 ) ;
  assign n3171 = ( n139 & ~n3167 ) | ( n139 & n3170 ) | ( ~n3167 & n3170 ) ;
  assign n3172 = ~n139 & n3171 ;
  assign n3173 = ( x2 & n3167 ) | ( x2 & n3172 ) | ( n3167 & n3172 ) ;
  assign n3174 = ( x2 & ~n3172 ) | ( x2 & n3167 ) | ( ~n3172 & n3167 ) ;
  assign n3175 = ( n3172 & ~n3173 ) | ( n3172 & n3174 ) | ( ~n3173 & n3174 ) ;
  assign n3176 = ( n3161 & ~n3162 ) | ( n3161 & n3175 ) | ( ~n3162 & n3175 ) ;
  assign n3177 = ( n3161 & ~n3175 ) | ( n3161 & n3162 ) | ( ~n3175 & n3162 ) ;
  assign n3178 = ( n3176 & ~n3161 ) | ( n3176 & n3177 ) | ( ~n3161 & n3177 ) ;
  assign n3179 = ( n3008 & n3018 ) | ( n3008 & n3158 ) | ( n3018 & n3158 ) ;
  assign n3183 = x94 &  n225 ;
  assign n3180 = ( x96 & ~n197 ) | ( x96 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n3181 = x95 &  n192 ;
  assign n3182 = n3180 | n3181 ;
  assign n3184 = ( x94 & ~n3183 ) | ( x94 & n3182 ) | ( ~n3183 & n3182 ) ;
  assign n3185 = ~n200 & n2836 ;
  assign n3186 = n3184 | n3185 ;
  assign n3187 = ( x5 & ~n3186 ) | ( x5 & 1'b0 ) | ( ~n3186 & 1'b0 ) ;
  assign n3188 = ~x5 & n3186 ;
  assign n3189 = n3187 | n3188 ;
  assign n3193 = x88 &  n503 ;
  assign n3190 = ( x90 & ~n450 ) | ( x90 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n3191 = x89 &  n445 ;
  assign n3192 = n3190 | n3191 ;
  assign n3194 = ( x88 & ~n3193 ) | ( x88 & n3192 ) | ( ~n3193 & n3192 ) ;
  assign n3195 = ~n453 & n1976 ;
  assign n3196 = n3194 | n3195 ;
  assign n3197 = ( x11 & ~n3196 ) | ( x11 & 1'b0 ) | ( ~n3196 & 1'b0 ) ;
  assign n3198 = ~x11 & n3196 ;
  assign n3199 = n3197 | n3198 ;
  assign n3200 = ( n3140 & n3141 ) | ( n3140 & n3151 ) | ( n3141 & n3151 ) ;
  assign n3287 = x82 &  n942 ;
  assign n3284 = ( x84 & ~n896 ) | ( x84 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n3285 = x83 &  n891 ;
  assign n3286 = n3284 | n3285 ;
  assign n3288 = ( x82 & ~n3287 ) | ( x82 & n3286 ) | ( ~n3287 & n3286 ) ;
  assign n3289 = ~n899 & n1199 ;
  assign n3290 = n3288 | n3289 ;
  assign n3291 = ( x17 & ~n3290 ) | ( x17 & 1'b0 ) | ( ~n3290 & 1'b0 ) ;
  assign n3292 = ~x17 & n3290 ;
  assign n3293 = n3291 | n3292 ;
  assign n3204 = x73 &  n1894 ;
  assign n3201 = ( x75 & ~n1816 ) | ( x75 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n3202 = x74 &  n1811 ;
  assign n3203 = n3201 | n3202 ;
  assign n3205 = ( x73 & ~n3204 ) | ( x73 & n3203 ) | ( ~n3204 & n3203 ) ;
  assign n3206 = ( n540 & ~n1819 ) | ( n540 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n3207 = n3205 | n3206 ;
  assign n3208 = ( x26 & ~n3207 ) | ( x26 & 1'b0 ) | ( ~n3207 & 1'b0 ) ;
  assign n3209 = ~x26 & n3207 ;
  assign n3210 = n3208 | n3209 ;
  assign n3211 = ( n3101 & n3111 ) | ( n3101 & n3112 ) | ( n3111 & n3112 ) ;
  assign n3230 = x67 &  n2718 ;
  assign n3227 = ( x69 & ~n2642 ) | ( x69 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n3228 = x68 &  n2637 ;
  assign n3229 = n3227 | n3228 ;
  assign n3231 = ( x67 & ~n3230 ) | ( x67 & n3229 ) | ( ~n3230 & n3229 ) ;
  assign n3232 = ( n246 & ~n2645 ) | ( n246 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n3233 = n3231 | n3232 ;
  assign n3234 = ( x32 & ~n3233 ) | ( x32 & 1'b0 ) | ( ~n3233 & 1'b0 ) ;
  assign n3235 = ~x32 & n3233 ;
  assign n3236 = n3234 | n3235 ;
  assign n3213 = ( x33 & ~x34 ) | ( x33 & n3086 ) | ( ~x34 & n3086 ) ;
  assign n3212 = ( x33 & ~x34 ) | ( x33 & n2858 ) | ( ~x34 & n2858 ) ;
  assign n3214 = ~n3213 |  n3212 ;
  assign n3218 = x64 &  n3214 ;
  assign n3215 = ( x66 & ~n3087 ) | ( x66 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n3216 = x65 &  n3082 ;
  assign n3217 = n3215 | n3216 ;
  assign n3219 = ( x64 & ~n3218 ) | ( x64 & n3217 ) | ( ~n3218 & n3217 ) ;
  assign n3220 = ( n157 & ~n3090 ) | ( n157 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n3221 = n3219 | n3220 ;
  assign n3222 = ( x35 & ~n2859 ) | ( x35 & n3092 ) | ( ~n2859 & n3092 ) ;
  assign n3223 = ~n3092 & n3222 ;
  assign n3224 = ( n3221 & ~x35 ) | ( n3221 & n3223 ) | ( ~x35 & n3223 ) ;
  assign n3225 = ( x35 & ~n3221 ) | ( x35 & n3223 ) | ( ~n3221 & n3223 ) ;
  assign n3226 = ( n3224 & ~n3223 ) | ( n3224 & n3225 ) | ( ~n3223 & n3225 ) ;
  assign n3237 = ( n3097 & ~n3236 ) | ( n3097 & n3226 ) | ( ~n3236 & n3226 ) ;
  assign n3238 = ( n3226 & ~n3097 ) | ( n3226 & n3236 ) | ( ~n3097 & n3236 ) ;
  assign n3239 = ( n3237 & ~n3226 ) | ( n3237 & n3238 ) | ( ~n3226 & n3238 ) ;
  assign n3243 = x70 &  n2312 ;
  assign n3240 = ( x72 & ~n2195 ) | ( x72 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n3241 = x71 &  n2190 ;
  assign n3242 = n3240 | n3241 ;
  assign n3244 = ( x70 & ~n3243 ) | ( x70 & n3242 ) | ( ~n3243 & n3242 ) ;
  assign n3245 = ( n345 & ~n2198 ) | ( n345 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n3246 = n3244 | n3245 ;
  assign n3247 = ( x29 & ~n3246 ) | ( x29 & 1'b0 ) | ( ~n3246 & 1'b0 ) ;
  assign n3248 = ~x29 & n3246 ;
  assign n3249 = n3247 | n3248 ;
  assign n3250 = ( n3239 & ~n3100 ) | ( n3239 & n3249 ) | ( ~n3100 & n3249 ) ;
  assign n3251 = ( n3100 & ~n3249 ) | ( n3100 & n3239 ) | ( ~n3249 & n3239 ) ;
  assign n3252 = ( n3250 & ~n3239 ) | ( n3250 & n3251 ) | ( ~n3239 & n3251 ) ;
  assign n3254 = ( n3210 & n3211 ) | ( n3210 & n3252 ) | ( n3211 & n3252 ) ;
  assign n3253 = ( n3211 & ~n3210 ) | ( n3211 & n3252 ) | ( ~n3210 & n3252 ) ;
  assign n3255 = ( n3210 & ~n3254 ) | ( n3210 & n3253 ) | ( ~n3254 & n3253 ) ;
  assign n3256 = ( n3115 & n3116 ) | ( n3115 & n3126 ) | ( n3116 & n3126 ) ;
  assign n3260 = x76 &  n1551 ;
  assign n3257 = ( x78 & ~n1451 ) | ( x78 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n3258 = x77 &  n1446 ;
  assign n3259 = n3257 | n3258 ;
  assign n3261 = ( x76 & ~n3260 ) | ( x76 & n3259 ) | ( ~n3260 & n3259 ) ;
  assign n3262 = ( n693 & ~n1454 ) | ( n693 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n3263 = n3261 | n3262 ;
  assign n3264 = ( x23 & ~n3263 ) | ( x23 & 1'b0 ) | ( ~n3263 & 1'b0 ) ;
  assign n3265 = ~x23 & n3263 ;
  assign n3266 = n3264 | n3265 ;
  assign n3267 = ( n3255 & ~n3256 ) | ( n3255 & n3266 ) | ( ~n3256 & n3266 ) ;
  assign n3268 = ( n3255 & ~n3266 ) | ( n3255 & n3256 ) | ( ~n3266 & n3256 ) ;
  assign n3269 = ( n3267 & ~n3255 ) | ( n3267 & n3268 ) | ( ~n3255 & n3268 ) ;
  assign n3280 = ( n2930 & n3058 ) | ( n2930 & n3129 ) | ( n3058 & n3129 ) ;
  assign n3273 = x79 &  n1227 ;
  assign n3270 = ( x81 & ~n1154 ) | ( x81 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n3271 = x80 &  n1149 ;
  assign n3272 = n3270 | n3271 ;
  assign n3274 = ( x79 & ~n3273 ) | ( x79 & n3272 ) | ( ~n3273 & n3272 ) ;
  assign n3275 = ( n994 & ~n1157 ) | ( n994 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n3276 = n3274 | n3275 ;
  assign n3277 = ( x20 & ~n3276 ) | ( x20 & 1'b0 ) | ( ~n3276 & 1'b0 ) ;
  assign n3278 = ~x20 & n3276 ;
  assign n3279 = n3277 | n3278 ;
  assign n3281 = ( n3269 & ~n3280 ) | ( n3269 & n3279 ) | ( ~n3280 & n3279 ) ;
  assign n3282 = ( n3269 & ~n3279 ) | ( n3269 & n3280 ) | ( ~n3279 & n3280 ) ;
  assign n3283 = ( n3281 & ~n3269 ) | ( n3281 & n3282 ) | ( ~n3269 & n3282 ) ;
  assign n3294 = ( n3134 & ~n3293 ) | ( n3134 & n3283 ) | ( ~n3293 & n3283 ) ;
  assign n3295 = ( n3283 & ~n3134 ) | ( n3283 & n3293 ) | ( ~n3134 & n3293 ) ;
  assign n3296 = ( n3294 & ~n3283 ) | ( n3294 & n3295 ) | ( ~n3283 & n3295 ) ;
  assign n3300 = x85 &  n713 ;
  assign n3297 = ( x87 & ~n641 ) | ( x87 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n3298 = x86 &  n636 ;
  assign n3299 = n3297 | n3298 ;
  assign n3301 = ( x85 & ~n3300 ) | ( x85 & n3299 ) | ( ~n3300 & n3299 ) ;
  assign n3302 = ~n644 & n1512 ;
  assign n3303 = n3301 | n3302 ;
  assign n3304 = ( x14 & ~n3303 ) | ( x14 & 1'b0 ) | ( ~n3303 & 1'b0 ) ;
  assign n3305 = ~x14 & n3303 ;
  assign n3306 = n3304 | n3305 ;
  assign n3307 = ( n3296 & ~n3138 ) | ( n3296 & n3306 ) | ( ~n3138 & n3306 ) ;
  assign n3308 = ( n3138 & ~n3306 ) | ( n3138 & n3296 ) | ( ~n3306 & n3296 ) ;
  assign n3309 = ( n3307 & ~n3296 ) | ( n3307 & n3308 ) | ( ~n3296 & n3308 ) ;
  assign n3311 = ( n3199 & n3200 ) | ( n3199 & n3309 ) | ( n3200 & n3309 ) ;
  assign n3310 = ( n3200 & ~n3199 ) | ( n3200 & n3309 ) | ( ~n3199 & n3309 ) ;
  assign n3312 = ( n3199 & ~n3311 ) | ( n3199 & n3310 ) | ( ~n3311 & n3310 ) ;
  assign n3316 = x91 &  n353 ;
  assign n3313 = ( x93 & ~n313 ) | ( x93 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n3314 = x92 &  n308 ;
  assign n3315 = n3313 | n3314 ;
  assign n3317 = ( x91 & ~n3316 ) | ( x91 & n3315 ) | ( ~n3316 & n3315 ) ;
  assign n3318 = n316 | n2264 ;
  assign n3319 = ~n3317 & n3318 ;
  assign n3320 = x8 &  n3319 ;
  assign n3321 = x8 | n3319 ;
  assign n3322 = ~n3320 & n3321 ;
  assign n3323 = ( n3028 & n3154 ) | ( n3028 & n3155 ) | ( n3154 & n3155 ) ;
  assign n3325 = ( n3312 & n3322 ) | ( n3312 & n3323 ) | ( n3322 & n3323 ) ;
  assign n3324 = ( n3322 & ~n3312 ) | ( n3322 & n3323 ) | ( ~n3312 & n3323 ) ;
  assign n3326 = ( n3312 & ~n3325 ) | ( n3312 & n3324 ) | ( ~n3325 & n3324 ) ;
  assign n3327 = ( n3179 & n3189 ) | ( n3179 & n3326 ) | ( n3189 & n3326 ) ;
  assign n3328 = ( n3189 & ~n3179 ) | ( n3189 & n3326 ) | ( ~n3179 & n3326 ) ;
  assign n3329 = ( n3179 & ~n3327 ) | ( n3179 & n3328 ) | ( ~n3327 & n3328 ) ;
  assign n3334 = ~n136 & x99 ;
  assign n3331 = ( x97 & ~n150 ) | ( x97 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n3332 = ( x98 & ~n131 ) | ( x98 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n3333 = n3331 | n3332 ;
  assign n3335 = ( x99 & ~n3334 ) | ( x99 & n3333 ) | ( ~n3334 & n3333 ) ;
  assign n3337 = ( x98 & x99 ) | ( x98 & n3169 ) | ( x99 & n3169 ) ;
  assign n3336 = ( x98 & ~x99 ) | ( x98 & n3169 ) | ( ~x99 & n3169 ) ;
  assign n3338 = ( x99 & ~n3337 ) | ( x99 & n3336 ) | ( ~n3337 & n3336 ) ;
  assign n3339 = ( n139 & ~n3335 ) | ( n139 & n3338 ) | ( ~n3335 & n3338 ) ;
  assign n3340 = ~n139 & n3339 ;
  assign n3341 = ( x2 & n3335 ) | ( x2 & n3340 ) | ( n3335 & n3340 ) ;
  assign n3342 = ( x2 & ~n3340 ) | ( x2 & n3335 ) | ( ~n3340 & n3335 ) ;
  assign n3343 = ( n3340 & ~n3341 ) | ( n3340 & n3342 ) | ( ~n3341 & n3342 ) ;
  assign n3330 = ( n3161 & n3162 ) | ( n3161 & n3175 ) | ( n3162 & n3175 ) ;
  assign n3344 = ( n3329 & ~n3343 ) | ( n3329 & n3330 ) | ( ~n3343 & n3330 ) ;
  assign n3345 = ( n3329 & ~n3330 ) | ( n3329 & n3343 ) | ( ~n3330 & n3343 ) ;
  assign n3346 = ( n3344 & ~n3329 ) | ( n3344 & n3345 ) | ( ~n3329 & n3345 ) ;
  assign n3350 = ~n136 & x100 ;
  assign n3347 = ( x98 & ~n150 ) | ( x98 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n3348 = ( x99 & ~n131 ) | ( x99 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n3349 = n3347 | n3348 ;
  assign n3351 = ( x100 & ~n3350 ) | ( x100 & n3349 ) | ( ~n3350 & n3349 ) ;
  assign n3352 = ( x99 & ~x100 ) | ( x99 & n3337 ) | ( ~x100 & n3337 ) ;
  assign n3353 = ( x99 & x100 ) | ( x99 & n3337 ) | ( x100 & n3337 ) ;
  assign n3354 = ( ~x100 & ~n3352 ) | ( ~x100 & n3353 ) | ( ~n3352 & n3353 ) ;
  assign n3355 = ( n3351 & ~n139 ) | ( n3351 & n3354 ) | ( ~n139 & n3354 ) ;
  assign n3356 = n139 | n3355 ;
  assign n3358 = ( x2 & n3351 ) | ( x2 & n3356 ) | ( n3351 & n3356 ) ;
  assign n3357 = ( x2 & ~n3356 ) | ( x2 & n3351 ) | ( ~n3356 & n3351 ) ;
  assign n3359 = ( n3356 & ~n3358 ) | ( n3356 & n3357 ) | ( ~n3358 & n3357 ) ;
  assign n3518 = ( n3330 & ~n3329 ) | ( n3330 & n3343 ) | ( ~n3329 & n3343 ) ;
  assign n3381 = ( x35 & ~x36 ) | ( x35 & 1'b0 ) | ( ~x36 & 1'b0 ) ;
  assign n3382 = ~x35 & x36 ;
  assign n3383 = n3381 | n3382 ;
  assign n3384 = x64 &  n3383 ;
  assign n3385 = ( n2859 & ~n3092 ) | ( n2859 & n3221 ) | ( ~n3092 & n3221 ) ;
  assign n3386 = ( x35 & n3092 ) | ( x35 & n3385 ) | ( n3092 & n3385 ) ;
  assign n3387 = ( x35 & ~n3386 ) | ( x35 & 1'b0 ) | ( ~n3386 & 1'b0 ) ;
  assign n3391 = x65 &  n3214 ;
  assign n3388 = ( x67 & ~n3087 ) | ( x67 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n3389 = x66 &  n3082 ;
  assign n3390 = n3388 | n3389 ;
  assign n3392 = ( x65 & ~n3391 ) | ( x65 & n3390 ) | ( ~n3391 & n3390 ) ;
  assign n3393 = n173 | n3090 ;
  assign n3394 = ~n3392 & n3393 ;
  assign n3395 = x35 &  n3394 ;
  assign n3396 = x35 | n3394 ;
  assign n3397 = ~n3395 & n3396 ;
  assign n3398 = ( n3384 & ~n3387 ) | ( n3384 & n3397 ) | ( ~n3387 & n3397 ) ;
  assign n3399 = ( n3384 & ~n3397 ) | ( n3384 & n3387 ) | ( ~n3397 & n3387 ) ;
  assign n3400 = ( n3398 & ~n3384 ) | ( n3398 & n3399 ) | ( ~n3384 & n3399 ) ;
  assign n3401 = ( n3097 & n3226 ) | ( n3097 & n3236 ) | ( n3226 & n3236 ) ;
  assign n3405 = x68 &  n2718 ;
  assign n3402 = ( x70 & ~n2642 ) | ( x70 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n3403 = x69 &  n2637 ;
  assign n3404 = n3402 | n3403 ;
  assign n3406 = ( x68 & ~n3405 ) | ( x68 & n3404 ) | ( ~n3405 & n3404 ) ;
  assign n3407 = ( n282 & ~n2645 ) | ( n282 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n3408 = n3406 | n3407 ;
  assign n3409 = ( x32 & ~n3408 ) | ( x32 & 1'b0 ) | ( ~n3408 & 1'b0 ) ;
  assign n3410 = ~x32 & n3408 ;
  assign n3411 = n3409 | n3410 ;
  assign n3412 = ( n3400 & ~n3401 ) | ( n3400 & n3411 ) | ( ~n3401 & n3411 ) ;
  assign n3413 = ( n3401 & ~n3400 ) | ( n3401 & n3411 ) | ( ~n3400 & n3411 ) ;
  assign n3414 = ( n3412 & ~n3411 ) | ( n3412 & n3413 ) | ( ~n3411 & n3413 ) ;
  assign n3419 = x71 &  n2312 ;
  assign n3416 = ( x73 & ~n2195 ) | ( x73 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n3417 = x72 &  n2190 ;
  assign n3418 = n3416 | n3417 ;
  assign n3420 = ( x71 & ~n3419 ) | ( x71 & n3418 ) | ( ~n3419 & n3418 ) ;
  assign n3421 = ( n389 & ~n2198 ) | ( n389 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n3422 = n3420 | n3421 ;
  assign n3423 = ( x29 & ~n3422 ) | ( x29 & 1'b0 ) | ( ~n3422 & 1'b0 ) ;
  assign n3424 = ~x29 & n3422 ;
  assign n3425 = n3423 | n3424 ;
  assign n3415 = ( n3100 & n3239 ) | ( n3100 & n3249 ) | ( n3239 & n3249 ) ;
  assign n3426 = ( n3414 & ~n3425 ) | ( n3414 & n3415 ) | ( ~n3425 & n3415 ) ;
  assign n3427 = ( n3414 & ~n3415 ) | ( n3414 & n3425 ) | ( ~n3415 & n3425 ) ;
  assign n3428 = ( n3426 & ~n3414 ) | ( n3426 & n3427 ) | ( ~n3414 & n3427 ) ;
  assign n3374 = x74 &  n1894 ;
  assign n3371 = ( x76 & ~n1816 ) | ( x76 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n3372 = x75 &  n1811 ;
  assign n3373 = n3371 | n3372 ;
  assign n3375 = ( x74 & ~n3374 ) | ( x74 & n3373 ) | ( ~n3374 & n3373 ) ;
  assign n3376 = ( n603 & ~n1819 ) | ( n603 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n3377 = n3375 | n3376 ;
  assign n3378 = ( x26 & ~n3377 ) | ( x26 & 1'b0 ) | ( ~n3377 & 1'b0 ) ;
  assign n3379 = ~x26 & n3377 ;
  assign n3380 = n3378 | n3379 ;
  assign n3429 = ( n3254 & ~n3428 ) | ( n3254 & n3380 ) | ( ~n3428 & n3380 ) ;
  assign n3430 = ( n3380 & ~n3254 ) | ( n3380 & n3428 ) | ( ~n3254 & n3428 ) ;
  assign n3431 = ( n3429 & ~n3380 ) | ( n3429 & n3430 ) | ( ~n3380 & n3430 ) ;
  assign n3432 = ( n3255 & n3256 ) | ( n3255 & n3266 ) | ( n3256 & n3266 ) ;
  assign n3436 = x77 &  n1551 ;
  assign n3433 = ( x79 & ~n1451 ) | ( x79 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n3434 = x78 &  n1446 ;
  assign n3435 = n3433 | n3434 ;
  assign n3437 = ( x77 & ~n3436 ) | ( x77 & n3435 ) | ( ~n3436 & n3435 ) ;
  assign n3438 = ( n766 & ~n1454 ) | ( n766 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n3439 = n3437 | n3438 ;
  assign n3440 = ( x23 & ~n3439 ) | ( x23 & 1'b0 ) | ( ~n3439 & 1'b0 ) ;
  assign n3441 = ~x23 & n3439 ;
  assign n3442 = n3440 | n3441 ;
  assign n3443 = ( n3431 & ~n3432 ) | ( n3431 & n3442 ) | ( ~n3432 & n3442 ) ;
  assign n3444 = ( n3432 & ~n3431 ) | ( n3432 & n3442 ) | ( ~n3431 & n3442 ) ;
  assign n3445 = ( n3443 & ~n3442 ) | ( n3443 & n3444 ) | ( ~n3442 & n3444 ) ;
  assign n3450 = x80 &  n1227 ;
  assign n3447 = ( x82 & ~n1154 ) | ( x82 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n3448 = x81 &  n1149 ;
  assign n3449 = n3447 | n3448 ;
  assign n3451 = ( x80 & ~n3450 ) | ( x80 & n3449 ) | ( ~n3450 & n3449 ) ;
  assign n3452 = ( n1084 & ~n1157 ) | ( n1084 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n3453 = n3451 | n3452 ;
  assign n3454 = ( x20 & ~n3453 ) | ( x20 & 1'b0 ) | ( ~n3453 & 1'b0 ) ;
  assign n3455 = ~x20 & n3453 ;
  assign n3456 = n3454 | n3455 ;
  assign n3446 = ( n3269 & n3279 ) | ( n3269 & n3280 ) | ( n3279 & n3280 ) ;
  assign n3457 = ( n3445 & ~n3456 ) | ( n3445 & n3446 ) | ( ~n3456 & n3446 ) ;
  assign n3458 = ( n3445 & ~n3446 ) | ( n3445 & n3456 ) | ( ~n3446 & n3456 ) ;
  assign n3459 = ( n3457 & ~n3445 ) | ( n3457 & n3458 ) | ( ~n3445 & n3458 ) ;
  assign n3460 = ( n3134 & n3283 ) | ( n3134 & n3293 ) | ( n3283 & n3293 ) ;
  assign n3464 = x83 &  n942 ;
  assign n3461 = ( x85 & ~n896 ) | ( x85 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n3462 = x84 &  n891 ;
  assign n3463 = n3461 | n3462 ;
  assign n3465 = ( x83 & ~n3464 ) | ( x83 & n3463 ) | ( ~n3464 & n3463 ) ;
  assign n3466 = ~n899 & n1295 ;
  assign n3467 = n3465 | n3466 ;
  assign n3468 = ( x17 & ~n3467 ) | ( x17 & 1'b0 ) | ( ~n3467 & 1'b0 ) ;
  assign n3469 = ~x17 & n3467 ;
  assign n3470 = n3468 | n3469 ;
  assign n3471 = ( n3459 & ~n3460 ) | ( n3459 & n3470 ) | ( ~n3460 & n3470 ) ;
  assign n3472 = ( n3459 & ~n3470 ) | ( n3459 & n3460 ) | ( ~n3470 & n3460 ) ;
  assign n3473 = ( n3471 & ~n3459 ) | ( n3471 & n3472 ) | ( ~n3459 & n3472 ) ;
  assign n3478 = x86 &  n713 ;
  assign n3475 = ( x88 & ~n641 ) | ( x88 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n3476 = x87 &  n636 ;
  assign n3477 = n3475 | n3476 ;
  assign n3479 = ( x86 & ~n3478 ) | ( x86 & n3477 ) | ( ~n3478 & n3477 ) ;
  assign n3480 = ~n644 & n1624 ;
  assign n3481 = n3479 | n3480 ;
  assign n3482 = ( x14 & ~n3481 ) | ( x14 & 1'b0 ) | ( ~n3481 & 1'b0 ) ;
  assign n3483 = ~x14 & n3481 ;
  assign n3484 = n3482 | n3483 ;
  assign n3474 = ( n3138 & n3296 ) | ( n3138 & n3306 ) | ( n3296 & n3306 ) ;
  assign n3485 = ( n3473 & ~n3484 ) | ( n3473 & n3474 ) | ( ~n3484 & n3474 ) ;
  assign n3486 = ( n3473 & ~n3474 ) | ( n3473 & n3484 ) | ( ~n3474 & n3484 ) ;
  assign n3487 = ( n3485 & ~n3473 ) | ( n3485 & n3486 ) | ( ~n3473 & n3486 ) ;
  assign n3491 = x89 &  n503 ;
  assign n3488 = ( x91 & ~n450 ) | ( x91 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n3489 = x90 &  n445 ;
  assign n3490 = n3488 | n3489 ;
  assign n3492 = ( x89 & ~n3491 ) | ( x89 & n3490 ) | ( ~n3491 & n3490 ) ;
  assign n3493 = ~n453 & n2108 ;
  assign n3494 = n3492 | n3493 ;
  assign n3495 = ( x11 & ~n3494 ) | ( x11 & 1'b0 ) | ( ~n3494 & 1'b0 ) ;
  assign n3496 = ~x11 & n3494 ;
  assign n3497 = n3495 | n3496 ;
  assign n3498 = ( n3487 & ~n3311 ) | ( n3487 & n3497 ) | ( ~n3311 & n3497 ) ;
  assign n3499 = ( n3311 & ~n3487 ) | ( n3311 & n3497 ) | ( ~n3487 & n3497 ) ;
  assign n3500 = ( n3498 & ~n3497 ) | ( n3498 & n3499 ) | ( ~n3497 & n3499 ) ;
  assign n3505 = x92 &  n353 ;
  assign n3502 = ( x94 & ~n313 ) | ( x94 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n3503 = x93 &  n308 ;
  assign n3504 = n3502 | n3503 ;
  assign n3506 = ( x92 & ~n3505 ) | ( x92 & n3504 ) | ( ~n3505 & n3504 ) ;
  assign n3507 = ~n316 & n2401 ;
  assign n3508 = n3506 | n3507 ;
  assign n3509 = ( x8 & ~n3508 ) | ( x8 & 1'b0 ) | ( ~n3508 & 1'b0 ) ;
  assign n3510 = ~x8 & n3508 ;
  assign n3511 = n3509 | n3510 ;
  assign n3501 = ( n3312 & ~n3322 ) | ( n3312 & n3323 ) | ( ~n3322 & n3323 ) ;
  assign n3512 = ( n3500 & ~n3511 ) | ( n3500 & n3501 ) | ( ~n3511 & n3501 ) ;
  assign n3513 = ( n3500 & ~n3501 ) | ( n3500 & n3511 ) | ( ~n3501 & n3511 ) ;
  assign n3514 = ( n3512 & ~n3500 ) | ( n3512 & n3513 ) | ( ~n3500 & n3513 ) ;
  assign n3363 = x95 &  n225 ;
  assign n3360 = ( x97 & ~n197 ) | ( x97 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n3361 = x96 &  n192 ;
  assign n3362 = n3360 | n3361 ;
  assign n3364 = ( x95 & ~n3363 ) | ( x95 & n3362 ) | ( ~n3363 & n3362 ) ;
  assign n3365 = ~n200 & n2999 ;
  assign n3366 = n3364 | n3365 ;
  assign n3367 = ( x5 & ~n3366 ) | ( x5 & 1'b0 ) | ( ~n3366 & 1'b0 ) ;
  assign n3368 = ~x5 & n3366 ;
  assign n3369 = n3367 | n3368 ;
  assign n3370 = ( n3179 & ~n3326 ) | ( n3179 & n3189 ) | ( ~n3326 & n3189 ) ;
  assign n3516 = ( n3369 & n3370 ) | ( n3369 & n3514 ) | ( n3370 & n3514 ) ;
  assign n3515 = ( n3369 & ~n3514 ) | ( n3369 & n3370 ) | ( ~n3514 & n3370 ) ;
  assign n3517 = ( n3514 & ~n3516 ) | ( n3514 & n3515 ) | ( ~n3516 & n3515 ) ;
  assign n3519 = ( n3359 & ~n3518 ) | ( n3359 & n3517 ) | ( ~n3518 & n3517 ) ;
  assign n3520 = ( n3359 & ~n3517 ) | ( n3359 & n3518 ) | ( ~n3517 & n3518 ) ;
  assign n3521 = ( n3519 & ~n3359 ) | ( n3519 & n3520 ) | ( ~n3359 & n3520 ) ;
  assign n3525 = x93 &  n353 ;
  assign n3522 = ( x95 & ~n313 ) | ( x95 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n3523 = x94 &  n308 ;
  assign n3524 = n3522 | n3523 ;
  assign n3526 = ( x93 & ~n3525 ) | ( x93 & n3524 ) | ( ~n3525 & n3524 ) ;
  assign n3527 = ~n316 & n2547 ;
  assign n3528 = n3526 | n3527 ;
  assign n3529 = ( x8 & ~n3528 ) | ( x8 & 1'b0 ) | ( ~n3528 & 1'b0 ) ;
  assign n3530 = ~x8 & n3528 ;
  assign n3531 = n3529 | n3530 ;
  assign n3532 = ( n3501 & ~n3500 ) | ( n3501 & n3511 ) | ( ~n3500 & n3511 ) ;
  assign n3536 = x84 &  n942 ;
  assign n3533 = ( x86 & ~n896 ) | ( x86 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n3534 = x85 &  n891 ;
  assign n3535 = n3533 | n3534 ;
  assign n3537 = ( x84 & ~n3536 ) | ( x84 & n3535 ) | ( ~n3536 & n3535 ) ;
  assign n3538 = ~n899 & n1496 ;
  assign n3539 = n3537 | n3538 ;
  assign n3540 = ( x17 & ~n3539 ) | ( x17 & 1'b0 ) | ( ~n3539 & 1'b0 ) ;
  assign n3541 = ~x17 & n3539 ;
  assign n3542 = n3540 | n3541 ;
  assign n3546 = x81 &  n1227 ;
  assign n3543 = ( x83 & ~n1154 ) | ( x83 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n3544 = x82 &  n1149 ;
  assign n3545 = n3543 | n3544 ;
  assign n3547 = ( x81 & ~n3546 ) | ( x81 & n3545 ) | ( ~n3546 & n3545 ) ;
  assign n3548 = ( n1100 & ~n1157 ) | ( n1100 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n3549 = n3547 | n3548 ;
  assign n3550 = ( x20 & ~n3549 ) | ( x20 & 1'b0 ) | ( ~n3549 & 1'b0 ) ;
  assign n3551 = ~x20 & n3549 ;
  assign n3552 = n3550 | n3551 ;
  assign n3556 = x75 &  n1894 ;
  assign n3553 = ( x77 & ~n1816 ) | ( x77 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n3554 = x76 &  n1811 ;
  assign n3555 = n3553 | n3554 ;
  assign n3557 = ( x75 & ~n3556 ) | ( x75 & n3555 ) | ( ~n3556 & n3555 ) ;
  assign n3558 = ( n677 & ~n1819 ) | ( n677 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n3559 = n3557 | n3558 ;
  assign n3560 = ( x26 & ~n3559 ) | ( x26 & 1'b0 ) | ( ~n3559 & 1'b0 ) ;
  assign n3561 = ~x26 & n3559 ;
  assign n3562 = n3560 | n3561 ;
  assign n3566 = x72 &  n2312 ;
  assign n3563 = ( x74 & ~n2195 ) | ( x74 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n3564 = x73 &  n2190 ;
  assign n3565 = n3563 | n3564 ;
  assign n3567 = ( x72 & ~n3566 ) | ( x72 & n3565 ) | ( ~n3566 & n3565 ) ;
  assign n3568 = ( n482 & ~n2198 ) | ( n482 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n3569 = n3567 | n3568 ;
  assign n3570 = ( x29 & ~n3569 ) | ( x29 & 1'b0 ) | ( ~n3569 & 1'b0 ) ;
  assign n3571 = ~x29 & n3569 ;
  assign n3572 = n3570 | n3571 ;
  assign n3573 = ( n3415 & ~n3414 ) | ( n3415 & n3425 ) | ( ~n3414 & n3425 ) ;
  assign n3577 = x69 &  n2718 ;
  assign n3574 = ( x71 & ~n2642 ) | ( x71 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n3575 = x70 &  n2637 ;
  assign n3576 = n3574 | n3575 ;
  assign n3578 = ( x69 & ~n3577 ) | ( x69 & n3576 ) | ( ~n3577 & n3576 ) ;
  assign n3579 = ( n298 & ~n2645 ) | ( n298 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n3580 = n3578 | n3579 ;
  assign n3581 = ( x32 & ~n3580 ) | ( x32 & 1'b0 ) | ( ~n3580 & 1'b0 ) ;
  assign n3582 = ~x32 & n3580 ;
  assign n3583 = n3581 | n3582 ;
  assign n3587 = x66 &  n3214 ;
  assign n3584 = ( x68 & ~n3087 ) | ( x68 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n3585 = x67 &  n3082 ;
  assign n3586 = n3584 | n3585 ;
  assign n3588 = ( x66 & ~n3587 ) | ( x66 & n3586 ) | ( ~n3587 & n3586 ) ;
  assign n3589 = ( n213 & ~n3090 ) | ( n213 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n3590 = n3588 | n3589 ;
  assign n3591 = ( x35 & ~n3590 ) | ( x35 & 1'b0 ) | ( ~n3590 & 1'b0 ) ;
  assign n3592 = ~x35 & n3590 ;
  assign n3593 = n3591 | n3592 ;
  assign n3594 = ( x38 & ~n3384 ) | ( x38 & 1'b0 ) | ( ~n3384 & 1'b0 ) ;
  assign n3595 = ( x36 & x37 ) | ( x36 & n3381 ) | ( x37 & n3381 ) ;
  assign n3596 = ( x36 & ~n3382 ) | ( x36 & x37 ) | ( ~n3382 & x37 ) ;
  assign n3597 = ~n3595 &  n3596 ;
  assign n3598 = x64 &  n3597 ;
  assign n3599 = ~x37 & x38 ;
  assign n3600 = ( x37 & ~x38 ) | ( x37 & 1'b0 ) | ( ~x38 & 1'b0 ) ;
  assign n3601 = n3599 | n3600 ;
  assign n3602 = ~n3383 |  n3601 ;
  assign n3603 = ( x65 & ~n3602 ) | ( x65 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n3604 = n3598 | n3603 ;
  assign n3605 = ~n3383 | ~n3601 ;
  assign n3606 = ( n142 & ~n3605 ) | ( n142 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n3607 = n3604 | n3606 ;
  assign n3609 = ( x38 & n3594 ) | ( x38 & n3607 ) | ( n3594 & n3607 ) ;
  assign n3608 = ( x38 & ~n3594 ) | ( x38 & n3607 ) | ( ~n3594 & n3607 ) ;
  assign n3610 = ( n3594 & ~n3609 ) | ( n3594 & n3608 ) | ( ~n3609 & n3608 ) ;
  assign n3612 = ( n3399 & n3593 ) | ( n3399 & n3610 ) | ( n3593 & n3610 ) ;
  assign n3611 = ( n3399 & ~n3593 ) | ( n3399 & n3610 ) | ( ~n3593 & n3610 ) ;
  assign n3613 = ( n3593 & ~n3612 ) | ( n3593 & n3611 ) | ( ~n3612 & n3611 ) ;
  assign n3615 = ( n3413 & n3583 ) | ( n3413 & n3613 ) | ( n3583 & n3613 ) ;
  assign n3614 = ( n3413 & ~n3583 ) | ( n3413 & n3613 ) | ( ~n3583 & n3613 ) ;
  assign n3616 = ( n3583 & ~n3615 ) | ( n3583 & n3614 ) | ( ~n3615 & n3614 ) ;
  assign n3618 = ( n3572 & n3573 ) | ( n3572 & n3616 ) | ( n3573 & n3616 ) ;
  assign n3617 = ( n3573 & ~n3572 ) | ( n3573 & n3616 ) | ( ~n3572 & n3616 ) ;
  assign n3619 = ( n3572 & ~n3618 ) | ( n3572 & n3617 ) | ( ~n3618 & n3617 ) ;
  assign n3621 = ( n3429 & n3562 ) | ( n3429 & n3619 ) | ( n3562 & n3619 ) ;
  assign n3620 = ( n3429 & ~n3562 ) | ( n3429 & n3619 ) | ( ~n3562 & n3619 ) ;
  assign n3622 = ( n3562 & ~n3621 ) | ( n3562 & n3620 ) | ( ~n3621 & n3620 ) ;
  assign n3626 = x78 &  n1551 ;
  assign n3623 = ( x80 & ~n1451 ) | ( x80 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n3624 = x79 &  n1446 ;
  assign n3625 = n3623 | n3624 ;
  assign n3627 = ( x78 & ~n3626 ) | ( x78 & n3625 ) | ( ~n3626 & n3625 ) ;
  assign n3628 = ( n842 & ~n1454 ) | ( n842 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n3629 = n3627 | n3628 ;
  assign n3630 = ( x23 & ~n3629 ) | ( x23 & 1'b0 ) | ( ~n3629 & 1'b0 ) ;
  assign n3631 = ~x23 & n3629 ;
  assign n3632 = n3630 | n3631 ;
  assign n3633 = ( n3622 & ~n3444 ) | ( n3622 & n3632 ) | ( ~n3444 & n3632 ) ;
  assign n3634 = ( n3444 & ~n3632 ) | ( n3444 & n3622 ) | ( ~n3632 & n3622 ) ;
  assign n3635 = ( n3633 & ~n3622 ) | ( n3633 & n3634 ) | ( ~n3622 & n3634 ) ;
  assign n3636 = ( n3446 & ~n3445 ) | ( n3446 & n3456 ) | ( ~n3445 & n3456 ) ;
  assign n3637 = ( n3552 & n3635 ) | ( n3552 & n3636 ) | ( n3635 & n3636 ) ;
  assign n3638 = ( n3635 & ~n3552 ) | ( n3635 & n3636 ) | ( ~n3552 & n3636 ) ;
  assign n3639 = ( n3552 & ~n3637 ) | ( n3552 & n3638 ) | ( ~n3637 & n3638 ) ;
  assign n3640 = ( n3460 & ~n3459 ) | ( n3460 & n3470 ) | ( ~n3459 & n3470 ) ;
  assign n3641 = ( n3542 & n3639 ) | ( n3542 & n3640 ) | ( n3639 & n3640 ) ;
  assign n3642 = ( n3639 & ~n3542 ) | ( n3639 & n3640 ) | ( ~n3542 & n3640 ) ;
  assign n3643 = ( n3542 & ~n3641 ) | ( n3542 & n3642 ) | ( ~n3641 & n3642 ) ;
  assign n3648 = x87 &  n713 ;
  assign n3645 = ( x89 & ~n641 ) | ( x89 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n3646 = x88 &  n636 ;
  assign n3647 = n3645 | n3646 ;
  assign n3649 = ( x87 & ~n3648 ) | ( x87 & n3647 ) | ( ~n3648 & n3647 ) ;
  assign n3650 = ~n644 & n1741 ;
  assign n3651 = n3649 | n3650 ;
  assign n3652 = ( x14 & ~n3651 ) | ( x14 & 1'b0 ) | ( ~n3651 & 1'b0 ) ;
  assign n3653 = ~x14 & n3651 ;
  assign n3654 = n3652 | n3653 ;
  assign n3644 = ( n3474 & ~n3473 ) | ( n3474 & n3484 ) | ( ~n3473 & n3484 ) ;
  assign n3655 = ( n3643 & ~n3654 ) | ( n3643 & n3644 ) | ( ~n3654 & n3644 ) ;
  assign n3656 = ( n3643 & ~n3644 ) | ( n3643 & n3654 ) | ( ~n3644 & n3654 ) ;
  assign n3657 = ( n3655 & ~n3643 ) | ( n3655 & n3656 ) | ( ~n3643 & n3656 ) ;
  assign n3661 = x90 &  n503 ;
  assign n3658 = ( x92 & ~n450 ) | ( x92 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n3659 = x91 &  n445 ;
  assign n3660 = n3658 | n3659 ;
  assign n3662 = ( x90 & ~n3661 ) | ( x90 & n3660 ) | ( ~n3661 & n3660 ) ;
  assign n3663 = ~n453 & n2248 ;
  assign n3664 = n3662 | n3663 ;
  assign n3665 = ( x11 & ~n3664 ) | ( x11 & 1'b0 ) | ( ~n3664 & 1'b0 ) ;
  assign n3666 = ~x11 & n3664 ;
  assign n3667 = n3665 | n3666 ;
  assign n3668 = ( n3657 & ~n3499 ) | ( n3657 & n3667 ) | ( ~n3499 & n3667 ) ;
  assign n3669 = ( n3499 & ~n3667 ) | ( n3499 & n3657 ) | ( ~n3667 & n3657 ) ;
  assign n3670 = ( n3668 & ~n3657 ) | ( n3668 & n3669 ) | ( ~n3657 & n3669 ) ;
  assign n3672 = ( n3531 & n3532 ) | ( n3531 & n3670 ) | ( n3532 & n3670 ) ;
  assign n3671 = ( n3532 & ~n3531 ) | ( n3532 & n3670 ) | ( ~n3531 & n3670 ) ;
  assign n3673 = ( n3531 & ~n3672 ) | ( n3531 & n3671 ) | ( ~n3672 & n3671 ) ;
  assign n3677 = x96 &  n225 ;
  assign n3674 = ( x98 & ~n197 ) | ( x98 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n3675 = x97 &  n192 ;
  assign n3676 = n3674 | n3675 ;
  assign n3678 = ( x96 & ~n3677 ) | ( x96 & n3676 ) | ( ~n3677 & n3676 ) ;
  assign n3679 = ~n200 & n3170 ;
  assign n3680 = n3678 | n3679 ;
  assign n3681 = ( x5 & ~n3680 ) | ( x5 & 1'b0 ) | ( ~n3680 & 1'b0 ) ;
  assign n3682 = ~x5 & n3680 ;
  assign n3683 = n3681 | n3682 ;
  assign n3684 = ( n3515 & n3673 ) | ( n3515 & n3683 ) | ( n3673 & n3683 ) ;
  assign n3685 = ( n3515 & ~n3673 ) | ( n3515 & n3683 ) | ( ~n3673 & n3683 ) ;
  assign n3686 = ( n3673 & ~n3684 ) | ( n3673 & n3685 ) | ( ~n3684 & n3685 ) ;
  assign n3690 = ~n136 & x101 ;
  assign n3687 = ( x99 & ~n150 ) | ( x99 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n3688 = ( x100 & ~n131 ) | ( x100 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n3689 = n3687 | n3688 ;
  assign n3691 = ( x101 & ~n3690 ) | ( x101 & n3689 ) | ( ~n3690 & n3689 ) ;
  assign n3692 = ( x100 & ~x101 ) | ( x100 & n3353 ) | ( ~x101 & n3353 ) ;
  assign n3693 = ( x100 & x101 ) | ( x100 & n3353 ) | ( x101 & n3353 ) ;
  assign n3694 = ( ~x101 & ~n3692 ) | ( ~x101 & n3693 ) | ( ~n3692 & n3693 ) ;
  assign n3695 = ( n3691 & ~n139 ) | ( n3691 & n3694 ) | ( ~n139 & n3694 ) ;
  assign n3696 = n139 | n3695 ;
  assign n3698 = ( x2 & n3691 ) | ( x2 & n3696 ) | ( n3691 & n3696 ) ;
  assign n3697 = ( x2 & ~n3696 ) | ( x2 & n3691 ) | ( ~n3696 & n3691 ) ;
  assign n3699 = ( n3696 & ~n3698 ) | ( n3696 & n3697 ) | ( ~n3698 & n3697 ) ;
  assign n3700 = ( n3686 & ~n3519 ) | ( n3686 & n3699 ) | ( ~n3519 & n3699 ) ;
  assign n3701 = ( n3519 & ~n3699 ) | ( n3519 & n3686 ) | ( ~n3699 & n3686 ) ;
  assign n3702 = ( n3700 & ~n3686 ) | ( n3700 & n3701 ) | ( ~n3686 & n3701 ) ;
  assign n3716 = x94 &  n353 ;
  assign n3713 = ( x96 & ~n313 ) | ( x96 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n3714 = x95 &  n308 ;
  assign n3715 = n3713 | n3714 ;
  assign n3717 = ( x94 & ~n3716 ) | ( x94 & n3715 ) | ( ~n3716 & n3715 ) ;
  assign n3718 = ~n316 & n2836 ;
  assign n3719 = n3717 | n3718 ;
  assign n3720 = ( x8 & ~n3719 ) | ( x8 & 1'b0 ) | ( ~n3719 & 1'b0 ) ;
  assign n3721 = ~x8 & n3719 ;
  assign n3722 = n3720 | n3721 ;
  assign n3726 = x91 &  n503 ;
  assign n3723 = ( x93 & ~n450 ) | ( x93 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n3724 = x92 &  n445 ;
  assign n3725 = n3723 | n3724 ;
  assign n3727 = ( x91 & ~n3726 ) | ( x91 & n3725 ) | ( ~n3726 & n3725 ) ;
  assign n3728 = n453 | n2264 ;
  assign n3729 = ~n3727 & n3728 ;
  assign n3730 = x11 &  n3729 ;
  assign n3731 = x11 | n3729 ;
  assign n3732 = ~n3730 & n3731 ;
  assign n3733 = ( n3499 & n3657 ) | ( n3499 & n3667 ) | ( n3657 & n3667 ) ;
  assign n3831 = x85 &  n942 ;
  assign n3828 = ( x87 & ~n896 ) | ( x87 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n3829 = x86 &  n891 ;
  assign n3830 = n3828 | n3829 ;
  assign n3832 = ( x85 & ~n3831 ) | ( x85 & n3830 ) | ( ~n3831 & n3830 ) ;
  assign n3833 = ~n899 & n1512 ;
  assign n3834 = n3832 | n3833 ;
  assign n3835 = ( x17 & ~n3834 ) | ( x17 & 1'b0 ) | ( ~n3834 & 1'b0 ) ;
  assign n3836 = ~x17 & n3834 ;
  assign n3837 = n3835 | n3836 ;
  assign n3737 = x82 &  n1227 ;
  assign n3734 = ( x84 & ~n1154 ) | ( x84 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n3735 = x83 &  n1149 ;
  assign n3736 = n3734 | n3735 ;
  assign n3738 = ( x82 & ~n3737 ) | ( x82 & n3736 ) | ( ~n3737 & n3736 ) ;
  assign n3739 = ~n1157 & n1199 ;
  assign n3740 = n3738 | n3739 ;
  assign n3741 = ( x20 & ~n3740 ) | ( x20 & 1'b0 ) | ( ~n3740 & 1'b0 ) ;
  assign n3742 = ~x20 & n3740 ;
  assign n3743 = n3741 | n3742 ;
  assign n3747 = x73 &  n2312 ;
  assign n3744 = ( x75 & ~n2195 ) | ( x75 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n3745 = x74 &  n2190 ;
  assign n3746 = n3744 | n3745 ;
  assign n3748 = ( x73 & ~n3747 ) | ( x73 & n3746 ) | ( ~n3747 & n3746 ) ;
  assign n3749 = ( n540 & ~n2198 ) | ( n540 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n3750 = n3748 | n3749 ;
  assign n3751 = ( x29 & ~n3750 ) | ( x29 & 1'b0 ) | ( ~n3750 & 1'b0 ) ;
  assign n3752 = ~x29 & n3750 ;
  assign n3753 = n3751 | n3752 ;
  assign n3772 = x67 &  n3214 ;
  assign n3769 = ( x69 & ~n3087 ) | ( x69 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n3770 = x68 &  n3082 ;
  assign n3771 = n3769 | n3770 ;
  assign n3773 = ( x67 & ~n3772 ) | ( x67 & n3771 ) | ( ~n3772 & n3771 ) ;
  assign n3774 = ( n246 & ~n3090 ) | ( n246 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n3775 = n3773 | n3774 ;
  assign n3776 = ( x35 & ~n3775 ) | ( x35 & 1'b0 ) | ( ~n3775 & 1'b0 ) ;
  assign n3777 = ~x35 & n3775 ;
  assign n3778 = n3776 | n3777 ;
  assign n3755 = ( x36 & ~x37 ) | ( x36 & n3601 ) | ( ~x37 & n3601 ) ;
  assign n3754 = ( x36 & ~x37 ) | ( x36 & n3383 ) | ( ~x37 & n3383 ) ;
  assign n3756 = ~n3755 |  n3754 ;
  assign n3760 = x64 &  n3756 ;
  assign n3757 = ( x66 & ~n3602 ) | ( x66 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n3758 = x65 &  n3597 ;
  assign n3759 = n3757 | n3758 ;
  assign n3761 = ( x64 & ~n3760 ) | ( x64 & n3759 ) | ( ~n3760 & n3759 ) ;
  assign n3762 = ( n157 & ~n3605 ) | ( n157 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n3763 = n3761 | n3762 ;
  assign n3764 = ( x38 & n3384 ) | ( x38 & n3607 ) | ( n3384 & n3607 ) ;
  assign n3765 = ( x38 & ~n3764 ) | ( x38 & 1'b0 ) | ( ~n3764 & 1'b0 ) ;
  assign n3767 = ( x38 & n3763 ) | ( x38 & n3765 ) | ( n3763 & n3765 ) ;
  assign n3766 = ( n3763 & ~x38 ) | ( n3763 & n3765 ) | ( ~x38 & n3765 ) ;
  assign n3768 = ( x38 & ~n3767 ) | ( x38 & n3766 ) | ( ~n3767 & n3766 ) ;
  assign n3779 = ( n3612 & ~n3778 ) | ( n3612 & n3768 ) | ( ~n3778 & n3768 ) ;
  assign n3780 = ( n3768 & ~n3612 ) | ( n3768 & n3778 ) | ( ~n3612 & n3778 ) ;
  assign n3781 = ( n3779 & ~n3768 ) | ( n3779 & n3780 ) | ( ~n3768 & n3780 ) ;
  assign n3785 = x70 &  n2718 ;
  assign n3782 = ( x72 & ~n2642 ) | ( x72 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n3783 = x71 &  n2637 ;
  assign n3784 = n3782 | n3783 ;
  assign n3786 = ( x70 & ~n3785 ) | ( x70 & n3784 ) | ( ~n3785 & n3784 ) ;
  assign n3787 = ( n345 & ~n2645 ) | ( n345 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n3788 = n3786 | n3787 ;
  assign n3789 = ( x32 & ~n3788 ) | ( x32 & 1'b0 ) | ( ~n3788 & 1'b0 ) ;
  assign n3790 = ~x32 & n3788 ;
  assign n3791 = n3789 | n3790 ;
  assign n3792 = ( n3781 & ~n3615 ) | ( n3781 & n3791 ) | ( ~n3615 & n3791 ) ;
  assign n3793 = ( n3615 & ~n3791 ) | ( n3615 & n3781 ) | ( ~n3791 & n3781 ) ;
  assign n3794 = ( n3792 & ~n3781 ) | ( n3792 & n3793 ) | ( ~n3781 & n3793 ) ;
  assign n3796 = ( n3618 & n3753 ) | ( n3618 & n3794 ) | ( n3753 & n3794 ) ;
  assign n3795 = ( n3618 & ~n3753 ) | ( n3618 & n3794 ) | ( ~n3753 & n3794 ) ;
  assign n3797 = ( n3753 & ~n3796 ) | ( n3753 & n3795 ) | ( ~n3796 & n3795 ) ;
  assign n3801 = x76 &  n1894 ;
  assign n3798 = ( x78 & ~n1816 ) | ( x78 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n3799 = x77 &  n1811 ;
  assign n3800 = n3798 | n3799 ;
  assign n3802 = ( x76 & ~n3801 ) | ( x76 & n3800 ) | ( ~n3801 & n3800 ) ;
  assign n3803 = ( n693 & ~n1819 ) | ( n693 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n3804 = n3802 | n3803 ;
  assign n3805 = ( x26 & ~n3804 ) | ( x26 & 1'b0 ) | ( ~n3804 & 1'b0 ) ;
  assign n3806 = ~x26 & n3804 ;
  assign n3807 = n3805 | n3806 ;
  assign n3808 = ( n3797 & ~n3621 ) | ( n3797 & n3807 ) | ( ~n3621 & n3807 ) ;
  assign n3809 = ( n3621 & ~n3807 ) | ( n3621 & n3797 ) | ( ~n3807 & n3797 ) ;
  assign n3810 = ( n3808 & ~n3797 ) | ( n3808 & n3809 ) | ( ~n3797 & n3809 ) ;
  assign n3821 = ( n3444 & n3622 ) | ( n3444 & n3632 ) | ( n3622 & n3632 ) ;
  assign n3814 = x79 &  n1551 ;
  assign n3811 = ( x81 & ~n1451 ) | ( x81 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n3812 = x80 &  n1446 ;
  assign n3813 = n3811 | n3812 ;
  assign n3815 = ( x79 & ~n3814 ) | ( x79 & n3813 ) | ( ~n3814 & n3813 ) ;
  assign n3816 = ( n994 & ~n1454 ) | ( n994 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n3817 = n3815 | n3816 ;
  assign n3818 = ( x23 & ~n3817 ) | ( x23 & 1'b0 ) | ( ~n3817 & 1'b0 ) ;
  assign n3819 = ~x23 & n3817 ;
  assign n3820 = n3818 | n3819 ;
  assign n3822 = ( n3810 & ~n3821 ) | ( n3810 & n3820 ) | ( ~n3821 & n3820 ) ;
  assign n3823 = ( n3810 & ~n3820 ) | ( n3810 & n3821 ) | ( ~n3820 & n3821 ) ;
  assign n3824 = ( n3822 & ~n3810 ) | ( n3822 & n3823 ) | ( ~n3810 & n3823 ) ;
  assign n3825 = ( n3637 & n3743 ) | ( n3637 & n3824 ) | ( n3743 & n3824 ) ;
  assign n3826 = ( n3637 & ~n3743 ) | ( n3637 & n3824 ) | ( ~n3743 & n3824 ) ;
  assign n3827 = ( n3743 & ~n3825 ) | ( n3743 & n3826 ) | ( ~n3825 & n3826 ) ;
  assign n3838 = ( n3641 & ~n3837 ) | ( n3641 & n3827 ) | ( ~n3837 & n3827 ) ;
  assign n3839 = ( n3827 & ~n3641 ) | ( n3827 & n3837 ) | ( ~n3641 & n3837 ) ;
  assign n3840 = ( n3838 & ~n3827 ) | ( n3838 & n3839 ) | ( ~n3827 & n3839 ) ;
  assign n3841 = ( n3643 & n3644 ) | ( n3643 & n3654 ) | ( n3644 & n3654 ) ;
  assign n3845 = x88 &  n713 ;
  assign n3842 = ( x90 & ~n641 ) | ( x90 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n3843 = x89 &  n636 ;
  assign n3844 = n3842 | n3843 ;
  assign n3846 = ( x88 & ~n3845 ) | ( x88 & n3844 ) | ( ~n3845 & n3844 ) ;
  assign n3847 = ~n644 & n1976 ;
  assign n3848 = n3846 | n3847 ;
  assign n3849 = ( x14 & ~n3848 ) | ( x14 & 1'b0 ) | ( ~n3848 & 1'b0 ) ;
  assign n3850 = ~x14 & n3848 ;
  assign n3851 = n3849 | n3850 ;
  assign n3852 = ( n3840 & ~n3841 ) | ( n3840 & n3851 ) | ( ~n3841 & n3851 ) ;
  assign n3853 = ( n3840 & ~n3851 ) | ( n3840 & n3841 ) | ( ~n3851 & n3841 ) ;
  assign n3854 = ( n3852 & ~n3840 ) | ( n3852 & n3853 ) | ( ~n3840 & n3853 ) ;
  assign n3855 = ( n3732 & n3733 ) | ( n3732 & n3854 ) | ( n3733 & n3854 ) ;
  assign n3856 = ( n3733 & ~n3732 ) | ( n3733 & n3854 ) | ( ~n3732 & n3854 ) ;
  assign n3857 = ( n3732 & ~n3855 ) | ( n3732 & n3856 ) | ( ~n3855 & n3856 ) ;
  assign n3858 = ( n3722 & ~n3672 ) | ( n3722 & n3857 ) | ( ~n3672 & n3857 ) ;
  assign n3859 = ( n3672 & ~n3857 ) | ( n3672 & n3722 ) | ( ~n3857 & n3722 ) ;
  assign n3860 = ( n3858 & ~n3722 ) | ( n3858 & n3859 ) | ( ~n3722 & n3859 ) ;
  assign n3706 = x97 &  n225 ;
  assign n3703 = ( x99 & ~n197 ) | ( x99 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n3704 = x98 &  n192 ;
  assign n3705 = n3703 | n3704 ;
  assign n3707 = ( x97 & ~n3706 ) | ( x97 & n3705 ) | ( ~n3706 & n3705 ) ;
  assign n3708 = ~n200 & n3338 ;
  assign n3709 = n3707 | n3708 ;
  assign n3710 = ( x5 & ~n3709 ) | ( x5 & 1'b0 ) | ( ~n3709 & 1'b0 ) ;
  assign n3711 = ~x5 & n3709 ;
  assign n3712 = n3710 | n3711 ;
  assign n3862 = ( n3684 & n3712 ) | ( n3684 & n3860 ) | ( n3712 & n3860 ) ;
  assign n3861 = ( n3684 & ~n3860 ) | ( n3684 & n3712 ) | ( ~n3860 & n3712 ) ;
  assign n3863 = ( n3860 & ~n3862 ) | ( n3860 & n3861 ) | ( ~n3862 & n3861 ) ;
  assign n3864 = ( n3519 & ~n3686 ) | ( n3519 & n3699 ) | ( ~n3686 & n3699 ) ;
  assign n3868 = ~n136 & x102 ;
  assign n3865 = ( x100 & ~n150 ) | ( x100 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n3866 = ( x101 & ~n131 ) | ( x101 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n3867 = n3865 | n3866 ;
  assign n3869 = ( x102 & ~n3868 ) | ( x102 & n3867 ) | ( ~n3868 & n3867 ) ;
  assign n3870 = ( x101 & ~x102 ) | ( x101 & n3693 ) | ( ~x102 & n3693 ) ;
  assign n3871 = ( x101 & x102 ) | ( x101 & n3693 ) | ( x102 & n3693 ) ;
  assign n3872 = ( ~x102 & ~n3870 ) | ( ~x102 & n3871 ) | ( ~n3870 & n3871 ) ;
  assign n3873 = ( n3869 & ~n139 ) | ( n3869 & n3872 ) | ( ~n139 & n3872 ) ;
  assign n3874 = n139 | n3873 ;
  assign n3875 = ( x2 & ~n3869 ) | ( x2 & n3874 ) | ( ~n3869 & n3874 ) ;
  assign n3876 = ( n3869 & ~x2 ) | ( n3869 & n3874 ) | ( ~x2 & n3874 ) ;
  assign n3877 = ( n3875 & ~n3874 ) | ( n3875 & n3876 ) | ( ~n3874 & n3876 ) ;
  assign n3878 = ( n3863 & n3864 ) | ( n3863 & n3877 ) | ( n3864 & n3877 ) ;
  assign n3879 = ( n3864 & ~n3863 ) | ( n3864 & n3877 ) | ( ~n3863 & n3877 ) ;
  assign n3880 = ( n3863 & ~n3878 ) | ( n3863 & n3879 ) | ( ~n3878 & n3879 ) ;
  assign n3884 = x98 &  n225 ;
  assign n3881 = ( x100 & ~n197 ) | ( x100 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n3882 = x99 &  n192 ;
  assign n3883 = n3881 | n3882 ;
  assign n3885 = ( x98 & ~n3884 ) | ( x98 & n3883 ) | ( ~n3884 & n3883 ) ;
  assign n3886 = n200 | n3354 ;
  assign n3887 = ~n3885 & n3886 ;
  assign n3888 = x5 &  n3887 ;
  assign n3889 = x5 | n3887 ;
  assign n3890 = ~n3888 & n3889 ;
  assign n4023 = x92 &  n503 ;
  assign n4020 = ( x94 & ~n450 ) | ( x94 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n4021 = x93 &  n445 ;
  assign n4022 = n4020 | n4021 ;
  assign n4024 = ( x92 & ~n4023 ) | ( x92 & n4022 ) | ( ~n4023 & n4022 ) ;
  assign n4025 = ~n453 & n2401 ;
  assign n4026 = n4024 | n4025 ;
  assign n4027 = ( x11 & ~n4026 ) | ( x11 & 1'b0 ) | ( ~n4026 & 1'b0 ) ;
  assign n4028 = ~x11 & n4026 ;
  assign n4029 = n4027 | n4028 ;
  assign n3914 = x71 &  n2718 ;
  assign n3911 = ( x73 & ~n2642 ) | ( x73 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n3912 = x72 &  n2637 ;
  assign n3913 = n3911 | n3912 ;
  assign n3915 = ( x71 & ~n3914 ) | ( x71 & n3913 ) | ( ~n3914 & n3913 ) ;
  assign n3916 = ( n389 & ~n2645 ) | ( n389 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n3917 = n3915 | n3916 ;
  assign n3918 = ( x32 & ~n3917 ) | ( x32 & 1'b0 ) | ( ~n3917 & 1'b0 ) ;
  assign n3919 = ~x32 & n3917 ;
  assign n3920 = n3918 | n3919 ;
  assign n3921 = ( x38 & ~x39 ) | ( x38 & 1'b0 ) | ( ~x39 & 1'b0 ) ;
  assign n3922 = ~x38 & x39 ;
  assign n3923 = n3921 | n3922 ;
  assign n3924 = x64 &  n3923 ;
  assign n3925 = ( x38 & n3763 ) | ( x38 & n3764 ) | ( n3763 & n3764 ) ;
  assign n3926 = ( x38 & ~n3925 ) | ( x38 & 1'b0 ) | ( ~n3925 & 1'b0 ) ;
  assign n3930 = x65 &  n3756 ;
  assign n3927 = ( x67 & ~n3602 ) | ( x67 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n3928 = x66 &  n3597 ;
  assign n3929 = n3927 | n3928 ;
  assign n3931 = ( x65 & ~n3930 ) | ( x65 & n3929 ) | ( ~n3930 & n3929 ) ;
  assign n3932 = n173 | n3605 ;
  assign n3933 = ~n3931 & n3932 ;
  assign n3934 = x38 &  n3933 ;
  assign n3935 = x38 | n3933 ;
  assign n3936 = ~n3934 & n3935 ;
  assign n3937 = ( n3924 & ~n3926 ) | ( n3924 & n3936 ) | ( ~n3926 & n3936 ) ;
  assign n3938 = ( n3924 & ~n3936 ) | ( n3924 & n3926 ) | ( ~n3936 & n3926 ) ;
  assign n3939 = ( n3937 & ~n3924 ) | ( n3937 & n3938 ) | ( ~n3924 & n3938 ) ;
  assign n3943 = x68 &  n3214 ;
  assign n3940 = ( x70 & ~n3087 ) | ( x70 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n3941 = x69 &  n3082 ;
  assign n3942 = n3940 | n3941 ;
  assign n3944 = ( x68 & ~n3943 ) | ( x68 & n3942 ) | ( ~n3943 & n3942 ) ;
  assign n3945 = ( n282 & ~n3090 ) | ( n282 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n3946 = n3944 | n3945 ;
  assign n3947 = ( x35 & ~n3946 ) | ( x35 & 1'b0 ) | ( ~n3946 & 1'b0 ) ;
  assign n3948 = ~x35 & n3946 ;
  assign n3949 = n3947 | n3948 ;
  assign n3950 = ( n3612 & n3768 ) | ( n3612 & n3778 ) | ( n3768 & n3778 ) ;
  assign n3951 = ( n3939 & ~n3949 ) | ( n3939 & n3950 ) | ( ~n3949 & n3950 ) ;
  assign n3952 = ( n3939 & ~n3950 ) | ( n3939 & n3949 ) | ( ~n3950 & n3949 ) ;
  assign n3953 = ( n3951 & ~n3939 ) | ( n3951 & n3952 ) | ( ~n3939 & n3952 ) ;
  assign n3954 = ( n3615 & n3781 ) | ( n3615 & n3791 ) | ( n3781 & n3791 ) ;
  assign n3955 = ( n3920 & ~n3953 ) | ( n3920 & n3954 ) | ( ~n3953 & n3954 ) ;
  assign n3956 = ( n3920 & ~n3954 ) | ( n3920 & n3953 ) | ( ~n3954 & n3953 ) ;
  assign n3957 = ( n3955 & ~n3920 ) | ( n3955 & n3956 ) | ( ~n3920 & n3956 ) ;
  assign n3904 = x74 &  n2312 ;
  assign n3901 = ( x76 & ~n2195 ) | ( x76 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n3902 = x75 &  n2190 ;
  assign n3903 = n3901 | n3902 ;
  assign n3905 = ( x74 & ~n3904 ) | ( x74 & n3903 ) | ( ~n3904 & n3903 ) ;
  assign n3906 = ( n603 & ~n2198 ) | ( n603 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n3907 = n3905 | n3906 ;
  assign n3908 = ( x29 & ~n3907 ) | ( x29 & 1'b0 ) | ( ~n3907 & 1'b0 ) ;
  assign n3909 = ~x29 & n3907 ;
  assign n3910 = n3908 | n3909 ;
  assign n3958 = ( n3796 & ~n3957 ) | ( n3796 & n3910 ) | ( ~n3957 & n3910 ) ;
  assign n3959 = ( n3910 & ~n3796 ) | ( n3910 & n3957 ) | ( ~n3796 & n3957 ) ;
  assign n3960 = ( n3958 & ~n3910 ) | ( n3958 & n3959 ) | ( ~n3910 & n3959 ) ;
  assign n3961 = ( n3621 & n3797 ) | ( n3621 & n3807 ) | ( n3797 & n3807 ) ;
  assign n3965 = x77 &  n1894 ;
  assign n3962 = ( x79 & ~n1816 ) | ( x79 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n3963 = x78 &  n1811 ;
  assign n3964 = n3962 | n3963 ;
  assign n3966 = ( x77 & ~n3965 ) | ( x77 & n3964 ) | ( ~n3965 & n3964 ) ;
  assign n3967 = ( n766 & ~n1819 ) | ( n766 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n3968 = n3966 | n3967 ;
  assign n3969 = ( x26 & ~n3968 ) | ( x26 & 1'b0 ) | ( ~n3968 & 1'b0 ) ;
  assign n3970 = ~x26 & n3968 ;
  assign n3971 = n3969 | n3970 ;
  assign n3972 = ( n3960 & ~n3961 ) | ( n3960 & n3971 ) | ( ~n3961 & n3971 ) ;
  assign n3973 = ( n3961 & ~n3960 ) | ( n3961 & n3971 ) | ( ~n3960 & n3971 ) ;
  assign n3974 = ( n3972 & ~n3971 ) | ( n3972 & n3973 ) | ( ~n3971 & n3973 ) ;
  assign n3979 = x80 &  n1551 ;
  assign n3976 = ( x82 & ~n1451 ) | ( x82 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n3977 = x81 &  n1446 ;
  assign n3978 = n3976 | n3977 ;
  assign n3980 = ( x80 & ~n3979 ) | ( x80 & n3978 ) | ( ~n3979 & n3978 ) ;
  assign n3981 = ( n1084 & ~n1454 ) | ( n1084 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n3982 = n3980 | n3981 ;
  assign n3983 = ( x23 & ~n3982 ) | ( x23 & 1'b0 ) | ( ~n3982 & 1'b0 ) ;
  assign n3984 = ~x23 & n3982 ;
  assign n3985 = n3983 | n3984 ;
  assign n3975 = ( n3810 & n3820 ) | ( n3810 & n3821 ) | ( n3820 & n3821 ) ;
  assign n3986 = ( n3974 & ~n3985 ) | ( n3974 & n3975 ) | ( ~n3985 & n3975 ) ;
  assign n3987 = ( n3974 & ~n3975 ) | ( n3974 & n3985 ) | ( ~n3975 & n3985 ) ;
  assign n3988 = ( n3986 & ~n3974 ) | ( n3986 & n3987 ) | ( ~n3974 & n3987 ) ;
  assign n3894 = x83 &  n1227 ;
  assign n3891 = ( x85 & ~n1154 ) | ( x85 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n3892 = x84 &  n1149 ;
  assign n3893 = n3891 | n3892 ;
  assign n3895 = ( x83 & ~n3894 ) | ( x83 & n3893 ) | ( ~n3894 & n3893 ) ;
  assign n3896 = ~n1157 & n1295 ;
  assign n3897 = n3895 | n3896 ;
  assign n3898 = ( x20 & ~n3897 ) | ( x20 & 1'b0 ) | ( ~n3897 & 1'b0 ) ;
  assign n3899 = ~x20 & n3897 ;
  assign n3900 = n3898 | n3899 ;
  assign n3989 = ( n3825 & ~n3988 ) | ( n3825 & n3900 ) | ( ~n3988 & n3900 ) ;
  assign n3990 = ( n3900 & ~n3825 ) | ( n3900 & n3988 ) | ( ~n3825 & n3988 ) ;
  assign n3991 = ( n3989 & ~n3900 ) | ( n3989 & n3990 ) | ( ~n3900 & n3990 ) ;
  assign n3992 = ( n3641 & n3827 ) | ( n3641 & n3837 ) | ( n3827 & n3837 ) ;
  assign n3996 = x86 &  n942 ;
  assign n3993 = ( x88 & ~n896 ) | ( x88 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n3994 = x87 &  n891 ;
  assign n3995 = n3993 | n3994 ;
  assign n3997 = ( x86 & ~n3996 ) | ( x86 & n3995 ) | ( ~n3996 & n3995 ) ;
  assign n3998 = ~n899 & n1624 ;
  assign n3999 = n3997 | n3998 ;
  assign n4000 = ( x17 & ~n3999 ) | ( x17 & 1'b0 ) | ( ~n3999 & 1'b0 ) ;
  assign n4001 = ~x17 & n3999 ;
  assign n4002 = n4000 | n4001 ;
  assign n4003 = ( n3991 & ~n3992 ) | ( n3991 & n4002 ) | ( ~n3992 & n4002 ) ;
  assign n4004 = ( n3991 & ~n4002 ) | ( n3991 & n3992 ) | ( ~n4002 & n3992 ) ;
  assign n4005 = ( n4003 & ~n3991 ) | ( n4003 & n4004 ) | ( ~n3991 & n4004 ) ;
  assign n4006 = ( n3840 & n3841 ) | ( n3840 & n3851 ) | ( n3841 & n3851 ) ;
  assign n4010 = x89 &  n713 ;
  assign n4007 = ( x91 & ~n641 ) | ( x91 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n4008 = x90 &  n636 ;
  assign n4009 = n4007 | n4008 ;
  assign n4011 = ( x89 & ~n4010 ) | ( x89 & n4009 ) | ( ~n4010 & n4009 ) ;
  assign n4012 = ~n644 & n2108 ;
  assign n4013 = n4011 | n4012 ;
  assign n4014 = ( x14 & ~n4013 ) | ( x14 & 1'b0 ) | ( ~n4013 & 1'b0 ) ;
  assign n4015 = ~x14 & n4013 ;
  assign n4016 = n4014 | n4015 ;
  assign n4017 = ( n4005 & ~n4006 ) | ( n4005 & n4016 ) | ( ~n4006 & n4016 ) ;
  assign n4018 = ( n4006 & ~n4005 ) | ( n4006 & n4016 ) | ( ~n4005 & n4016 ) ;
  assign n4019 = ( n4017 & ~n4016 ) | ( n4017 & n4018 ) | ( ~n4016 & n4018 ) ;
  assign n4030 = ( n3856 & ~n4029 ) | ( n3856 & n4019 ) | ( ~n4029 & n4019 ) ;
  assign n4031 = ( n4019 & ~n3856 ) | ( n4019 & n4029 ) | ( ~n3856 & n4029 ) ;
  assign n4032 = ( n4030 & ~n4019 ) | ( n4030 & n4031 ) | ( ~n4019 & n4031 ) ;
  assign n4036 = x95 &  n353 ;
  assign n4033 = ( x97 & ~n313 ) | ( x97 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n4034 = x96 &  n308 ;
  assign n4035 = n4033 | n4034 ;
  assign n4037 = ( x95 & ~n4036 ) | ( x95 & n4035 ) | ( ~n4036 & n4035 ) ;
  assign n4038 = ~n316 & n2999 ;
  assign n4039 = n4037 | n4038 ;
  assign n4040 = ( x8 & ~n4039 ) | ( x8 & 1'b0 ) | ( ~n4039 & 1'b0 ) ;
  assign n4041 = ~x8 & n4039 ;
  assign n4042 = n4040 | n4041 ;
  assign n4043 = ( n4032 & ~n3859 ) | ( n4032 & n4042 ) | ( ~n3859 & n4042 ) ;
  assign n4044 = ( n3859 & ~n4032 ) | ( n3859 & n4042 ) | ( ~n4032 & n4042 ) ;
  assign n4045 = ( n4043 & ~n4042 ) | ( n4043 & n4044 ) | ( ~n4042 & n4044 ) ;
  assign n4047 = ( n3861 & n3890 ) | ( n3861 & n4045 ) | ( n3890 & n4045 ) ;
  assign n4046 = ( n3890 & ~n3861 ) | ( n3890 & n4045 ) | ( ~n3861 & n4045 ) ;
  assign n4048 = ( n3861 & ~n4047 ) | ( n3861 & n4046 ) | ( ~n4047 & n4046 ) ;
  assign n4052 = ~n136 & x103 ;
  assign n4049 = ( x101 & ~n150 ) | ( x101 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n4050 = ( x102 & ~n131 ) | ( x102 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n4051 = n4049 | n4050 ;
  assign n4053 = ( x103 & ~n4052 ) | ( x103 & n4051 ) | ( ~n4052 & n4051 ) ;
  assign n4054 = ( x102 & ~x103 ) | ( x102 & n3871 ) | ( ~x103 & n3871 ) ;
  assign n4055 = ( x102 & x103 ) | ( x102 & n3871 ) | ( x103 & n3871 ) ;
  assign n4056 = ( ~x103 & ~n4054 ) | ( ~x103 & n4055 ) | ( ~n4054 & n4055 ) ;
  assign n4057 = ( n4053 & ~n139 ) | ( n4053 & n4056 ) | ( ~n139 & n4056 ) ;
  assign n4058 = n139 | n4057 ;
  assign n4059 = ( x2 & ~n4053 ) | ( x2 & n4058 ) | ( ~n4053 & n4058 ) ;
  assign n4060 = ( n4053 & ~x2 ) | ( n4053 & n4058 ) | ( ~x2 & n4058 ) ;
  assign n4061 = ( n4059 & ~n4058 ) | ( n4059 & n4060 ) | ( ~n4058 & n4060 ) ;
  assign n4063 = ( n3878 & n4048 ) | ( n3878 & n4061 ) | ( n4048 & n4061 ) ;
  assign n4062 = ( n3878 & ~n4048 ) | ( n3878 & n4061 ) | ( ~n4048 & n4061 ) ;
  assign n4064 = ( n4048 & ~n4063 ) | ( n4048 & n4062 ) | ( ~n4063 & n4062 ) ;
  assign n4245 = ~n136 & x104 ;
  assign n4242 = ( x102 & ~n150 ) | ( x102 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n4243 = ( x103 & ~n131 ) | ( x103 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n4244 = n4242 | n4243 ;
  assign n4246 = ( x104 & ~n4245 ) | ( x104 & n4244 ) | ( ~n4245 & n4244 ) ;
  assign n4247 = ( x103 & ~x104 ) | ( x103 & n4055 ) | ( ~x104 & n4055 ) ;
  assign n4248 = ( x103 & x104 ) | ( x103 & n4055 ) | ( x104 & n4055 ) ;
  assign n4249 = ( ~x104 & ~n4247 ) | ( ~x104 & n4248 ) | ( ~n4247 & n4248 ) ;
  assign n4250 = ( n4246 & ~n139 ) | ( n4246 & n4249 ) | ( ~n139 & n4249 ) ;
  assign n4251 = n139 | n4250 ;
  assign n4253 = ( x2 & n4246 ) | ( x2 & n4251 ) | ( n4246 & n4251 ) ;
  assign n4252 = ( x2 & ~n4251 ) | ( x2 & n4246 ) | ( ~n4251 & n4246 ) ;
  assign n4254 = ( n4251 & ~n4253 ) | ( n4251 & n4252 ) | ( ~n4253 & n4252 ) ;
  assign n4078 = x96 &  n353 ;
  assign n4075 = ( x98 & ~n313 ) | ( x98 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n4076 = x97 &  n308 ;
  assign n4077 = n4075 | n4076 ;
  assign n4079 = ( x96 & ~n4078 ) | ( x96 & n4077 ) | ( ~n4078 & n4077 ) ;
  assign n4080 = ~n316 & n3170 ;
  assign n4081 = n4079 | n4080 ;
  assign n4082 = ( x8 & ~n4081 ) | ( x8 & 1'b0 ) | ( ~n4081 & 1'b0 ) ;
  assign n4083 = ~x8 & n4081 ;
  assign n4084 = n4082 | n4083 ;
  assign n4088 = x90 &  n713 ;
  assign n4085 = ( x92 & ~n641 ) | ( x92 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n4086 = x91 &  n636 ;
  assign n4087 = n4085 | n4086 ;
  assign n4089 = ( x90 & ~n4088 ) | ( x90 & n4087 ) | ( ~n4088 & n4087 ) ;
  assign n4090 = ~n644 & n2248 ;
  assign n4091 = n4089 | n4090 ;
  assign n4092 = ( x14 & ~n4091 ) | ( x14 & 1'b0 ) | ( ~n4091 & 1'b0 ) ;
  assign n4093 = ~x14 & n4091 ;
  assign n4094 = n4092 | n4093 ;
  assign n4098 = x87 &  n942 ;
  assign n4095 = ( x89 & ~n896 ) | ( x89 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n4096 = x88 &  n891 ;
  assign n4097 = n4095 | n4096 ;
  assign n4099 = ( x87 & ~n4098 ) | ( x87 & n4097 ) | ( ~n4098 & n4097 ) ;
  assign n4100 = ~n899 & n1741 ;
  assign n4101 = n4099 | n4100 ;
  assign n4102 = ( x17 & ~n4101 ) | ( x17 & 1'b0 ) | ( ~n4101 & 1'b0 ) ;
  assign n4103 = ~x17 & n4101 ;
  assign n4104 = n4102 | n4103 ;
  assign n4108 = x84 &  n1227 ;
  assign n4105 = ( x86 & ~n1154 ) | ( x86 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n4106 = x85 &  n1149 ;
  assign n4107 = n4105 | n4106 ;
  assign n4109 = ( x84 & ~n4108 ) | ( x84 & n4107 ) | ( ~n4108 & n4107 ) ;
  assign n4110 = ~n1157 & n1496 ;
  assign n4111 = n4109 | n4110 ;
  assign n4112 = ( x20 & ~n4111 ) | ( x20 & 1'b0 ) | ( ~n4111 & 1'b0 ) ;
  assign n4113 = ~x20 & n4111 ;
  assign n4114 = n4112 | n4113 ;
  assign n4118 = x81 &  n1551 ;
  assign n4115 = ( x83 & ~n1451 ) | ( x83 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n4116 = x82 &  n1446 ;
  assign n4117 = n4115 | n4116 ;
  assign n4119 = ( x81 & ~n4118 ) | ( x81 & n4117 ) | ( ~n4118 & n4117 ) ;
  assign n4120 = ( n1100 & ~n1454 ) | ( n1100 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n4121 = n4119 | n4120 ;
  assign n4122 = ( x23 & ~n4121 ) | ( x23 & 1'b0 ) | ( ~n4121 & 1'b0 ) ;
  assign n4123 = ~x23 & n4121 ;
  assign n4124 = n4122 | n4123 ;
  assign n4172 = x72 &  n2718 ;
  assign n4169 = ( x74 & ~n2642 ) | ( x74 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n4170 = x73 &  n2637 ;
  assign n4171 = n4169 | n4170 ;
  assign n4173 = ( x72 & ~n4172 ) | ( x72 & n4171 ) | ( ~n4172 & n4171 ) ;
  assign n4174 = ( n482 & ~n2645 ) | ( n482 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n4175 = n4173 | n4174 ;
  assign n4176 = ( x32 & ~n4175 ) | ( x32 & 1'b0 ) | ( ~n4175 & 1'b0 ) ;
  assign n4177 = ~x32 & n4175 ;
  assign n4178 = n4176 | n4177 ;
  assign n4128 = x66 &  n3756 ;
  assign n4125 = ( x68 & ~n3602 ) | ( x68 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n4126 = x67 &  n3597 ;
  assign n4127 = n4125 | n4126 ;
  assign n4129 = ( x66 & ~n4128 ) | ( x66 & n4127 ) | ( ~n4128 & n4127 ) ;
  assign n4130 = ( n213 & ~n3605 ) | ( n213 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n4131 = n4129 | n4130 ;
  assign n4132 = ( x38 & ~n4131 ) | ( x38 & 1'b0 ) | ( ~n4131 & 1'b0 ) ;
  assign n4133 = ~x38 & n4131 ;
  assign n4134 = n4132 | n4133 ;
  assign n4135 = ( x41 & ~n3924 ) | ( x41 & 1'b0 ) | ( ~n3924 & 1'b0 ) ;
  assign n4136 = ( x39 & x40 ) | ( x39 & n3921 ) | ( x40 & n3921 ) ;
  assign n4137 = ( x39 & ~n3922 ) | ( x39 & x40 ) | ( ~n3922 & x40 ) ;
  assign n4138 = ~n4136 &  n4137 ;
  assign n4139 = x64 &  n4138 ;
  assign n4140 = ~x40 & x41 ;
  assign n4141 = ( x40 & ~x41 ) | ( x40 & 1'b0 ) | ( ~x41 & 1'b0 ) ;
  assign n4142 = n4140 | n4141 ;
  assign n4143 = ~n3923 |  n4142 ;
  assign n4144 = ( x65 & ~n4143 ) | ( x65 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n4145 = n4139 | n4144 ;
  assign n4146 = ~n3923 | ~n4142 ;
  assign n4147 = ( n142 & ~n4146 ) | ( n142 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n4148 = n4145 | n4147 ;
  assign n4150 = ( x41 & n4135 ) | ( x41 & n4148 ) | ( n4135 & n4148 ) ;
  assign n4149 = ( x41 & ~n4135 ) | ( x41 & n4148 ) | ( ~n4135 & n4148 ) ;
  assign n4151 = ( n4135 & ~n4150 ) | ( n4135 & n4149 ) | ( ~n4150 & n4149 ) ;
  assign n4153 = ( n3938 & n4134 ) | ( n3938 & n4151 ) | ( n4134 & n4151 ) ;
  assign n4152 = ( n3938 & ~n4134 ) | ( n3938 & n4151 ) | ( ~n4134 & n4151 ) ;
  assign n4154 = ( n4134 & ~n4153 ) | ( n4134 & n4152 ) | ( ~n4153 & n4152 ) ;
  assign n4165 = ( n3949 & ~n3939 ) | ( n3949 & n3950 ) | ( ~n3939 & n3950 ) ;
  assign n4158 = x69 &  n3214 ;
  assign n4155 = ( x71 & ~n3087 ) | ( x71 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n4156 = x70 &  n3082 ;
  assign n4157 = n4155 | n4156 ;
  assign n4159 = ( x69 & ~n4158 ) | ( x69 & n4157 ) | ( ~n4158 & n4157 ) ;
  assign n4160 = ( n298 & ~n3090 ) | ( n298 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n4161 = n4159 | n4160 ;
  assign n4162 = ( x35 & ~n4161 ) | ( x35 & 1'b0 ) | ( ~n4161 & 1'b0 ) ;
  assign n4163 = ~x35 & n4161 ;
  assign n4164 = n4162 | n4163 ;
  assign n4166 = ( n4154 & ~n4165 ) | ( n4154 & n4164 ) | ( ~n4165 & n4164 ) ;
  assign n4167 = ( n4154 & ~n4164 ) | ( n4154 & n4165 ) | ( ~n4164 & n4165 ) ;
  assign n4168 = ( n4166 & ~n4154 ) | ( n4166 & n4167 ) | ( ~n4154 & n4167 ) ;
  assign n4179 = ( n3955 & ~n4178 ) | ( n3955 & n4168 ) | ( ~n4178 & n4168 ) ;
  assign n4180 = ( n4168 & ~n3955 ) | ( n4168 & n4178 ) | ( ~n3955 & n4178 ) ;
  assign n4181 = ( n4179 & ~n4168 ) | ( n4179 & n4180 ) | ( ~n4168 & n4180 ) ;
  assign n4185 = x75 &  n2312 ;
  assign n4182 = ( x77 & ~n2195 ) | ( x77 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n4183 = x76 &  n2190 ;
  assign n4184 = n4182 | n4183 ;
  assign n4186 = ( x75 & ~n4185 ) | ( x75 & n4184 ) | ( ~n4185 & n4184 ) ;
  assign n4187 = ( n677 & ~n2198 ) | ( n677 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n4188 = n4186 | n4187 ;
  assign n4189 = ( x29 & ~n4188 ) | ( x29 & 1'b0 ) | ( ~n4188 & 1'b0 ) ;
  assign n4190 = ~x29 & n4188 ;
  assign n4191 = n4189 | n4190 ;
  assign n4192 = ( n4181 & ~n3958 ) | ( n4181 & n4191 ) | ( ~n3958 & n4191 ) ;
  assign n4193 = ( n3958 & ~n4191 ) | ( n3958 & n4181 ) | ( ~n4191 & n4181 ) ;
  assign n4194 = ( n4192 & ~n4181 ) | ( n4192 & n4193 ) | ( ~n4181 & n4193 ) ;
  assign n4198 = x78 &  n1894 ;
  assign n4195 = ( x80 & ~n1816 ) | ( x80 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n4196 = x79 &  n1811 ;
  assign n4197 = n4195 | n4196 ;
  assign n4199 = ( x78 & ~n4198 ) | ( x78 & n4197 ) | ( ~n4198 & n4197 ) ;
  assign n4200 = ( n842 & ~n1819 ) | ( n842 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n4201 = n4199 | n4200 ;
  assign n4202 = ( x26 & ~n4201 ) | ( x26 & 1'b0 ) | ( ~n4201 & 1'b0 ) ;
  assign n4203 = ~x26 & n4201 ;
  assign n4204 = n4202 | n4203 ;
  assign n4205 = ( n4194 & ~n3973 ) | ( n4194 & n4204 ) | ( ~n3973 & n4204 ) ;
  assign n4206 = ( n3973 & ~n4204 ) | ( n3973 & n4194 ) | ( ~n4204 & n4194 ) ;
  assign n4207 = ( n4205 & ~n4194 ) | ( n4205 & n4206 ) | ( ~n4194 & n4206 ) ;
  assign n4208 = ( n3975 & ~n3974 ) | ( n3975 & n3985 ) | ( ~n3974 & n3985 ) ;
  assign n4209 = ( n4124 & n4207 ) | ( n4124 & n4208 ) | ( n4207 & n4208 ) ;
  assign n4210 = ( n4207 & ~n4124 ) | ( n4207 & n4208 ) | ( ~n4124 & n4208 ) ;
  assign n4211 = ( n4124 & ~n4209 ) | ( n4124 & n4210 ) | ( ~n4209 & n4210 ) ;
  assign n4212 = ( n3989 & n4114 ) | ( n3989 & n4211 ) | ( n4114 & n4211 ) ;
  assign n4213 = ( n3989 & ~n4114 ) | ( n3989 & n4211 ) | ( ~n4114 & n4211 ) ;
  assign n4214 = ( n4114 & ~n4212 ) | ( n4114 & n4213 ) | ( ~n4212 & n4213 ) ;
  assign n4215 = ( n3992 & ~n3991 ) | ( n3992 & n4002 ) | ( ~n3991 & n4002 ) ;
  assign n4216 = ( n4104 & n4214 ) | ( n4104 & n4215 ) | ( n4214 & n4215 ) ;
  assign n4217 = ( n4214 & ~n4104 ) | ( n4214 & n4215 ) | ( ~n4104 & n4215 ) ;
  assign n4218 = ( n4104 & ~n4216 ) | ( n4104 & n4217 ) | ( ~n4216 & n4217 ) ;
  assign n4220 = ( n4018 & n4094 ) | ( n4018 & n4218 ) | ( n4094 & n4218 ) ;
  assign n4219 = ( n4018 & ~n4094 ) | ( n4018 & n4218 ) | ( ~n4094 & n4218 ) ;
  assign n4221 = ( n4094 & ~n4220 ) | ( n4094 & n4219 ) | ( ~n4220 & n4219 ) ;
  assign n4222 = ( n3856 & ~n4019 ) | ( n3856 & n4029 ) | ( ~n4019 & n4029 ) ;
  assign n4226 = x93 &  n503 ;
  assign n4223 = ( x95 & ~n450 ) | ( x95 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n4224 = x94 &  n445 ;
  assign n4225 = n4223 | n4224 ;
  assign n4227 = ( x93 & ~n4226 ) | ( x93 & n4225 ) | ( ~n4226 & n4225 ) ;
  assign n4228 = ~n453 & n2547 ;
  assign n4229 = n4227 | n4228 ;
  assign n4230 = ( x11 & ~n4229 ) | ( x11 & 1'b0 ) | ( ~n4229 & 1'b0 ) ;
  assign n4231 = ~x11 & n4229 ;
  assign n4232 = n4230 | n4231 ;
  assign n4233 = ( n4221 & ~n4222 ) | ( n4221 & n4232 ) | ( ~n4222 & n4232 ) ;
  assign n4234 = ( n4221 & ~n4232 ) | ( n4221 & n4222 ) | ( ~n4232 & n4222 ) ;
  assign n4235 = ( n4233 & ~n4221 ) | ( n4233 & n4234 ) | ( ~n4221 & n4234 ) ;
  assign n4237 = ( n4044 & n4084 ) | ( n4044 & n4235 ) | ( n4084 & n4235 ) ;
  assign n4236 = ( n4044 & ~n4084 ) | ( n4044 & n4235 ) | ( ~n4084 & n4235 ) ;
  assign n4238 = ( n4084 & ~n4237 ) | ( n4084 & n4236 ) | ( ~n4237 & n4236 ) ;
  assign n4068 = x99 &  n225 ;
  assign n4065 = ( x101 & ~n197 ) | ( x101 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n4066 = x100 &  n192 ;
  assign n4067 = n4065 | n4066 ;
  assign n4069 = ( x99 & ~n4068 ) | ( x99 & n4067 ) | ( ~n4068 & n4067 ) ;
  assign n4070 = n200 | n3694 ;
  assign n4071 = ~n4069 & n4070 ;
  assign n4072 = x5 &  n4071 ;
  assign n4073 = x5 | n4071 ;
  assign n4074 = ~n4072 & n4073 ;
  assign n4239 = ( n4046 & n4074 ) | ( n4046 & n4238 ) | ( n4074 & n4238 ) ;
  assign n4240 = ( n4046 & ~n4238 ) | ( n4046 & n4074 ) | ( ~n4238 & n4074 ) ;
  assign n4241 = ( n4238 & ~n4239 ) | ( n4238 & n4240 ) | ( ~n4239 & n4240 ) ;
  assign n4255 = ( n4062 & ~n4254 ) | ( n4062 & n4241 ) | ( ~n4254 & n4241 ) ;
  assign n4256 = ( n4241 & ~n4062 ) | ( n4241 & n4254 ) | ( ~n4062 & n4254 ) ;
  assign n4257 = ( n4255 & ~n4241 ) | ( n4255 & n4256 ) | ( ~n4241 & n4256 ) ;
  assign n4261 = x100 &  n225 ;
  assign n4258 = ( x102 & ~n197 ) | ( x102 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n4259 = x101 &  n192 ;
  assign n4260 = n4258 | n4259 ;
  assign n4262 = ( x100 & ~n4261 ) | ( x100 & n4260 ) | ( ~n4261 & n4260 ) ;
  assign n4263 = n200 | n3872 ;
  assign n4264 = ~n4262 & n4263 ;
  assign n4265 = x5 &  n4264 ;
  assign n4266 = x5 | n4264 ;
  assign n4267 = ~n4265 & n4266 ;
  assign n4281 = x94 &  n503 ;
  assign n4278 = ( x96 & ~n450 ) | ( x96 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n4279 = x95 &  n445 ;
  assign n4280 = n4278 | n4279 ;
  assign n4282 = ( x94 & ~n4281 ) | ( x94 & n4280 ) | ( ~n4281 & n4280 ) ;
  assign n4283 = ~n453 & n2836 ;
  assign n4284 = n4282 | n4283 ;
  assign n4285 = ( x11 & ~n4284 ) | ( x11 & 1'b0 ) | ( ~n4284 & 1'b0 ) ;
  assign n4286 = ~x11 & n4284 ;
  assign n4287 = n4285 | n4286 ;
  assign n4288 = ( n4221 & n4222 ) | ( n4221 & n4232 ) | ( n4222 & n4232 ) ;
  assign n4292 = x91 &  n713 ;
  assign n4289 = ( x93 & ~n641 ) | ( x93 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n4290 = x92 &  n636 ;
  assign n4291 = n4289 | n4290 ;
  assign n4293 = ( x91 & ~n4292 ) | ( x91 & n4291 ) | ( ~n4292 & n4291 ) ;
  assign n4294 = n644 | n2264 ;
  assign n4295 = ~n4293 & n4294 ;
  assign n4296 = x14 &  n4295 ;
  assign n4297 = x14 | n4295 ;
  assign n4298 = ~n4296 & n4297 ;
  assign n4302 = x88 &  n942 ;
  assign n4299 = ( x90 & ~n896 ) | ( x90 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n4300 = x89 &  n891 ;
  assign n4301 = n4299 | n4300 ;
  assign n4303 = ( x88 & ~n4302 ) | ( x88 & n4301 ) | ( ~n4302 & n4301 ) ;
  assign n4304 = ~n899 & n1976 ;
  assign n4305 = n4303 | n4304 ;
  assign n4306 = ( x17 & ~n4305 ) | ( x17 & 1'b0 ) | ( ~n4305 & 1'b0 ) ;
  assign n4307 = ~x17 & n4305 ;
  assign n4308 = n4306 | n4307 ;
  assign n4409 = x85 &  n1227 ;
  assign n4406 = ( x87 & ~n1154 ) | ( x87 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n4407 = x86 &  n1149 ;
  assign n4408 = n4406 | n4407 ;
  assign n4410 = ( x85 & ~n4409 ) | ( x85 & n4408 ) | ( ~n4409 & n4408 ) ;
  assign n4411 = ~n1157 & n1512 ;
  assign n4412 = n4410 | n4411 ;
  assign n4413 = ( x20 & ~n4412 ) | ( x20 & 1'b0 ) | ( ~n4412 & 1'b0 ) ;
  assign n4414 = ~x20 & n4412 ;
  assign n4415 = n4413 | n4414 ;
  assign n4312 = x79 &  n1894 ;
  assign n4309 = ( x81 & ~n1816 ) | ( x81 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n4310 = x80 &  n1811 ;
  assign n4311 = n4309 | n4310 ;
  assign n4313 = ( x79 & ~n4312 ) | ( x79 & n4311 ) | ( ~n4312 & n4311 ) ;
  assign n4314 = ( n994 & ~n1819 ) | ( n994 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n4315 = n4313 | n4314 ;
  assign n4316 = ( x26 & ~n4315 ) | ( x26 & 1'b0 ) | ( ~n4315 & 1'b0 ) ;
  assign n4317 = ~x26 & n4315 ;
  assign n4318 = n4316 | n4317 ;
  assign n4319 = ( n3973 & n4194 ) | ( n3973 & n4204 ) | ( n4194 & n4204 ) ;
  assign n4323 = x76 &  n2312 ;
  assign n4320 = ( x78 & ~n2195 ) | ( x78 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n4321 = x77 &  n2190 ;
  assign n4322 = n4320 | n4321 ;
  assign n4324 = ( x76 & ~n4323 ) | ( x76 & n4322 ) | ( ~n4323 & n4322 ) ;
  assign n4325 = ( n693 & ~n2198 ) | ( n693 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n4326 = n4324 | n4325 ;
  assign n4327 = ( x29 & ~n4326 ) | ( x29 & 1'b0 ) | ( ~n4326 & 1'b0 ) ;
  assign n4328 = ~x29 & n4326 ;
  assign n4329 = n4327 | n4328 ;
  assign n4330 = ( n3958 & n4181 ) | ( n3958 & n4191 ) | ( n4181 & n4191 ) ;
  assign n4334 = x70 &  n3214 ;
  assign n4331 = ( x72 & ~n3087 ) | ( x72 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n4332 = x71 &  n3082 ;
  assign n4333 = n4331 | n4332 ;
  assign n4335 = ( x70 & ~n4334 ) | ( x70 & n4333 ) | ( ~n4334 & n4333 ) ;
  assign n4336 = ( n345 & ~n3090 ) | ( n345 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n4337 = n4335 | n4336 ;
  assign n4339 = x35 &  n4337 ;
  assign n4338 = ~x35 & n4337 ;
  assign n4340 = ( x35 & ~n4339 ) | ( x35 & n4338 ) | ( ~n4339 & n4338 ) ;
  assign n4341 = ( n4154 & n4164 ) | ( n4154 & n4165 ) | ( n4164 & n4165 ) ;
  assign n4360 = x67 &  n3756 ;
  assign n4357 = ( x69 & ~n3602 ) | ( x69 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n4358 = x68 &  n3597 ;
  assign n4359 = n4357 | n4358 ;
  assign n4361 = ( x67 & ~n4360 ) | ( x67 & n4359 ) | ( ~n4360 & n4359 ) ;
  assign n4362 = ( n246 & ~n3605 ) | ( n246 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n4363 = n4361 | n4362 ;
  assign n4364 = ( x38 & ~n4363 ) | ( x38 & 1'b0 ) | ( ~n4363 & 1'b0 ) ;
  assign n4365 = ~x38 & n4363 ;
  assign n4366 = n4364 | n4365 ;
  assign n4343 = ( x39 & ~x40 ) | ( x39 & n4142 ) | ( ~x40 & n4142 ) ;
  assign n4342 = ( x39 & ~x40 ) | ( x39 & n3923 ) | ( ~x40 & n3923 ) ;
  assign n4344 = ~n4343 |  n4342 ;
  assign n4348 = x64 &  n4344 ;
  assign n4345 = ( x66 & ~n4143 ) | ( x66 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n4346 = x65 &  n4138 ;
  assign n4347 = n4345 | n4346 ;
  assign n4349 = ( x64 & ~n4348 ) | ( x64 & n4347 ) | ( ~n4348 & n4347 ) ;
  assign n4350 = ( n157 & ~n4146 ) | ( n157 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n4351 = n4349 | n4350 ;
  assign n4352 = ( x41 & n3924 ) | ( x41 & n4148 ) | ( n3924 & n4148 ) ;
  assign n4353 = ( x41 & ~n4352 ) | ( x41 & 1'b0 ) | ( ~n4352 & 1'b0 ) ;
  assign n4355 = ( x41 & n4351 ) | ( x41 & n4353 ) | ( n4351 & n4353 ) ;
  assign n4354 = ( n4351 & ~x41 ) | ( n4351 & n4353 ) | ( ~x41 & n4353 ) ;
  assign n4356 = ( x41 & ~n4355 ) | ( x41 & n4354 ) | ( ~n4355 & n4354 ) ;
  assign n4367 = ( n4153 & ~n4366 ) | ( n4153 & n4356 ) | ( ~n4366 & n4356 ) ;
  assign n4368 = ( n4356 & ~n4153 ) | ( n4356 & n4366 ) | ( ~n4153 & n4366 ) ;
  assign n4369 = ( n4367 & ~n4356 ) | ( n4367 & n4368 ) | ( ~n4356 & n4368 ) ;
  assign n4371 = ( n4340 & n4341 ) | ( n4340 & n4369 ) | ( n4341 & n4369 ) ;
  assign n4370 = ( n4341 & ~n4340 ) | ( n4341 & n4369 ) | ( ~n4340 & n4369 ) ;
  assign n4372 = ( n4340 & ~n4371 ) | ( n4340 & n4370 ) | ( ~n4371 & n4370 ) ;
  assign n4373 = ( n3955 & n4168 ) | ( n3955 & n4178 ) | ( n4168 & n4178 ) ;
  assign n4377 = x73 &  n2718 ;
  assign n4374 = ( x75 & ~n2642 ) | ( x75 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n4375 = x74 &  n2637 ;
  assign n4376 = n4374 | n4375 ;
  assign n4378 = ( x73 & ~n4377 ) | ( x73 & n4376 ) | ( ~n4377 & n4376 ) ;
  assign n4379 = ( n540 & ~n2645 ) | ( n540 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n4380 = n4378 | n4379 ;
  assign n4381 = ( x32 & ~n4380 ) | ( x32 & 1'b0 ) | ( ~n4380 & 1'b0 ) ;
  assign n4382 = ~x32 & n4380 ;
  assign n4383 = n4381 | n4382 ;
  assign n4384 = ( n4372 & ~n4373 ) | ( n4372 & n4383 ) | ( ~n4373 & n4383 ) ;
  assign n4385 = ( n4372 & ~n4383 ) | ( n4372 & n4373 ) | ( ~n4383 & n4373 ) ;
  assign n4386 = ( n4384 & ~n4372 ) | ( n4384 & n4385 ) | ( ~n4372 & n4385 ) ;
  assign n4388 = ( n4329 & n4330 ) | ( n4329 & n4386 ) | ( n4330 & n4386 ) ;
  assign n4387 = ( n4330 & ~n4329 ) | ( n4330 & n4386 ) | ( ~n4329 & n4386 ) ;
  assign n4389 = ( n4329 & ~n4388 ) | ( n4329 & n4387 ) | ( ~n4388 & n4387 ) ;
  assign n4391 = ( n4318 & n4319 ) | ( n4318 & n4389 ) | ( n4319 & n4389 ) ;
  assign n4390 = ( n4319 & ~n4318 ) | ( n4319 & n4389 ) | ( ~n4318 & n4389 ) ;
  assign n4392 = ( n4318 & ~n4391 ) | ( n4318 & n4390 ) | ( ~n4391 & n4390 ) ;
  assign n4396 = x82 &  n1551 ;
  assign n4393 = ( x84 & ~n1451 ) | ( x84 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n4394 = x83 &  n1446 ;
  assign n4395 = n4393 | n4394 ;
  assign n4397 = ( x82 & ~n4396 ) | ( x82 & n4395 ) | ( ~n4396 & n4395 ) ;
  assign n4398 = ( n1199 & ~n1454 ) | ( n1199 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n4399 = n4397 | n4398 ;
  assign n4400 = ( x23 & ~n4399 ) | ( x23 & 1'b0 ) | ( ~n4399 & 1'b0 ) ;
  assign n4401 = ~x23 & n4399 ;
  assign n4402 = n4400 | n4401 ;
  assign n4403 = ( n4392 & ~n4209 ) | ( n4392 & n4402 ) | ( ~n4209 & n4402 ) ;
  assign n4404 = ( n4209 & ~n4402 ) | ( n4209 & n4392 ) | ( ~n4402 & n4392 ) ;
  assign n4405 = ( n4403 & ~n4392 ) | ( n4403 & n4404 ) | ( ~n4392 & n4404 ) ;
  assign n4416 = ( n4212 & ~n4415 ) | ( n4212 & n4405 ) | ( ~n4415 & n4405 ) ;
  assign n4417 = ( n4405 & ~n4212 ) | ( n4405 & n4415 ) | ( ~n4212 & n4415 ) ;
  assign n4418 = ( n4416 & ~n4405 ) | ( n4416 & n4417 ) | ( ~n4405 & n4417 ) ;
  assign n4419 = ( n4216 & n4308 ) | ( n4216 & n4418 ) | ( n4308 & n4418 ) ;
  assign n4420 = ( n4308 & ~n4216 ) | ( n4308 & n4418 ) | ( ~n4216 & n4418 ) ;
  assign n4421 = ( n4216 & ~n4419 ) | ( n4216 & n4420 ) | ( ~n4419 & n4420 ) ;
  assign n4422 = ( n4220 & n4298 ) | ( n4220 & n4421 ) | ( n4298 & n4421 ) ;
  assign n4423 = ( n4220 & ~n4298 ) | ( n4220 & n4421 ) | ( ~n4298 & n4421 ) ;
  assign n4424 = ( n4298 & ~n4422 ) | ( n4298 & n4423 ) | ( ~n4422 & n4423 ) ;
  assign n4425 = ( n4287 & ~n4288 ) | ( n4287 & n4424 ) | ( ~n4288 & n4424 ) ;
  assign n4426 = ( n4287 & ~n4424 ) | ( n4287 & n4288 ) | ( ~n4424 & n4288 ) ;
  assign n4427 = ( n4425 & ~n4287 ) | ( n4425 & n4426 ) | ( ~n4287 & n4426 ) ;
  assign n4271 = x97 &  n353 ;
  assign n4268 = ( x99 & ~n313 ) | ( x99 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n4269 = x98 &  n308 ;
  assign n4270 = n4268 | n4269 ;
  assign n4272 = ( x97 & ~n4271 ) | ( x97 & n4270 ) | ( ~n4271 & n4270 ) ;
  assign n4273 = ~n316 & n3338 ;
  assign n4274 = n4272 | n4273 ;
  assign n4275 = ( x8 & ~n4274 ) | ( x8 & 1'b0 ) | ( ~n4274 & 1'b0 ) ;
  assign n4276 = ~x8 & n4274 ;
  assign n4277 = n4275 | n4276 ;
  assign n4428 = ( n4237 & n4277 ) | ( n4237 & n4427 ) | ( n4277 & n4427 ) ;
  assign n4429 = ( n4237 & ~n4427 ) | ( n4237 & n4277 ) | ( ~n4427 & n4277 ) ;
  assign n4430 = ( n4427 & ~n4428 ) | ( n4427 & n4429 ) | ( ~n4428 & n4429 ) ;
  assign n4431 = ( n4240 & n4267 ) | ( n4240 & n4430 ) | ( n4267 & n4430 ) ;
  assign n4432 = ( n4267 & ~n4240 ) | ( n4267 & n4430 ) | ( ~n4240 & n4430 ) ;
  assign n4433 = ( n4240 & ~n4431 ) | ( n4240 & n4432 ) | ( ~n4431 & n4432 ) ;
  assign n4434 = ( n4062 & ~n4241 ) | ( n4062 & n4254 ) | ( ~n4241 & n4254 ) ;
  assign n4438 = ~n136 & x105 ;
  assign n4435 = ( x103 & ~n150 ) | ( x103 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n4436 = ( x104 & ~n131 ) | ( x104 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n4437 = n4435 | n4436 ;
  assign n4439 = ( x105 & ~n4438 ) | ( x105 & n4437 ) | ( ~n4438 & n4437 ) ;
  assign n4441 = ( x104 & x105 ) | ( x104 & n4248 ) | ( x105 & n4248 ) ;
  assign n4440 = ( x104 & ~x105 ) | ( x104 & n4248 ) | ( ~x105 & n4248 ) ;
  assign n4442 = ( x105 & ~n4441 ) | ( x105 & n4440 ) | ( ~n4441 & n4440 ) ;
  assign n4443 = ( n139 & ~n4439 ) | ( n139 & n4442 ) | ( ~n4439 & n4442 ) ;
  assign n4444 = ~n139 & n4443 ;
  assign n4445 = ( x2 & n4439 ) | ( x2 & n4444 ) | ( n4439 & n4444 ) ;
  assign n4446 = ( x2 & ~n4444 ) | ( x2 & n4439 ) | ( ~n4444 & n4439 ) ;
  assign n4447 = ( n4444 & ~n4445 ) | ( n4444 & n4446 ) | ( ~n4445 & n4446 ) ;
  assign n4448 = ( n4433 & n4434 ) | ( n4433 & n4447 ) | ( n4434 & n4447 ) ;
  assign n4449 = ( n4434 & ~n4433 ) | ( n4434 & n4447 ) | ( ~n4433 & n4447 ) ;
  assign n4450 = ( n4433 & ~n4448 ) | ( n4433 & n4449 ) | ( ~n4448 & n4449 ) ;
  assign n4454 = ~n136 & x106 ;
  assign n4451 = ( x104 & ~n150 ) | ( x104 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n4452 = ( x105 & ~n131 ) | ( x105 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n4453 = n4451 | n4452 ;
  assign n4455 = ( x106 & ~n4454 ) | ( x106 & n4453 ) | ( ~n4454 & n4453 ) ;
  assign n4457 = ( x105 & x106 ) | ( x105 & n4441 ) | ( x106 & n4441 ) ;
  assign n4456 = ( x105 & ~x106 ) | ( x105 & n4441 ) | ( ~x106 & n4441 ) ;
  assign n4458 = ( x106 & ~n4457 ) | ( x106 & n4456 ) | ( ~n4457 & n4456 ) ;
  assign n4459 = ( n139 & ~n4455 ) | ( n139 & n4458 ) | ( ~n4455 & n4458 ) ;
  assign n4460 = ~n139 & n4459 ;
  assign n4461 = ( x2 & n4455 ) | ( x2 & n4460 ) | ( n4455 & n4460 ) ;
  assign n4462 = ( x2 & ~n4460 ) | ( x2 & n4455 ) | ( ~n4460 & n4455 ) ;
  assign n4463 = ( n4460 & ~n4461 ) | ( n4460 & n4462 ) | ( ~n4461 & n4462 ) ;
  assign n4477 = x98 &  n353 ;
  assign n4474 = ( x100 & ~n313 ) | ( x100 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n4475 = x99 &  n308 ;
  assign n4476 = n4474 | n4475 ;
  assign n4478 = ( x98 & ~n4477 ) | ( x98 & n4476 ) | ( ~n4477 & n4476 ) ;
  assign n4479 = n316 | n3354 ;
  assign n4480 = ~n4478 & n4479 ;
  assign n4481 = x8 &  n4480 ;
  assign n4482 = x8 | n4480 ;
  assign n4483 = ~n4481 & n4482 ;
  assign n4614 = x92 &  n713 ;
  assign n4611 = ( x94 & ~n641 ) | ( x94 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n4612 = x93 &  n636 ;
  assign n4613 = n4611 | n4612 ;
  assign n4615 = ( x92 & ~n4614 ) | ( x92 & n4613 ) | ( ~n4614 & n4613 ) ;
  assign n4616 = ~n644 & n2401 ;
  assign n4617 = n4615 | n4616 ;
  assign n4618 = ( x14 & ~n4617 ) | ( x14 & 1'b0 ) | ( ~n4617 & 1'b0 ) ;
  assign n4619 = ~x14 & n4617 ;
  assign n4620 = n4618 | n4619 ;
  assign n4570 = x80 &  n1894 ;
  assign n4567 = ( x82 & ~n1816 ) | ( x82 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n4568 = x81 &  n1811 ;
  assign n4569 = n4567 | n4568 ;
  assign n4571 = ( x80 & ~n4570 ) | ( x80 & n4569 ) | ( ~n4570 & n4569 ) ;
  assign n4572 = ( n1084 & ~n1819 ) | ( n1084 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n4573 = n4571 | n4572 ;
  assign n4574 = ( x26 & ~n4573 ) | ( x26 & 1'b0 ) | ( ~n4573 & 1'b0 ) ;
  assign n4575 = ~x26 & n4573 ;
  assign n4576 = n4574 | n4575 ;
  assign n4557 = x77 &  n2312 ;
  assign n4554 = ( x79 & ~n2195 ) | ( x79 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n4555 = x78 &  n2190 ;
  assign n4556 = n4554 | n4555 ;
  assign n4558 = ( x77 & ~n4557 ) | ( x77 & n4556 ) | ( ~n4557 & n4556 ) ;
  assign n4559 = ( n766 & ~n2198 ) | ( n766 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n4560 = n4558 | n4559 ;
  assign n4561 = ( x29 & ~n4560 ) | ( x29 & 1'b0 ) | ( ~n4560 & 1'b0 ) ;
  assign n4562 = ~x29 & n4560 ;
  assign n4563 = n4561 | n4562 ;
  assign n4497 = x74 &  n2718 ;
  assign n4494 = ( x76 & ~n2642 ) | ( x76 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n4495 = x75 &  n2637 ;
  assign n4496 = n4494 | n4495 ;
  assign n4498 = ( x74 & ~n4497 ) | ( x74 & n4496 ) | ( ~n4497 & n4496 ) ;
  assign n4499 = ( n603 & ~n2645 ) | ( n603 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n4500 = n4498 | n4499 ;
  assign n4501 = ( x32 & ~n4500 ) | ( x32 & 1'b0 ) | ( ~n4500 & 1'b0 ) ;
  assign n4502 = ~x32 & n4500 ;
  assign n4503 = n4501 | n4502 ;
  assign n4504 = ( n4372 & n4373 ) | ( n4372 & n4383 ) | ( n4373 & n4383 ) ;
  assign n4505 = ( x41 & ~x42 ) | ( x41 & 1'b0 ) | ( ~x42 & 1'b0 ) ;
  assign n4506 = ~x41 & x42 ;
  assign n4507 = n4505 | n4506 ;
  assign n4508 = x64 &  n4507 ;
  assign n4509 = ( x41 & n4351 ) | ( x41 & n4352 ) | ( n4351 & n4352 ) ;
  assign n4510 = ( x41 & ~n4509 ) | ( x41 & 1'b0 ) | ( ~n4509 & 1'b0 ) ;
  assign n4514 = x65 &  n4344 ;
  assign n4511 = ( x67 & ~n4143 ) | ( x67 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n4512 = x66 &  n4138 ;
  assign n4513 = n4511 | n4512 ;
  assign n4515 = ( x65 & ~n4514 ) | ( x65 & n4513 ) | ( ~n4514 & n4513 ) ;
  assign n4516 = n173 | n4146 ;
  assign n4517 = ~n4515 & n4516 ;
  assign n4518 = x41 &  n4517 ;
  assign n4519 = x41 | n4517 ;
  assign n4520 = ~n4518 & n4519 ;
  assign n4521 = ( n4508 & ~n4510 ) | ( n4508 & n4520 ) | ( ~n4510 & n4520 ) ;
  assign n4522 = ( n4508 & ~n4520 ) | ( n4508 & n4510 ) | ( ~n4520 & n4510 ) ;
  assign n4523 = ( n4521 & ~n4508 ) | ( n4521 & n4522 ) | ( ~n4508 & n4522 ) ;
  assign n4527 = x68 &  n3756 ;
  assign n4524 = ( x70 & ~n3602 ) | ( x70 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n4525 = x69 &  n3597 ;
  assign n4526 = n4524 | n4525 ;
  assign n4528 = ( x68 & ~n4527 ) | ( x68 & n4526 ) | ( ~n4527 & n4526 ) ;
  assign n4529 = ( n282 & ~n3605 ) | ( n282 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n4530 = n4528 | n4529 ;
  assign n4531 = ( x38 & ~n4530 ) | ( x38 & 1'b0 ) | ( ~n4530 & 1'b0 ) ;
  assign n4532 = ~x38 & n4530 ;
  assign n4533 = n4531 | n4532 ;
  assign n4534 = ( n4153 & n4356 ) | ( n4153 & n4366 ) | ( n4356 & n4366 ) ;
  assign n4535 = ( n4523 & ~n4533 ) | ( n4523 & n4534 ) | ( ~n4533 & n4534 ) ;
  assign n4536 = ( n4523 & ~n4534 ) | ( n4523 & n4533 ) | ( ~n4534 & n4533 ) ;
  assign n4537 = ( n4535 & ~n4523 ) | ( n4535 & n4536 ) | ( ~n4523 & n4536 ) ;
  assign n4541 = x71 &  n3214 ;
  assign n4538 = ( x73 & ~n3087 ) | ( x73 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n4539 = x72 &  n3082 ;
  assign n4540 = n4538 | n4539 ;
  assign n4542 = ( x71 & ~n4541 ) | ( x71 & n4540 ) | ( ~n4541 & n4540 ) ;
  assign n4543 = ( n389 & ~n3090 ) | ( n389 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n4544 = n4542 | n4543 ;
  assign n4545 = ( x35 & ~n4544 ) | ( x35 & 1'b0 ) | ( ~n4544 & 1'b0 ) ;
  assign n4546 = ~x35 & n4544 ;
  assign n4547 = n4545 | n4546 ;
  assign n4548 = ( n4537 & ~n4371 ) | ( n4537 & n4547 ) | ( ~n4371 & n4547 ) ;
  assign n4549 = ( n4371 & ~n4547 ) | ( n4371 & n4537 ) | ( ~n4547 & n4537 ) ;
  assign n4550 = ( n4548 & ~n4537 ) | ( n4548 & n4549 ) | ( ~n4537 & n4549 ) ;
  assign n4551 = ( n4503 & ~n4504 ) | ( n4503 & n4550 ) | ( ~n4504 & n4550 ) ;
  assign n4552 = ( n4503 & ~n4550 ) | ( n4503 & n4504 ) | ( ~n4550 & n4504 ) ;
  assign n4553 = ( n4551 & ~n4503 ) | ( n4551 & n4552 ) | ( ~n4503 & n4552 ) ;
  assign n4564 = ( n4388 & ~n4563 ) | ( n4388 & n4553 ) | ( ~n4563 & n4553 ) ;
  assign n4565 = ( n4553 & ~n4388 ) | ( n4553 & n4563 ) | ( ~n4388 & n4563 ) ;
  assign n4566 = ( n4564 & ~n4553 ) | ( n4564 & n4565 ) | ( ~n4553 & n4565 ) ;
  assign n4577 = ( n4391 & ~n4576 ) | ( n4391 & n4566 ) | ( ~n4576 & n4566 ) ;
  assign n4578 = ( n4566 & ~n4391 ) | ( n4566 & n4576 ) | ( ~n4391 & n4576 ) ;
  assign n4579 = ( n4577 & ~n4566 ) | ( n4577 & n4578 ) | ( ~n4566 & n4578 ) ;
  assign n4583 = x83 &  n1551 ;
  assign n4580 = ( x85 & ~n1451 ) | ( x85 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n4581 = x84 &  n1446 ;
  assign n4582 = n4580 | n4581 ;
  assign n4584 = ( x83 & ~n4583 ) | ( x83 & n4582 ) | ( ~n4583 & n4582 ) ;
  assign n4585 = ( n1295 & ~n1454 ) | ( n1295 & 1'b0 ) | ( ~n1454 & 1'b0 ) ;
  assign n4586 = n4584 | n4585 ;
  assign n4587 = ( x23 & ~n4586 ) | ( x23 & 1'b0 ) | ( ~n4586 & 1'b0 ) ;
  assign n4588 = ~x23 & n4586 ;
  assign n4589 = n4587 | n4588 ;
  assign n4590 = ( n4209 & n4392 ) | ( n4209 & n4402 ) | ( n4392 & n4402 ) ;
  assign n4591 = ( n4579 & ~n4589 ) | ( n4579 & n4590 ) | ( ~n4589 & n4590 ) ;
  assign n4592 = ( n4579 & ~n4590 ) | ( n4579 & n4589 ) | ( ~n4590 & n4589 ) ;
  assign n4593 = ( n4591 & ~n4579 ) | ( n4591 & n4592 ) | ( ~n4579 & n4592 ) ;
  assign n4594 = ( n4212 & n4405 ) | ( n4212 & n4415 ) | ( n4405 & n4415 ) ;
  assign n4598 = x86 &  n1227 ;
  assign n4595 = ( x88 & ~n1154 ) | ( x88 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n4596 = x87 &  n1149 ;
  assign n4597 = n4595 | n4596 ;
  assign n4599 = ( x86 & ~n4598 ) | ( x86 & n4597 ) | ( ~n4598 & n4597 ) ;
  assign n4600 = ~n1157 & n1624 ;
  assign n4601 = n4599 | n4600 ;
  assign n4602 = ( x20 & ~n4601 ) | ( x20 & 1'b0 ) | ( ~n4601 & 1'b0 ) ;
  assign n4603 = ~x20 & n4601 ;
  assign n4604 = n4602 | n4603 ;
  assign n4605 = ( n4593 & ~n4594 ) | ( n4593 & n4604 ) | ( ~n4594 & n4604 ) ;
  assign n4606 = ( n4593 & ~n4604 ) | ( n4593 & n4594 ) | ( ~n4604 & n4594 ) ;
  assign n4607 = ( n4605 & ~n4593 ) | ( n4605 & n4606 ) | ( ~n4593 & n4606 ) ;
  assign n4487 = x89 &  n942 ;
  assign n4484 = ( x91 & ~n896 ) | ( x91 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n4485 = x90 &  n891 ;
  assign n4486 = n4484 | n4485 ;
  assign n4488 = ( x89 & ~n4487 ) | ( x89 & n4486 ) | ( ~n4487 & n4486 ) ;
  assign n4489 = ~n899 & n2108 ;
  assign n4490 = n4488 | n4489 ;
  assign n4491 = ( x17 & ~n4490 ) | ( x17 & 1'b0 ) | ( ~n4490 & 1'b0 ) ;
  assign n4492 = ~x17 & n4490 ;
  assign n4493 = n4491 | n4492 ;
  assign n4608 = ( n4419 & n4493 ) | ( n4419 & n4607 ) | ( n4493 & n4607 ) ;
  assign n4609 = ( n4419 & ~n4607 ) | ( n4419 & n4493 ) | ( ~n4607 & n4493 ) ;
  assign n4610 = ( n4607 & ~n4608 ) | ( n4607 & n4609 ) | ( ~n4608 & n4609 ) ;
  assign n4621 = ( n4423 & ~n4620 ) | ( n4423 & n4610 ) | ( ~n4620 & n4610 ) ;
  assign n4622 = ( n4610 & ~n4423 ) | ( n4610 & n4620 ) | ( ~n4423 & n4620 ) ;
  assign n4623 = ( n4621 & ~n4610 ) | ( n4621 & n4622 ) | ( ~n4610 & n4622 ) ;
  assign n4627 = x95 &  n503 ;
  assign n4624 = ( x97 & ~n450 ) | ( x97 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n4625 = x96 &  n445 ;
  assign n4626 = n4624 | n4625 ;
  assign n4628 = ( x95 & ~n4627 ) | ( x95 & n4626 ) | ( ~n4627 & n4626 ) ;
  assign n4629 = ~n453 & n2999 ;
  assign n4630 = n4628 | n4629 ;
  assign n4631 = ( x11 & ~n4630 ) | ( x11 & 1'b0 ) | ( ~n4630 & 1'b0 ) ;
  assign n4632 = ~x11 & n4630 ;
  assign n4633 = n4631 | n4632 ;
  assign n4634 = ( n4623 & ~n4426 ) | ( n4623 & n4633 ) | ( ~n4426 & n4633 ) ;
  assign n4635 = ( n4426 & ~n4623 ) | ( n4426 & n4633 ) | ( ~n4623 & n4633 ) ;
  assign n4636 = ( n4634 & ~n4633 ) | ( n4634 & n4635 ) | ( ~n4633 & n4635 ) ;
  assign n4638 = ( n4429 & n4483 ) | ( n4429 & n4636 ) | ( n4483 & n4636 ) ;
  assign n4637 = ( n4483 & ~n4429 ) | ( n4483 & n4636 ) | ( ~n4429 & n4636 ) ;
  assign n4639 = ( n4429 & ~n4638 ) | ( n4429 & n4637 ) | ( ~n4638 & n4637 ) ;
  assign n4467 = x101 &  n225 ;
  assign n4464 = ( x103 & ~n197 ) | ( x103 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n4465 = x102 &  n192 ;
  assign n4466 = n4464 | n4465 ;
  assign n4468 = ( x101 & ~n4467 ) | ( x101 & n4466 ) | ( ~n4467 & n4466 ) ;
  assign n4469 = n200 | n4056 ;
  assign n4470 = ~n4468 & n4469 ;
  assign n4471 = x5 &  n4470 ;
  assign n4472 = x5 | n4470 ;
  assign n4473 = ~n4471 & n4472 ;
  assign n4641 = ( n4431 & n4473 ) | ( n4431 & n4639 ) | ( n4473 & n4639 ) ;
  assign n4640 = ( n4431 & ~n4639 ) | ( n4431 & n4473 ) | ( ~n4639 & n4473 ) ;
  assign n4642 = ( n4639 & ~n4641 ) | ( n4639 & n4640 ) | ( ~n4641 & n4640 ) ;
  assign n4643 = ( n4433 & ~n4447 ) | ( n4433 & n4434 ) | ( ~n4447 & n4434 ) ;
  assign n4645 = ( n4463 & n4642 ) | ( n4463 & n4643 ) | ( n4642 & n4643 ) ;
  assign n4644 = ( n4642 & ~n4463 ) | ( n4642 & n4643 ) | ( ~n4463 & n4643 ) ;
  assign n4646 = ( n4463 & ~n4645 ) | ( n4463 & n4644 ) | ( ~n4645 & n4644 ) ;
  assign n4660 = x99 &  n353 ;
  assign n4657 = ( x101 & ~n313 ) | ( x101 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n4658 = x100 &  n308 ;
  assign n4659 = n4657 | n4658 ;
  assign n4661 = ( x99 & ~n4660 ) | ( x99 & n4659 ) | ( ~n4660 & n4659 ) ;
  assign n4662 = n316 | n3694 ;
  assign n4663 = ~n4661 & n4662 ;
  assign n4664 = x8 &  n4663 ;
  assign n4665 = x8 | n4663 ;
  assign n4666 = ~n4664 & n4665 ;
  assign n4680 = x87 &  n1227 ;
  assign n4677 = ( x89 & ~n1154 ) | ( x89 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n4678 = x88 &  n1149 ;
  assign n4679 = n4677 | n4678 ;
  assign n4681 = ( x87 & ~n4680 ) | ( x87 & n4679 ) | ( ~n4680 & n4679 ) ;
  assign n4682 = ~n1157 & n1741 ;
  assign n4683 = n4681 | n4682 ;
  assign n4684 = ( x20 & ~n4683 ) | ( x20 & 1'b0 ) | ( ~n4683 & 1'b0 ) ;
  assign n4685 = ~x20 & n4683 ;
  assign n4686 = n4684 | n4685 ;
  assign n4690 = x84 &  n1551 ;
  assign n4687 = ( x86 & ~n1451 ) | ( x86 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n4688 = x85 &  n1446 ;
  assign n4689 = n4687 | n4688 ;
  assign n4691 = ( x84 & ~n4690 ) | ( x84 & n4689 ) | ( ~n4690 & n4689 ) ;
  assign n4692 = ~n1454 & n1496 ;
  assign n4693 = n4691 | n4692 ;
  assign n4694 = ( x23 & ~n4693 ) | ( x23 & 1'b0 ) | ( ~n4693 & 1'b0 ) ;
  assign n4695 = ~x23 & n4693 ;
  assign n4696 = n4694 | n4695 ;
  assign n4700 = x81 &  n1894 ;
  assign n4697 = ( x83 & ~n1816 ) | ( x83 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n4698 = x82 &  n1811 ;
  assign n4699 = n4697 | n4698 ;
  assign n4701 = ( x81 & ~n4700 ) | ( x81 & n4699 ) | ( ~n4700 & n4699 ) ;
  assign n4702 = ( n1100 & ~n1819 ) | ( n1100 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n4703 = n4701 | n4702 ;
  assign n4704 = ( x26 & ~n4703 ) | ( x26 & 1'b0 ) | ( ~n4703 & 1'b0 ) ;
  assign n4705 = ~x26 & n4703 ;
  assign n4706 = n4704 | n4705 ;
  assign n4710 = x66 &  n4344 ;
  assign n4707 = ( x68 & ~n4143 ) | ( x68 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n4708 = x67 &  n4138 ;
  assign n4709 = n4707 | n4708 ;
  assign n4711 = ( x66 & ~n4710 ) | ( x66 & n4709 ) | ( ~n4710 & n4709 ) ;
  assign n4712 = ( n213 & ~n4146 ) | ( n213 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n4713 = n4711 | n4712 ;
  assign n4714 = ( x41 & ~n4713 ) | ( x41 & 1'b0 ) | ( ~n4713 & 1'b0 ) ;
  assign n4715 = ~x41 & n4713 ;
  assign n4716 = n4714 | n4715 ;
  assign n4717 = ( x44 & ~n4508 ) | ( x44 & 1'b0 ) | ( ~n4508 & 1'b0 ) ;
  assign n4718 = ( x42 & x43 ) | ( x42 & n4505 ) | ( x43 & n4505 ) ;
  assign n4719 = ( x42 & ~n4506 ) | ( x42 & x43 ) | ( ~n4506 & x43 ) ;
  assign n4720 = ~n4718 &  n4719 ;
  assign n4721 = x64 &  n4720 ;
  assign n4722 = ~x43 & x44 ;
  assign n4723 = ( x43 & ~x44 ) | ( x43 & 1'b0 ) | ( ~x44 & 1'b0 ) ;
  assign n4724 = n4722 | n4723 ;
  assign n4725 = ~n4507 |  n4724 ;
  assign n4726 = ( x65 & ~n4725 ) | ( x65 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n4727 = n4721 | n4726 ;
  assign n4728 = ~n4507 | ~n4724 ;
  assign n4729 = ( n142 & ~n4728 ) | ( n142 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n4730 = n4727 | n4729 ;
  assign n4732 = ( x44 & n4717 ) | ( x44 & n4730 ) | ( n4717 & n4730 ) ;
  assign n4731 = ( x44 & ~n4717 ) | ( x44 & n4730 ) | ( ~n4717 & n4730 ) ;
  assign n4733 = ( n4717 & ~n4732 ) | ( n4717 & n4731 ) | ( ~n4732 & n4731 ) ;
  assign n4735 = ( n4522 & n4716 ) | ( n4522 & n4733 ) | ( n4716 & n4733 ) ;
  assign n4734 = ( n4522 & ~n4716 ) | ( n4522 & n4733 ) | ( ~n4716 & n4733 ) ;
  assign n4736 = ( n4716 & ~n4735 ) | ( n4716 & n4734 ) | ( ~n4735 & n4734 ) ;
  assign n4747 = ( n4533 & ~n4523 ) | ( n4533 & n4534 ) | ( ~n4523 & n4534 ) ;
  assign n4740 = x69 &  n3756 ;
  assign n4737 = ( x71 & ~n3602 ) | ( x71 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n4738 = x70 &  n3597 ;
  assign n4739 = n4737 | n4738 ;
  assign n4741 = ( x69 & ~n4740 ) | ( x69 & n4739 ) | ( ~n4740 & n4739 ) ;
  assign n4742 = ( n298 & ~n3605 ) | ( n298 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n4743 = n4741 | n4742 ;
  assign n4744 = ( x38 & ~n4743 ) | ( x38 & 1'b0 ) | ( ~n4743 & 1'b0 ) ;
  assign n4745 = ~x38 & n4743 ;
  assign n4746 = n4744 | n4745 ;
  assign n4748 = ( n4736 & ~n4747 ) | ( n4736 & n4746 ) | ( ~n4747 & n4746 ) ;
  assign n4749 = ( n4736 & ~n4746 ) | ( n4736 & n4747 ) | ( ~n4746 & n4747 ) ;
  assign n4750 = ( n4748 & ~n4736 ) | ( n4748 & n4749 ) | ( ~n4736 & n4749 ) ;
  assign n4755 = x72 &  n3214 ;
  assign n4752 = ( x74 & ~n3087 ) | ( x74 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n4753 = x73 &  n3082 ;
  assign n4754 = n4752 | n4753 ;
  assign n4756 = ( x72 & ~n4755 ) | ( x72 & n4754 ) | ( ~n4755 & n4754 ) ;
  assign n4757 = ( n482 & ~n3090 ) | ( n482 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n4758 = n4756 | n4757 ;
  assign n4759 = ( x35 & ~n4758 ) | ( x35 & 1'b0 ) | ( ~n4758 & 1'b0 ) ;
  assign n4760 = ~x35 & n4758 ;
  assign n4761 = n4759 | n4760 ;
  assign n4751 = ( n4371 & ~n4537 ) | ( n4371 & n4547 ) | ( ~n4537 & n4547 ) ;
  assign n4762 = ( n4750 & ~n4761 ) | ( n4750 & n4751 ) | ( ~n4761 & n4751 ) ;
  assign n4763 = ( n4750 & ~n4751 ) | ( n4750 & n4761 ) | ( ~n4751 & n4761 ) ;
  assign n4764 = ( n4762 & ~n4750 ) | ( n4762 & n4763 ) | ( ~n4750 & n4763 ) ;
  assign n4768 = x75 &  n2718 ;
  assign n4765 = ( x77 & ~n2642 ) | ( x77 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n4766 = x76 &  n2637 ;
  assign n4767 = n4765 | n4766 ;
  assign n4769 = ( x75 & ~n4768 ) | ( x75 & n4767 ) | ( ~n4768 & n4767 ) ;
  assign n4770 = ( n677 & ~n2645 ) | ( n677 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n4771 = n4769 | n4770 ;
  assign n4772 = ( x32 & ~n4771 ) | ( x32 & 1'b0 ) | ( ~n4771 & 1'b0 ) ;
  assign n4773 = ~x32 & n4771 ;
  assign n4774 = n4772 | n4773 ;
  assign n4775 = ( n4764 & ~n4552 ) | ( n4764 & n4774 ) | ( ~n4552 & n4774 ) ;
  assign n4776 = ( n4552 & ~n4774 ) | ( n4552 & n4764 ) | ( ~n4774 & n4764 ) ;
  assign n4777 = ( n4775 & ~n4764 ) | ( n4775 & n4776 ) | ( ~n4764 & n4776 ) ;
  assign n4788 = ( n4388 & ~n4553 ) | ( n4388 & n4563 ) | ( ~n4553 & n4563 ) ;
  assign n4781 = x78 &  n2312 ;
  assign n4778 = ( x80 & ~n2195 ) | ( x80 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n4779 = x79 &  n2190 ;
  assign n4780 = n4778 | n4779 ;
  assign n4782 = ( x78 & ~n4781 ) | ( x78 & n4780 ) | ( ~n4781 & n4780 ) ;
  assign n4783 = ( n842 & ~n2198 ) | ( n842 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n4784 = n4782 | n4783 ;
  assign n4785 = ( x29 & ~n4784 ) | ( x29 & 1'b0 ) | ( ~n4784 & 1'b0 ) ;
  assign n4786 = ~x29 & n4784 ;
  assign n4787 = n4785 | n4786 ;
  assign n4789 = ( n4777 & ~n4788 ) | ( n4777 & n4787 ) | ( ~n4788 & n4787 ) ;
  assign n4790 = ( n4777 & ~n4787 ) | ( n4777 & n4788 ) | ( ~n4787 & n4788 ) ;
  assign n4791 = ( n4789 & ~n4777 ) | ( n4789 & n4790 ) | ( ~n4777 & n4790 ) ;
  assign n4792 = ( n4391 & ~n4566 ) | ( n4391 & n4576 ) | ( ~n4566 & n4576 ) ;
  assign n4793 = ( n4706 & n4791 ) | ( n4706 & n4792 ) | ( n4791 & n4792 ) ;
  assign n4794 = ( n4791 & ~n4706 ) | ( n4791 & n4792 ) | ( ~n4706 & n4792 ) ;
  assign n4795 = ( n4706 & ~n4793 ) | ( n4706 & n4794 ) | ( ~n4793 & n4794 ) ;
  assign n4796 = ( n4589 & ~n4579 ) | ( n4589 & n4590 ) | ( ~n4579 & n4590 ) ;
  assign n4797 = ( n4696 & n4795 ) | ( n4696 & n4796 ) | ( n4795 & n4796 ) ;
  assign n4798 = ( n4795 & ~n4696 ) | ( n4795 & n4796 ) | ( ~n4696 & n4796 ) ;
  assign n4799 = ( n4696 & ~n4797 ) | ( n4696 & n4798 ) | ( ~n4797 & n4798 ) ;
  assign n4800 = ( n4594 & ~n4593 ) | ( n4594 & n4604 ) | ( ~n4593 & n4604 ) ;
  assign n4801 = ( n4686 & n4799 ) | ( n4686 & n4800 ) | ( n4799 & n4800 ) ;
  assign n4802 = ( n4799 & ~n4686 ) | ( n4799 & n4800 ) | ( ~n4686 & n4800 ) ;
  assign n4803 = ( n4686 & ~n4801 ) | ( n4686 & n4802 ) | ( ~n4801 & n4802 ) ;
  assign n4670 = x90 &  n942 ;
  assign n4667 = ( x92 & ~n896 ) | ( x92 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n4668 = x91 &  n891 ;
  assign n4669 = n4667 | n4668 ;
  assign n4671 = ( x90 & ~n4670 ) | ( x90 & n4669 ) | ( ~n4670 & n4669 ) ;
  assign n4672 = ~n899 & n2248 ;
  assign n4673 = n4671 | n4672 ;
  assign n4674 = ( x17 & ~n4673 ) | ( x17 & 1'b0 ) | ( ~n4673 & 1'b0 ) ;
  assign n4675 = ~x17 & n4673 ;
  assign n4676 = n4674 | n4675 ;
  assign n4804 = ( n4609 & n4676 ) | ( n4609 & n4803 ) | ( n4676 & n4803 ) ;
  assign n4805 = ( n4609 & ~n4803 ) | ( n4609 & n4676 ) | ( ~n4803 & n4676 ) ;
  assign n4806 = ( n4803 & ~n4804 ) | ( n4803 & n4805 ) | ( ~n4804 & n4805 ) ;
  assign n4807 = ( n4423 & ~n4610 ) | ( n4423 & n4620 ) | ( ~n4610 & n4620 ) ;
  assign n4811 = x93 &  n713 ;
  assign n4808 = ( x95 & ~n641 ) | ( x95 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n4809 = x94 &  n636 ;
  assign n4810 = n4808 | n4809 ;
  assign n4812 = ( x93 & ~n4811 ) | ( x93 & n4810 ) | ( ~n4811 & n4810 ) ;
  assign n4813 = ~n644 & n2547 ;
  assign n4814 = n4812 | n4813 ;
  assign n4815 = ( x14 & ~n4814 ) | ( x14 & 1'b0 ) | ( ~n4814 & 1'b0 ) ;
  assign n4816 = ~x14 & n4814 ;
  assign n4817 = n4815 | n4816 ;
  assign n4818 = ( n4806 & ~n4807 ) | ( n4806 & n4817 ) | ( ~n4807 & n4817 ) ;
  assign n4819 = ( n4806 & ~n4817 ) | ( n4806 & n4807 ) | ( ~n4817 & n4807 ) ;
  assign n4820 = ( n4818 & ~n4806 ) | ( n4818 & n4819 ) | ( ~n4806 & n4819 ) ;
  assign n4824 = x96 &  n503 ;
  assign n4821 = ( x98 & ~n450 ) | ( x98 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n4822 = x97 &  n445 ;
  assign n4823 = n4821 | n4822 ;
  assign n4825 = ( x96 & ~n4824 ) | ( x96 & n4823 ) | ( ~n4824 & n4823 ) ;
  assign n4826 = ~n453 & n3170 ;
  assign n4827 = n4825 | n4826 ;
  assign n4828 = ( x11 & ~n4827 ) | ( x11 & 1'b0 ) | ( ~n4827 & 1'b0 ) ;
  assign n4829 = ~x11 & n4827 ;
  assign n4830 = n4828 | n4829 ;
  assign n4831 = ( n4820 & ~n4635 ) | ( n4820 & n4830 ) | ( ~n4635 & n4830 ) ;
  assign n4832 = ( n4635 & ~n4830 ) | ( n4635 & n4820 ) | ( ~n4830 & n4820 ) ;
  assign n4833 = ( n4831 & ~n4820 ) | ( n4831 & n4832 ) | ( ~n4820 & n4832 ) ;
  assign n4834 = ( n4637 & n4666 ) | ( n4637 & n4833 ) | ( n4666 & n4833 ) ;
  assign n4835 = ( n4666 & ~n4637 ) | ( n4666 & n4833 ) | ( ~n4637 & n4833 ) ;
  assign n4836 = ( n4637 & ~n4834 ) | ( n4637 & n4835 ) | ( ~n4834 & n4835 ) ;
  assign n4650 = x102 &  n225 ;
  assign n4647 = ( x104 & ~n197 ) | ( x104 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n4648 = x103 &  n192 ;
  assign n4649 = n4647 | n4648 ;
  assign n4651 = ( x102 & ~n4650 ) | ( x102 & n4649 ) | ( ~n4650 & n4649 ) ;
  assign n4652 = n200 | n4249 ;
  assign n4653 = ~n4651 & n4652 ;
  assign n4654 = x5 &  n4653 ;
  assign n4655 = x5 | n4653 ;
  assign n4656 = ~n4654 & n4655 ;
  assign n4837 = ( n4640 & ~n4836 ) | ( n4640 & n4656 ) | ( ~n4836 & n4656 ) ;
  assign n4838 = ( n4640 & ~n4656 ) | ( n4640 & n4836 ) | ( ~n4656 & n4836 ) ;
  assign n4839 = ( n4837 & ~n4640 ) | ( n4837 & n4838 ) | ( ~n4640 & n4838 ) ;
  assign n4840 = ( n4463 & ~n4643 ) | ( n4463 & n4642 ) | ( ~n4643 & n4642 ) ;
  assign n4844 = ~n136 & x107 ;
  assign n4841 = ( x105 & ~n150 ) | ( x105 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n4842 = ( x106 & ~n131 ) | ( x106 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n4843 = n4841 | n4842 ;
  assign n4845 = ( x107 & ~n4844 ) | ( x107 & n4843 ) | ( ~n4844 & n4843 ) ;
  assign n4847 = ( x106 & x107 ) | ( x106 & n4457 ) | ( x107 & n4457 ) ;
  assign n4846 = ( x106 & ~x107 ) | ( x106 & n4457 ) | ( ~x107 & n4457 ) ;
  assign n4848 = ( x107 & ~n4847 ) | ( x107 & n4846 ) | ( ~n4847 & n4846 ) ;
  assign n4849 = ( n139 & ~n4845 ) | ( n139 & n4848 ) | ( ~n4845 & n4848 ) ;
  assign n4850 = ~n139 & n4849 ;
  assign n4851 = ( n4845 & ~x2 ) | ( n4845 & n4850 ) | ( ~x2 & n4850 ) ;
  assign n4852 = ( x2 & ~n4845 ) | ( x2 & n4850 ) | ( ~n4845 & n4850 ) ;
  assign n4853 = ( n4851 & ~n4850 ) | ( n4851 & n4852 ) | ( ~n4850 & n4852 ) ;
  assign n4854 = ( n4839 & n4840 ) | ( n4839 & n4853 ) | ( n4840 & n4853 ) ;
  assign n4855 = ( n4840 & ~n4839 ) | ( n4840 & n4853 ) | ( ~n4839 & n4853 ) ;
  assign n4856 = ( n4839 & ~n4854 ) | ( n4839 & n4855 ) | ( ~n4854 & n4855 ) ;
  assign n4860 = x103 &  n225 ;
  assign n4857 = ( x105 & ~n197 ) | ( x105 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n4858 = x104 &  n192 ;
  assign n4859 = n4857 | n4858 ;
  assign n4861 = ( x103 & ~n4860 ) | ( x103 & n4859 ) | ( ~n4860 & n4859 ) ;
  assign n4862 = ~n200 & n4442 ;
  assign n4863 = n4861 | n4862 ;
  assign n4864 = ( x5 & ~n4863 ) | ( x5 & 1'b0 ) | ( ~n4863 & 1'b0 ) ;
  assign n4865 = ~x5 & n4863 ;
  assign n4866 = n4864 | n4865 ;
  assign n4867 = ( n4637 & ~n4833 ) | ( n4637 & n4666 ) | ( ~n4833 & n4666 ) ;
  assign n4881 = x94 &  n713 ;
  assign n4878 = ( x96 & ~n641 ) | ( x96 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n4879 = x95 &  n636 ;
  assign n4880 = n4878 | n4879 ;
  assign n4882 = ( x94 & ~n4881 ) | ( x94 & n4880 ) | ( ~n4881 & n4880 ) ;
  assign n4883 = ~n644 & n2836 ;
  assign n4884 = n4882 | n4883 ;
  assign n4885 = ( x14 & ~n4884 ) | ( x14 & 1'b0 ) | ( ~n4884 & 1'b0 ) ;
  assign n4886 = ~x14 & n4884 ;
  assign n4887 = n4885 | n4886 ;
  assign n4888 = ( n4806 & n4807 ) | ( n4806 & n4817 ) | ( n4807 & n4817 ) ;
  assign n4892 = x91 &  n942 ;
  assign n4889 = ( x93 & ~n896 ) | ( x93 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n4890 = x92 &  n891 ;
  assign n4891 = n4889 | n4890 ;
  assign n4893 = ( x91 & ~n4892 ) | ( x91 & n4891 ) | ( ~n4892 & n4891 ) ;
  assign n4894 = n899 | n2264 ;
  assign n4895 = ~n4893 & n4894 ;
  assign n4896 = x17 &  n4895 ;
  assign n4897 = x17 | n4895 ;
  assign n4898 = ~n4896 & n4897 ;
  assign n4999 = x85 &  n1551 ;
  assign n4996 = ( x87 & ~n1451 ) | ( x87 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n4997 = x86 &  n1446 ;
  assign n4998 = n4996 | n4997 ;
  assign n5000 = ( x85 & ~n4999 ) | ( x85 & n4998 ) | ( ~n4999 & n4998 ) ;
  assign n5001 = ~n1454 & n1512 ;
  assign n5002 = n5000 | n5001 ;
  assign n5003 = ( x23 & ~n5002 ) | ( x23 & 1'b0 ) | ( ~n5002 & 1'b0 ) ;
  assign n5004 = ~x23 & n5002 ;
  assign n5005 = n5003 | n5004 ;
  assign n4902 = x79 &  n2312 ;
  assign n4899 = ( x81 & ~n2195 ) | ( x81 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n4900 = x80 &  n2190 ;
  assign n4901 = n4899 | n4900 ;
  assign n4903 = ( x79 & ~n4902 ) | ( x79 & n4901 ) | ( ~n4902 & n4901 ) ;
  assign n4904 = ( n994 & ~n2198 ) | ( n994 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n4905 = n4903 | n4904 ;
  assign n4906 = ( x29 & ~n4905 ) | ( x29 & 1'b0 ) | ( ~n4905 & 1'b0 ) ;
  assign n4907 = ~x29 & n4905 ;
  assign n4908 = n4906 | n4907 ;
  assign n4909 = ( n4777 & n4787 ) | ( n4777 & n4788 ) | ( n4787 & n4788 ) ;
  assign n4913 = x76 &  n2718 ;
  assign n4910 = ( x78 & ~n2642 ) | ( x78 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n4911 = x77 &  n2637 ;
  assign n4912 = n4910 | n4911 ;
  assign n4914 = ( x76 & ~n4913 ) | ( x76 & n4912 ) | ( ~n4913 & n4912 ) ;
  assign n4915 = ( n693 & ~n2645 ) | ( n693 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n4916 = n4914 | n4915 ;
  assign n4917 = ( x32 & ~n4916 ) | ( x32 & 1'b0 ) | ( ~n4916 & 1'b0 ) ;
  assign n4918 = ~x32 & n4916 ;
  assign n4919 = n4917 | n4918 ;
  assign n4920 = ( n4552 & n4764 ) | ( n4552 & n4774 ) | ( n4764 & n4774 ) ;
  assign n4924 = x70 &  n3756 ;
  assign n4921 = ( x72 & ~n3602 ) | ( x72 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n4922 = x71 &  n3597 ;
  assign n4923 = n4921 | n4922 ;
  assign n4925 = ( x70 & ~n4924 ) | ( x70 & n4923 ) | ( ~n4924 & n4923 ) ;
  assign n4926 = ( n345 & ~n3605 ) | ( n345 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n4927 = n4925 | n4926 ;
  assign n4929 = x38 &  n4927 ;
  assign n4928 = ~x38 & n4927 ;
  assign n4930 = ( x38 & ~n4929 ) | ( x38 & n4928 ) | ( ~n4929 & n4928 ) ;
  assign n4931 = ( n4736 & n4746 ) | ( n4736 & n4747 ) | ( n4746 & n4747 ) ;
  assign n4950 = x67 &  n4344 ;
  assign n4947 = ( x69 & ~n4143 ) | ( x69 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n4948 = x68 &  n4138 ;
  assign n4949 = n4947 | n4948 ;
  assign n4951 = ( x67 & ~n4950 ) | ( x67 & n4949 ) | ( ~n4950 & n4949 ) ;
  assign n4952 = ( n246 & ~n4146 ) | ( n246 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n4953 = n4951 | n4952 ;
  assign n4954 = ( x41 & ~n4953 ) | ( x41 & 1'b0 ) | ( ~n4953 & 1'b0 ) ;
  assign n4955 = ~x41 & n4953 ;
  assign n4956 = n4954 | n4955 ;
  assign n4933 = ( x42 & ~x43 ) | ( x42 & n4724 ) | ( ~x43 & n4724 ) ;
  assign n4932 = ( x42 & ~x43 ) | ( x42 & n4507 ) | ( ~x43 & n4507 ) ;
  assign n4934 = ~n4933 |  n4932 ;
  assign n4938 = x64 &  n4934 ;
  assign n4935 = ( x66 & ~n4725 ) | ( x66 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n4936 = x65 &  n4720 ;
  assign n4937 = n4935 | n4936 ;
  assign n4939 = ( x64 & ~n4938 ) | ( x64 & n4937 ) | ( ~n4938 & n4937 ) ;
  assign n4940 = ( n157 & ~n4728 ) | ( n157 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n4941 = n4939 | n4940 ;
  assign n4942 = ( x44 & n4508 ) | ( x44 & n4730 ) | ( n4508 & n4730 ) ;
  assign n4943 = ( x44 & ~n4942 ) | ( x44 & 1'b0 ) | ( ~n4942 & 1'b0 ) ;
  assign n4945 = ( x44 & n4941 ) | ( x44 & n4943 ) | ( n4941 & n4943 ) ;
  assign n4944 = ( n4941 & ~x44 ) | ( n4941 & n4943 ) | ( ~x44 & n4943 ) ;
  assign n4946 = ( x44 & ~n4945 ) | ( x44 & n4944 ) | ( ~n4945 & n4944 ) ;
  assign n4957 = ( n4735 & ~n4956 ) | ( n4735 & n4946 ) | ( ~n4956 & n4946 ) ;
  assign n4958 = ( n4946 & ~n4735 ) | ( n4946 & n4956 ) | ( ~n4735 & n4956 ) ;
  assign n4959 = ( n4957 & ~n4946 ) | ( n4957 & n4958 ) | ( ~n4946 & n4958 ) ;
  assign n4961 = ( n4930 & n4931 ) | ( n4930 & n4959 ) | ( n4931 & n4959 ) ;
  assign n4960 = ( n4931 & ~n4930 ) | ( n4931 & n4959 ) | ( ~n4930 & n4959 ) ;
  assign n4962 = ( n4930 & ~n4961 ) | ( n4930 & n4960 ) | ( ~n4961 & n4960 ) ;
  assign n4963 = ( n4750 & n4751 ) | ( n4750 & n4761 ) | ( n4751 & n4761 ) ;
  assign n4967 = x73 &  n3214 ;
  assign n4964 = ( x75 & ~n3087 ) | ( x75 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n4965 = x74 &  n3082 ;
  assign n4966 = n4964 | n4965 ;
  assign n4968 = ( x73 & ~n4967 ) | ( x73 & n4966 ) | ( ~n4967 & n4966 ) ;
  assign n4969 = ( n540 & ~n3090 ) | ( n540 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n4970 = n4968 | n4969 ;
  assign n4971 = ( x35 & ~n4970 ) | ( x35 & 1'b0 ) | ( ~n4970 & 1'b0 ) ;
  assign n4972 = ~x35 & n4970 ;
  assign n4973 = n4971 | n4972 ;
  assign n4974 = ( n4962 & ~n4963 ) | ( n4962 & n4973 ) | ( ~n4963 & n4973 ) ;
  assign n4975 = ( n4962 & ~n4973 ) | ( n4962 & n4963 ) | ( ~n4973 & n4963 ) ;
  assign n4976 = ( n4974 & ~n4962 ) | ( n4974 & n4975 ) | ( ~n4962 & n4975 ) ;
  assign n4978 = ( n4919 & n4920 ) | ( n4919 & n4976 ) | ( n4920 & n4976 ) ;
  assign n4977 = ( n4920 & ~n4919 ) | ( n4920 & n4976 ) | ( ~n4919 & n4976 ) ;
  assign n4979 = ( n4919 & ~n4978 ) | ( n4919 & n4977 ) | ( ~n4978 & n4977 ) ;
  assign n4981 = ( n4908 & n4909 ) | ( n4908 & n4979 ) | ( n4909 & n4979 ) ;
  assign n4980 = ( n4909 & ~n4908 ) | ( n4909 & n4979 ) | ( ~n4908 & n4979 ) ;
  assign n4982 = ( n4908 & ~n4981 ) | ( n4908 & n4980 ) | ( ~n4981 & n4980 ) ;
  assign n4986 = x82 &  n1894 ;
  assign n4983 = ( x84 & ~n1816 ) | ( x84 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n4984 = x83 &  n1811 ;
  assign n4985 = n4983 | n4984 ;
  assign n4987 = ( x82 & ~n4986 ) | ( x82 & n4985 ) | ( ~n4986 & n4985 ) ;
  assign n4988 = ( n1199 & ~n1819 ) | ( n1199 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n4989 = n4987 | n4988 ;
  assign n4990 = ( x26 & ~n4989 ) | ( x26 & 1'b0 ) | ( ~n4989 & 1'b0 ) ;
  assign n4991 = ~x26 & n4989 ;
  assign n4992 = n4990 | n4991 ;
  assign n4993 = ( n4982 & ~n4793 ) | ( n4982 & n4992 ) | ( ~n4793 & n4992 ) ;
  assign n4994 = ( n4793 & ~n4992 ) | ( n4793 & n4982 ) | ( ~n4992 & n4982 ) ;
  assign n4995 = ( n4993 & ~n4982 ) | ( n4993 & n4994 ) | ( ~n4982 & n4994 ) ;
  assign n5006 = ( n4797 & ~n5005 ) | ( n4797 & n4995 ) | ( ~n5005 & n4995 ) ;
  assign n5007 = ( n4995 & ~n4797 ) | ( n4995 & n5005 ) | ( ~n4797 & n5005 ) ;
  assign n5008 = ( n5006 & ~n4995 ) | ( n5006 & n5007 ) | ( ~n4995 & n5007 ) ;
  assign n5012 = x88 &  n1227 ;
  assign n5009 = ( x90 & ~n1154 ) | ( x90 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n5010 = x89 &  n1149 ;
  assign n5011 = n5009 | n5010 ;
  assign n5013 = ( x88 & ~n5012 ) | ( x88 & n5011 ) | ( ~n5012 & n5011 ) ;
  assign n5014 = ~n1157 & n1976 ;
  assign n5015 = n5013 | n5014 ;
  assign n5016 = ( x20 & ~n5015 ) | ( x20 & 1'b0 ) | ( ~n5015 & 1'b0 ) ;
  assign n5017 = ~x20 & n5015 ;
  assign n5018 = n5016 | n5017 ;
  assign n5019 = ( n5008 & ~n4801 ) | ( n5008 & n5018 ) | ( ~n4801 & n5018 ) ;
  assign n5020 = ( n4801 & ~n5018 ) | ( n4801 & n5008 ) | ( ~n5018 & n5008 ) ;
  assign n5021 = ( n5019 & ~n5008 ) | ( n5019 & n5020 ) | ( ~n5008 & n5020 ) ;
  assign n5022 = ( n4804 & ~n4898 ) | ( n4804 & n5021 ) | ( ~n4898 & n5021 ) ;
  assign n5023 = ( n4898 & ~n4804 ) | ( n4898 & n5021 ) | ( ~n4804 & n5021 ) ;
  assign n5024 = ( n5022 & ~n5021 ) | ( n5022 & n5023 ) | ( ~n5021 & n5023 ) ;
  assign n5025 = ( n4887 & ~n4888 ) | ( n4887 & n5024 ) | ( ~n4888 & n5024 ) ;
  assign n5026 = ( n4887 & ~n5024 ) | ( n4887 & n4888 ) | ( ~n5024 & n4888 ) ;
  assign n5027 = ( n5025 & ~n4887 ) | ( n5025 & n5026 ) | ( ~n4887 & n5026 ) ;
  assign n5031 = x97 &  n503 ;
  assign n5028 = ( x99 & ~n450 ) | ( x99 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n5029 = x98 &  n445 ;
  assign n5030 = n5028 | n5029 ;
  assign n5032 = ( x97 & ~n5031 ) | ( x97 & n5030 ) | ( ~n5031 & n5030 ) ;
  assign n5033 = ~n453 & n3338 ;
  assign n5034 = n5032 | n5033 ;
  assign n5035 = ( x11 & ~n5034 ) | ( x11 & 1'b0 ) | ( ~n5034 & 1'b0 ) ;
  assign n5036 = ~x11 & n5034 ;
  assign n5037 = n5035 | n5036 ;
  assign n5038 = ( n4635 & n4820 ) | ( n4635 & n4830 ) | ( n4820 & n4830 ) ;
  assign n5039 = ( n5027 & ~n5037 ) | ( n5027 & n5038 ) | ( ~n5037 & n5038 ) ;
  assign n5040 = ( n5027 & ~n5038 ) | ( n5027 & n5037 ) | ( ~n5038 & n5037 ) ;
  assign n5041 = ( n5039 & ~n5027 ) | ( n5039 & n5040 ) | ( ~n5027 & n5040 ) ;
  assign n4871 = x100 &  n353 ;
  assign n4868 = ( x102 & ~n313 ) | ( x102 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n4869 = x101 &  n308 ;
  assign n4870 = n4868 | n4869 ;
  assign n4872 = ( x100 & ~n4871 ) | ( x100 & n4870 ) | ( ~n4871 & n4870 ) ;
  assign n4873 = n316 | n3872 ;
  assign n4874 = ~n4872 & n4873 ;
  assign n4875 = x8 &  n4874 ;
  assign n4876 = x8 | n4874 ;
  assign n4877 = ~n4875 & n4876 ;
  assign n5042 = ( n4867 & ~n5041 ) | ( n4867 & n4877 ) | ( ~n5041 & n4877 ) ;
  assign n5043 = ( n4867 & ~n4877 ) | ( n4867 & n5041 ) | ( ~n4877 & n5041 ) ;
  assign n5044 = ( n5042 & ~n4867 ) | ( n5042 & n5043 ) | ( ~n4867 & n5043 ) ;
  assign n5045 = ( n4837 & ~n4866 ) | ( n4837 & n5044 ) | ( ~n4866 & n5044 ) ;
  assign n5046 = ( n4866 & ~n4837 ) | ( n4866 & n5044 ) | ( ~n4837 & n5044 ) ;
  assign n5047 = ( n5045 & ~n5044 ) | ( n5045 & n5046 ) | ( ~n5044 & n5046 ) ;
  assign n5051 = ~n136 & x108 ;
  assign n5048 = ( x106 & ~n150 ) | ( x106 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n5049 = ( x107 & ~n131 ) | ( x107 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n5050 = n5048 | n5049 ;
  assign n5052 = ( x108 & ~n5051 ) | ( x108 & n5050 ) | ( ~n5051 & n5050 ) ;
  assign n5053 = ( x107 & ~x108 ) | ( x107 & n4847 ) | ( ~x108 & n4847 ) ;
  assign n5054 = ( x107 & x108 ) | ( x107 & n4847 ) | ( x108 & n4847 ) ;
  assign n5055 = ( ~x108 & ~n5053 ) | ( ~x108 & n5054 ) | ( ~n5053 & n5054 ) ;
  assign n5056 = ( n5052 & ~n139 ) | ( n5052 & n5055 ) | ( ~n139 & n5055 ) ;
  assign n5057 = n139 | n5056 ;
  assign n5059 = ( x2 & n5052 ) | ( x2 & n5057 ) | ( n5052 & n5057 ) ;
  assign n5058 = ( x2 & ~n5057 ) | ( x2 & n5052 ) | ( ~n5057 & n5052 ) ;
  assign n5060 = ( n5057 & ~n5059 ) | ( n5057 & n5058 ) | ( ~n5059 & n5058 ) ;
  assign n5062 = ( n4854 & n5047 ) | ( n4854 & n5060 ) | ( n5047 & n5060 ) ;
  assign n5061 = ( n4854 & ~n5047 ) | ( n4854 & n5060 ) | ( ~n5047 & n5060 ) ;
  assign n5063 = ( n5047 & ~n5062 ) | ( n5047 & n5061 ) | ( ~n5062 & n5061 ) ;
  assign n5249 = x104 &  n225 ;
  assign n5246 = ( x106 & ~n197 ) | ( x106 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n5247 = x105 &  n192 ;
  assign n5248 = n5246 | n5247 ;
  assign n5250 = ( x104 & ~n5249 ) | ( x104 & n5248 ) | ( ~n5249 & n5248 ) ;
  assign n5251 = ~n200 & n4458 ;
  assign n5252 = n5250 | n5251 ;
  assign n5253 = ( x5 & ~n5252 ) | ( x5 & 1'b0 ) | ( ~n5252 & 1'b0 ) ;
  assign n5254 = ~x5 & n5252 ;
  assign n5255 = n5253 | n5254 ;
  assign n5242 = ( n4867 & n4877 ) | ( n4867 & n5041 ) | ( n4877 & n5041 ) ;
  assign n5150 = x80 &  n2312 ;
  assign n5147 = ( x82 & ~n2195 ) | ( x82 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n5148 = x81 &  n2190 ;
  assign n5149 = n5147 | n5148 ;
  assign n5151 = ( x80 & ~n5150 ) | ( x80 & n5149 ) | ( ~n5150 & n5149 ) ;
  assign n5152 = ( n1084 & ~n2198 ) | ( n1084 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n5153 = n5151 | n5152 ;
  assign n5154 = ( x29 & ~n5153 ) | ( x29 & 1'b0 ) | ( ~n5153 & 1'b0 ) ;
  assign n5155 = ~x29 & n5153 ;
  assign n5156 = n5154 | n5155 ;
  assign n5137 = x77 &  n2718 ;
  assign n5134 = ( x79 & ~n2642 ) | ( x79 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n5135 = x78 &  n2637 ;
  assign n5136 = n5134 | n5135 ;
  assign n5138 = ( x77 & ~n5137 ) | ( x77 & n5136 ) | ( ~n5137 & n5136 ) ;
  assign n5139 = ( n766 & ~n2645 ) | ( n766 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n5140 = n5138 | n5139 ;
  assign n5141 = ( x32 & ~n5140 ) | ( x32 & 1'b0 ) | ( ~n5140 & 1'b0 ) ;
  assign n5142 = ~x32 & n5140 ;
  assign n5143 = n5141 | n5142 ;
  assign n5077 = x74 &  n3214 ;
  assign n5074 = ( x76 & ~n3087 ) | ( x76 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n5075 = x75 &  n3082 ;
  assign n5076 = n5074 | n5075 ;
  assign n5078 = ( x74 & ~n5077 ) | ( x74 & n5076 ) | ( ~n5077 & n5076 ) ;
  assign n5079 = ( n603 & ~n3090 ) | ( n603 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n5080 = n5078 | n5079 ;
  assign n5081 = ( x35 & ~n5080 ) | ( x35 & 1'b0 ) | ( ~n5080 & 1'b0 ) ;
  assign n5082 = ~x35 & n5080 ;
  assign n5083 = n5081 | n5082 ;
  assign n5084 = ( n4962 & n4963 ) | ( n4962 & n4973 ) | ( n4963 & n4973 ) ;
  assign n5085 = ( x44 & ~x45 ) | ( x44 & 1'b0 ) | ( ~x45 & 1'b0 ) ;
  assign n5086 = ~x44 & x45 ;
  assign n5087 = n5085 | n5086 ;
  assign n5088 = x64 &  n5087 ;
  assign n5089 = ( x44 & n4941 ) | ( x44 & n4942 ) | ( n4941 & n4942 ) ;
  assign n5090 = ( x44 & ~n5089 ) | ( x44 & 1'b0 ) | ( ~n5089 & 1'b0 ) ;
  assign n5094 = x65 &  n4934 ;
  assign n5091 = ( x67 & ~n4725 ) | ( x67 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n5092 = x66 &  n4720 ;
  assign n5093 = n5091 | n5092 ;
  assign n5095 = ( x65 & ~n5094 ) | ( x65 & n5093 ) | ( ~n5094 & n5093 ) ;
  assign n5096 = n173 | n4728 ;
  assign n5097 = ~n5095 & n5096 ;
  assign n5098 = x44 &  n5097 ;
  assign n5099 = x44 | n5097 ;
  assign n5100 = ~n5098 & n5099 ;
  assign n5101 = ( n5088 & ~n5090 ) | ( n5088 & n5100 ) | ( ~n5090 & n5100 ) ;
  assign n5102 = ( n5088 & ~n5100 ) | ( n5088 & n5090 ) | ( ~n5100 & n5090 ) ;
  assign n5103 = ( n5101 & ~n5088 ) | ( n5101 & n5102 ) | ( ~n5088 & n5102 ) ;
  assign n5107 = x68 &  n4344 ;
  assign n5104 = ( x70 & ~n4143 ) | ( x70 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n5105 = x69 &  n4138 ;
  assign n5106 = n5104 | n5105 ;
  assign n5108 = ( x68 & ~n5107 ) | ( x68 & n5106 ) | ( ~n5107 & n5106 ) ;
  assign n5109 = ( n282 & ~n4146 ) | ( n282 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n5110 = n5108 | n5109 ;
  assign n5111 = ( x41 & ~n5110 ) | ( x41 & 1'b0 ) | ( ~n5110 & 1'b0 ) ;
  assign n5112 = ~x41 & n5110 ;
  assign n5113 = n5111 | n5112 ;
  assign n5114 = ( n4735 & n4946 ) | ( n4735 & n4956 ) | ( n4946 & n4956 ) ;
  assign n5115 = ( n5103 & ~n5113 ) | ( n5103 & n5114 ) | ( ~n5113 & n5114 ) ;
  assign n5116 = ( n5103 & ~n5114 ) | ( n5103 & n5113 ) | ( ~n5114 & n5113 ) ;
  assign n5117 = ( n5115 & ~n5103 ) | ( n5115 & n5116 ) | ( ~n5103 & n5116 ) ;
  assign n5121 = x71 &  n3756 ;
  assign n5118 = ( x73 & ~n3602 ) | ( x73 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n5119 = x72 &  n3597 ;
  assign n5120 = n5118 | n5119 ;
  assign n5122 = ( x71 & ~n5121 ) | ( x71 & n5120 ) | ( ~n5121 & n5120 ) ;
  assign n5123 = ( n389 & ~n3605 ) | ( n389 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n5124 = n5122 | n5123 ;
  assign n5125 = ( x38 & ~n5124 ) | ( x38 & 1'b0 ) | ( ~n5124 & 1'b0 ) ;
  assign n5126 = ~x38 & n5124 ;
  assign n5127 = n5125 | n5126 ;
  assign n5128 = ( n5117 & ~n4961 ) | ( n5117 & n5127 ) | ( ~n4961 & n5127 ) ;
  assign n5129 = ( n4961 & ~n5127 ) | ( n4961 & n5117 ) | ( ~n5127 & n5117 ) ;
  assign n5130 = ( n5128 & ~n5117 ) | ( n5128 & n5129 ) | ( ~n5117 & n5129 ) ;
  assign n5131 = ( n5083 & ~n5084 ) | ( n5083 & n5130 ) | ( ~n5084 & n5130 ) ;
  assign n5132 = ( n5083 & ~n5130 ) | ( n5083 & n5084 ) | ( ~n5130 & n5084 ) ;
  assign n5133 = ( n5131 & ~n5083 ) | ( n5131 & n5132 ) | ( ~n5083 & n5132 ) ;
  assign n5144 = ( n4978 & ~n5143 ) | ( n4978 & n5133 ) | ( ~n5143 & n5133 ) ;
  assign n5145 = ( n5133 & ~n4978 ) | ( n5133 & n5143 ) | ( ~n4978 & n5143 ) ;
  assign n5146 = ( n5144 & ~n5133 ) | ( n5144 & n5145 ) | ( ~n5133 & n5145 ) ;
  assign n5157 = ( n4981 & ~n5156 ) | ( n4981 & n5146 ) | ( ~n5156 & n5146 ) ;
  assign n5158 = ( n5146 & ~n4981 ) | ( n5146 & n5156 ) | ( ~n4981 & n5156 ) ;
  assign n5159 = ( n5157 & ~n5146 ) | ( n5157 & n5158 ) | ( ~n5146 & n5158 ) ;
  assign n5163 = x83 &  n1894 ;
  assign n5160 = ( x85 & ~n1816 ) | ( x85 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n5161 = x84 &  n1811 ;
  assign n5162 = n5160 | n5161 ;
  assign n5164 = ( x83 & ~n5163 ) | ( x83 & n5162 ) | ( ~n5163 & n5162 ) ;
  assign n5165 = ( n1295 & ~n1819 ) | ( n1295 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n5166 = n5164 | n5165 ;
  assign n5167 = ( x26 & ~n5166 ) | ( x26 & 1'b0 ) | ( ~n5166 & 1'b0 ) ;
  assign n5168 = ~x26 & n5166 ;
  assign n5169 = n5167 | n5168 ;
  assign n5170 = ( n4793 & n4982 ) | ( n4793 & n4992 ) | ( n4982 & n4992 ) ;
  assign n5171 = ( n5159 & ~n5169 ) | ( n5159 & n5170 ) | ( ~n5169 & n5170 ) ;
  assign n5172 = ( n5159 & ~n5170 ) | ( n5159 & n5169 ) | ( ~n5170 & n5169 ) ;
  assign n5173 = ( n5171 & ~n5159 ) | ( n5171 & n5172 ) | ( ~n5159 & n5172 ) ;
  assign n5174 = ( n4797 & n4995 ) | ( n4797 & n5005 ) | ( n4995 & n5005 ) ;
  assign n5178 = x86 &  n1551 ;
  assign n5175 = ( x88 & ~n1451 ) | ( x88 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n5176 = x87 &  n1446 ;
  assign n5177 = n5175 | n5176 ;
  assign n5179 = ( x86 & ~n5178 ) | ( x86 & n5177 ) | ( ~n5178 & n5177 ) ;
  assign n5180 = ~n1454 & n1624 ;
  assign n5181 = n5179 | n5180 ;
  assign n5182 = ( x23 & ~n5181 ) | ( x23 & 1'b0 ) | ( ~n5181 & 1'b0 ) ;
  assign n5183 = ~x23 & n5181 ;
  assign n5184 = n5182 | n5183 ;
  assign n5185 = ( n5173 & ~n5174 ) | ( n5173 & n5184 ) | ( ~n5174 & n5184 ) ;
  assign n5186 = ( n5173 & ~n5184 ) | ( n5173 & n5174 ) | ( ~n5184 & n5174 ) ;
  assign n5187 = ( n5185 & ~n5173 ) | ( n5185 & n5186 ) | ( ~n5173 & n5186 ) ;
  assign n5188 = ( n4801 & n5008 ) | ( n4801 & n5018 ) | ( n5008 & n5018 ) ;
  assign n5192 = x89 &  n1227 ;
  assign n5189 = ( x91 & ~n1154 ) | ( x91 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n5190 = x90 &  n1149 ;
  assign n5191 = n5189 | n5190 ;
  assign n5193 = ( x89 & ~n5192 ) | ( x89 & n5191 ) | ( ~n5192 & n5191 ) ;
  assign n5194 = ~n1157 & n2108 ;
  assign n5195 = n5193 | n5194 ;
  assign n5196 = ( x20 & ~n5195 ) | ( x20 & 1'b0 ) | ( ~n5195 & 1'b0 ) ;
  assign n5197 = ~x20 & n5195 ;
  assign n5198 = n5196 | n5197 ;
  assign n5199 = ( n5187 & ~n5188 ) | ( n5187 & n5198 ) | ( ~n5188 & n5198 ) ;
  assign n5200 = ( n5188 & ~n5187 ) | ( n5188 & n5198 ) | ( ~n5187 & n5198 ) ;
  assign n5201 = ( n5199 & ~n5198 ) | ( n5199 & n5200 ) | ( ~n5198 & n5200 ) ;
  assign n5067 = x92 &  n942 ;
  assign n5064 = ( x94 & ~n896 ) | ( x94 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n5065 = x93 &  n891 ;
  assign n5066 = n5064 | n5065 ;
  assign n5068 = ( x92 & ~n5067 ) | ( x92 & n5066 ) | ( ~n5067 & n5066 ) ;
  assign n5069 = ~n899 & n2401 ;
  assign n5070 = n5068 | n5069 ;
  assign n5071 = ( x17 & ~n5070 ) | ( x17 & 1'b0 ) | ( ~n5070 & 1'b0 ) ;
  assign n5072 = ~x17 & n5070 ;
  assign n5073 = n5071 | n5072 ;
  assign n5202 = ( n5022 & ~n5201 ) | ( n5022 & n5073 ) | ( ~n5201 & n5073 ) ;
  assign n5203 = ( n5022 & ~n5073 ) | ( n5022 & n5201 ) | ( ~n5073 & n5201 ) ;
  assign n5204 = ( n5202 & ~n5022 ) | ( n5202 & n5203 ) | ( ~n5022 & n5203 ) ;
  assign n5208 = x95 &  n713 ;
  assign n5205 = ( x97 & ~n641 ) | ( x97 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n5206 = x96 &  n636 ;
  assign n5207 = n5205 | n5206 ;
  assign n5209 = ( x95 & ~n5208 ) | ( x95 & n5207 ) | ( ~n5208 & n5207 ) ;
  assign n5210 = ~n644 & n2999 ;
  assign n5211 = n5209 | n5210 ;
  assign n5212 = ( x14 & ~n5211 ) | ( x14 & 1'b0 ) | ( ~n5211 & 1'b0 ) ;
  assign n5213 = ~x14 & n5211 ;
  assign n5214 = n5212 | n5213 ;
  assign n5215 = ( n5204 & ~n5026 ) | ( n5204 & n5214 ) | ( ~n5026 & n5214 ) ;
  assign n5216 = ( n5026 & ~n5204 ) | ( n5026 & n5214 ) | ( ~n5204 & n5214 ) ;
  assign n5217 = ( n5215 & ~n5214 ) | ( n5215 & n5216 ) | ( ~n5214 & n5216 ) ;
  assign n5218 = ( n5037 & ~n5027 ) | ( n5037 & n5038 ) | ( ~n5027 & n5038 ) ;
  assign n5222 = x98 &  n503 ;
  assign n5219 = ( x100 & ~n450 ) | ( x100 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n5220 = x99 &  n445 ;
  assign n5221 = n5219 | n5220 ;
  assign n5223 = ( x98 & ~n5222 ) | ( x98 & n5221 ) | ( ~n5222 & n5221 ) ;
  assign n5224 = n453 | n3354 ;
  assign n5225 = ~n5223 & n5224 ;
  assign n5226 = x11 &  n5225 ;
  assign n5227 = x11 | n5225 ;
  assign n5228 = ~n5226 & n5227 ;
  assign n5229 = ( n5217 & n5218 ) | ( n5217 & n5228 ) | ( n5218 & n5228 ) ;
  assign n5230 = ( n5218 & ~n5217 ) | ( n5218 & n5228 ) | ( ~n5217 & n5228 ) ;
  assign n5231 = ( n5217 & ~n5229 ) | ( n5217 & n5230 ) | ( ~n5229 & n5230 ) ;
  assign n5235 = x101 &  n353 ;
  assign n5232 = ( x103 & ~n313 ) | ( x103 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n5233 = x102 &  n308 ;
  assign n5234 = n5232 | n5233 ;
  assign n5236 = ( x101 & ~n5235 ) | ( x101 & n5234 ) | ( ~n5235 & n5234 ) ;
  assign n5237 = n316 | n4056 ;
  assign n5238 = ~n5236 & n5237 ;
  assign n5239 = x8 &  n5238 ;
  assign n5240 = x8 | n5238 ;
  assign n5241 = ~n5239 & n5240 ;
  assign n5243 = ( n5231 & n5241 ) | ( n5231 & n5242 ) | ( n5241 & n5242 ) ;
  assign n5244 = ( n5231 & ~n5242 ) | ( n5231 & n5241 ) | ( ~n5242 & n5241 ) ;
  assign n5245 = ( n5242 & ~n5243 ) | ( n5242 & n5244 ) | ( ~n5243 & n5244 ) ;
  assign n5256 = ( n5045 & ~n5255 ) | ( n5045 & n5245 ) | ( ~n5255 & n5245 ) ;
  assign n5257 = ( n5045 & ~n5245 ) | ( n5045 & n5255 ) | ( ~n5245 & n5255 ) ;
  assign n5258 = ( n5256 & ~n5045 ) | ( n5256 & n5257 ) | ( ~n5045 & n5257 ) ;
  assign n5259 = ( n4854 & ~n5060 ) | ( n4854 & n5047 ) | ( ~n5060 & n5047 ) ;
  assign n5263 = ~n136 & x109 ;
  assign n5260 = ( x107 & ~n150 ) | ( x107 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n5261 = ( x108 & ~n131 ) | ( x108 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n5262 = n5260 | n5261 ;
  assign n5264 = ( x109 & ~n5263 ) | ( x109 & n5262 ) | ( ~n5263 & n5262 ) ;
  assign n5266 = ( x108 & x109 ) | ( x108 & n5054 ) | ( x109 & n5054 ) ;
  assign n5265 = ( x108 & ~x109 ) | ( x108 & n5054 ) | ( ~x109 & n5054 ) ;
  assign n5267 = ( x109 & ~n5266 ) | ( x109 & n5265 ) | ( ~n5266 & n5265 ) ;
  assign n5268 = ( n139 & ~n5264 ) | ( n139 & n5267 ) | ( ~n5264 & n5267 ) ;
  assign n5269 = ~n139 & n5268 ;
  assign n5270 = ( x2 & n5264 ) | ( x2 & n5269 ) | ( n5264 & n5269 ) ;
  assign n5271 = ( x2 & ~n5269 ) | ( x2 & n5264 ) | ( ~n5269 & n5264 ) ;
  assign n5272 = ( n5269 & ~n5270 ) | ( n5269 & n5271 ) | ( ~n5270 & n5271 ) ;
  assign n5273 = ( n5258 & ~n5259 ) | ( n5258 & n5272 ) | ( ~n5259 & n5272 ) ;
  assign n5274 = ( n5258 & ~n5272 ) | ( n5258 & n5259 ) | ( ~n5272 & n5259 ) ;
  assign n5275 = ( n5273 & ~n5258 ) | ( n5273 & n5274 ) | ( ~n5258 & n5274 ) ;
  assign n5279 = ~n136 & x110 ;
  assign n5276 = ( x108 & ~n150 ) | ( x108 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n5277 = ( x109 & ~n131 ) | ( x109 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n5278 = n5276 | n5277 ;
  assign n5280 = ( x110 & ~n5279 ) | ( x110 & n5278 ) | ( ~n5279 & n5278 ) ;
  assign n5281 = ( x109 & ~x110 ) | ( x109 & n5266 ) | ( ~x110 & n5266 ) ;
  assign n5282 = ( x109 & x110 ) | ( x109 & n5266 ) | ( x110 & n5266 ) ;
  assign n5283 = ( ~x110 & ~n5281 ) | ( ~x110 & n5282 ) | ( ~n5281 & n5282 ) ;
  assign n5284 = ( n5280 & ~n139 ) | ( n5280 & n5283 ) | ( ~n139 & n5283 ) ;
  assign n5285 = n139 | n5284 ;
  assign n5287 = ( x2 & n5280 ) | ( x2 & n5285 ) | ( n5280 & n5285 ) ;
  assign n5286 = ( x2 & ~n5285 ) | ( x2 & n5280 ) | ( ~n5285 & n5280 ) ;
  assign n5288 = ( n5285 & ~n5287 ) | ( n5285 & n5286 ) | ( ~n5287 & n5286 ) ;
  assign n5289 = ( n5245 & ~n5045 ) | ( n5245 & n5255 ) | ( ~n5045 & n5255 ) ;
  assign n5293 = x105 &  n225 ;
  assign n5290 = ( x107 & ~n197 ) | ( x107 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n5291 = x106 &  n192 ;
  assign n5292 = n5290 | n5291 ;
  assign n5294 = ( x105 & ~n5293 ) | ( x105 & n5292 ) | ( ~n5293 & n5292 ) ;
  assign n5295 = ~n200 & n4848 ;
  assign n5296 = n5294 | n5295 ;
  assign n5297 = ( x5 & ~n5296 ) | ( x5 & 1'b0 ) | ( ~n5296 & 1'b0 ) ;
  assign n5298 = ~x5 & n5296 ;
  assign n5299 = n5297 | n5298 ;
  assign n5300 = ( n5241 & ~n5231 ) | ( n5241 & n5242 ) | ( ~n5231 & n5242 ) ;
  assign n5304 = x102 &  n353 ;
  assign n5301 = ( x104 & ~n313 ) | ( x104 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n5302 = x103 &  n308 ;
  assign n5303 = n5301 | n5302 ;
  assign n5305 = ( x102 & ~n5304 ) | ( x102 & n5303 ) | ( ~n5304 & n5303 ) ;
  assign n5306 = n316 | n4249 ;
  assign n5307 = ~n5305 & n5306 ;
  assign n5308 = x8 &  n5307 ;
  assign n5309 = x8 | n5307 ;
  assign n5310 = ~n5308 & n5309 ;
  assign n5314 = x99 &  n503 ;
  assign n5311 = ( x101 & ~n450 ) | ( x101 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n5312 = x100 &  n445 ;
  assign n5313 = n5311 | n5312 ;
  assign n5315 = ( x99 & ~n5314 ) | ( x99 & n5313 ) | ( ~n5314 & n5313 ) ;
  assign n5316 = n453 | n3694 ;
  assign n5317 = ~n5315 & n5316 ;
  assign n5318 = x11 &  n5317 ;
  assign n5319 = x11 | n5317 ;
  assign n5320 = ~n5318 & n5319 ;
  assign n5324 = x93 &  n942 ;
  assign n5321 = ( x95 & ~n896 ) | ( x95 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n5322 = x94 &  n891 ;
  assign n5323 = n5321 | n5322 ;
  assign n5325 = ( x93 & ~n5324 ) | ( x93 & n5323 ) | ( ~n5324 & n5323 ) ;
  assign n5326 = ~n899 & n2547 ;
  assign n5327 = n5325 | n5326 ;
  assign n5328 = ( x17 & ~n5327 ) | ( x17 & 1'b0 ) | ( ~n5327 & 1'b0 ) ;
  assign n5329 = ~x17 & n5327 ;
  assign n5330 = n5328 | n5329 ;
  assign n5334 = x90 &  n1227 ;
  assign n5331 = ( x92 & ~n1154 ) | ( x92 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n5332 = x91 &  n1149 ;
  assign n5333 = n5331 | n5332 ;
  assign n5335 = ( x90 & ~n5334 ) | ( x90 & n5333 ) | ( ~n5334 & n5333 ) ;
  assign n5336 = ~n1157 & n2248 ;
  assign n5337 = n5335 | n5336 ;
  assign n5338 = ( x20 & ~n5337 ) | ( x20 & 1'b0 ) | ( ~n5337 & 1'b0 ) ;
  assign n5339 = ~x20 & n5337 ;
  assign n5340 = n5338 | n5339 ;
  assign n5344 = x87 &  n1551 ;
  assign n5341 = ( x89 & ~n1451 ) | ( x89 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n5342 = x88 &  n1446 ;
  assign n5343 = n5341 | n5342 ;
  assign n5345 = ( x87 & ~n5344 ) | ( x87 & n5343 ) | ( ~n5344 & n5343 ) ;
  assign n5346 = ~n1454 & n1741 ;
  assign n5347 = n5345 | n5346 ;
  assign n5348 = ( x23 & ~n5347 ) | ( x23 & 1'b0 ) | ( ~n5347 & 1'b0 ) ;
  assign n5349 = ~x23 & n5347 ;
  assign n5350 = n5348 | n5349 ;
  assign n5354 = x84 &  n1894 ;
  assign n5351 = ( x86 & ~n1816 ) | ( x86 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n5352 = x85 &  n1811 ;
  assign n5353 = n5351 | n5352 ;
  assign n5355 = ( x84 & ~n5354 ) | ( x84 & n5353 ) | ( ~n5354 & n5353 ) ;
  assign n5356 = ( n1496 & ~n1819 ) | ( n1496 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n5357 = n5355 | n5356 ;
  assign n5358 = ( x26 & ~n5357 ) | ( x26 & 1'b0 ) | ( ~n5357 & 1'b0 ) ;
  assign n5359 = ~x26 & n5357 ;
  assign n5360 = n5358 | n5359 ;
  assign n5364 = x81 &  n2312 ;
  assign n5361 = ( x83 & ~n2195 ) | ( x83 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n5362 = x82 &  n2190 ;
  assign n5363 = n5361 | n5362 ;
  assign n5365 = ( x81 & ~n5364 ) | ( x81 & n5363 ) | ( ~n5364 & n5363 ) ;
  assign n5366 = ( n1100 & ~n2198 ) | ( n1100 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n5367 = n5365 | n5366 ;
  assign n5368 = ( x29 & ~n5367 ) | ( x29 & 1'b0 ) | ( ~n5367 & 1'b0 ) ;
  assign n5369 = ~x29 & n5367 ;
  assign n5370 = n5368 | n5369 ;
  assign n5374 = x66 &  n4934 ;
  assign n5371 = ( x68 & ~n4725 ) | ( x68 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n5372 = x67 &  n4720 ;
  assign n5373 = n5371 | n5372 ;
  assign n5375 = ( x66 & ~n5374 ) | ( x66 & n5373 ) | ( ~n5374 & n5373 ) ;
  assign n5376 = ( n213 & ~n4728 ) | ( n213 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n5377 = n5375 | n5376 ;
  assign n5378 = ( x44 & ~n5377 ) | ( x44 & 1'b0 ) | ( ~n5377 & 1'b0 ) ;
  assign n5379 = ~x44 & n5377 ;
  assign n5380 = n5378 | n5379 ;
  assign n5381 = ( x47 & ~n5088 ) | ( x47 & 1'b0 ) | ( ~n5088 & 1'b0 ) ;
  assign n5382 = ( x45 & x46 ) | ( x45 & n5085 ) | ( x46 & n5085 ) ;
  assign n5383 = ( x45 & ~n5086 ) | ( x45 & x46 ) | ( ~n5086 & x46 ) ;
  assign n5384 = ~n5382 &  n5383 ;
  assign n5385 = x64 &  n5384 ;
  assign n5386 = ~x46 & x47 ;
  assign n5387 = ( x46 & ~x47 ) | ( x46 & 1'b0 ) | ( ~x47 & 1'b0 ) ;
  assign n5388 = n5386 | n5387 ;
  assign n5389 = ~n5087 |  n5388 ;
  assign n5390 = ( x65 & ~n5389 ) | ( x65 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n5391 = n5385 | n5390 ;
  assign n5392 = ~n5087 | ~n5388 ;
  assign n5393 = ( n142 & ~n5392 ) | ( n142 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n5394 = n5391 | n5393 ;
  assign n5396 = ( x47 & n5381 ) | ( x47 & n5394 ) | ( n5381 & n5394 ) ;
  assign n5395 = ( x47 & ~n5381 ) | ( x47 & n5394 ) | ( ~n5381 & n5394 ) ;
  assign n5397 = ( n5381 & ~n5396 ) | ( n5381 & n5395 ) | ( ~n5396 & n5395 ) ;
  assign n5399 = ( n5102 & n5380 ) | ( n5102 & n5397 ) | ( n5380 & n5397 ) ;
  assign n5398 = ( n5102 & ~n5380 ) | ( n5102 & n5397 ) | ( ~n5380 & n5397 ) ;
  assign n5400 = ( n5380 & ~n5399 ) | ( n5380 & n5398 ) | ( ~n5399 & n5398 ) ;
  assign n5411 = ( n5113 & ~n5103 ) | ( n5113 & n5114 ) | ( ~n5103 & n5114 ) ;
  assign n5404 = x69 &  n4344 ;
  assign n5401 = ( x71 & ~n4143 ) | ( x71 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n5402 = x70 &  n4138 ;
  assign n5403 = n5401 | n5402 ;
  assign n5405 = ( x69 & ~n5404 ) | ( x69 & n5403 ) | ( ~n5404 & n5403 ) ;
  assign n5406 = ( n298 & ~n4146 ) | ( n298 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n5407 = n5405 | n5406 ;
  assign n5408 = ( x41 & ~n5407 ) | ( x41 & 1'b0 ) | ( ~n5407 & 1'b0 ) ;
  assign n5409 = ~x41 & n5407 ;
  assign n5410 = n5408 | n5409 ;
  assign n5412 = ( n5400 & ~n5411 ) | ( n5400 & n5410 ) | ( ~n5411 & n5410 ) ;
  assign n5413 = ( n5400 & ~n5410 ) | ( n5400 & n5411 ) | ( ~n5410 & n5411 ) ;
  assign n5414 = ( n5412 & ~n5400 ) | ( n5412 & n5413 ) | ( ~n5400 & n5413 ) ;
  assign n5419 = x72 &  n3756 ;
  assign n5416 = ( x74 & ~n3602 ) | ( x74 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n5417 = x73 &  n3597 ;
  assign n5418 = n5416 | n5417 ;
  assign n5420 = ( x72 & ~n5419 ) | ( x72 & n5418 ) | ( ~n5419 & n5418 ) ;
  assign n5421 = ( n482 & ~n3605 ) | ( n482 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n5422 = n5420 | n5421 ;
  assign n5423 = ( x38 & ~n5422 ) | ( x38 & 1'b0 ) | ( ~n5422 & 1'b0 ) ;
  assign n5424 = ~x38 & n5422 ;
  assign n5425 = n5423 | n5424 ;
  assign n5415 = ( n4961 & ~n5117 ) | ( n4961 & n5127 ) | ( ~n5117 & n5127 ) ;
  assign n5426 = ( n5414 & ~n5425 ) | ( n5414 & n5415 ) | ( ~n5425 & n5415 ) ;
  assign n5427 = ( n5414 & ~n5415 ) | ( n5414 & n5425 ) | ( ~n5415 & n5425 ) ;
  assign n5428 = ( n5426 & ~n5414 ) | ( n5426 & n5427 ) | ( ~n5414 & n5427 ) ;
  assign n5432 = x75 &  n3214 ;
  assign n5429 = ( x77 & ~n3087 ) | ( x77 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n5430 = x76 &  n3082 ;
  assign n5431 = n5429 | n5430 ;
  assign n5433 = ( x75 & ~n5432 ) | ( x75 & n5431 ) | ( ~n5432 & n5431 ) ;
  assign n5434 = ( n677 & ~n3090 ) | ( n677 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n5435 = n5433 | n5434 ;
  assign n5436 = ( x35 & ~n5435 ) | ( x35 & 1'b0 ) | ( ~n5435 & 1'b0 ) ;
  assign n5437 = ~x35 & n5435 ;
  assign n5438 = n5436 | n5437 ;
  assign n5439 = ( n5428 & ~n5132 ) | ( n5428 & n5438 ) | ( ~n5132 & n5438 ) ;
  assign n5440 = ( n5132 & ~n5438 ) | ( n5132 & n5428 ) | ( ~n5438 & n5428 ) ;
  assign n5441 = ( n5439 & ~n5428 ) | ( n5439 & n5440 ) | ( ~n5428 & n5440 ) ;
  assign n5452 = ( n4978 & ~n5133 ) | ( n4978 & n5143 ) | ( ~n5133 & n5143 ) ;
  assign n5445 = x78 &  n2718 ;
  assign n5442 = ( x80 & ~n2642 ) | ( x80 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n5443 = x79 &  n2637 ;
  assign n5444 = n5442 | n5443 ;
  assign n5446 = ( x78 & ~n5445 ) | ( x78 & n5444 ) | ( ~n5445 & n5444 ) ;
  assign n5447 = ( n842 & ~n2645 ) | ( n842 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n5448 = n5446 | n5447 ;
  assign n5449 = ( x32 & ~n5448 ) | ( x32 & 1'b0 ) | ( ~n5448 & 1'b0 ) ;
  assign n5450 = ~x32 & n5448 ;
  assign n5451 = n5449 | n5450 ;
  assign n5453 = ( n5441 & ~n5452 ) | ( n5441 & n5451 ) | ( ~n5452 & n5451 ) ;
  assign n5454 = ( n5441 & ~n5451 ) | ( n5441 & n5452 ) | ( ~n5451 & n5452 ) ;
  assign n5455 = ( n5453 & ~n5441 ) | ( n5453 & n5454 ) | ( ~n5441 & n5454 ) ;
  assign n5456 = ( n4981 & ~n5146 ) | ( n4981 & n5156 ) | ( ~n5146 & n5156 ) ;
  assign n5457 = ( n5370 & n5455 ) | ( n5370 & n5456 ) | ( n5455 & n5456 ) ;
  assign n5458 = ( n5455 & ~n5370 ) | ( n5455 & n5456 ) | ( ~n5370 & n5456 ) ;
  assign n5459 = ( n5370 & ~n5457 ) | ( n5370 & n5458 ) | ( ~n5457 & n5458 ) ;
  assign n5460 = ( n5169 & ~n5159 ) | ( n5169 & n5170 ) | ( ~n5159 & n5170 ) ;
  assign n5461 = ( n5360 & n5459 ) | ( n5360 & n5460 ) | ( n5459 & n5460 ) ;
  assign n5462 = ( n5459 & ~n5360 ) | ( n5459 & n5460 ) | ( ~n5360 & n5460 ) ;
  assign n5463 = ( n5360 & ~n5461 ) | ( n5360 & n5462 ) | ( ~n5461 & n5462 ) ;
  assign n5464 = ( n5174 & ~n5173 ) | ( n5174 & n5184 ) | ( ~n5173 & n5184 ) ;
  assign n5465 = ( n5350 & n5463 ) | ( n5350 & n5464 ) | ( n5463 & n5464 ) ;
  assign n5466 = ( n5463 & ~n5350 ) | ( n5463 & n5464 ) | ( ~n5350 & n5464 ) ;
  assign n5467 = ( n5350 & ~n5465 ) | ( n5350 & n5466 ) | ( ~n5465 & n5466 ) ;
  assign n5469 = ( n5200 & n5340 ) | ( n5200 & n5467 ) | ( n5340 & n5467 ) ;
  assign n5468 = ( n5200 & ~n5340 ) | ( n5200 & n5467 ) | ( ~n5340 & n5467 ) ;
  assign n5470 = ( n5340 & ~n5469 ) | ( n5340 & n5468 ) | ( ~n5469 & n5468 ) ;
  assign n5471 = ( n5202 & n5330 ) | ( n5202 & n5470 ) | ( n5330 & n5470 ) ;
  assign n5472 = ( n5330 & ~n5202 ) | ( n5330 & n5470 ) | ( ~n5202 & n5470 ) ;
  assign n5473 = ( n5202 & ~n5471 ) | ( n5202 & n5472 ) | ( ~n5471 & n5472 ) ;
  assign n5477 = x96 &  n713 ;
  assign n5474 = ( x98 & ~n641 ) | ( x98 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n5475 = x97 &  n636 ;
  assign n5476 = n5474 | n5475 ;
  assign n5478 = ( x96 & ~n5477 ) | ( x96 & n5476 ) | ( ~n5477 & n5476 ) ;
  assign n5479 = ~n644 & n3170 ;
  assign n5480 = n5478 | n5479 ;
  assign n5481 = ( x14 & ~n5480 ) | ( x14 & 1'b0 ) | ( ~n5480 & 1'b0 ) ;
  assign n5482 = ~x14 & n5480 ;
  assign n5483 = n5481 | n5482 ;
  assign n5484 = ( n5473 & ~n5216 ) | ( n5473 & n5483 ) | ( ~n5216 & n5483 ) ;
  assign n5485 = ( n5216 & ~n5483 ) | ( n5216 & n5473 ) | ( ~n5483 & n5473 ) ;
  assign n5486 = ( n5484 & ~n5473 ) | ( n5484 & n5485 ) | ( ~n5473 & n5485 ) ;
  assign n5487 = ( n5217 & ~n5218 ) | ( n5217 & n5228 ) | ( ~n5218 & n5228 ) ;
  assign n5488 = ( n5320 & ~n5486 ) | ( n5320 & n5487 ) | ( ~n5486 & n5487 ) ;
  assign n5489 = ( n5320 & ~n5487 ) | ( n5320 & n5486 ) | ( ~n5487 & n5486 ) ;
  assign n5490 = ( n5488 & ~n5320 ) | ( n5488 & n5489 ) | ( ~n5320 & n5489 ) ;
  assign n5491 = ( n5300 & n5310 ) | ( n5300 & n5490 ) | ( n5310 & n5490 ) ;
  assign n5492 = ( n5310 & ~n5300 ) | ( n5310 & n5490 ) | ( ~n5300 & n5490 ) ;
  assign n5493 = ( n5300 & ~n5491 ) | ( n5300 & n5492 ) | ( ~n5491 & n5492 ) ;
  assign n5494 = ( n5289 & n5299 ) | ( n5289 & n5493 ) | ( n5299 & n5493 ) ;
  assign n5495 = ( n5299 & ~n5289 ) | ( n5299 & n5493 ) | ( ~n5289 & n5493 ) ;
  assign n5496 = ( n5289 & ~n5494 ) | ( n5289 & n5495 ) | ( ~n5494 & n5495 ) ;
  assign n5497 = ( n5259 & ~n5258 ) | ( n5259 & n5272 ) | ( ~n5258 & n5272 ) ;
  assign n5499 = ( n5288 & n5496 ) | ( n5288 & n5497 ) | ( n5496 & n5497 ) ;
  assign n5498 = ( n5496 & ~n5288 ) | ( n5496 & n5497 ) | ( ~n5288 & n5497 ) ;
  assign n5500 = ( n5288 & ~n5499 ) | ( n5288 & n5498 ) | ( ~n5499 & n5498 ) ;
  assign n5504 = x106 &  n225 ;
  assign n5501 = ( x108 & ~n197 ) | ( x108 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n5502 = x107 &  n192 ;
  assign n5503 = n5501 | n5502 ;
  assign n5505 = ( x106 & ~n5504 ) | ( x106 & n5503 ) | ( ~n5504 & n5503 ) ;
  assign n5506 = n200 | n5055 ;
  assign n5507 = ~n5505 & n5506 ;
  assign n5508 = x5 &  n5507 ;
  assign n5509 = x5 | n5507 ;
  assign n5510 = ~n5508 & n5509 ;
  assign n5511 = ( n5300 & ~n5490 ) | ( n5300 & n5310 ) | ( ~n5490 & n5310 ) ;
  assign n5515 = x103 &  n353 ;
  assign n5512 = ( x105 & ~n313 ) | ( x105 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n5513 = x104 &  n308 ;
  assign n5514 = n5512 | n5513 ;
  assign n5516 = ( x103 & ~n5515 ) | ( x103 & n5514 ) | ( ~n5515 & n5514 ) ;
  assign n5517 = ~n316 & n4442 ;
  assign n5518 = n5516 | n5517 ;
  assign n5519 = ( x8 & ~n5518 ) | ( x8 & 1'b0 ) | ( ~n5518 & 1'b0 ) ;
  assign n5520 = ~x8 & n5518 ;
  assign n5521 = n5519 | n5520 ;
  assign n5525 = x100 &  n503 ;
  assign n5522 = ( x102 & ~n450 ) | ( x102 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n5523 = x101 &  n445 ;
  assign n5524 = n5522 | n5523 ;
  assign n5526 = ( x100 & ~n5525 ) | ( x100 & n5524 ) | ( ~n5525 & n5524 ) ;
  assign n5527 = n453 | n3872 ;
  assign n5528 = ~n5526 & n5527 ;
  assign n5529 = x11 &  n5528 ;
  assign n5530 = x11 | n5528 ;
  assign n5531 = ~n5529 & n5530 ;
  assign n5545 = x91 &  n1227 ;
  assign n5542 = ( x93 & ~n1154 ) | ( x93 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n5543 = x92 &  n1149 ;
  assign n5544 = n5542 | n5543 ;
  assign n5546 = ( x91 & ~n5545 ) | ( x91 & n5544 ) | ( ~n5545 & n5544 ) ;
  assign n5547 = n1157 | n2264 ;
  assign n5548 = ~n5546 & n5547 ;
  assign n5549 = x20 &  n5548 ;
  assign n5550 = x20 | n5548 ;
  assign n5551 = ~n5549 & n5550 ;
  assign n5652 = x85 &  n1894 ;
  assign n5649 = ( x87 & ~n1816 ) | ( x87 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n5650 = x86 &  n1811 ;
  assign n5651 = n5649 | n5650 ;
  assign n5653 = ( x85 & ~n5652 ) | ( x85 & n5651 ) | ( ~n5652 & n5651 ) ;
  assign n5654 = ( n1512 & ~n1819 ) | ( n1512 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n5655 = n5653 | n5654 ;
  assign n5656 = ( x26 & ~n5655 ) | ( x26 & 1'b0 ) | ( ~n5655 & 1'b0 ) ;
  assign n5657 = ~x26 & n5655 ;
  assign n5658 = n5656 | n5657 ;
  assign n5565 = x79 &  n2718 ;
  assign n5562 = ( x81 & ~n2642 ) | ( x81 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n5563 = x80 &  n2637 ;
  assign n5564 = n5562 | n5563 ;
  assign n5566 = ( x79 & ~n5565 ) | ( x79 & n5564 ) | ( ~n5565 & n5564 ) ;
  assign n5567 = ( n994 & ~n2645 ) | ( n994 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n5568 = n5566 | n5567 ;
  assign n5569 = ( x32 & ~n5568 ) | ( x32 & 1'b0 ) | ( ~n5568 & 1'b0 ) ;
  assign n5570 = ~x32 & n5568 ;
  assign n5571 = n5569 | n5570 ;
  assign n5572 = ( n5441 & n5451 ) | ( n5441 & n5452 ) | ( n5451 & n5452 ) ;
  assign n5633 = x76 &  n3214 ;
  assign n5630 = ( x78 & ~n3087 ) | ( x78 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n5631 = x77 &  n3082 ;
  assign n5632 = n5630 | n5631 ;
  assign n5634 = ( x76 & ~n5633 ) | ( x76 & n5632 ) | ( ~n5633 & n5632 ) ;
  assign n5635 = ( n693 & ~n3090 ) | ( n693 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n5636 = n5634 | n5635 ;
  assign n5637 = ( x35 & ~n5636 ) | ( x35 & 1'b0 ) | ( ~n5636 & 1'b0 ) ;
  assign n5638 = ~x35 & n5636 ;
  assign n5639 = n5637 | n5638 ;
  assign n5576 = x70 &  n4344 ;
  assign n5573 = ( x72 & ~n4143 ) | ( x72 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n5574 = x71 &  n4138 ;
  assign n5575 = n5573 | n5574 ;
  assign n5577 = ( x70 & ~n5576 ) | ( x70 & n5575 ) | ( ~n5576 & n5575 ) ;
  assign n5578 = ( n345 & ~n4146 ) | ( n345 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n5579 = n5577 | n5578 ;
  assign n5581 = x41 &  n5579 ;
  assign n5580 = ~x41 & n5579 ;
  assign n5582 = ( x41 & ~n5581 ) | ( x41 & n5580 ) | ( ~n5581 & n5580 ) ;
  assign n5583 = ( n5400 & n5410 ) | ( n5400 & n5411 ) | ( n5410 & n5411 ) ;
  assign n5602 = x67 &  n4934 ;
  assign n5599 = ( x69 & ~n4725 ) | ( x69 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n5600 = x68 &  n4720 ;
  assign n5601 = n5599 | n5600 ;
  assign n5603 = ( x67 & ~n5602 ) | ( x67 & n5601 ) | ( ~n5602 & n5601 ) ;
  assign n5604 = ( n246 & ~n4728 ) | ( n246 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n5605 = n5603 | n5604 ;
  assign n5606 = ( x44 & ~n5605 ) | ( x44 & 1'b0 ) | ( ~n5605 & 1'b0 ) ;
  assign n5607 = ~x44 & n5605 ;
  assign n5608 = n5606 | n5607 ;
  assign n5585 = ( x45 & ~x46 ) | ( x45 & n5388 ) | ( ~x46 & n5388 ) ;
  assign n5584 = ( x45 & ~x46 ) | ( x45 & n5087 ) | ( ~x46 & n5087 ) ;
  assign n5586 = ~n5585 |  n5584 ;
  assign n5590 = x64 &  n5586 ;
  assign n5587 = ( x66 & ~n5389 ) | ( x66 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n5588 = x65 &  n5384 ;
  assign n5589 = n5587 | n5588 ;
  assign n5591 = ( x64 & ~n5590 ) | ( x64 & n5589 ) | ( ~n5590 & n5589 ) ;
  assign n5592 = ( n157 & ~n5392 ) | ( n157 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n5593 = n5591 | n5592 ;
  assign n5594 = ( x47 & n5088 ) | ( x47 & n5394 ) | ( n5088 & n5394 ) ;
  assign n5595 = ( x47 & ~n5594 ) | ( x47 & 1'b0 ) | ( ~n5594 & 1'b0 ) ;
  assign n5597 = ( x47 & n5593 ) | ( x47 & n5595 ) | ( n5593 & n5595 ) ;
  assign n5596 = ( n5593 & ~x47 ) | ( n5593 & n5595 ) | ( ~x47 & n5595 ) ;
  assign n5598 = ( x47 & ~n5597 ) | ( x47 & n5596 ) | ( ~n5597 & n5596 ) ;
  assign n5609 = ( n5399 & ~n5608 ) | ( n5399 & n5598 ) | ( ~n5608 & n5598 ) ;
  assign n5610 = ( n5598 & ~n5399 ) | ( n5598 & n5608 ) | ( ~n5399 & n5608 ) ;
  assign n5611 = ( n5609 & ~n5598 ) | ( n5609 & n5610 ) | ( ~n5598 & n5610 ) ;
  assign n5613 = ( n5582 & n5583 ) | ( n5582 & n5611 ) | ( n5583 & n5611 ) ;
  assign n5612 = ( n5583 & ~n5582 ) | ( n5583 & n5611 ) | ( ~n5582 & n5611 ) ;
  assign n5614 = ( n5582 & ~n5613 ) | ( n5582 & n5612 ) | ( ~n5613 & n5612 ) ;
  assign n5615 = ( n5414 & n5415 ) | ( n5414 & n5425 ) | ( n5415 & n5425 ) ;
  assign n5619 = x73 &  n3756 ;
  assign n5616 = ( x75 & ~n3602 ) | ( x75 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n5617 = x74 &  n3597 ;
  assign n5618 = n5616 | n5617 ;
  assign n5620 = ( x73 & ~n5619 ) | ( x73 & n5618 ) | ( ~n5619 & n5618 ) ;
  assign n5621 = ( n540 & ~n3605 ) | ( n540 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n5622 = n5620 | n5621 ;
  assign n5623 = ( x38 & ~n5622 ) | ( x38 & 1'b0 ) | ( ~n5622 & 1'b0 ) ;
  assign n5624 = ~x38 & n5622 ;
  assign n5625 = n5623 | n5624 ;
  assign n5626 = ( n5614 & ~n5615 ) | ( n5614 & n5625 ) | ( ~n5615 & n5625 ) ;
  assign n5627 = ( n5614 & ~n5625 ) | ( n5614 & n5615 ) | ( ~n5625 & n5615 ) ;
  assign n5628 = ( n5626 & ~n5614 ) | ( n5626 & n5627 ) | ( ~n5614 & n5627 ) ;
  assign n5629 = ( n5132 & n5428 ) | ( n5132 & n5438 ) | ( n5428 & n5438 ) ;
  assign n5641 = ( n5628 & n5629 ) | ( n5628 & n5639 ) | ( n5629 & n5639 ) ;
  assign n5640 = ( n5628 & ~n5639 ) | ( n5628 & n5629 ) | ( ~n5639 & n5629 ) ;
  assign n5642 = ( n5639 & ~n5641 ) | ( n5639 & n5640 ) | ( ~n5641 & n5640 ) ;
  assign n5644 = ( n5571 & n5572 ) | ( n5571 & n5642 ) | ( n5572 & n5642 ) ;
  assign n5643 = ( n5572 & ~n5571 ) | ( n5572 & n5642 ) | ( ~n5571 & n5642 ) ;
  assign n5645 = ( n5571 & ~n5644 ) | ( n5571 & n5643 ) | ( ~n5644 & n5643 ) ;
  assign n5555 = x82 &  n2312 ;
  assign n5552 = ( x84 & ~n2195 ) | ( x84 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n5553 = x83 &  n2190 ;
  assign n5554 = n5552 | n5553 ;
  assign n5556 = ( x82 & ~n5555 ) | ( x82 & n5554 ) | ( ~n5555 & n5554 ) ;
  assign n5557 = ( n1199 & ~n2198 ) | ( n1199 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n5558 = n5556 | n5557 ;
  assign n5559 = ( x29 & ~n5558 ) | ( x29 & 1'b0 ) | ( ~n5558 & 1'b0 ) ;
  assign n5560 = ~x29 & n5558 ;
  assign n5561 = n5559 | n5560 ;
  assign n5646 = ( n5457 & ~n5645 ) | ( n5457 & n5561 ) | ( ~n5645 & n5561 ) ;
  assign n5647 = ( n5561 & ~n5457 ) | ( n5561 & n5645 ) | ( ~n5457 & n5645 ) ;
  assign n5648 = ( n5646 & ~n5561 ) | ( n5646 & n5647 ) | ( ~n5561 & n5647 ) ;
  assign n5659 = ( n5461 & ~n5658 ) | ( n5461 & n5648 ) | ( ~n5658 & n5648 ) ;
  assign n5660 = ( n5648 & ~n5461 ) | ( n5648 & n5658 ) | ( ~n5461 & n5658 ) ;
  assign n5661 = ( n5659 & ~n5648 ) | ( n5659 & n5660 ) | ( ~n5648 & n5660 ) ;
  assign n5665 = x88 &  n1551 ;
  assign n5662 = ( x90 & ~n1451 ) | ( x90 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n5663 = x89 &  n1446 ;
  assign n5664 = n5662 | n5663 ;
  assign n5666 = ( x88 & ~n5665 ) | ( x88 & n5664 ) | ( ~n5665 & n5664 ) ;
  assign n5667 = ~n1454 & n1976 ;
  assign n5668 = n5666 | n5667 ;
  assign n5669 = ( x23 & ~n5668 ) | ( x23 & 1'b0 ) | ( ~n5668 & 1'b0 ) ;
  assign n5670 = ~x23 & n5668 ;
  assign n5671 = n5669 | n5670 ;
  assign n5672 = ( n5661 & ~n5465 ) | ( n5661 & n5671 ) | ( ~n5465 & n5671 ) ;
  assign n5673 = ( n5465 & ~n5671 ) | ( n5465 & n5661 ) | ( ~n5671 & n5661 ) ;
  assign n5674 = ( n5672 & ~n5661 ) | ( n5672 & n5673 ) | ( ~n5661 & n5673 ) ;
  assign n5675 = ( n5469 & n5551 ) | ( n5469 & n5674 ) | ( n5551 & n5674 ) ;
  assign n5676 = ( n5469 & ~n5551 ) | ( n5469 & n5674 ) | ( ~n5551 & n5674 ) ;
  assign n5677 = ( n5551 & ~n5675 ) | ( n5551 & n5676 ) | ( ~n5675 & n5676 ) ;
  assign n5535 = x94 &  n942 ;
  assign n5532 = ( x96 & ~n896 ) | ( x96 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n5533 = x95 &  n891 ;
  assign n5534 = n5532 | n5533 ;
  assign n5536 = ( x94 & ~n5535 ) | ( x94 & n5534 ) | ( ~n5535 & n5534 ) ;
  assign n5537 = ~n899 & n2836 ;
  assign n5538 = n5536 | n5537 ;
  assign n5539 = ( x17 & ~n5538 ) | ( x17 & 1'b0 ) | ( ~n5538 & 1'b0 ) ;
  assign n5540 = ~x17 & n5538 ;
  assign n5541 = n5539 | n5540 ;
  assign n5679 = ( n5471 & n5541 ) | ( n5471 & n5677 ) | ( n5541 & n5677 ) ;
  assign n5678 = ( n5471 & ~n5677 ) | ( n5471 & n5541 ) | ( ~n5677 & n5541 ) ;
  assign n5680 = ( n5677 & ~n5679 ) | ( n5677 & n5678 ) | ( ~n5679 & n5678 ) ;
  assign n5684 = x97 &  n713 ;
  assign n5681 = ( x99 & ~n641 ) | ( x99 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n5682 = x98 &  n636 ;
  assign n5683 = n5681 | n5682 ;
  assign n5685 = ( x97 & ~n5684 ) | ( x97 & n5683 ) | ( ~n5684 & n5683 ) ;
  assign n5686 = ~n644 & n3338 ;
  assign n5687 = n5685 | n5686 ;
  assign n5688 = ( x14 & ~n5687 ) | ( x14 & 1'b0 ) | ( ~n5687 & 1'b0 ) ;
  assign n5689 = ~x14 & n5687 ;
  assign n5690 = n5688 | n5689 ;
  assign n5691 = ( n5216 & n5473 ) | ( n5216 & n5483 ) | ( n5473 & n5483 ) ;
  assign n5692 = ( n5680 & ~n5690 ) | ( n5680 & n5691 ) | ( ~n5690 & n5691 ) ;
  assign n5693 = ( n5680 & ~n5691 ) | ( n5680 & n5690 ) | ( ~n5691 & n5690 ) ;
  assign n5694 = ( n5692 & ~n5680 ) | ( n5692 & n5693 ) | ( ~n5680 & n5693 ) ;
  assign n5695 = ( n5488 & n5531 ) | ( n5488 & n5694 ) | ( n5531 & n5694 ) ;
  assign n5696 = ( n5488 & ~n5531 ) | ( n5488 & n5694 ) | ( ~n5531 & n5694 ) ;
  assign n5697 = ( n5531 & ~n5695 ) | ( n5531 & n5696 ) | ( ~n5695 & n5696 ) ;
  assign n5699 = ( n5511 & n5521 ) | ( n5511 & n5697 ) | ( n5521 & n5697 ) ;
  assign n5698 = ( n5521 & ~n5511 ) | ( n5521 & n5697 ) | ( ~n5511 & n5697 ) ;
  assign n5700 = ( n5511 & ~n5699 ) | ( n5511 & n5698 ) | ( ~n5699 & n5698 ) ;
  assign n5701 = ( n5494 & ~n5510 ) | ( n5494 & n5700 ) | ( ~n5510 & n5700 ) ;
  assign n5702 = ( n5494 & ~n5700 ) | ( n5494 & n5510 ) | ( ~n5700 & n5510 ) ;
  assign n5703 = ( n5701 & ~n5494 ) | ( n5701 & n5702 ) | ( ~n5494 & n5702 ) ;
  assign n5707 = ~n136 & x111 ;
  assign n5704 = ( x109 & ~n150 ) | ( x109 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n5705 = ( x110 & ~n131 ) | ( x110 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n5706 = n5704 | n5705 ;
  assign n5708 = ( x111 & ~n5707 ) | ( x111 & n5706 ) | ( ~n5707 & n5706 ) ;
  assign n5709 = ( x110 & ~x111 ) | ( x110 & n5282 ) | ( ~x111 & n5282 ) ;
  assign n5710 = ( x110 & x111 ) | ( x110 & n5282 ) | ( x111 & n5282 ) ;
  assign n5711 = ( ~x111 & ~n5709 ) | ( ~x111 & n5710 ) | ( ~n5709 & n5710 ) ;
  assign n5712 = ( n5708 & ~n139 ) | ( n5708 & n5711 ) | ( ~n139 & n5711 ) ;
  assign n5713 = n139 | n5712 ;
  assign n5714 = ( x2 & ~n5708 ) | ( x2 & n5713 ) | ( ~n5708 & n5713 ) ;
  assign n5715 = ( n5708 & ~x2 ) | ( n5708 & n5713 ) | ( ~x2 & n5713 ) ;
  assign n5716 = ( n5714 & ~n5713 ) | ( n5714 & n5715 ) | ( ~n5713 & n5715 ) ;
  assign n5717 = ( n5703 & ~n5498 ) | ( n5703 & n5716 ) | ( ~n5498 & n5716 ) ;
  assign n5718 = ( n5498 & ~n5716 ) | ( n5498 & n5703 ) | ( ~n5716 & n5703 ) ;
  assign n5719 = ( n5717 & ~n5703 ) | ( n5717 & n5718 ) | ( ~n5703 & n5718 ) ;
  assign n5723 = ~n136 & x112 ;
  assign n5720 = ( x110 & ~n150 ) | ( x110 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n5721 = ( x111 & ~n131 ) | ( x111 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n5722 = n5720 | n5721 ;
  assign n5724 = ( x112 & ~n5723 ) | ( x112 & n5722 ) | ( ~n5723 & n5722 ) ;
  assign n5726 = ( x111 & x112 ) | ( x111 & n5710 ) | ( x112 & n5710 ) ;
  assign n5725 = ( x111 & ~x112 ) | ( x111 & n5710 ) | ( ~x112 & n5710 ) ;
  assign n5727 = ( x112 & ~n5726 ) | ( x112 & n5725 ) | ( ~n5726 & n5725 ) ;
  assign n5728 = ( n139 & ~n5724 ) | ( n139 & n5727 ) | ( ~n5724 & n5727 ) ;
  assign n5729 = ~n139 & n5728 ;
  assign n5730 = ( x2 & n5724 ) | ( x2 & n5729 ) | ( n5724 & n5729 ) ;
  assign n5731 = ( x2 & ~n5729 ) | ( x2 & n5724 ) | ( ~n5729 & n5724 ) ;
  assign n5732 = ( n5729 & ~n5730 ) | ( n5729 & n5731 ) | ( ~n5730 & n5731 ) ;
  assign n5743 = ( n5511 & ~n5521 ) | ( n5511 & n5697 ) | ( ~n5521 & n5697 ) ;
  assign n5747 = x104 &  n353 ;
  assign n5744 = ( x106 & ~n313 ) | ( x106 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n5745 = x105 &  n308 ;
  assign n5746 = n5744 | n5745 ;
  assign n5748 = ( x104 & ~n5747 ) | ( x104 & n5746 ) | ( ~n5747 & n5746 ) ;
  assign n5749 = ~n316 & n4458 ;
  assign n5750 = n5748 | n5749 ;
  assign n5751 = ( x8 & ~n5750 ) | ( x8 & 1'b0 ) | ( ~n5750 & 1'b0 ) ;
  assign n5752 = ~x8 & n5750 ;
  assign n5753 = n5751 | n5752 ;
  assign n5905 = x92 &  n1227 ;
  assign n5902 = ( x94 & ~n1154 ) | ( x94 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n5903 = x93 &  n1149 ;
  assign n5904 = n5902 | n5903 ;
  assign n5906 = ( x92 & ~n5905 ) | ( x92 & n5904 ) | ( ~n5905 & n5904 ) ;
  assign n5907 = ~n1157 & n2401 ;
  assign n5908 = n5906 | n5907 ;
  assign n5909 = ( x20 & ~n5908 ) | ( x20 & 1'b0 ) | ( ~n5908 & 1'b0 ) ;
  assign n5910 = ~x20 & n5908 ;
  assign n5911 = n5909 | n5910 ;
  assign n5777 = x83 &  n2312 ;
  assign n5774 = ( x85 & ~n2195 ) | ( x85 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n5775 = x84 &  n2190 ;
  assign n5776 = n5774 | n5775 ;
  assign n5778 = ( x83 & ~n5777 ) | ( x83 & n5776 ) | ( ~n5777 & n5776 ) ;
  assign n5779 = ( n1295 & ~n2198 ) | ( n1295 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n5780 = n5778 | n5779 ;
  assign n5781 = ( x29 & ~n5780 ) | ( x29 & 1'b0 ) | ( ~n5780 & 1'b0 ) ;
  assign n5782 = ~x29 & n5780 ;
  assign n5783 = n5781 | n5782 ;
  assign n5797 = x77 &  n3214 ;
  assign n5794 = ( x79 & ~n3087 ) | ( x79 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n5795 = x78 &  n3082 ;
  assign n5796 = n5794 | n5795 ;
  assign n5798 = ( x77 & ~n5797 ) | ( x77 & n5796 ) | ( ~n5797 & n5796 ) ;
  assign n5799 = ( n766 & ~n3090 ) | ( n766 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n5800 = n5798 | n5799 ;
  assign n5801 = ( x35 & ~n5800 ) | ( x35 & 1'b0 ) | ( ~n5800 & 1'b0 ) ;
  assign n5802 = ~x35 & n5800 ;
  assign n5803 = n5801 | n5802 ;
  assign n5807 = x74 &  n3756 ;
  assign n5804 = ( x76 & ~n3602 ) | ( x76 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n5805 = x75 &  n3597 ;
  assign n5806 = n5804 | n5805 ;
  assign n5808 = ( x74 & ~n5807 ) | ( x74 & n5806 ) | ( ~n5807 & n5806 ) ;
  assign n5809 = ( n603 & ~n3605 ) | ( n603 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n5810 = n5808 | n5809 ;
  assign n5811 = ( x38 & ~n5810 ) | ( x38 & 1'b0 ) | ( ~n5810 & 1'b0 ) ;
  assign n5812 = ~x38 & n5810 ;
  assign n5813 = n5811 | n5812 ;
  assign n5814 = ( n5614 & n5615 ) | ( n5614 & n5625 ) | ( n5615 & n5625 ) ;
  assign n5815 = ( x47 & ~x48 ) | ( x47 & 1'b0 ) | ( ~x48 & 1'b0 ) ;
  assign n5816 = ~x47 & x48 ;
  assign n5817 = n5815 | n5816 ;
  assign n5818 = x64 &  n5817 ;
  assign n5819 = ( x47 & n5593 ) | ( x47 & n5594 ) | ( n5593 & n5594 ) ;
  assign n5820 = ( x47 & ~n5819 ) | ( x47 & 1'b0 ) | ( ~n5819 & 1'b0 ) ;
  assign n5824 = x65 &  n5586 ;
  assign n5821 = ( x67 & ~n5389 ) | ( x67 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n5822 = x66 &  n5384 ;
  assign n5823 = n5821 | n5822 ;
  assign n5825 = ( x65 & ~n5824 ) | ( x65 & n5823 ) | ( ~n5824 & n5823 ) ;
  assign n5826 = n173 | n5392 ;
  assign n5827 = ~n5825 & n5826 ;
  assign n5828 = x47 &  n5827 ;
  assign n5829 = x47 | n5827 ;
  assign n5830 = ~n5828 & n5829 ;
  assign n5831 = ( n5818 & ~n5820 ) | ( n5818 & n5830 ) | ( ~n5820 & n5830 ) ;
  assign n5832 = ( n5818 & ~n5830 ) | ( n5818 & n5820 ) | ( ~n5830 & n5820 ) ;
  assign n5833 = ( n5831 & ~n5818 ) | ( n5831 & n5832 ) | ( ~n5818 & n5832 ) ;
  assign n5837 = x68 &  n4934 ;
  assign n5834 = ( x70 & ~n4725 ) | ( x70 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n5835 = x69 &  n4720 ;
  assign n5836 = n5834 | n5835 ;
  assign n5838 = ( x68 & ~n5837 ) | ( x68 & n5836 ) | ( ~n5837 & n5836 ) ;
  assign n5839 = ( n282 & ~n4728 ) | ( n282 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n5840 = n5838 | n5839 ;
  assign n5841 = ( x44 & ~n5840 ) | ( x44 & 1'b0 ) | ( ~n5840 & 1'b0 ) ;
  assign n5842 = ~x44 & n5840 ;
  assign n5843 = n5841 | n5842 ;
  assign n5844 = ( n5399 & n5598 ) | ( n5399 & n5608 ) | ( n5598 & n5608 ) ;
  assign n5845 = ( n5833 & ~n5843 ) | ( n5833 & n5844 ) | ( ~n5843 & n5844 ) ;
  assign n5846 = ( n5833 & ~n5844 ) | ( n5833 & n5843 ) | ( ~n5844 & n5843 ) ;
  assign n5847 = ( n5845 & ~n5833 ) | ( n5845 & n5846 ) | ( ~n5833 & n5846 ) ;
  assign n5851 = x71 &  n4344 ;
  assign n5848 = ( x73 & ~n4143 ) | ( x73 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n5849 = x72 &  n4138 ;
  assign n5850 = n5848 | n5849 ;
  assign n5852 = ( x71 & ~n5851 ) | ( x71 & n5850 ) | ( ~n5851 & n5850 ) ;
  assign n5853 = ( n389 & ~n4146 ) | ( n389 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n5854 = n5852 | n5853 ;
  assign n5855 = ( x41 & ~n5854 ) | ( x41 & 1'b0 ) | ( ~n5854 & 1'b0 ) ;
  assign n5856 = ~x41 & n5854 ;
  assign n5857 = n5855 | n5856 ;
  assign n5858 = ( n5847 & ~n5613 ) | ( n5847 & n5857 ) | ( ~n5613 & n5857 ) ;
  assign n5859 = ( n5613 & ~n5857 ) | ( n5613 & n5847 ) | ( ~n5857 & n5847 ) ;
  assign n5860 = ( n5858 & ~n5847 ) | ( n5858 & n5859 ) | ( ~n5847 & n5859 ) ;
  assign n5861 = ( n5813 & ~n5814 ) | ( n5813 & n5860 ) | ( ~n5814 & n5860 ) ;
  assign n5862 = ( n5813 & ~n5860 ) | ( n5813 & n5814 ) | ( ~n5860 & n5814 ) ;
  assign n5863 = ( n5861 & ~n5813 ) | ( n5861 & n5862 ) | ( ~n5813 & n5862 ) ;
  assign n5864 = ( n5803 & ~n5641 ) | ( n5803 & n5863 ) | ( ~n5641 & n5863 ) ;
  assign n5865 = ( n5641 & ~n5863 ) | ( n5641 & n5803 ) | ( ~n5863 & n5803 ) ;
  assign n5866 = ( n5864 & ~n5803 ) | ( n5864 & n5865 ) | ( ~n5803 & n5865 ) ;
  assign n5787 = x80 &  n2718 ;
  assign n5784 = ( x82 & ~n2642 ) | ( x82 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n5785 = x81 &  n2637 ;
  assign n5786 = n5784 | n5785 ;
  assign n5788 = ( x80 & ~n5787 ) | ( x80 & n5786 ) | ( ~n5787 & n5786 ) ;
  assign n5789 = ( n1084 & ~n2645 ) | ( n1084 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n5790 = n5788 | n5789 ;
  assign n5791 = ( x32 & ~n5790 ) | ( x32 & 1'b0 ) | ( ~n5790 & 1'b0 ) ;
  assign n5792 = ~x32 & n5790 ;
  assign n5793 = n5791 | n5792 ;
  assign n5867 = ( n5644 & ~n5866 ) | ( n5644 & n5793 ) | ( ~n5866 & n5793 ) ;
  assign n5868 = ( n5793 & ~n5644 ) | ( n5793 & n5866 ) | ( ~n5644 & n5866 ) ;
  assign n5869 = ( n5867 & ~n5793 ) | ( n5867 & n5868 ) | ( ~n5793 & n5868 ) ;
  assign n5870 = ( n5457 & n5561 ) | ( n5457 & n5645 ) | ( n5561 & n5645 ) ;
  assign n5871 = ( n5783 & ~n5869 ) | ( n5783 & n5870 ) | ( ~n5869 & n5870 ) ;
  assign n5872 = ( n5783 & ~n5870 ) | ( n5783 & n5869 ) | ( ~n5870 & n5869 ) ;
  assign n5873 = ( n5871 & ~n5783 ) | ( n5871 & n5872 ) | ( ~n5783 & n5872 ) ;
  assign n5874 = ( n5461 & n5648 ) | ( n5461 & n5658 ) | ( n5648 & n5658 ) ;
  assign n5878 = x86 &  n1894 ;
  assign n5875 = ( x88 & ~n1816 ) | ( x88 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n5876 = x87 &  n1811 ;
  assign n5877 = n5875 | n5876 ;
  assign n5879 = ( x86 & ~n5878 ) | ( x86 & n5877 ) | ( ~n5878 & n5877 ) ;
  assign n5880 = ( n1624 & ~n1819 ) | ( n1624 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n5881 = n5879 | n5880 ;
  assign n5882 = ( x26 & ~n5881 ) | ( x26 & 1'b0 ) | ( ~n5881 & 1'b0 ) ;
  assign n5883 = ~x26 & n5881 ;
  assign n5884 = n5882 | n5883 ;
  assign n5885 = ( n5873 & ~n5874 ) | ( n5873 & n5884 ) | ( ~n5874 & n5884 ) ;
  assign n5886 = ( n5873 & ~n5884 ) | ( n5873 & n5874 ) | ( ~n5884 & n5874 ) ;
  assign n5887 = ( n5885 & ~n5873 ) | ( n5885 & n5886 ) | ( ~n5873 & n5886 ) ;
  assign n5888 = ( n5465 & n5661 ) | ( n5465 & n5671 ) | ( n5661 & n5671 ) ;
  assign n5892 = x89 &  n1551 ;
  assign n5889 = ( x91 & ~n1451 ) | ( x91 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n5890 = x90 &  n1446 ;
  assign n5891 = n5889 | n5890 ;
  assign n5893 = ( x89 & ~n5892 ) | ( x89 & n5891 ) | ( ~n5892 & n5891 ) ;
  assign n5894 = ~n1454 & n2108 ;
  assign n5895 = n5893 | n5894 ;
  assign n5896 = ( x23 & ~n5895 ) | ( x23 & 1'b0 ) | ( ~n5895 & 1'b0 ) ;
  assign n5897 = ~x23 & n5895 ;
  assign n5898 = n5896 | n5897 ;
  assign n5899 = ( n5887 & ~n5888 ) | ( n5887 & n5898 ) | ( ~n5888 & n5898 ) ;
  assign n5900 = ( n5888 & ~n5887 ) | ( n5888 & n5898 ) | ( ~n5887 & n5898 ) ;
  assign n5901 = ( n5899 & ~n5898 ) | ( n5899 & n5900 ) | ( ~n5898 & n5900 ) ;
  assign n5912 = ( n5676 & ~n5911 ) | ( n5676 & n5901 ) | ( ~n5911 & n5901 ) ;
  assign n5913 = ( n5901 & ~n5676 ) | ( n5901 & n5911 ) | ( ~n5676 & n5911 ) ;
  assign n5914 = ( n5912 & ~n5901 ) | ( n5912 & n5913 ) | ( ~n5901 & n5913 ) ;
  assign n5767 = x95 &  n942 ;
  assign n5764 = ( x97 & ~n896 ) | ( x97 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n5765 = x96 &  n891 ;
  assign n5766 = n5764 | n5765 ;
  assign n5768 = ( x95 & ~n5767 ) | ( x95 & n5766 ) | ( ~n5767 & n5766 ) ;
  assign n5769 = ~n899 & n2999 ;
  assign n5770 = n5768 | n5769 ;
  assign n5771 = ( x17 & ~n5770 ) | ( x17 & 1'b0 ) | ( ~n5770 & 1'b0 ) ;
  assign n5772 = ~x17 & n5770 ;
  assign n5773 = n5771 | n5772 ;
  assign n5915 = ( n5678 & n5773 ) | ( n5678 & n5914 ) | ( n5773 & n5914 ) ;
  assign n5916 = ( n5678 & ~n5914 ) | ( n5678 & n5773 ) | ( ~n5914 & n5773 ) ;
  assign n5917 = ( n5914 & ~n5915 ) | ( n5914 & n5916 ) | ( ~n5915 & n5916 ) ;
  assign n5918 = ( n5690 & ~n5680 ) | ( n5690 & n5691 ) | ( ~n5680 & n5691 ) ;
  assign n5922 = x98 &  n713 ;
  assign n5919 = ( x100 & ~n641 ) | ( x100 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n5920 = x99 &  n636 ;
  assign n5921 = n5919 | n5920 ;
  assign n5923 = ( x98 & ~n5922 ) | ( x98 & n5921 ) | ( ~n5922 & n5921 ) ;
  assign n5924 = n644 | n3354 ;
  assign n5925 = ~n5923 & n5924 ;
  assign n5926 = x14 &  n5925 ;
  assign n5927 = x14 | n5925 ;
  assign n5928 = ~n5926 & n5927 ;
  assign n5929 = ( n5917 & n5918 ) | ( n5917 & n5928 ) | ( n5918 & n5928 ) ;
  assign n5930 = ( n5918 & ~n5917 ) | ( n5918 & n5928 ) | ( ~n5917 & n5928 ) ;
  assign n5931 = ( n5917 & ~n5929 ) | ( n5917 & n5930 ) | ( ~n5929 & n5930 ) ;
  assign n5757 = x101 &  n503 ;
  assign n5754 = ( x103 & ~n450 ) | ( x103 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n5755 = x102 &  n445 ;
  assign n5756 = n5754 | n5755 ;
  assign n5758 = ( x101 & ~n5757 ) | ( x101 & n5756 ) | ( ~n5757 & n5756 ) ;
  assign n5759 = n453 | n4056 ;
  assign n5760 = ~n5758 & n5759 ;
  assign n5761 = x11 &  n5760 ;
  assign n5762 = x11 | n5760 ;
  assign n5763 = ~n5761 & n5762 ;
  assign n5932 = ( n5695 & ~n5931 ) | ( n5695 & n5763 ) | ( ~n5931 & n5763 ) ;
  assign n5933 = ( n5763 & ~n5695 ) | ( n5763 & n5931 ) | ( ~n5695 & n5931 ) ;
  assign n5934 = ( n5932 & ~n5763 ) | ( n5932 & n5933 ) | ( ~n5763 & n5933 ) ;
  assign n5935 = ( n5743 & ~n5753 ) | ( n5743 & n5934 ) | ( ~n5753 & n5934 ) ;
  assign n5936 = ( n5743 & ~n5934 ) | ( n5743 & n5753 ) | ( ~n5934 & n5753 ) ;
  assign n5937 = ( n5935 & ~n5743 ) | ( n5935 & n5936 ) | ( ~n5743 & n5936 ) ;
  assign n5736 = x107 &  n225 ;
  assign n5733 = ( x109 & ~n197 ) | ( x109 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n5734 = x108 &  n192 ;
  assign n5735 = n5733 | n5734 ;
  assign n5737 = ( x107 & ~n5736 ) | ( x107 & n5735 ) | ( ~n5736 & n5735 ) ;
  assign n5738 = ~n200 & n5267 ;
  assign n5739 = n5737 | n5738 ;
  assign n5740 = ( x5 & ~n5739 ) | ( x5 & 1'b0 ) | ( ~n5739 & 1'b0 ) ;
  assign n5741 = ~x5 & n5739 ;
  assign n5742 = n5740 | n5741 ;
  assign n5938 = ( n5701 & ~n5937 ) | ( n5701 & n5742 ) | ( ~n5937 & n5742 ) ;
  assign n5939 = ( n5701 & ~n5742 ) | ( n5701 & n5937 ) | ( ~n5742 & n5937 ) ;
  assign n5940 = ( n5938 & ~n5701 ) | ( n5938 & n5939 ) | ( ~n5701 & n5939 ) ;
  assign n5941 = ( n5717 & n5732 ) | ( n5717 & n5940 ) | ( n5732 & n5940 ) ;
  assign n5942 = ( n5717 & ~n5732 ) | ( n5717 & n5940 ) | ( ~n5732 & n5940 ) ;
  assign n5943 = ( n5732 & ~n5941 ) | ( n5732 & n5942 ) | ( ~n5941 & n5942 ) ;
  assign n6165 = ~n136 & x113 ;
  assign n6162 = ( x111 & ~n150 ) | ( x111 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n6163 = ( x112 & ~n131 ) | ( x112 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n6164 = n6162 | n6163 ;
  assign n6166 = ( x113 & ~n6165 ) | ( x113 & n6164 ) | ( ~n6165 & n6164 ) ;
  assign n6167 = ( x112 & ~x113 ) | ( x112 & n5726 ) | ( ~x113 & n5726 ) ;
  assign n6168 = ( x112 & x113 ) | ( x112 & n5726 ) | ( x113 & n5726 ) ;
  assign n6169 = ( ~x113 & ~n6167 ) | ( ~x113 & n6168 ) | ( ~n6167 & n6168 ) ;
  assign n6170 = ( n6166 & ~n139 ) | ( n6166 & n6169 ) | ( ~n139 & n6169 ) ;
  assign n6171 = n139 | n6170 ;
  assign n6173 = ( x2 & n6166 ) | ( x2 & n6171 ) | ( n6166 & n6171 ) ;
  assign n6172 = ( x2 & ~n6171 ) | ( x2 & n6166 ) | ( ~n6171 & n6166 ) ;
  assign n6174 = ( n6171 & ~n6173 ) | ( n6171 & n6172 ) | ( ~n6173 & n6172 ) ;
  assign n6138 = x105 &  n353 ;
  assign n6135 = ( x107 & ~n313 ) | ( x107 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n6136 = x106 &  n308 ;
  assign n6137 = n6135 | n6136 ;
  assign n6139 = ( x105 & ~n6138 ) | ( x105 & n6137 ) | ( ~n6138 & n6137 ) ;
  assign n6140 = ~n316 & n4848 ;
  assign n6141 = n6139 | n6140 ;
  assign n6142 = ( x8 & ~n6141 ) | ( x8 & 1'b0 ) | ( ~n6141 & 1'b0 ) ;
  assign n6143 = ~x8 & n6141 ;
  assign n6144 = n6142 | n6143 ;
  assign n5957 = x99 &  n713 ;
  assign n5954 = ( x101 & ~n641 ) | ( x101 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n5955 = x100 &  n636 ;
  assign n5956 = n5954 | n5955 ;
  assign n5958 = ( x99 & ~n5957 ) | ( x99 & n5956 ) | ( ~n5957 & n5956 ) ;
  assign n5959 = n644 | n3694 ;
  assign n5960 = ~n5958 & n5959 ;
  assign n5961 = x14 &  n5960 ;
  assign n5962 = x14 | n5960 ;
  assign n5963 = ~n5961 & n5962 ;
  assign n5967 = x93 &  n1227 ;
  assign n5964 = ( x95 & ~n1154 ) | ( x95 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n5965 = x94 &  n1149 ;
  assign n5966 = n5964 | n5965 ;
  assign n5968 = ( x93 & ~n5967 ) | ( x93 & n5966 ) | ( ~n5967 & n5966 ) ;
  assign n5969 = ~n1157 & n2547 ;
  assign n5970 = n5968 | n5969 ;
  assign n5971 = ( x20 & ~n5970 ) | ( x20 & 1'b0 ) | ( ~n5970 & 1'b0 ) ;
  assign n5972 = ~x20 & n5970 ;
  assign n5973 = n5971 | n5972 ;
  assign n5977 = x90 &  n1551 ;
  assign n5974 = ( x92 & ~n1451 ) | ( x92 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n5975 = x91 &  n1446 ;
  assign n5976 = n5974 | n5975 ;
  assign n5978 = ( x90 & ~n5977 ) | ( x90 & n5976 ) | ( ~n5977 & n5976 ) ;
  assign n5979 = ~n1454 & n2248 ;
  assign n5980 = n5978 | n5979 ;
  assign n5981 = ( x23 & ~n5980 ) | ( x23 & 1'b0 ) | ( ~n5980 & 1'b0 ) ;
  assign n5982 = ~x23 & n5980 ;
  assign n5983 = n5981 | n5982 ;
  assign n5987 = x87 &  n1894 ;
  assign n5984 = ( x89 & ~n1816 ) | ( x89 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n5985 = x88 &  n1811 ;
  assign n5986 = n5984 | n5985 ;
  assign n5988 = ( x87 & ~n5987 ) | ( x87 & n5986 ) | ( ~n5987 & n5986 ) ;
  assign n5989 = ( n1741 & ~n1819 ) | ( n1741 & 1'b0 ) | ( ~n1819 & 1'b0 ) ;
  assign n5990 = n5988 | n5989 ;
  assign n5991 = ( x26 & ~n5990 ) | ( x26 & 1'b0 ) | ( ~n5990 & 1'b0 ) ;
  assign n5992 = ~x26 & n5990 ;
  assign n5993 = n5991 | n5992 ;
  assign n5997 = x84 &  n2312 ;
  assign n5994 = ( x86 & ~n2195 ) | ( x86 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n5995 = x85 &  n2190 ;
  assign n5996 = n5994 | n5995 ;
  assign n5998 = ( x84 & ~n5997 ) | ( x84 & n5996 ) | ( ~n5997 & n5996 ) ;
  assign n5999 = ( n1496 & ~n2198 ) | ( n1496 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n6000 = n5998 | n5999 ;
  assign n6001 = ( x29 & ~n6000 ) | ( x29 & 1'b0 ) | ( ~n6000 & 1'b0 ) ;
  assign n6002 = ~x29 & n6000 ;
  assign n6003 = n6001 | n6002 ;
  assign n6007 = x81 &  n2718 ;
  assign n6004 = ( x83 & ~n2642 ) | ( x83 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n6005 = x82 &  n2637 ;
  assign n6006 = n6004 | n6005 ;
  assign n6008 = ( x81 & ~n6007 ) | ( x81 & n6006 ) | ( ~n6007 & n6006 ) ;
  assign n6009 = ( n1100 & ~n2645 ) | ( n1100 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n6010 = n6008 | n6009 ;
  assign n6011 = ( x32 & ~n6010 ) | ( x32 & 1'b0 ) | ( ~n6010 & 1'b0 ) ;
  assign n6012 = ~x32 & n6010 ;
  assign n6013 = n6011 | n6012 ;
  assign n6017 = x66 &  n5586 ;
  assign n6014 = ( x68 & ~n5389 ) | ( x68 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n6015 = x67 &  n5384 ;
  assign n6016 = n6014 | n6015 ;
  assign n6018 = ( x66 & ~n6017 ) | ( x66 & n6016 ) | ( ~n6017 & n6016 ) ;
  assign n6019 = ( n213 & ~n5392 ) | ( n213 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n6020 = n6018 | n6019 ;
  assign n6021 = ( x47 & ~n6020 ) | ( x47 & 1'b0 ) | ( ~n6020 & 1'b0 ) ;
  assign n6022 = ~x47 & n6020 ;
  assign n6023 = n6021 | n6022 ;
  assign n6024 = ( x50 & ~n5818 ) | ( x50 & 1'b0 ) | ( ~n5818 & 1'b0 ) ;
  assign n6025 = ( x48 & x49 ) | ( x48 & n5815 ) | ( x49 & n5815 ) ;
  assign n6026 = ( x48 & ~n5816 ) | ( x48 & x49 ) | ( ~n5816 & x49 ) ;
  assign n6027 = ~n6025 &  n6026 ;
  assign n6028 = x64 &  n6027 ;
  assign n6029 = ~x49 & x50 ;
  assign n6030 = ( x49 & ~x50 ) | ( x49 & 1'b0 ) | ( ~x50 & 1'b0 ) ;
  assign n6031 = n6029 | n6030 ;
  assign n6032 = ~n5817 |  n6031 ;
  assign n6033 = ( x65 & ~n6032 ) | ( x65 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n6034 = n6028 | n6033 ;
  assign n6035 = ~n5817 | ~n6031 ;
  assign n6036 = ( n142 & ~n6035 ) | ( n142 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n6037 = n6034 | n6036 ;
  assign n6039 = ( x50 & n6024 ) | ( x50 & n6037 ) | ( n6024 & n6037 ) ;
  assign n6038 = ( x50 & ~n6024 ) | ( x50 & n6037 ) | ( ~n6024 & n6037 ) ;
  assign n6040 = ( n6024 & ~n6039 ) | ( n6024 & n6038 ) | ( ~n6039 & n6038 ) ;
  assign n6042 = ( n5832 & n6023 ) | ( n5832 & n6040 ) | ( n6023 & n6040 ) ;
  assign n6041 = ( n5832 & ~n6023 ) | ( n5832 & n6040 ) | ( ~n6023 & n6040 ) ;
  assign n6043 = ( n6023 & ~n6042 ) | ( n6023 & n6041 ) | ( ~n6042 & n6041 ) ;
  assign n6054 = ( n5843 & ~n5833 ) | ( n5843 & n5844 ) | ( ~n5833 & n5844 ) ;
  assign n6047 = x69 &  n4934 ;
  assign n6044 = ( x71 & ~n4725 ) | ( x71 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n6045 = x70 &  n4720 ;
  assign n6046 = n6044 | n6045 ;
  assign n6048 = ( x69 & ~n6047 ) | ( x69 & n6046 ) | ( ~n6047 & n6046 ) ;
  assign n6049 = ( n298 & ~n4728 ) | ( n298 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n6050 = n6048 | n6049 ;
  assign n6051 = ( x44 & ~n6050 ) | ( x44 & 1'b0 ) | ( ~n6050 & 1'b0 ) ;
  assign n6052 = ~x44 & n6050 ;
  assign n6053 = n6051 | n6052 ;
  assign n6055 = ( n6043 & ~n6054 ) | ( n6043 & n6053 ) | ( ~n6054 & n6053 ) ;
  assign n6056 = ( n6043 & ~n6053 ) | ( n6043 & n6054 ) | ( ~n6053 & n6054 ) ;
  assign n6057 = ( n6055 & ~n6043 ) | ( n6055 & n6056 ) | ( ~n6043 & n6056 ) ;
  assign n6062 = x72 &  n4344 ;
  assign n6059 = ( x74 & ~n4143 ) | ( x74 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n6060 = x73 &  n4138 ;
  assign n6061 = n6059 | n6060 ;
  assign n6063 = ( x72 & ~n6062 ) | ( x72 & n6061 ) | ( ~n6062 & n6061 ) ;
  assign n6064 = ( n482 & ~n4146 ) | ( n482 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n6065 = n6063 | n6064 ;
  assign n6066 = ( x41 & ~n6065 ) | ( x41 & 1'b0 ) | ( ~n6065 & 1'b0 ) ;
  assign n6067 = ~x41 & n6065 ;
  assign n6068 = n6066 | n6067 ;
  assign n6058 = ( n5613 & ~n5847 ) | ( n5613 & n5857 ) | ( ~n5847 & n5857 ) ;
  assign n6069 = ( n6057 & ~n6068 ) | ( n6057 & n6058 ) | ( ~n6068 & n6058 ) ;
  assign n6070 = ( n6057 & ~n6058 ) | ( n6057 & n6068 ) | ( ~n6058 & n6068 ) ;
  assign n6071 = ( n6069 & ~n6057 ) | ( n6069 & n6070 ) | ( ~n6057 & n6070 ) ;
  assign n6075 = x75 &  n3756 ;
  assign n6072 = ( x77 & ~n3602 ) | ( x77 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n6073 = x76 &  n3597 ;
  assign n6074 = n6072 | n6073 ;
  assign n6076 = ( x75 & ~n6075 ) | ( x75 & n6074 ) | ( ~n6075 & n6074 ) ;
  assign n6077 = ( n677 & ~n3605 ) | ( n677 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n6078 = n6076 | n6077 ;
  assign n6079 = ( x38 & ~n6078 ) | ( x38 & 1'b0 ) | ( ~n6078 & 1'b0 ) ;
  assign n6080 = ~x38 & n6078 ;
  assign n6081 = n6079 | n6080 ;
  assign n6082 = ( n6071 & ~n5862 ) | ( n6071 & n6081 ) | ( ~n5862 & n6081 ) ;
  assign n6083 = ( n5862 & ~n6081 ) | ( n5862 & n6071 ) | ( ~n6081 & n6071 ) ;
  assign n6084 = ( n6082 & ~n6071 ) | ( n6082 & n6083 ) | ( ~n6071 & n6083 ) ;
  assign n6088 = x78 &  n3214 ;
  assign n6085 = ( x80 & ~n3087 ) | ( x80 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n6086 = x79 &  n3082 ;
  assign n6087 = n6085 | n6086 ;
  assign n6089 = ( x78 & ~n6088 ) | ( x78 & n6087 ) | ( ~n6088 & n6087 ) ;
  assign n6090 = ( n842 & ~n3090 ) | ( n842 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n6091 = n6089 | n6090 ;
  assign n6092 = ( x35 & ~n6091 ) | ( x35 & 1'b0 ) | ( ~n6091 & 1'b0 ) ;
  assign n6093 = ~x35 & n6091 ;
  assign n6094 = n6092 | n6093 ;
  assign n6095 = ( n6084 & ~n5865 ) | ( n6084 & n6094 ) | ( ~n5865 & n6094 ) ;
  assign n6096 = ( n5865 & ~n6094 ) | ( n5865 & n6084 ) | ( ~n6094 & n6084 ) ;
  assign n6097 = ( n6095 & ~n6084 ) | ( n6095 & n6096 ) | ( ~n6084 & n6096 ) ;
  assign n6098 = ( n5867 & n6013 ) | ( n5867 & n6097 ) | ( n6013 & n6097 ) ;
  assign n6099 = ( n5867 & ~n6013 ) | ( n5867 & n6097 ) | ( ~n6013 & n6097 ) ;
  assign n6100 = ( n6013 & ~n6098 ) | ( n6013 & n6099 ) | ( ~n6098 & n6099 ) ;
  assign n6101 = ( n5871 & n6003 ) | ( n5871 & n6100 ) | ( n6003 & n6100 ) ;
  assign n6102 = ( n5871 & ~n6003 ) | ( n5871 & n6100 ) | ( ~n6003 & n6100 ) ;
  assign n6103 = ( n6003 & ~n6101 ) | ( n6003 & n6102 ) | ( ~n6101 & n6102 ) ;
  assign n6104 = ( n5874 & ~n5873 ) | ( n5874 & n5884 ) | ( ~n5873 & n5884 ) ;
  assign n6105 = ( n5993 & n6103 ) | ( n5993 & n6104 ) | ( n6103 & n6104 ) ;
  assign n6106 = ( n6103 & ~n5993 ) | ( n6103 & n6104 ) | ( ~n5993 & n6104 ) ;
  assign n6107 = ( n5993 & ~n6105 ) | ( n5993 & n6106 ) | ( ~n6105 & n6106 ) ;
  assign n6109 = ( n5900 & n5983 ) | ( n5900 & n6107 ) | ( n5983 & n6107 ) ;
  assign n6108 = ( n5900 & ~n5983 ) | ( n5900 & n6107 ) | ( ~n5983 & n6107 ) ;
  assign n6110 = ( n5983 & ~n6109 ) | ( n5983 & n6108 ) | ( ~n6109 & n6108 ) ;
  assign n6111 = ( n5676 & ~n5901 ) | ( n5676 & n5911 ) | ( ~n5901 & n5911 ) ;
  assign n6112 = ( n5973 & ~n6110 ) | ( n5973 & n6111 ) | ( ~n6110 & n6111 ) ;
  assign n6113 = ( n5973 & ~n6111 ) | ( n5973 & n6110 ) | ( ~n6111 & n6110 ) ;
  assign n6114 = ( n6112 & ~n5973 ) | ( n6112 & n6113 ) | ( ~n5973 & n6113 ) ;
  assign n6118 = x96 &  n942 ;
  assign n6115 = ( x98 & ~n896 ) | ( x98 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n6116 = x97 &  n891 ;
  assign n6117 = n6115 | n6116 ;
  assign n6119 = ( x96 & ~n6118 ) | ( x96 & n6117 ) | ( ~n6118 & n6117 ) ;
  assign n6120 = ~n899 & n3170 ;
  assign n6121 = n6119 | n6120 ;
  assign n6122 = ( x17 & ~n6121 ) | ( x17 & 1'b0 ) | ( ~n6121 & 1'b0 ) ;
  assign n6123 = ~x17 & n6121 ;
  assign n6124 = n6122 | n6123 ;
  assign n6125 = ( n5916 & ~n6114 ) | ( n5916 & n6124 ) | ( ~n6114 & n6124 ) ;
  assign n6126 = ( n5916 & ~n6124 ) | ( n5916 & n6114 ) | ( ~n6124 & n6114 ) ;
  assign n6127 = ( n6125 & ~n5916 ) | ( n6125 & n6126 ) | ( ~n5916 & n6126 ) ;
  assign n6128 = ( n5917 & ~n5918 ) | ( n5917 & n5928 ) | ( ~n5918 & n5928 ) ;
  assign n6129 = ( n5963 & ~n6127 ) | ( n5963 & n6128 ) | ( ~n6127 & n6128 ) ;
  assign n6130 = ( n5963 & ~n6128 ) | ( n5963 & n6127 ) | ( ~n6128 & n6127 ) ;
  assign n6131 = ( n6129 & ~n5963 ) | ( n6129 & n6130 ) | ( ~n5963 & n6130 ) ;
  assign n5947 = x102 &  n503 ;
  assign n5944 = ( x104 & ~n450 ) | ( x104 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n5945 = x103 &  n445 ;
  assign n5946 = n5944 | n5945 ;
  assign n5948 = ( x102 & ~n5947 ) | ( x102 & n5946 ) | ( ~n5947 & n5946 ) ;
  assign n5949 = n453 | n4249 ;
  assign n5950 = ~n5948 & n5949 ;
  assign n5951 = x11 &  n5950 ;
  assign n5952 = x11 | n5950 ;
  assign n5953 = ~n5951 & n5952 ;
  assign n6132 = ( n5932 & ~n6131 ) | ( n5932 & n5953 ) | ( ~n6131 & n5953 ) ;
  assign n6133 = ( n5953 & ~n5932 ) | ( n5953 & n6131 ) | ( ~n5932 & n6131 ) ;
  assign n6134 = ( n6132 & ~n5953 ) | ( n6132 & n6133 ) | ( ~n5953 & n6133 ) ;
  assign n6145 = ( n5753 & ~n5743 ) | ( n5753 & n5934 ) | ( ~n5743 & n5934 ) ;
  assign n6146 = ( n6144 & ~n6134 ) | ( n6144 & n6145 ) | ( ~n6134 & n6145 ) ;
  assign n6147 = ( n6134 & ~n6144 ) | ( n6134 & n6145 ) | ( ~n6144 & n6145 ) ;
  assign n6148 = ( n6146 & ~n6145 ) | ( n6146 & n6147 ) | ( ~n6145 & n6147 ) ;
  assign n6152 = x108 &  n225 ;
  assign n6149 = ( x110 & ~n197 ) | ( x110 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n6150 = x109 &  n192 ;
  assign n6151 = n6149 | n6150 ;
  assign n6153 = ( x108 & ~n6152 ) | ( x108 & n6151 ) | ( ~n6152 & n6151 ) ;
  assign n6154 = n200 | n5283 ;
  assign n6155 = ~n6153 & n6154 ;
  assign n6156 = x5 &  n6155 ;
  assign n6157 = x5 | n6155 ;
  assign n6158 = ~n6156 & n6157 ;
  assign n6160 = ( n5938 & n6148 ) | ( n5938 & n6158 ) | ( n6148 & n6158 ) ;
  assign n6159 = ( n6148 & ~n5938 ) | ( n6148 & n6158 ) | ( ~n5938 & n6158 ) ;
  assign n6161 = ( n5938 & ~n6160 ) | ( n5938 & n6159 ) | ( ~n6160 & n6159 ) ;
  assign n6175 = ( n5942 & ~n6174 ) | ( n5942 & n6161 ) | ( ~n6174 & n6161 ) ;
  assign n6176 = ( n6161 & ~n5942 ) | ( n6161 & n6174 ) | ( ~n5942 & n6174 ) ;
  assign n6177 = ( n6175 & ~n6161 ) | ( n6175 & n6176 ) | ( ~n6161 & n6176 ) ;
  assign n6181 = ~n136 & x114 ;
  assign n6178 = ( x112 & ~n150 ) | ( x112 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n6179 = ( x113 & ~n131 ) | ( x113 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n6180 = n6178 | n6179 ;
  assign n6182 = ( x114 & ~n6181 ) | ( x114 & n6180 ) | ( ~n6181 & n6180 ) ;
  assign n6183 = ( x113 & ~x114 ) | ( x113 & n6168 ) | ( ~x114 & n6168 ) ;
  assign n6184 = ( x113 & x114 ) | ( x113 & n6168 ) | ( x114 & n6168 ) ;
  assign n6185 = ( ~x114 & ~n6183 ) | ( ~x114 & n6184 ) | ( ~n6183 & n6184 ) ;
  assign n6186 = ( n6182 & ~n139 ) | ( n6182 & n6185 ) | ( ~n139 & n6185 ) ;
  assign n6187 = n139 | n6186 ;
  assign n6189 = ( x2 & n6182 ) | ( x2 & n6187 ) | ( n6182 & n6187 ) ;
  assign n6188 = ( x2 & ~n6187 ) | ( x2 & n6182 ) | ( ~n6187 & n6182 ) ;
  assign n6190 = ( n6187 & ~n6189 ) | ( n6187 & n6188 ) | ( ~n6189 & n6188 ) ;
  assign n6191 = ( n5938 & ~n6158 ) | ( n5938 & n6148 ) | ( ~n6158 & n6148 ) ;
  assign n6195 = x109 &  n225 ;
  assign n6192 = ( x111 & ~n197 ) | ( x111 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n6193 = x110 &  n192 ;
  assign n6194 = n6192 | n6193 ;
  assign n6196 = ( x109 & ~n6195 ) | ( x109 & n6194 ) | ( ~n6195 & n6194 ) ;
  assign n6197 = n200 | n5711 ;
  assign n6198 = ~n6196 & n6197 ;
  assign n6199 = x5 &  n6198 ;
  assign n6200 = x5 | n6198 ;
  assign n6201 = ~n6199 & n6200 ;
  assign n6202 = ( n6134 & n6144 ) | ( n6134 & n6145 ) | ( n6144 & n6145 ) ;
  assign n6206 = x106 &  n353 ;
  assign n6203 = ( x108 & ~n313 ) | ( x108 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n6204 = x107 &  n308 ;
  assign n6205 = n6203 | n6204 ;
  assign n6207 = ( x106 & ~n6206 ) | ( x106 & n6205 ) | ( ~n6206 & n6205 ) ;
  assign n6208 = n316 | n5055 ;
  assign n6209 = ~n6207 & n6208 ;
  assign n6210 = x8 &  n6209 ;
  assign n6211 = x8 | n6209 ;
  assign n6212 = ~n6210 & n6211 ;
  assign n6216 = x103 &  n503 ;
  assign n6213 = ( x105 & ~n450 ) | ( x105 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n6214 = x104 &  n445 ;
  assign n6215 = n6213 | n6214 ;
  assign n6217 = ( x103 & ~n6216 ) | ( x103 & n6215 ) | ( ~n6216 & n6215 ) ;
  assign n6218 = ~n453 & n4442 ;
  assign n6219 = n6217 | n6218 ;
  assign n6220 = ( x11 & ~n6219 ) | ( x11 & 1'b0 ) | ( ~n6219 & 1'b0 ) ;
  assign n6221 = ~x11 & n6219 ;
  assign n6222 = n6220 | n6221 ;
  assign n6226 = x100 &  n713 ;
  assign n6223 = ( x102 & ~n641 ) | ( x102 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n6224 = x101 &  n636 ;
  assign n6225 = n6223 | n6224 ;
  assign n6227 = ( x100 & ~n6226 ) | ( x100 & n6225 ) | ( ~n6226 & n6225 ) ;
  assign n6228 = n644 | n3872 ;
  assign n6229 = ~n6227 & n6228 ;
  assign n6230 = x14 &  n6229 ;
  assign n6231 = x14 | n6229 ;
  assign n6232 = ~n6230 & n6231 ;
  assign n6236 = x94 &  n1227 ;
  assign n6233 = ( x96 & ~n1154 ) | ( x96 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n6234 = x95 &  n1149 ;
  assign n6235 = n6233 | n6234 ;
  assign n6237 = ( x94 & ~n6236 ) | ( x94 & n6235 ) | ( ~n6236 & n6235 ) ;
  assign n6238 = ~n1157 & n2836 ;
  assign n6239 = n6237 | n6238 ;
  assign n6240 = ( x20 & ~n6239 ) | ( x20 & 1'b0 ) | ( ~n6239 & 1'b0 ) ;
  assign n6241 = ~x20 & n6239 ;
  assign n6242 = n6240 | n6241 ;
  assign n6243 = ( n5973 & n6110 ) | ( n5973 & n6111 ) | ( n6110 & n6111 ) ;
  assign n6247 = x91 &  n1551 ;
  assign n6244 = ( x93 & ~n1451 ) | ( x93 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n6245 = x92 &  n1446 ;
  assign n6246 = n6244 | n6245 ;
  assign n6248 = ( x91 & ~n6247 ) | ( x91 & n6246 ) | ( ~n6247 & n6246 ) ;
  assign n6249 = n1454 | n2264 ;
  assign n6250 = ~n6248 & n6249 ;
  assign n6251 = x23 &  n6250 ;
  assign n6252 = x23 | n6250 ;
  assign n6253 = ~n6251 & n6252 ;
  assign n6354 = x85 &  n2312 ;
  assign n6351 = ( x87 & ~n2195 ) | ( x87 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n6352 = x86 &  n2190 ;
  assign n6353 = n6351 | n6352 ;
  assign n6355 = ( x85 & ~n6354 ) | ( x85 & n6353 ) | ( ~n6354 & n6353 ) ;
  assign n6356 = ( n1512 & ~n2198 ) | ( n1512 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n6357 = n6355 | n6356 ;
  assign n6358 = ( x29 & ~n6357 ) | ( x29 & 1'b0 ) | ( ~n6357 & 1'b0 ) ;
  assign n6359 = ~x29 & n6357 ;
  assign n6360 = n6358 | n6359 ;
  assign n6267 = x79 &  n3214 ;
  assign n6264 = ( x81 & ~n3087 ) | ( x81 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n6265 = x80 &  n3082 ;
  assign n6266 = n6264 | n6265 ;
  assign n6268 = ( x79 & ~n6267 ) | ( x79 & n6266 ) | ( ~n6267 & n6266 ) ;
  assign n6269 = ( n994 & ~n3090 ) | ( n994 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n6270 = n6268 | n6269 ;
  assign n6271 = ( x35 & ~n6270 ) | ( x35 & 1'b0 ) | ( ~n6270 & 1'b0 ) ;
  assign n6272 = ~x35 & n6270 ;
  assign n6273 = n6271 | n6272 ;
  assign n6274 = ( n5865 & n6084 ) | ( n5865 & n6094 ) | ( n6084 & n6094 ) ;
  assign n6335 = x76 &  n3756 ;
  assign n6332 = ( x78 & ~n3602 ) | ( x78 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n6333 = x77 &  n3597 ;
  assign n6334 = n6332 | n6333 ;
  assign n6336 = ( x76 & ~n6335 ) | ( x76 & n6334 ) | ( ~n6335 & n6334 ) ;
  assign n6337 = ( n693 & ~n3605 ) | ( n693 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n6338 = n6336 | n6337 ;
  assign n6339 = ( x38 & ~n6338 ) | ( x38 & 1'b0 ) | ( ~n6338 & 1'b0 ) ;
  assign n6340 = ~x38 & n6338 ;
  assign n6341 = n6339 | n6340 ;
  assign n6278 = x70 &  n4934 ;
  assign n6275 = ( x72 & ~n4725 ) | ( x72 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n6276 = x71 &  n4720 ;
  assign n6277 = n6275 | n6276 ;
  assign n6279 = ( x70 & ~n6278 ) | ( x70 & n6277 ) | ( ~n6278 & n6277 ) ;
  assign n6280 = ( n345 & ~n4728 ) | ( n345 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n6281 = n6279 | n6280 ;
  assign n6283 = x44 &  n6281 ;
  assign n6282 = ~x44 & n6281 ;
  assign n6284 = ( x44 & ~n6283 ) | ( x44 & n6282 ) | ( ~n6283 & n6282 ) ;
  assign n6285 = ( n6043 & n6053 ) | ( n6043 & n6054 ) | ( n6053 & n6054 ) ;
  assign n6304 = x67 &  n5586 ;
  assign n6301 = ( x69 & ~n5389 ) | ( x69 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n6302 = x68 &  n5384 ;
  assign n6303 = n6301 | n6302 ;
  assign n6305 = ( x67 & ~n6304 ) | ( x67 & n6303 ) | ( ~n6304 & n6303 ) ;
  assign n6306 = ( n246 & ~n5392 ) | ( n246 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n6307 = n6305 | n6306 ;
  assign n6308 = ( x47 & ~n6307 ) | ( x47 & 1'b0 ) | ( ~n6307 & 1'b0 ) ;
  assign n6309 = ~x47 & n6307 ;
  assign n6310 = n6308 | n6309 ;
  assign n6287 = ( x48 & ~x49 ) | ( x48 & n6031 ) | ( ~x49 & n6031 ) ;
  assign n6286 = ( x48 & ~x49 ) | ( x48 & n5817 ) | ( ~x49 & n5817 ) ;
  assign n6288 = ~n6287 |  n6286 ;
  assign n6292 = x64 &  n6288 ;
  assign n6289 = ( x66 & ~n6032 ) | ( x66 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n6290 = x65 &  n6027 ;
  assign n6291 = n6289 | n6290 ;
  assign n6293 = ( x64 & ~n6292 ) | ( x64 & n6291 ) | ( ~n6292 & n6291 ) ;
  assign n6294 = ( n157 & ~n6035 ) | ( n157 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n6295 = n6293 | n6294 ;
  assign n6296 = ( x50 & n5818 ) | ( x50 & n6037 ) | ( n5818 & n6037 ) ;
  assign n6297 = ( x50 & ~n6296 ) | ( x50 & 1'b0 ) | ( ~n6296 & 1'b0 ) ;
  assign n6299 = ( x50 & n6295 ) | ( x50 & n6297 ) | ( n6295 & n6297 ) ;
  assign n6298 = ( n6295 & ~x50 ) | ( n6295 & n6297 ) | ( ~x50 & n6297 ) ;
  assign n6300 = ( x50 & ~n6299 ) | ( x50 & n6298 ) | ( ~n6299 & n6298 ) ;
  assign n6311 = ( n6042 & ~n6310 ) | ( n6042 & n6300 ) | ( ~n6310 & n6300 ) ;
  assign n6312 = ( n6300 & ~n6042 ) | ( n6300 & n6310 ) | ( ~n6042 & n6310 ) ;
  assign n6313 = ( n6311 & ~n6300 ) | ( n6311 & n6312 ) | ( ~n6300 & n6312 ) ;
  assign n6315 = ( n6284 & n6285 ) | ( n6284 & n6313 ) | ( n6285 & n6313 ) ;
  assign n6314 = ( n6285 & ~n6284 ) | ( n6285 & n6313 ) | ( ~n6284 & n6313 ) ;
  assign n6316 = ( n6284 & ~n6315 ) | ( n6284 & n6314 ) | ( ~n6315 & n6314 ) ;
  assign n6317 = ( n6057 & n6058 ) | ( n6057 & n6068 ) | ( n6058 & n6068 ) ;
  assign n6321 = x73 &  n4344 ;
  assign n6318 = ( x75 & ~n4143 ) | ( x75 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n6319 = x74 &  n4138 ;
  assign n6320 = n6318 | n6319 ;
  assign n6322 = ( x73 & ~n6321 ) | ( x73 & n6320 ) | ( ~n6321 & n6320 ) ;
  assign n6323 = ( n540 & ~n4146 ) | ( n540 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n6324 = n6322 | n6323 ;
  assign n6325 = ( x41 & ~n6324 ) | ( x41 & 1'b0 ) | ( ~n6324 & 1'b0 ) ;
  assign n6326 = ~x41 & n6324 ;
  assign n6327 = n6325 | n6326 ;
  assign n6328 = ( n6316 & ~n6317 ) | ( n6316 & n6327 ) | ( ~n6317 & n6327 ) ;
  assign n6329 = ( n6316 & ~n6327 ) | ( n6316 & n6317 ) | ( ~n6327 & n6317 ) ;
  assign n6330 = ( n6328 & ~n6316 ) | ( n6328 & n6329 ) | ( ~n6316 & n6329 ) ;
  assign n6331 = ( n5862 & n6071 ) | ( n5862 & n6081 ) | ( n6071 & n6081 ) ;
  assign n6343 = ( n6330 & n6331 ) | ( n6330 & n6341 ) | ( n6331 & n6341 ) ;
  assign n6342 = ( n6330 & ~n6341 ) | ( n6330 & n6331 ) | ( ~n6341 & n6331 ) ;
  assign n6344 = ( n6341 & ~n6343 ) | ( n6341 & n6342 ) | ( ~n6343 & n6342 ) ;
  assign n6346 = ( n6273 & n6274 ) | ( n6273 & n6344 ) | ( n6274 & n6344 ) ;
  assign n6345 = ( n6274 & ~n6273 ) | ( n6274 & n6344 ) | ( ~n6273 & n6344 ) ;
  assign n6347 = ( n6273 & ~n6346 ) | ( n6273 & n6345 ) | ( ~n6346 & n6345 ) ;
  assign n6257 = x82 &  n2718 ;
  assign n6254 = ( x84 & ~n2642 ) | ( x84 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n6255 = x83 &  n2637 ;
  assign n6256 = n6254 | n6255 ;
  assign n6258 = ( x82 & ~n6257 ) | ( x82 & n6256 ) | ( ~n6257 & n6256 ) ;
  assign n6259 = ( n1199 & ~n2645 ) | ( n1199 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n6260 = n6258 | n6259 ;
  assign n6261 = ( x32 & ~n6260 ) | ( x32 & 1'b0 ) | ( ~n6260 & 1'b0 ) ;
  assign n6262 = ~x32 & n6260 ;
  assign n6263 = n6261 | n6262 ;
  assign n6348 = ( n6098 & ~n6347 ) | ( n6098 & n6263 ) | ( ~n6347 & n6263 ) ;
  assign n6349 = ( n6263 & ~n6098 ) | ( n6263 & n6347 ) | ( ~n6098 & n6347 ) ;
  assign n6350 = ( n6348 & ~n6263 ) | ( n6348 & n6349 ) | ( ~n6263 & n6349 ) ;
  assign n6361 = ( n6101 & ~n6360 ) | ( n6101 & n6350 ) | ( ~n6360 & n6350 ) ;
  assign n6362 = ( n6350 & ~n6101 ) | ( n6350 & n6360 ) | ( ~n6101 & n6360 ) ;
  assign n6363 = ( n6361 & ~n6350 ) | ( n6361 & n6362 ) | ( ~n6350 & n6362 ) ;
  assign n6367 = x88 &  n1894 ;
  assign n6364 = ( x90 & ~n1816 ) | ( x90 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n6365 = x89 &  n1811 ;
  assign n6366 = n6364 | n6365 ;
  assign n6368 = ( x88 & ~n6367 ) | ( x88 & n6366 ) | ( ~n6367 & n6366 ) ;
  assign n6369 = ~n1819 & n1976 ;
  assign n6370 = n6368 | n6369 ;
  assign n6371 = ( x26 & ~n6370 ) | ( x26 & 1'b0 ) | ( ~n6370 & 1'b0 ) ;
  assign n6372 = ~x26 & n6370 ;
  assign n6373 = n6371 | n6372 ;
  assign n6374 = ( n6363 & ~n6105 ) | ( n6363 & n6373 ) | ( ~n6105 & n6373 ) ;
  assign n6375 = ( n6105 & ~n6373 ) | ( n6105 & n6363 ) | ( ~n6373 & n6363 ) ;
  assign n6376 = ( n6374 & ~n6363 ) | ( n6374 & n6375 ) | ( ~n6363 & n6375 ) ;
  assign n6377 = ( n6109 & n6253 ) | ( n6109 & n6376 ) | ( n6253 & n6376 ) ;
  assign n6378 = ( n6109 & ~n6253 ) | ( n6109 & n6376 ) | ( ~n6253 & n6376 ) ;
  assign n6379 = ( n6253 & ~n6377 ) | ( n6253 & n6378 ) | ( ~n6377 & n6378 ) ;
  assign n6380 = ( n6242 & ~n6243 ) | ( n6242 & n6379 ) | ( ~n6243 & n6379 ) ;
  assign n6381 = ( n6242 & ~n6379 ) | ( n6242 & n6243 ) | ( ~n6379 & n6243 ) ;
  assign n6382 = ( n6380 & ~n6242 ) | ( n6380 & n6381 ) | ( ~n6242 & n6381 ) ;
  assign n6383 = ( n5916 & n6114 ) | ( n5916 & n6124 ) | ( n6114 & n6124 ) ;
  assign n6387 = x97 &  n942 ;
  assign n6384 = ( x99 & ~n896 ) | ( x99 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n6385 = x98 &  n891 ;
  assign n6386 = n6384 | n6385 ;
  assign n6388 = ( x97 & ~n6387 ) | ( x97 & n6386 ) | ( ~n6387 & n6386 ) ;
  assign n6389 = ~n899 & n3338 ;
  assign n6390 = n6388 | n6389 ;
  assign n6391 = ( x17 & ~n6390 ) | ( x17 & 1'b0 ) | ( ~n6390 & 1'b0 ) ;
  assign n6392 = ~x17 & n6390 ;
  assign n6393 = n6391 | n6392 ;
  assign n6395 = ( n6382 & n6383 ) | ( n6382 & n6393 ) | ( n6383 & n6393 ) ;
  assign n6394 = ( n6383 & ~n6382 ) | ( n6383 & n6393 ) | ( ~n6382 & n6393 ) ;
  assign n6396 = ( n6382 & ~n6395 ) | ( n6382 & n6394 ) | ( ~n6395 & n6394 ) ;
  assign n6397 = ( n6129 & n6232 ) | ( n6129 & n6396 ) | ( n6232 & n6396 ) ;
  assign n6398 = ( n6129 & ~n6232 ) | ( n6129 & n6396 ) | ( ~n6232 & n6396 ) ;
  assign n6399 = ( n6232 & ~n6397 ) | ( n6232 & n6398 ) | ( ~n6397 & n6398 ) ;
  assign n6401 = ( n6132 & n6222 ) | ( n6132 & n6399 ) | ( n6222 & n6399 ) ;
  assign n6400 = ( n6132 & ~n6222 ) | ( n6132 & n6399 ) | ( ~n6222 & n6399 ) ;
  assign n6402 = ( n6222 & ~n6401 ) | ( n6222 & n6400 ) | ( ~n6401 & n6400 ) ;
  assign n6404 = ( n6202 & n6212 ) | ( n6202 & n6402 ) | ( n6212 & n6402 ) ;
  assign n6403 = ( n6212 & ~n6202 ) | ( n6212 & n6402 ) | ( ~n6202 & n6402 ) ;
  assign n6405 = ( n6202 & ~n6404 ) | ( n6202 & n6403 ) | ( ~n6404 & n6403 ) ;
  assign n6407 = ( n6191 & n6201 ) | ( n6191 & n6405 ) | ( n6201 & n6405 ) ;
  assign n6406 = ( n6201 & ~n6191 ) | ( n6201 & n6405 ) | ( ~n6191 & n6405 ) ;
  assign n6408 = ( n6191 & ~n6407 ) | ( n6191 & n6406 ) | ( ~n6407 & n6406 ) ;
  assign n6409 = ( n5942 & n6161 ) | ( n5942 & n6174 ) | ( n6161 & n6174 ) ;
  assign n6410 = ( n6190 & ~n6408 ) | ( n6190 & n6409 ) | ( ~n6408 & n6409 ) ;
  assign n6411 = ( n6190 & ~n6409 ) | ( n6190 & n6408 ) | ( ~n6409 & n6408 ) ;
  assign n6412 = ( n6410 & ~n6190 ) | ( n6410 & n6411 ) | ( ~n6190 & n6411 ) ;
  assign n6429 = x110 &  n225 ;
  assign n6426 = ( x112 & ~n197 ) | ( x112 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n6427 = x111 &  n192 ;
  assign n6428 = n6426 | n6427 ;
  assign n6430 = ( x110 & ~n6429 ) | ( x110 & n6428 ) | ( ~n6429 & n6428 ) ;
  assign n6431 = ~n200 & n5727 ;
  assign n6432 = n6430 | n6431 ;
  assign n6433 = ( x5 & ~n6432 ) | ( x5 & 1'b0 ) | ( ~n6432 & 1'b0 ) ;
  assign n6434 = ~x5 & n6432 ;
  assign n6435 = n6433 | n6434 ;
  assign n6450 = x104 &  n503 ;
  assign n6447 = ( x106 & ~n450 ) | ( x106 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n6448 = x105 &  n445 ;
  assign n6449 = n6447 | n6448 ;
  assign n6451 = ( x104 & ~n6450 ) | ( x104 & n6449 ) | ( ~n6450 & n6449 ) ;
  assign n6452 = ~n453 & n4458 ;
  assign n6453 = n6451 | n6452 ;
  assign n6454 = ( x11 & ~n6453 ) | ( x11 & 1'b0 ) | ( ~n6453 & 1'b0 ) ;
  assign n6455 = ~x11 & n6453 ;
  assign n6456 = n6454 | n6455 ;
  assign n6470 = x98 &  n942 ;
  assign n6467 = ( x100 & ~n896 ) | ( x100 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n6468 = x99 &  n891 ;
  assign n6469 = n6467 | n6468 ;
  assign n6471 = ( x98 & ~n6470 ) | ( x98 & n6469 ) | ( ~n6470 & n6469 ) ;
  assign n6472 = n899 | n3354 ;
  assign n6473 = ~n6471 & n6472 ;
  assign n6474 = x17 &  n6473 ;
  assign n6475 = x17 | n6473 ;
  assign n6476 = ~n6474 & n6475 ;
  assign n6608 = x92 &  n1551 ;
  assign n6605 = ( x94 & ~n1451 ) | ( x94 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n6606 = x93 &  n1446 ;
  assign n6607 = n6605 | n6606 ;
  assign n6609 = ( x92 & ~n6608 ) | ( x92 & n6607 ) | ( ~n6608 & n6607 ) ;
  assign n6610 = ~n1454 & n2401 ;
  assign n6611 = n6609 | n6610 ;
  assign n6612 = ( x23 & ~n6611 ) | ( x23 & 1'b0 ) | ( ~n6611 & 1'b0 ) ;
  assign n6613 = ~x23 & n6611 ;
  assign n6614 = n6612 | n6613 ;
  assign n6480 = x83 &  n2718 ;
  assign n6477 = ( x85 & ~n2642 ) | ( x85 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n6478 = x84 &  n2637 ;
  assign n6479 = n6477 | n6478 ;
  assign n6481 = ( x83 & ~n6480 ) | ( x83 & n6479 ) | ( ~n6480 & n6479 ) ;
  assign n6482 = ( n1295 & ~n2645 ) | ( n1295 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n6483 = n6481 | n6482 ;
  assign n6484 = ( x32 & ~n6483 ) | ( x32 & 1'b0 ) | ( ~n6483 & 1'b0 ) ;
  assign n6485 = ~x32 & n6483 ;
  assign n6486 = n6484 | n6485 ;
  assign n6490 = x80 &  n3214 ;
  assign n6487 = ( x82 & ~n3087 ) | ( x82 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n6488 = x81 &  n3082 ;
  assign n6489 = n6487 | n6488 ;
  assign n6491 = ( x80 & ~n6490 ) | ( x80 & n6489 ) | ( ~n6490 & n6489 ) ;
  assign n6492 = ( n1084 & ~n3090 ) | ( n1084 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n6493 = n6491 | n6492 ;
  assign n6494 = ( x35 & ~n6493 ) | ( x35 & 1'b0 ) | ( ~n6493 & 1'b0 ) ;
  assign n6495 = ~x35 & n6493 ;
  assign n6496 = n6494 | n6495 ;
  assign n6500 = x77 &  n3756 ;
  assign n6497 = ( x79 & ~n3602 ) | ( x79 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n6498 = x78 &  n3597 ;
  assign n6499 = n6497 | n6498 ;
  assign n6501 = ( x77 & ~n6500 ) | ( x77 & n6499 ) | ( ~n6500 & n6499 ) ;
  assign n6502 = ( n766 & ~n3605 ) | ( n766 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n6503 = n6501 | n6502 ;
  assign n6504 = ( x38 & ~n6503 ) | ( x38 & 1'b0 ) | ( ~n6503 & 1'b0 ) ;
  assign n6505 = ~x38 & n6503 ;
  assign n6506 = n6504 | n6505 ;
  assign n6510 = x74 &  n4344 ;
  assign n6507 = ( x76 & ~n4143 ) | ( x76 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n6508 = x75 &  n4138 ;
  assign n6509 = n6507 | n6508 ;
  assign n6511 = ( x74 & ~n6510 ) | ( x74 & n6509 ) | ( ~n6510 & n6509 ) ;
  assign n6512 = ( n603 & ~n4146 ) | ( n603 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n6513 = n6511 | n6512 ;
  assign n6514 = ( x41 & ~n6513 ) | ( x41 & 1'b0 ) | ( ~n6513 & 1'b0 ) ;
  assign n6515 = ~x41 & n6513 ;
  assign n6516 = n6514 | n6515 ;
  assign n6517 = ( n6316 & n6317 ) | ( n6316 & n6327 ) | ( n6317 & n6327 ) ;
  assign n6518 = ( x50 & ~x51 ) | ( x50 & 1'b0 ) | ( ~x51 & 1'b0 ) ;
  assign n6519 = ~x50 & x51 ;
  assign n6520 = n6518 | n6519 ;
  assign n6521 = x64 &  n6520 ;
  assign n6522 = ( x50 & n6295 ) | ( x50 & n6296 ) | ( n6295 & n6296 ) ;
  assign n6523 = ( x50 & ~n6522 ) | ( x50 & 1'b0 ) | ( ~n6522 & 1'b0 ) ;
  assign n6527 = x65 &  n6288 ;
  assign n6524 = ( x67 & ~n6032 ) | ( x67 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n6525 = x66 &  n6027 ;
  assign n6526 = n6524 | n6525 ;
  assign n6528 = ( x65 & ~n6527 ) | ( x65 & n6526 ) | ( ~n6527 & n6526 ) ;
  assign n6529 = n173 | n6035 ;
  assign n6530 = ~n6528 & n6529 ;
  assign n6531 = x50 &  n6530 ;
  assign n6532 = x50 | n6530 ;
  assign n6533 = ~n6531 & n6532 ;
  assign n6534 = ( n6521 & ~n6523 ) | ( n6521 & n6533 ) | ( ~n6523 & n6533 ) ;
  assign n6535 = ( n6521 & ~n6533 ) | ( n6521 & n6523 ) | ( ~n6533 & n6523 ) ;
  assign n6536 = ( n6534 & ~n6521 ) | ( n6534 & n6535 ) | ( ~n6521 & n6535 ) ;
  assign n6540 = x68 &  n5586 ;
  assign n6537 = ( x70 & ~n5389 ) | ( x70 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n6538 = x69 &  n5384 ;
  assign n6539 = n6537 | n6538 ;
  assign n6541 = ( x68 & ~n6540 ) | ( x68 & n6539 ) | ( ~n6540 & n6539 ) ;
  assign n6542 = ( n282 & ~n5392 ) | ( n282 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n6543 = n6541 | n6542 ;
  assign n6544 = ( x47 & ~n6543 ) | ( x47 & 1'b0 ) | ( ~n6543 & 1'b0 ) ;
  assign n6545 = ~x47 & n6543 ;
  assign n6546 = n6544 | n6545 ;
  assign n6547 = ( n6042 & n6300 ) | ( n6042 & n6310 ) | ( n6300 & n6310 ) ;
  assign n6548 = ( n6536 & ~n6546 ) | ( n6536 & n6547 ) | ( ~n6546 & n6547 ) ;
  assign n6549 = ( n6536 & ~n6547 ) | ( n6536 & n6546 ) | ( ~n6547 & n6546 ) ;
  assign n6550 = ( n6548 & ~n6536 ) | ( n6548 & n6549 ) | ( ~n6536 & n6549 ) ;
  assign n6554 = x71 &  n4934 ;
  assign n6551 = ( x73 & ~n4725 ) | ( x73 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n6552 = x72 &  n4720 ;
  assign n6553 = n6551 | n6552 ;
  assign n6555 = ( x71 & ~n6554 ) | ( x71 & n6553 ) | ( ~n6554 & n6553 ) ;
  assign n6556 = ( n389 & ~n4728 ) | ( n389 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n6557 = n6555 | n6556 ;
  assign n6558 = ( x44 & ~n6557 ) | ( x44 & 1'b0 ) | ( ~n6557 & 1'b0 ) ;
  assign n6559 = ~x44 & n6557 ;
  assign n6560 = n6558 | n6559 ;
  assign n6561 = ( n6550 & ~n6315 ) | ( n6550 & n6560 ) | ( ~n6315 & n6560 ) ;
  assign n6562 = ( n6315 & ~n6560 ) | ( n6315 & n6550 ) | ( ~n6560 & n6550 ) ;
  assign n6563 = ( n6561 & ~n6550 ) | ( n6561 & n6562 ) | ( ~n6550 & n6562 ) ;
  assign n6564 = ( n6516 & ~n6517 ) | ( n6516 & n6563 ) | ( ~n6517 & n6563 ) ;
  assign n6565 = ( n6516 & ~n6563 ) | ( n6516 & n6517 ) | ( ~n6563 & n6517 ) ;
  assign n6566 = ( n6564 & ~n6516 ) | ( n6564 & n6565 ) | ( ~n6516 & n6565 ) ;
  assign n6567 = ( n6506 & ~n6343 ) | ( n6506 & n6566 ) | ( ~n6343 & n6566 ) ;
  assign n6568 = ( n6343 & ~n6566 ) | ( n6343 & n6506 ) | ( ~n6566 & n6506 ) ;
  assign n6569 = ( n6567 & ~n6506 ) | ( n6567 & n6568 ) | ( ~n6506 & n6568 ) ;
  assign n6570 = ( n6496 & ~n6346 ) | ( n6496 & n6569 ) | ( ~n6346 & n6569 ) ;
  assign n6571 = ( n6346 & ~n6569 ) | ( n6346 & n6496 ) | ( ~n6569 & n6496 ) ;
  assign n6572 = ( n6570 & ~n6496 ) | ( n6570 & n6571 ) | ( ~n6496 & n6571 ) ;
  assign n6573 = ( n6098 & n6263 ) | ( n6098 & n6347 ) | ( n6263 & n6347 ) ;
  assign n6574 = ( n6486 & ~n6572 ) | ( n6486 & n6573 ) | ( ~n6572 & n6573 ) ;
  assign n6575 = ( n6486 & ~n6573 ) | ( n6486 & n6572 ) | ( ~n6573 & n6572 ) ;
  assign n6576 = ( n6574 & ~n6486 ) | ( n6574 & n6575 ) | ( ~n6486 & n6575 ) ;
  assign n6577 = ( n6101 & n6350 ) | ( n6101 & n6360 ) | ( n6350 & n6360 ) ;
  assign n6581 = x86 &  n2312 ;
  assign n6578 = ( x88 & ~n2195 ) | ( x88 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n6579 = x87 &  n2190 ;
  assign n6580 = n6578 | n6579 ;
  assign n6582 = ( x86 & ~n6581 ) | ( x86 & n6580 ) | ( ~n6581 & n6580 ) ;
  assign n6583 = ( n1624 & ~n2198 ) | ( n1624 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n6584 = n6582 | n6583 ;
  assign n6585 = ( x29 & ~n6584 ) | ( x29 & 1'b0 ) | ( ~n6584 & 1'b0 ) ;
  assign n6586 = ~x29 & n6584 ;
  assign n6587 = n6585 | n6586 ;
  assign n6588 = ( n6576 & ~n6577 ) | ( n6576 & n6587 ) | ( ~n6577 & n6587 ) ;
  assign n6589 = ( n6576 & ~n6587 ) | ( n6576 & n6577 ) | ( ~n6587 & n6577 ) ;
  assign n6590 = ( n6588 & ~n6576 ) | ( n6588 & n6589 ) | ( ~n6576 & n6589 ) ;
  assign n6591 = ( n6105 & n6363 ) | ( n6105 & n6373 ) | ( n6363 & n6373 ) ;
  assign n6595 = x89 &  n1894 ;
  assign n6592 = ( x91 & ~n1816 ) | ( x91 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n6593 = x90 &  n1811 ;
  assign n6594 = n6592 | n6593 ;
  assign n6596 = ( x89 & ~n6595 ) | ( x89 & n6594 ) | ( ~n6595 & n6594 ) ;
  assign n6597 = ~n1819 & n2108 ;
  assign n6598 = n6596 | n6597 ;
  assign n6599 = ( x26 & ~n6598 ) | ( x26 & 1'b0 ) | ( ~n6598 & 1'b0 ) ;
  assign n6600 = ~x26 & n6598 ;
  assign n6601 = n6599 | n6600 ;
  assign n6602 = ( n6590 & ~n6591 ) | ( n6590 & n6601 ) | ( ~n6591 & n6601 ) ;
  assign n6603 = ( n6591 & ~n6590 ) | ( n6591 & n6601 ) | ( ~n6590 & n6601 ) ;
  assign n6604 = ( n6602 & ~n6601 ) | ( n6602 & n6603 ) | ( ~n6601 & n6603 ) ;
  assign n6615 = ( n6378 & ~n6614 ) | ( n6378 & n6604 ) | ( ~n6614 & n6604 ) ;
  assign n6616 = ( n6604 & ~n6378 ) | ( n6604 & n6614 ) | ( ~n6378 & n6614 ) ;
  assign n6617 = ( n6615 & ~n6604 ) | ( n6615 & n6616 ) | ( ~n6604 & n6616 ) ;
  assign n6621 = x95 &  n1227 ;
  assign n6618 = ( x97 & ~n1154 ) | ( x97 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n6619 = x96 &  n1149 ;
  assign n6620 = n6618 | n6619 ;
  assign n6622 = ( x95 & ~n6621 ) | ( x95 & n6620 ) | ( ~n6621 & n6620 ) ;
  assign n6623 = ~n1157 & n2999 ;
  assign n6624 = n6622 | n6623 ;
  assign n6625 = ( x20 & ~n6624 ) | ( x20 & 1'b0 ) | ( ~n6624 & 1'b0 ) ;
  assign n6626 = ~x20 & n6624 ;
  assign n6627 = n6625 | n6626 ;
  assign n6628 = ( n6617 & ~n6381 ) | ( n6617 & n6627 ) | ( ~n6381 & n6627 ) ;
  assign n6629 = ( n6381 & ~n6617 ) | ( n6381 & n6627 ) | ( ~n6617 & n6627 ) ;
  assign n6630 = ( n6628 & ~n6627 ) | ( n6628 & n6629 ) | ( ~n6627 & n6629 ) ;
  assign n6632 = ( n6394 & n6476 ) | ( n6394 & n6630 ) | ( n6476 & n6630 ) ;
  assign n6631 = ( n6476 & ~n6394 ) | ( n6476 & n6630 ) | ( ~n6394 & n6630 ) ;
  assign n6633 = ( n6394 & ~n6632 ) | ( n6394 & n6631 ) | ( ~n6632 & n6631 ) ;
  assign n6460 = x101 &  n713 ;
  assign n6457 = ( x103 & ~n641 ) | ( x103 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n6458 = x102 &  n636 ;
  assign n6459 = n6457 | n6458 ;
  assign n6461 = ( x101 & ~n6460 ) | ( x101 & n6459 ) | ( ~n6460 & n6459 ) ;
  assign n6462 = n644 | n4056 ;
  assign n6463 = ~n6461 & n6462 ;
  assign n6464 = x14 &  n6463 ;
  assign n6465 = x14 | n6463 ;
  assign n6466 = ~n6464 & n6465 ;
  assign n6634 = ( n6397 & ~n6633 ) | ( n6397 & n6466 ) | ( ~n6633 & n6466 ) ;
  assign n6635 = ( n6466 & ~n6397 ) | ( n6466 & n6633 ) | ( ~n6397 & n6633 ) ;
  assign n6636 = ( n6634 & ~n6466 ) | ( n6634 & n6635 ) | ( ~n6466 & n6635 ) ;
  assign n6637 = ( n6456 & ~n6400 ) | ( n6456 & n6636 ) | ( ~n6400 & n6636 ) ;
  assign n6638 = ( n6400 & ~n6636 ) | ( n6400 & n6456 ) | ( ~n6636 & n6456 ) ;
  assign n6639 = ( n6637 & ~n6456 ) | ( n6637 & n6638 ) | ( ~n6456 & n6638 ) ;
  assign n6436 = ( n6202 & ~n6212 ) | ( n6202 & n6402 ) | ( ~n6212 & n6402 ) ;
  assign n6440 = x107 &  n353 ;
  assign n6437 = ( x109 & ~n313 ) | ( x109 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n6438 = x108 &  n308 ;
  assign n6439 = n6437 | n6438 ;
  assign n6441 = ( x107 & ~n6440 ) | ( x107 & n6439 ) | ( ~n6440 & n6439 ) ;
  assign n6442 = ~n316 & n5267 ;
  assign n6443 = n6441 | n6442 ;
  assign n6444 = ( x8 & ~n6443 ) | ( x8 & 1'b0 ) | ( ~n6443 & 1'b0 ) ;
  assign n6445 = ~x8 & n6443 ;
  assign n6446 = n6444 | n6445 ;
  assign n6640 = ( n6436 & n6446 ) | ( n6436 & n6639 ) | ( n6446 & n6639 ) ;
  assign n6641 = ( n6436 & ~n6639 ) | ( n6436 & n6446 ) | ( ~n6639 & n6446 ) ;
  assign n6642 = ( n6639 & ~n6640 ) | ( n6639 & n6641 ) | ( ~n6640 & n6641 ) ;
  assign n6643 = ( n6406 & ~n6435 ) | ( n6406 & n6642 ) | ( ~n6435 & n6642 ) ;
  assign n6644 = ( n6406 & ~n6642 ) | ( n6406 & n6435 ) | ( ~n6642 & n6435 ) ;
  assign n6645 = ( n6643 & ~n6406 ) | ( n6643 & n6644 ) | ( ~n6406 & n6644 ) ;
  assign n6416 = ~n136 & x115 ;
  assign n6413 = ( x113 & ~n150 ) | ( x113 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n6414 = ( x114 & ~n131 ) | ( x114 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n6415 = n6413 | n6414 ;
  assign n6417 = ( x115 & ~n6416 ) | ( x115 & n6415 ) | ( ~n6416 & n6415 ) ;
  assign n6419 = ( x114 & x115 ) | ( x114 & n6184 ) | ( x115 & n6184 ) ;
  assign n6418 = ( x114 & ~x115 ) | ( x114 & n6184 ) | ( ~x115 & n6184 ) ;
  assign n6420 = ( x115 & ~n6419 ) | ( x115 & n6418 ) | ( ~n6419 & n6418 ) ;
  assign n6421 = ( n139 & ~n6417 ) | ( n139 & n6420 ) | ( ~n6417 & n6420 ) ;
  assign n6422 = ~n139 & n6421 ;
  assign n6423 = ( x2 & n6417 ) | ( x2 & n6422 ) | ( n6417 & n6422 ) ;
  assign n6424 = ( x2 & ~n6422 ) | ( x2 & n6417 ) | ( ~n6422 & n6417 ) ;
  assign n6425 = ( n6422 & ~n6423 ) | ( n6422 & n6424 ) | ( ~n6423 & n6424 ) ;
  assign n6646 = ( n6410 & ~n6645 ) | ( n6410 & n6425 ) | ( ~n6645 & n6425 ) ;
  assign n6647 = ( n6425 & ~n6410 ) | ( n6425 & n6645 ) | ( ~n6410 & n6645 ) ;
  assign n6648 = ( n6646 & ~n6425 ) | ( n6646 & n6647 ) | ( ~n6425 & n6647 ) ;
  assign n6662 = x108 &  n353 ;
  assign n6659 = ( x110 & ~n313 ) | ( x110 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n6660 = x109 &  n308 ;
  assign n6661 = n6659 | n6660 ;
  assign n6663 = ( x108 & ~n6662 ) | ( x108 & n6661 ) | ( ~n6662 & n6661 ) ;
  assign n6664 = n316 | n5283 ;
  assign n6665 = ~n6663 & n6664 ;
  assign n6666 = x8 &  n6665 ;
  assign n6667 = x8 | n6665 ;
  assign n6668 = ~n6666 & n6667 ;
  assign n6862 = x105 &  n503 ;
  assign n6859 = ( x107 & ~n450 ) | ( x107 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n6860 = x106 &  n445 ;
  assign n6861 = n6859 | n6860 ;
  assign n6863 = ( x105 & ~n6862 ) | ( x105 & n6861 ) | ( ~n6862 & n6861 ) ;
  assign n6864 = ~n453 & n4848 ;
  assign n6865 = n6863 | n6864 ;
  assign n6866 = ( x11 & ~n6865 ) | ( x11 & 1'b0 ) | ( ~n6865 & 1'b0 ) ;
  assign n6867 = ~x11 & n6865 ;
  assign n6868 = n6866 | n6867 ;
  assign n6682 = x96 &  n1227 ;
  assign n6679 = ( x98 & ~n1154 ) | ( x98 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n6680 = x97 &  n1149 ;
  assign n6681 = n6679 | n6680 ;
  assign n6683 = ( x96 & ~n6682 ) | ( x96 & n6681 ) | ( ~n6682 & n6681 ) ;
  assign n6684 = ~n1157 & n3170 ;
  assign n6685 = n6683 | n6684 ;
  assign n6686 = ( x20 & ~n6685 ) | ( x20 & 1'b0 ) | ( ~n6685 & 1'b0 ) ;
  assign n6687 = ~x20 & n6685 ;
  assign n6688 = n6686 | n6687 ;
  assign n6692 = x93 &  n1551 ;
  assign n6689 = ( x95 & ~n1451 ) | ( x95 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n6690 = x94 &  n1446 ;
  assign n6691 = n6689 | n6690 ;
  assign n6693 = ( x93 & ~n6692 ) | ( x93 & n6691 ) | ( ~n6692 & n6691 ) ;
  assign n6694 = ~n1454 & n2547 ;
  assign n6695 = n6693 | n6694 ;
  assign n6696 = ( x23 & ~n6695 ) | ( x23 & 1'b0 ) | ( ~n6695 & 1'b0 ) ;
  assign n6697 = ~x23 & n6695 ;
  assign n6698 = n6696 | n6697 ;
  assign n6796 = x81 &  n3214 ;
  assign n6793 = ( x83 & ~n3087 ) | ( x83 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n6794 = x82 &  n3082 ;
  assign n6795 = n6793 | n6794 ;
  assign n6797 = ( x81 & ~n6796 ) | ( x81 & n6795 ) | ( ~n6796 & n6795 ) ;
  assign n6798 = ( n1100 & ~n3090 ) | ( n1100 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n6799 = n6797 | n6798 ;
  assign n6800 = ( x35 & ~n6799 ) | ( x35 & 1'b0 ) | ( ~n6799 & 1'b0 ) ;
  assign n6801 = ~x35 & n6799 ;
  assign n6802 = n6800 | n6801 ;
  assign n6712 = x66 &  n6288 ;
  assign n6709 = ( x68 & ~n6032 ) | ( x68 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n6710 = x67 &  n6027 ;
  assign n6711 = n6709 | n6710 ;
  assign n6713 = ( x66 & ~n6712 ) | ( x66 & n6711 ) | ( ~n6712 & n6711 ) ;
  assign n6714 = ( n213 & ~n6035 ) | ( n213 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n6715 = n6713 | n6714 ;
  assign n6716 = ( x50 & ~n6715 ) | ( x50 & 1'b0 ) | ( ~n6715 & 1'b0 ) ;
  assign n6717 = ~x50 & n6715 ;
  assign n6718 = n6716 | n6717 ;
  assign n6719 = ( x53 & ~n6521 ) | ( x53 & 1'b0 ) | ( ~n6521 & 1'b0 ) ;
  assign n6720 = ( x51 & x52 ) | ( x51 & n6518 ) | ( x52 & n6518 ) ;
  assign n6721 = ( x51 & ~n6519 ) | ( x51 & x52 ) | ( ~n6519 & x52 ) ;
  assign n6722 = ~n6720 &  n6721 ;
  assign n6723 = x64 &  n6722 ;
  assign n6724 = ~x52 & x53 ;
  assign n6725 = ( x52 & ~x53 ) | ( x52 & 1'b0 ) | ( ~x53 & 1'b0 ) ;
  assign n6726 = n6724 | n6725 ;
  assign n6727 = ~n6520 |  n6726 ;
  assign n6728 = ( x65 & ~n6727 ) | ( x65 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n6729 = n6723 | n6728 ;
  assign n6730 = ~n6520 | ~n6726 ;
  assign n6731 = ( n142 & ~n6730 ) | ( n142 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n6732 = n6729 | n6731 ;
  assign n6734 = ( x53 & n6719 ) | ( x53 & n6732 ) | ( n6719 & n6732 ) ;
  assign n6733 = ( x53 & ~n6719 ) | ( x53 & n6732 ) | ( ~n6719 & n6732 ) ;
  assign n6735 = ( n6719 & ~n6734 ) | ( n6719 & n6733 ) | ( ~n6734 & n6733 ) ;
  assign n6737 = ( n6535 & n6718 ) | ( n6535 & n6735 ) | ( n6718 & n6735 ) ;
  assign n6736 = ( n6535 & ~n6718 ) | ( n6535 & n6735 ) | ( ~n6718 & n6735 ) ;
  assign n6738 = ( n6718 & ~n6737 ) | ( n6718 & n6736 ) | ( ~n6737 & n6736 ) ;
  assign n6749 = ( n6546 & ~n6536 ) | ( n6546 & n6547 ) | ( ~n6536 & n6547 ) ;
  assign n6742 = x69 &  n5586 ;
  assign n6739 = ( x71 & ~n5389 ) | ( x71 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n6740 = x70 &  n5384 ;
  assign n6741 = n6739 | n6740 ;
  assign n6743 = ( x69 & ~n6742 ) | ( x69 & n6741 ) | ( ~n6742 & n6741 ) ;
  assign n6744 = ( n298 & ~n5392 ) | ( n298 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n6745 = n6743 | n6744 ;
  assign n6746 = ( x47 & ~n6745 ) | ( x47 & 1'b0 ) | ( ~n6745 & 1'b0 ) ;
  assign n6747 = ~x47 & n6745 ;
  assign n6748 = n6746 | n6747 ;
  assign n6750 = ( n6738 & ~n6749 ) | ( n6738 & n6748 ) | ( ~n6749 & n6748 ) ;
  assign n6751 = ( n6738 & ~n6748 ) | ( n6738 & n6749 ) | ( ~n6748 & n6749 ) ;
  assign n6752 = ( n6750 & ~n6738 ) | ( n6750 & n6751 ) | ( ~n6738 & n6751 ) ;
  assign n6757 = x72 &  n4934 ;
  assign n6754 = ( x74 & ~n4725 ) | ( x74 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n6755 = x73 &  n4720 ;
  assign n6756 = n6754 | n6755 ;
  assign n6758 = ( x72 & ~n6757 ) | ( x72 & n6756 ) | ( ~n6757 & n6756 ) ;
  assign n6759 = ( n482 & ~n4728 ) | ( n482 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n6760 = n6758 | n6759 ;
  assign n6761 = ( x44 & ~n6760 ) | ( x44 & 1'b0 ) | ( ~n6760 & 1'b0 ) ;
  assign n6762 = ~x44 & n6760 ;
  assign n6763 = n6761 | n6762 ;
  assign n6753 = ( n6315 & ~n6550 ) | ( n6315 & n6560 ) | ( ~n6550 & n6560 ) ;
  assign n6764 = ( n6752 & ~n6763 ) | ( n6752 & n6753 ) | ( ~n6763 & n6753 ) ;
  assign n6765 = ( n6752 & ~n6753 ) | ( n6752 & n6763 ) | ( ~n6753 & n6763 ) ;
  assign n6766 = ( n6764 & ~n6752 ) | ( n6764 & n6765 ) | ( ~n6752 & n6765 ) ;
  assign n6770 = x75 &  n4344 ;
  assign n6767 = ( x77 & ~n4143 ) | ( x77 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n6768 = x76 &  n4138 ;
  assign n6769 = n6767 | n6768 ;
  assign n6771 = ( x75 & ~n6770 ) | ( x75 & n6769 ) | ( ~n6770 & n6769 ) ;
  assign n6772 = ( n677 & ~n4146 ) | ( n677 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n6773 = n6771 | n6772 ;
  assign n6774 = ( x41 & ~n6773 ) | ( x41 & 1'b0 ) | ( ~n6773 & 1'b0 ) ;
  assign n6775 = ~x41 & n6773 ;
  assign n6776 = n6774 | n6775 ;
  assign n6777 = ( n6766 & ~n6565 ) | ( n6766 & n6776 ) | ( ~n6565 & n6776 ) ;
  assign n6778 = ( n6565 & ~n6776 ) | ( n6565 & n6766 ) | ( ~n6776 & n6766 ) ;
  assign n6779 = ( n6777 & ~n6766 ) | ( n6777 & n6778 ) | ( ~n6766 & n6778 ) ;
  assign n6783 = x78 &  n3756 ;
  assign n6780 = ( x80 & ~n3602 ) | ( x80 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n6781 = x79 &  n3597 ;
  assign n6782 = n6780 | n6781 ;
  assign n6784 = ( x78 & ~n6783 ) | ( x78 & n6782 ) | ( ~n6783 & n6782 ) ;
  assign n6785 = ( n842 & ~n3605 ) | ( n842 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n6786 = n6784 | n6785 ;
  assign n6787 = ( x38 & ~n6786 ) | ( x38 & 1'b0 ) | ( ~n6786 & 1'b0 ) ;
  assign n6788 = ~x38 & n6786 ;
  assign n6789 = n6787 | n6788 ;
  assign n6790 = ( n6779 & ~n6568 ) | ( n6779 & n6789 ) | ( ~n6568 & n6789 ) ;
  assign n6791 = ( n6568 & ~n6789 ) | ( n6568 & n6779 ) | ( ~n6789 & n6779 ) ;
  assign n6792 = ( n6790 & ~n6779 ) | ( n6790 & n6791 ) | ( ~n6779 & n6791 ) ;
  assign n6803 = ( n6571 & ~n6802 ) | ( n6571 & n6792 ) | ( ~n6802 & n6792 ) ;
  assign n6804 = ( n6792 & ~n6571 ) | ( n6792 & n6802 ) | ( ~n6571 & n6802 ) ;
  assign n6805 = ( n6803 & ~n6792 ) | ( n6803 & n6804 ) | ( ~n6792 & n6804 ) ;
  assign n6702 = x84 &  n2718 ;
  assign n6699 = ( x86 & ~n2642 ) | ( x86 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n6700 = x85 &  n2637 ;
  assign n6701 = n6699 | n6700 ;
  assign n6703 = ( x84 & ~n6702 ) | ( x84 & n6701 ) | ( ~n6702 & n6701 ) ;
  assign n6704 = ( n1496 & ~n2645 ) | ( n1496 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n6705 = n6703 | n6704 ;
  assign n6706 = ( x32 & ~n6705 ) | ( x32 & 1'b0 ) | ( ~n6705 & 1'b0 ) ;
  assign n6707 = ~x32 & n6705 ;
  assign n6708 = n6706 | n6707 ;
  assign n6806 = ( n6574 & ~n6805 ) | ( n6574 & n6708 ) | ( ~n6805 & n6708 ) ;
  assign n6807 = ( n6708 & ~n6574 ) | ( n6708 & n6805 ) | ( ~n6574 & n6805 ) ;
  assign n6808 = ( n6806 & ~n6708 ) | ( n6806 & n6807 ) | ( ~n6708 & n6807 ) ;
  assign n6813 = x87 &  n2312 ;
  assign n6810 = ( x89 & ~n2195 ) | ( x89 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n6811 = x88 &  n2190 ;
  assign n6812 = n6810 | n6811 ;
  assign n6814 = ( x87 & ~n6813 ) | ( x87 & n6812 ) | ( ~n6813 & n6812 ) ;
  assign n6815 = ( n1741 & ~n2198 ) | ( n1741 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n6816 = n6814 | n6815 ;
  assign n6817 = ( x29 & ~n6816 ) | ( x29 & 1'b0 ) | ( ~n6816 & 1'b0 ) ;
  assign n6818 = ~x29 & n6816 ;
  assign n6819 = n6817 | n6818 ;
  assign n6809 = ( n6577 & ~n6576 ) | ( n6577 & n6587 ) | ( ~n6576 & n6587 ) ;
  assign n6820 = ( n6808 & ~n6819 ) | ( n6808 & n6809 ) | ( ~n6819 & n6809 ) ;
  assign n6821 = ( n6808 & ~n6809 ) | ( n6808 & n6819 ) | ( ~n6809 & n6819 ) ;
  assign n6822 = ( n6820 & ~n6808 ) | ( n6820 & n6821 ) | ( ~n6808 & n6821 ) ;
  assign n6826 = x90 &  n1894 ;
  assign n6823 = ( x92 & ~n1816 ) | ( x92 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n6824 = x91 &  n1811 ;
  assign n6825 = n6823 | n6824 ;
  assign n6827 = ( x90 & ~n6826 ) | ( x90 & n6825 ) | ( ~n6826 & n6825 ) ;
  assign n6828 = ~n1819 & n2248 ;
  assign n6829 = n6827 | n6828 ;
  assign n6830 = ( x26 & ~n6829 ) | ( x26 & 1'b0 ) | ( ~n6829 & 1'b0 ) ;
  assign n6831 = ~x26 & n6829 ;
  assign n6832 = n6830 | n6831 ;
  assign n6833 = ( n6822 & ~n6603 ) | ( n6822 & n6832 ) | ( ~n6603 & n6832 ) ;
  assign n6834 = ( n6603 & ~n6832 ) | ( n6603 & n6822 ) | ( ~n6832 & n6822 ) ;
  assign n6835 = ( n6833 & ~n6822 ) | ( n6833 & n6834 ) | ( ~n6822 & n6834 ) ;
  assign n6836 = ( n6378 & ~n6604 ) | ( n6378 & n6614 ) | ( ~n6604 & n6614 ) ;
  assign n6837 = ( n6698 & n6835 ) | ( n6698 & n6836 ) | ( n6835 & n6836 ) ;
  assign n6838 = ( n6835 & ~n6698 ) | ( n6835 & n6836 ) | ( ~n6698 & n6836 ) ;
  assign n6839 = ( n6698 & ~n6837 ) | ( n6698 & n6838 ) | ( ~n6837 & n6838 ) ;
  assign n6840 = ( n6629 & n6688 ) | ( n6629 & n6839 ) | ( n6688 & n6839 ) ;
  assign n6841 = ( n6629 & ~n6688 ) | ( n6629 & n6839 ) | ( ~n6688 & n6839 ) ;
  assign n6842 = ( n6688 & ~n6840 ) | ( n6688 & n6841 ) | ( ~n6840 & n6841 ) ;
  assign n6846 = x99 &  n942 ;
  assign n6843 = ( x101 & ~n896 ) | ( x101 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n6844 = x100 &  n891 ;
  assign n6845 = n6843 | n6844 ;
  assign n6847 = ( x99 & ~n6846 ) | ( x99 & n6845 ) | ( ~n6846 & n6845 ) ;
  assign n6848 = n899 | n3694 ;
  assign n6849 = ~n6847 & n6848 ;
  assign n6850 = x17 &  n6849 ;
  assign n6851 = x17 | n6849 ;
  assign n6852 = ~n6850 & n6851 ;
  assign n6853 = ( n6631 & n6842 ) | ( n6631 & n6852 ) | ( n6842 & n6852 ) ;
  assign n6854 = ( n6842 & ~n6631 ) | ( n6842 & n6852 ) | ( ~n6631 & n6852 ) ;
  assign n6855 = ( n6631 & ~n6853 ) | ( n6631 & n6854 ) | ( ~n6853 & n6854 ) ;
  assign n6672 = x102 &  n713 ;
  assign n6669 = ( x104 & ~n641 ) | ( x104 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n6670 = x103 &  n636 ;
  assign n6671 = n6669 | n6670 ;
  assign n6673 = ( x102 & ~n6672 ) | ( x102 & n6671 ) | ( ~n6672 & n6671 ) ;
  assign n6674 = n644 | n4249 ;
  assign n6675 = ~n6673 & n6674 ;
  assign n6676 = x14 &  n6675 ;
  assign n6677 = x14 | n6675 ;
  assign n6678 = ~n6676 & n6677 ;
  assign n6856 = ( n6634 & ~n6855 ) | ( n6634 & n6678 ) | ( ~n6855 & n6678 ) ;
  assign n6857 = ( n6678 & ~n6634 ) | ( n6678 & n6855 ) | ( ~n6634 & n6855 ) ;
  assign n6858 = ( n6856 & ~n6678 ) | ( n6856 & n6857 ) | ( ~n6678 & n6857 ) ;
  assign n6869 = ( n6637 & ~n6868 ) | ( n6637 & n6858 ) | ( ~n6868 & n6858 ) ;
  assign n6870 = ( n6858 & ~n6637 ) | ( n6858 & n6868 ) | ( ~n6637 & n6868 ) ;
  assign n6871 = ( n6869 & ~n6858 ) | ( n6869 & n6870 ) | ( ~n6858 & n6870 ) ;
  assign n6872 = ( n6641 & ~n6668 ) | ( n6641 & n6871 ) | ( ~n6668 & n6871 ) ;
  assign n6873 = ( n6641 & ~n6871 ) | ( n6641 & n6668 ) | ( ~n6871 & n6668 ) ;
  assign n6874 = ( n6872 & ~n6641 ) | ( n6872 & n6873 ) | ( ~n6641 & n6873 ) ;
  assign n6652 = x111 &  n225 ;
  assign n6649 = ( x113 & ~n197 ) | ( x113 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n6650 = x112 &  n192 ;
  assign n6651 = n6649 | n6650 ;
  assign n6653 = ( x111 & ~n6652 ) | ( x111 & n6651 ) | ( ~n6652 & n6651 ) ;
  assign n6654 = n200 | n6169 ;
  assign n6655 = ~n6653 & n6654 ;
  assign n6656 = x5 &  n6655 ;
  assign n6657 = x5 | n6655 ;
  assign n6658 = ~n6656 & n6657 ;
  assign n6875 = ( n6643 & ~n6874 ) | ( n6643 & n6658 ) | ( ~n6874 & n6658 ) ;
  assign n6876 = ( n6643 & ~n6658 ) | ( n6643 & n6874 ) | ( ~n6658 & n6874 ) ;
  assign n6877 = ( n6875 & ~n6643 ) | ( n6875 & n6876 ) | ( ~n6643 & n6876 ) ;
  assign n6881 = ~n136 & x116 ;
  assign n6878 = ( x114 & ~n150 ) | ( x114 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n6879 = ( x115 & ~n131 ) | ( x115 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n6880 = n6878 | n6879 ;
  assign n6882 = ( x116 & ~n6881 ) | ( x116 & n6880 ) | ( ~n6881 & n6880 ) ;
  assign n6883 = ( x115 & ~x116 ) | ( x115 & n6419 ) | ( ~x116 & n6419 ) ;
  assign n6884 = ( x115 & x116 ) | ( x115 & n6419 ) | ( x116 & n6419 ) ;
  assign n6885 = ( ~x116 & ~n6883 ) | ( ~x116 & n6884 ) | ( ~n6883 & n6884 ) ;
  assign n6886 = ( n6882 & ~n139 ) | ( n6882 & n6885 ) | ( ~n139 & n6885 ) ;
  assign n6887 = n139 | n6886 ;
  assign n6889 = ( x2 & n6882 ) | ( x2 & n6887 ) | ( n6882 & n6887 ) ;
  assign n6888 = ( x2 & ~n6887 ) | ( x2 & n6882 ) | ( ~n6887 & n6882 ) ;
  assign n6890 = ( n6887 & ~n6889 ) | ( n6887 & n6888 ) | ( ~n6889 & n6888 ) ;
  assign n6891 = ( n6647 & n6877 ) | ( n6647 & n6890 ) | ( n6877 & n6890 ) ;
  assign n6892 = ( n6647 & ~n6877 ) | ( n6647 & n6890 ) | ( ~n6877 & n6890 ) ;
  assign n6893 = ( n6877 & ~n6891 ) | ( n6877 & n6892 ) | ( ~n6891 & n6892 ) ;
  assign n6894 = ( n6643 & n6658 ) | ( n6643 & n6874 ) | ( n6658 & n6874 ) ;
  assign n6898 = x112 &  n225 ;
  assign n6895 = ( x114 & ~n197 ) | ( x114 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n6896 = x113 &  n192 ;
  assign n6897 = n6895 | n6896 ;
  assign n6899 = ( x112 & ~n6898 ) | ( x112 & n6897 ) | ( ~n6898 & n6897 ) ;
  assign n6900 = n200 | n6185 ;
  assign n6901 = ~n6899 & n6900 ;
  assign n6902 = x5 &  n6901 ;
  assign n6903 = x5 | n6901 ;
  assign n6904 = ~n6902 & n6903 ;
  assign n6908 = x103 &  n713 ;
  assign n6905 = ( x105 & ~n641 ) | ( x105 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n6906 = x104 &  n636 ;
  assign n6907 = n6905 | n6906 ;
  assign n6909 = ( x103 & ~n6908 ) | ( x103 & n6907 ) | ( ~n6908 & n6907 ) ;
  assign n6910 = ~n644 & n4442 ;
  assign n6911 = n6909 | n6910 ;
  assign n6912 = ( x14 & ~n6911 ) | ( x14 & 1'b0 ) | ( ~n6911 & 1'b0 ) ;
  assign n6913 = ~x14 & n6911 ;
  assign n6914 = n6912 | n6913 ;
  assign n6915 = ( n6631 & ~n6842 ) | ( n6631 & n6852 ) | ( ~n6842 & n6852 ) ;
  assign n7082 = x97 &  n1227 ;
  assign n7079 = ( x99 & ~n1154 ) | ( x99 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n7080 = x98 &  n1149 ;
  assign n7081 = n7079 | n7080 ;
  assign n7083 = ( x97 & ~n7082 ) | ( x97 & n7081 ) | ( ~n7082 & n7081 ) ;
  assign n7084 = ~n1157 & n3338 ;
  assign n7085 = n7083 | n7084 ;
  assign n7086 = ( x20 & ~n7085 ) | ( x20 & 1'b0 ) | ( ~n7085 & 1'b0 ) ;
  assign n7087 = ~x20 & n7085 ;
  assign n7088 = n7086 | n7087 ;
  assign n6929 = x94 &  n1551 ;
  assign n6926 = ( x96 & ~n1451 ) | ( x96 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n6927 = x95 &  n1446 ;
  assign n6928 = n6926 | n6927 ;
  assign n6930 = ( x94 & ~n6929 ) | ( x94 & n6928 ) | ( ~n6929 & n6928 ) ;
  assign n6931 = ~n1454 & n2836 ;
  assign n6932 = n6930 | n6931 ;
  assign n6933 = ( x23 & ~n6932 ) | ( x23 & 1'b0 ) | ( ~n6932 & 1'b0 ) ;
  assign n6934 = ~x23 & n6932 ;
  assign n6935 = n6933 | n6934 ;
  assign n6939 = x91 &  n1894 ;
  assign n6936 = ( x93 & ~n1816 ) | ( x93 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n6937 = x92 &  n1811 ;
  assign n6938 = n6936 | n6937 ;
  assign n6940 = ( x91 & ~n6939 ) | ( x91 & n6938 ) | ( ~n6939 & n6938 ) ;
  assign n6941 = n1819 | n2264 ;
  assign n6942 = ~n6940 & n6941 ;
  assign n6943 = x26 &  n6942 ;
  assign n6944 = x26 | n6942 ;
  assign n6945 = ~n6943 & n6944 ;
  assign n6946 = ( n6603 & n6822 ) | ( n6603 & n6832 ) | ( n6822 & n6832 ) ;
  assign n6950 = x85 &  n2718 ;
  assign n6947 = ( x87 & ~n2642 ) | ( x87 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n6948 = x86 &  n2637 ;
  assign n6949 = n6947 | n6948 ;
  assign n6951 = ( x85 & ~n6950 ) | ( x85 & n6949 ) | ( ~n6950 & n6949 ) ;
  assign n6952 = ( n1512 & ~n2645 ) | ( n1512 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n6953 = n6951 | n6952 ;
  assign n6954 = ( x32 & ~n6953 ) | ( x32 & 1'b0 ) | ( ~n6953 & 1'b0 ) ;
  assign n6955 = ~x32 & n6953 ;
  assign n6956 = n6954 | n6955 ;
  assign n6957 = ( n6574 & n6708 ) | ( n6574 & n6805 ) | ( n6708 & n6805 ) ;
  assign n6961 = x79 &  n3756 ;
  assign n6958 = ( x81 & ~n3602 ) | ( x81 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n6959 = x80 &  n3597 ;
  assign n6960 = n6958 | n6959 ;
  assign n6962 = ( x79 & ~n6961 ) | ( x79 & n6960 ) | ( ~n6961 & n6960 ) ;
  assign n6963 = ( n994 & ~n3605 ) | ( n994 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n6964 = n6962 | n6963 ;
  assign n6965 = ( x38 & ~n6964 ) | ( x38 & 1'b0 ) | ( ~n6964 & 1'b0 ) ;
  assign n6966 = ~x38 & n6964 ;
  assign n6967 = n6965 | n6966 ;
  assign n6968 = ( n6568 & n6779 ) | ( n6568 & n6789 ) | ( n6779 & n6789 ) ;
  assign n7029 = x76 &  n4344 ;
  assign n7026 = ( x78 & ~n4143 ) | ( x78 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n7027 = x77 &  n4138 ;
  assign n7028 = n7026 | n7027 ;
  assign n7030 = ( x76 & ~n7029 ) | ( x76 & n7028 ) | ( ~n7029 & n7028 ) ;
  assign n7031 = ( n693 & ~n4146 ) | ( n693 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n7032 = n7030 | n7031 ;
  assign n7033 = ( x41 & ~n7032 ) | ( x41 & 1'b0 ) | ( ~n7032 & 1'b0 ) ;
  assign n7034 = ~x41 & n7032 ;
  assign n7035 = n7033 | n7034 ;
  assign n6972 = x73 &  n4934 ;
  assign n6969 = ( x75 & ~n4725 ) | ( x75 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n6970 = x74 &  n4720 ;
  assign n6971 = n6969 | n6970 ;
  assign n6973 = ( x73 & ~n6972 ) | ( x73 & n6971 ) | ( ~n6972 & n6971 ) ;
  assign n6974 = ( n540 & ~n4728 ) | ( n540 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n6975 = n6973 | n6974 ;
  assign n6976 = ( x44 & ~n6975 ) | ( x44 & 1'b0 ) | ( ~n6975 & 1'b0 ) ;
  assign n6977 = ~x44 & n6975 ;
  assign n6978 = n6976 | n6977 ;
  assign n6979 = ( n6752 & n6753 ) | ( n6752 & n6763 ) | ( n6753 & n6763 ) ;
  assign n6998 = x67 &  n6288 ;
  assign n6995 = ( x69 & ~n6032 ) | ( x69 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n6996 = x68 &  n6027 ;
  assign n6997 = n6995 | n6996 ;
  assign n6999 = ( x67 & ~n6998 ) | ( x67 & n6997 ) | ( ~n6998 & n6997 ) ;
  assign n7000 = ( n246 & ~n6035 ) | ( n246 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n7001 = n6999 | n7000 ;
  assign n7002 = ( x50 & ~n7001 ) | ( x50 & 1'b0 ) | ( ~n7001 & 1'b0 ) ;
  assign n7003 = ~x50 & n7001 ;
  assign n7004 = n7002 | n7003 ;
  assign n6981 = ( x51 & ~x52 ) | ( x51 & n6726 ) | ( ~x52 & n6726 ) ;
  assign n6980 = ( x51 & ~x52 ) | ( x51 & n6520 ) | ( ~x52 & n6520 ) ;
  assign n6982 = ~n6981 |  n6980 ;
  assign n6986 = x64 &  n6982 ;
  assign n6983 = ( x66 & ~n6727 ) | ( x66 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n6984 = x65 &  n6722 ;
  assign n6985 = n6983 | n6984 ;
  assign n6987 = ( x64 & ~n6986 ) | ( x64 & n6985 ) | ( ~n6986 & n6985 ) ;
  assign n6988 = ( n157 & ~n6730 ) | ( n157 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n6989 = n6987 | n6988 ;
  assign n6990 = ( x53 & ~n6521 ) | ( x53 & n6732 ) | ( ~n6521 & n6732 ) ;
  assign n6991 = ~n6732 & n6990 ;
  assign n6992 = ( n6989 & ~x53 ) | ( n6989 & n6991 ) | ( ~x53 & n6991 ) ;
  assign n6993 = ( x53 & ~n6989 ) | ( x53 & n6991 ) | ( ~n6989 & n6991 ) ;
  assign n6994 = ( n6992 & ~n6991 ) | ( n6992 & n6993 ) | ( ~n6991 & n6993 ) ;
  assign n7005 = ( n6737 & ~n7004 ) | ( n6737 & n6994 ) | ( ~n7004 & n6994 ) ;
  assign n7006 = ( n6994 & ~n6737 ) | ( n6994 & n7004 ) | ( ~n6737 & n7004 ) ;
  assign n7007 = ( n7005 & ~n6994 ) | ( n7005 & n7006 ) | ( ~n6994 & n7006 ) ;
  assign n7008 = ( n6738 & n6748 ) | ( n6738 & n6749 ) | ( n6748 & n6749 ) ;
  assign n7012 = x70 &  n5586 ;
  assign n7009 = ( x72 & ~n5389 ) | ( x72 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n7010 = x71 &  n5384 ;
  assign n7011 = n7009 | n7010 ;
  assign n7013 = ( x70 & ~n7012 ) | ( x70 & n7011 ) | ( ~n7012 & n7011 ) ;
  assign n7014 = ( n345 & ~n5392 ) | ( n345 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n7015 = n7013 | n7014 ;
  assign n7016 = ( x47 & ~n7015 ) | ( x47 & 1'b0 ) | ( ~n7015 & 1'b0 ) ;
  assign n7017 = ~x47 & n7015 ;
  assign n7018 = n7016 | n7017 ;
  assign n7019 = ( n7007 & ~n7008 ) | ( n7007 & n7018 ) | ( ~n7008 & n7018 ) ;
  assign n7020 = ( n7007 & ~n7018 ) | ( n7007 & n7008 ) | ( ~n7018 & n7008 ) ;
  assign n7021 = ( n7019 & ~n7007 ) | ( n7019 & n7020 ) | ( ~n7007 & n7020 ) ;
  assign n7023 = ( n6978 & n6979 ) | ( n6978 & n7021 ) | ( n6979 & n7021 ) ;
  assign n7022 = ( n6979 & ~n6978 ) | ( n6979 & n7021 ) | ( ~n6978 & n7021 ) ;
  assign n7024 = ( n6978 & ~n7023 ) | ( n6978 & n7022 ) | ( ~n7023 & n7022 ) ;
  assign n7025 = ( n6565 & n6766 ) | ( n6565 & n6776 ) | ( n6766 & n6776 ) ;
  assign n7037 = ( n7024 & n7025 ) | ( n7024 & n7035 ) | ( n7025 & n7035 ) ;
  assign n7036 = ( n7024 & ~n7035 ) | ( n7024 & n7025 ) | ( ~n7035 & n7025 ) ;
  assign n7038 = ( n7035 & ~n7037 ) | ( n7035 & n7036 ) | ( ~n7037 & n7036 ) ;
  assign n7040 = ( n6967 & n6968 ) | ( n6967 & n7038 ) | ( n6968 & n7038 ) ;
  assign n7039 = ( n6968 & ~n6967 ) | ( n6968 & n7038 ) | ( ~n6967 & n7038 ) ;
  assign n7041 = ( n6967 & ~n7040 ) | ( n6967 & n7039 ) | ( ~n7040 & n7039 ) ;
  assign n7042 = ( n6571 & n6792 ) | ( n6571 & n6802 ) | ( n6792 & n6802 ) ;
  assign n7046 = x82 &  n3214 ;
  assign n7043 = ( x84 & ~n3087 ) | ( x84 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n7044 = x83 &  n3082 ;
  assign n7045 = n7043 | n7044 ;
  assign n7047 = ( x82 & ~n7046 ) | ( x82 & n7045 ) | ( ~n7046 & n7045 ) ;
  assign n7048 = ( n1199 & ~n3090 ) | ( n1199 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n7049 = n7047 | n7048 ;
  assign n7050 = ( x35 & ~n7049 ) | ( x35 & 1'b0 ) | ( ~n7049 & 1'b0 ) ;
  assign n7051 = ~x35 & n7049 ;
  assign n7052 = n7050 | n7051 ;
  assign n7053 = ( n7041 & ~n7042 ) | ( n7041 & n7052 ) | ( ~n7042 & n7052 ) ;
  assign n7054 = ( n7041 & ~n7052 ) | ( n7041 & n7042 ) | ( ~n7052 & n7042 ) ;
  assign n7055 = ( n7053 & ~n7041 ) | ( n7053 & n7054 ) | ( ~n7041 & n7054 ) ;
  assign n7057 = ( n6956 & n6957 ) | ( n6956 & n7055 ) | ( n6957 & n7055 ) ;
  assign n7056 = ( n6957 & ~n6956 ) | ( n6957 & n7055 ) | ( ~n6956 & n7055 ) ;
  assign n7058 = ( n6956 & ~n7057 ) | ( n6956 & n7056 ) | ( ~n7057 & n7056 ) ;
  assign n7059 = ( n6808 & n6809 ) | ( n6808 & n6819 ) | ( n6809 & n6819 ) ;
  assign n7063 = x88 &  n2312 ;
  assign n7060 = ( x90 & ~n2195 ) | ( x90 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n7061 = x89 &  n2190 ;
  assign n7062 = n7060 | n7061 ;
  assign n7064 = ( x88 & ~n7063 ) | ( x88 & n7062 ) | ( ~n7063 & n7062 ) ;
  assign n7065 = ( n1976 & ~n2198 ) | ( n1976 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n7066 = n7064 | n7065 ;
  assign n7067 = ( x29 & ~n7066 ) | ( x29 & 1'b0 ) | ( ~n7066 & 1'b0 ) ;
  assign n7068 = ~x29 & n7066 ;
  assign n7069 = n7067 | n7068 ;
  assign n7070 = ( n7058 & ~n7059 ) | ( n7058 & n7069 ) | ( ~n7059 & n7069 ) ;
  assign n7071 = ( n7058 & ~n7069 ) | ( n7058 & n7059 ) | ( ~n7069 & n7059 ) ;
  assign n7072 = ( n7070 & ~n7058 ) | ( n7070 & n7071 ) | ( ~n7058 & n7071 ) ;
  assign n7073 = ( n6945 & n6946 ) | ( n6945 & n7072 ) | ( n6946 & n7072 ) ;
  assign n7074 = ( n6946 & ~n6945 ) | ( n6946 & n7072 ) | ( ~n6945 & n7072 ) ;
  assign n7075 = ( n6945 & ~n7073 ) | ( n6945 & n7074 ) | ( ~n7073 & n7074 ) ;
  assign n7076 = ( n6935 & ~n6837 ) | ( n6935 & n7075 ) | ( ~n6837 & n7075 ) ;
  assign n7077 = ( n6837 & ~n7075 ) | ( n6837 & n6935 ) | ( ~n7075 & n6935 ) ;
  assign n7078 = ( n7076 & ~n6935 ) | ( n7076 & n7077 ) | ( ~n6935 & n7077 ) ;
  assign n7089 = ( n6840 & ~n7088 ) | ( n6840 & n7078 ) | ( ~n7088 & n7078 ) ;
  assign n7090 = ( n7078 & ~n6840 ) | ( n7078 & n7088 ) | ( ~n6840 & n7088 ) ;
  assign n7091 = ( n7089 & ~n7078 ) | ( n7089 & n7090 ) | ( ~n7078 & n7090 ) ;
  assign n6919 = x100 &  n942 ;
  assign n6916 = ( x102 & ~n896 ) | ( x102 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n6917 = x101 &  n891 ;
  assign n6918 = n6916 | n6917 ;
  assign n6920 = ( x100 & ~n6919 ) | ( x100 & n6918 ) | ( ~n6919 & n6918 ) ;
  assign n6921 = n899 | n3872 ;
  assign n6922 = ~n6920 & n6921 ;
  assign n6923 = x17 &  n6922 ;
  assign n6924 = x17 | n6922 ;
  assign n6925 = ~n6923 & n6924 ;
  assign n7092 = ( n6915 & ~n7091 ) | ( n6915 & n6925 ) | ( ~n7091 & n6925 ) ;
  assign n7093 = ( n6915 & ~n6925 ) | ( n6915 & n7091 ) | ( ~n6925 & n7091 ) ;
  assign n7094 = ( n7092 & ~n6915 ) | ( n7092 & n7093 ) | ( ~n6915 & n7093 ) ;
  assign n7096 = ( n6856 & n6914 ) | ( n6856 & n7094 ) | ( n6914 & n7094 ) ;
  assign n7095 = ( n6856 & ~n6914 ) | ( n6856 & n7094 ) | ( ~n6914 & n7094 ) ;
  assign n7097 = ( n6914 & ~n7096 ) | ( n6914 & n7095 ) | ( ~n7096 & n7095 ) ;
  assign n7098 = ( n6637 & n6858 ) | ( n6637 & n6868 ) | ( n6858 & n6868 ) ;
  assign n7102 = x106 &  n503 ;
  assign n7099 = ( x108 & ~n450 ) | ( x108 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n7100 = x107 &  n445 ;
  assign n7101 = n7099 | n7100 ;
  assign n7103 = ( x106 & ~n7102 ) | ( x106 & n7101 ) | ( ~n7102 & n7101 ) ;
  assign n7104 = n453 | n5055 ;
  assign n7105 = ~n7103 & n7104 ;
  assign n7106 = x11 &  n7105 ;
  assign n7107 = x11 | n7105 ;
  assign n7108 = ~n7106 & n7107 ;
  assign n7109 = ( n7097 & n7098 ) | ( n7097 & n7108 ) | ( n7098 & n7108 ) ;
  assign n7110 = ( n7098 & ~n7097 ) | ( n7098 & n7108 ) | ( ~n7097 & n7108 ) ;
  assign n7111 = ( n7097 & ~n7109 ) | ( n7097 & n7110 ) | ( ~n7109 & n7110 ) ;
  assign n7115 = x109 &  n353 ;
  assign n7112 = ( x111 & ~n313 ) | ( x111 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n7113 = x110 &  n308 ;
  assign n7114 = n7112 | n7113 ;
  assign n7116 = ( x109 & ~n7115 ) | ( x109 & n7114 ) | ( ~n7115 & n7114 ) ;
  assign n7117 = n316 | n5711 ;
  assign n7118 = ~n7116 & n7117 ;
  assign n7119 = x8 &  n7118 ;
  assign n7120 = x8 | n7118 ;
  assign n7121 = ~n7119 & n7120 ;
  assign n7123 = ( n6872 & n7111 ) | ( n6872 & n7121 ) | ( n7111 & n7121 ) ;
  assign n7122 = ( n7111 & ~n6872 ) | ( n7111 & n7121 ) | ( ~n6872 & n7121 ) ;
  assign n7124 = ( n6872 & ~n7123 ) | ( n6872 & n7122 ) | ( ~n7123 & n7122 ) ;
  assign n7125 = ( n6894 & n6904 ) | ( n6894 & n7124 ) | ( n6904 & n7124 ) ;
  assign n7126 = ( n6904 & ~n6894 ) | ( n6904 & n7124 ) | ( ~n6894 & n7124 ) ;
  assign n7127 = ( n6894 & ~n7125 ) | ( n6894 & n7126 ) | ( ~n7125 & n7126 ) ;
  assign n7132 = ~n136 & x117 ;
  assign n7129 = ( x115 & ~n150 ) | ( x115 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n7130 = ( x116 & ~n131 ) | ( x116 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n7131 = n7129 | n7130 ;
  assign n7133 = ( x117 & ~n7132 ) | ( x117 & n7131 ) | ( ~n7132 & n7131 ) ;
  assign n7134 = ( x116 & ~x117 ) | ( x116 & n6884 ) | ( ~x117 & n6884 ) ;
  assign n7135 = ( x116 & x117 ) | ( x116 & n6884 ) | ( x117 & n6884 ) ;
  assign n7136 = ( ~x117 & ~n7134 ) | ( ~x117 & n7135 ) | ( ~n7134 & n7135 ) ;
  assign n7137 = ( n7133 & ~n139 ) | ( n7133 & n7136 ) | ( ~n139 & n7136 ) ;
  assign n7138 = n139 | n7137 ;
  assign n7140 = ( x2 & n7133 ) | ( x2 & n7138 ) | ( n7133 & n7138 ) ;
  assign n7139 = ( x2 & ~n7138 ) | ( x2 & n7133 ) | ( ~n7138 & n7133 ) ;
  assign n7141 = ( n7138 & ~n7140 ) | ( n7138 & n7139 ) | ( ~n7140 & n7139 ) ;
  assign n7128 = ( n6877 & ~n6647 ) | ( n6877 & n6890 ) | ( ~n6647 & n6890 ) ;
  assign n7142 = ( n7127 & ~n7141 ) | ( n7127 & n7128 ) | ( ~n7141 & n7128 ) ;
  assign n7143 = ( n7127 & ~n7128 ) | ( n7127 & n7141 ) | ( ~n7128 & n7141 ) ;
  assign n7144 = ( n7142 & ~n7127 ) | ( n7142 & n7143 ) | ( ~n7127 & n7143 ) ;
  assign n7148 = ~n136 & x118 ;
  assign n7145 = ( x116 & ~n150 ) | ( x116 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n7146 = ( x117 & ~n131 ) | ( x117 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n7147 = n7145 | n7146 ;
  assign n7149 = ( x118 & ~n7148 ) | ( x118 & n7147 ) | ( ~n7148 & n7147 ) ;
  assign n7150 = ( x117 & ~x118 ) | ( x117 & n7135 ) | ( ~x118 & n7135 ) ;
  assign n7151 = ( x117 & x118 ) | ( x117 & n7135 ) | ( x118 & n7135 ) ;
  assign n7152 = ( ~x118 & ~n7150 ) | ( ~x118 & n7151 ) | ( ~n7150 & n7151 ) ;
  assign n7153 = ( n7149 & ~n139 ) | ( n7149 & n7152 ) | ( ~n139 & n7152 ) ;
  assign n7154 = n139 | n7153 ;
  assign n7156 = ( x2 & n7149 ) | ( x2 & n7154 ) | ( n7149 & n7154 ) ;
  assign n7155 = ( x2 & ~n7154 ) | ( x2 & n7149 ) | ( ~n7154 & n7149 ) ;
  assign n7157 = ( n7154 & ~n7156 ) | ( n7154 & n7155 ) | ( ~n7156 & n7155 ) ;
  assign n7158 = ( n7128 & ~n7127 ) | ( n7128 & n7141 ) | ( ~n7127 & n7141 ) ;
  assign n7159 = ( n6894 & ~n7124 ) | ( n6894 & n6904 ) | ( ~n7124 & n6904 ) ;
  assign n7163 = x113 &  n225 ;
  assign n7160 = ( x115 & ~n197 ) | ( x115 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n7161 = x114 &  n192 ;
  assign n7162 = n7160 | n7161 ;
  assign n7164 = ( x113 & ~n7163 ) | ( x113 & n7162 ) | ( ~n7163 & n7162 ) ;
  assign n7165 = ~n200 & n6420 ;
  assign n7166 = n7164 | n7165 ;
  assign n7167 = ( x5 & ~n7166 ) | ( x5 & 1'b0 ) | ( ~n7166 & 1'b0 ) ;
  assign n7168 = ~x5 & n7166 ;
  assign n7169 = n7167 | n7168 ;
  assign n7382 = x110 &  n353 ;
  assign n7379 = ( x112 & ~n313 ) | ( x112 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n7380 = x111 &  n308 ;
  assign n7381 = n7379 | n7380 ;
  assign n7383 = ( x110 & ~n7382 ) | ( x110 & n7381 ) | ( ~n7382 & n7381 ) ;
  assign n7384 = ~n316 & n5727 ;
  assign n7385 = n7383 | n7384 ;
  assign n7386 = ( x8 & ~n7385 ) | ( x8 & 1'b0 ) | ( ~n7385 & 1'b0 ) ;
  assign n7387 = ~x8 & n7385 ;
  assign n7388 = n7386 | n7387 ;
  assign n7173 = x107 &  n503 ;
  assign n7170 = ( x109 & ~n450 ) | ( x109 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n7171 = x108 &  n445 ;
  assign n7172 = n7170 | n7171 ;
  assign n7174 = ( x107 & ~n7173 ) | ( x107 & n7172 ) | ( ~n7173 & n7172 ) ;
  assign n7175 = ~n453 & n5267 ;
  assign n7176 = n7174 | n7175 ;
  assign n7177 = ( x11 & ~n7176 ) | ( x11 & 1'b0 ) | ( ~n7176 & 1'b0 ) ;
  assign n7178 = ~x11 & n7176 ;
  assign n7179 = n7177 | n7178 ;
  assign n7180 = ( n7097 & ~n7108 ) | ( n7097 & n7098 ) | ( ~n7108 & n7098 ) ;
  assign n7181 = ( n6915 & n6925 ) | ( n6915 & n7091 ) | ( n6925 & n7091 ) ;
  assign n7185 = x101 &  n942 ;
  assign n7182 = ( x103 & ~n896 ) | ( x103 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n7183 = x102 &  n891 ;
  assign n7184 = n7182 | n7183 ;
  assign n7186 = ( x101 & ~n7185 ) | ( x101 & n7184 ) | ( ~n7185 & n7184 ) ;
  assign n7187 = n899 | n4056 ;
  assign n7188 = ~n7186 & n7187 ;
  assign n7189 = x17 &  n7188 ;
  assign n7190 = x17 | n7188 ;
  assign n7191 = ~n7189 & n7190 ;
  assign n7195 = x92 &  n1894 ;
  assign n7192 = ( x94 & ~n1816 ) | ( x94 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n7193 = x93 &  n1811 ;
  assign n7194 = n7192 | n7193 ;
  assign n7196 = ( x92 & ~n7195 ) | ( x92 & n7194 ) | ( ~n7195 & n7194 ) ;
  assign n7197 = ~n1819 & n2401 ;
  assign n7198 = n7196 | n7197 ;
  assign n7199 = ( x26 & ~n7198 ) | ( x26 & 1'b0 ) | ( ~n7198 & 1'b0 ) ;
  assign n7200 = ~x26 & n7198 ;
  assign n7201 = n7199 | n7200 ;
  assign n7205 = x89 &  n2312 ;
  assign n7202 = ( x91 & ~n2195 ) | ( x91 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n7203 = x90 &  n2190 ;
  assign n7204 = n7202 | n7203 ;
  assign n7206 = ( x89 & ~n7205 ) | ( x89 & n7204 ) | ( ~n7205 & n7204 ) ;
  assign n7207 = ( n2108 & ~n2198 ) | ( n2108 & 1'b0 ) | ( ~n2198 & 1'b0 ) ;
  assign n7208 = n7206 | n7207 ;
  assign n7209 = ( x29 & ~n7208 ) | ( x29 & 1'b0 ) | ( ~n7208 & 1'b0 ) ;
  assign n7210 = ~x29 & n7208 ;
  assign n7211 = n7209 | n7210 ;
  assign n7212 = ( n7058 & n7059 ) | ( n7058 & n7069 ) | ( n7059 & n7069 ) ;
  assign n7216 = x86 &  n2718 ;
  assign n7213 = ( x88 & ~n2642 ) | ( x88 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n7214 = x87 &  n2637 ;
  assign n7215 = n7213 | n7214 ;
  assign n7217 = ( x86 & ~n7216 ) | ( x86 & n7215 ) | ( ~n7216 & n7215 ) ;
  assign n7218 = ( n1624 & ~n2645 ) | ( n1624 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n7219 = n7217 | n7218 ;
  assign n7220 = ( x32 & ~n7219 ) | ( x32 & 1'b0 ) | ( ~n7219 & 1'b0 ) ;
  assign n7221 = ~x32 & n7219 ;
  assign n7222 = n7220 | n7221 ;
  assign n7226 = x83 &  n3214 ;
  assign n7223 = ( x85 & ~n3087 ) | ( x85 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n7224 = x84 &  n3082 ;
  assign n7225 = n7223 | n7224 ;
  assign n7227 = ( x83 & ~n7226 ) | ( x83 & n7225 ) | ( ~n7226 & n7225 ) ;
  assign n7228 = ( n1295 & ~n3090 ) | ( n1295 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n7229 = n7227 | n7228 ;
  assign n7230 = ( x35 & ~n7229 ) | ( x35 & 1'b0 ) | ( ~n7229 & 1'b0 ) ;
  assign n7231 = ~x35 & n7229 ;
  assign n7232 = n7230 | n7231 ;
  assign n7233 = ( n7041 & n7042 ) | ( n7041 & n7052 ) | ( n7042 & n7052 ) ;
  assign n7237 = x80 &  n3756 ;
  assign n7234 = ( x82 & ~n3602 ) | ( x82 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n7235 = x81 &  n3597 ;
  assign n7236 = n7234 | n7235 ;
  assign n7238 = ( x80 & ~n7237 ) | ( x80 & n7236 ) | ( ~n7237 & n7236 ) ;
  assign n7239 = ( n1084 & ~n3605 ) | ( n1084 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n7240 = n7238 | n7239 ;
  assign n7241 = ( x38 & ~n7240 ) | ( x38 & 1'b0 ) | ( ~n7240 & 1'b0 ) ;
  assign n7242 = ~x38 & n7240 ;
  assign n7243 = n7241 | n7242 ;
  assign n7247 = x77 &  n4344 ;
  assign n7244 = ( x79 & ~n4143 ) | ( x79 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n7245 = x78 &  n4138 ;
  assign n7246 = n7244 | n7245 ;
  assign n7248 = ( x77 & ~n7247 ) | ( x77 & n7246 ) | ( ~n7247 & n7246 ) ;
  assign n7249 = ( n766 & ~n4146 ) | ( n766 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n7250 = n7248 | n7249 ;
  assign n7251 = ( x41 & ~n7250 ) | ( x41 & 1'b0 ) | ( ~n7250 & 1'b0 ) ;
  assign n7252 = ~x41 & n7250 ;
  assign n7253 = n7251 | n7252 ;
  assign n7257 = x74 &  n4934 ;
  assign n7254 = ( x76 & ~n4725 ) | ( x76 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n7255 = x75 &  n4720 ;
  assign n7256 = n7254 | n7255 ;
  assign n7258 = ( x74 & ~n7257 ) | ( x74 & n7256 ) | ( ~n7257 & n7256 ) ;
  assign n7259 = ( n603 & ~n4728 ) | ( n603 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n7260 = n7258 | n7259 ;
  assign n7261 = ( x44 & ~n7260 ) | ( x44 & 1'b0 ) | ( ~n7260 & 1'b0 ) ;
  assign n7262 = ~x44 & n7260 ;
  assign n7263 = n7261 | n7262 ;
  assign n7267 = x71 &  n5586 ;
  assign n7264 = ( x73 & ~n5389 ) | ( x73 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n7265 = x72 &  n5384 ;
  assign n7266 = n7264 | n7265 ;
  assign n7268 = ( x71 & ~n7267 ) | ( x71 & n7266 ) | ( ~n7267 & n7266 ) ;
  assign n7269 = ( n389 & ~n5392 ) | ( n389 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n7270 = n7268 | n7269 ;
  assign n7271 = ( x47 & ~n7270 ) | ( x47 & 1'b0 ) | ( ~n7270 & 1'b0 ) ;
  assign n7272 = ~x47 & n7270 ;
  assign n7273 = n7271 | n7272 ;
  assign n7274 = ( n7007 & n7008 ) | ( n7007 & n7018 ) | ( n7008 & n7018 ) ;
  assign n7275 = ( x53 & ~x54 ) | ( x53 & 1'b0 ) | ( ~x54 & 1'b0 ) ;
  assign n7276 = ~x53 & x54 ;
  assign n7277 = n7275 | n7276 ;
  assign n7278 = x64 &  n7277 ;
  assign n7279 = ( n6521 & ~n6732 ) | ( n6521 & n6989 ) | ( ~n6732 & n6989 ) ;
  assign n7280 = ( x53 & n6732 ) | ( x53 & n7279 ) | ( n6732 & n7279 ) ;
  assign n7281 = ( x53 & ~n7280 ) | ( x53 & 1'b0 ) | ( ~n7280 & 1'b0 ) ;
  assign n7285 = x65 &  n6982 ;
  assign n7282 = ( x67 & ~n6727 ) | ( x67 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n7283 = x66 &  n6722 ;
  assign n7284 = n7282 | n7283 ;
  assign n7286 = ( x65 & ~n7285 ) | ( x65 & n7284 ) | ( ~n7285 & n7284 ) ;
  assign n7287 = n173 | n6730 ;
  assign n7288 = ~n7286 & n7287 ;
  assign n7289 = x53 &  n7288 ;
  assign n7290 = x53 | n7288 ;
  assign n7291 = ~n7289 & n7290 ;
  assign n7292 = ( n7278 & ~n7281 ) | ( n7278 & n7291 ) | ( ~n7281 & n7291 ) ;
  assign n7293 = ( n7278 & ~n7291 ) | ( n7278 & n7281 ) | ( ~n7291 & n7281 ) ;
  assign n7294 = ( n7292 & ~n7278 ) | ( n7292 & n7293 ) | ( ~n7278 & n7293 ) ;
  assign n7295 = ( n6737 & n6994 ) | ( n6737 & n7004 ) | ( n6994 & n7004 ) ;
  assign n7299 = x68 &  n6288 ;
  assign n7296 = ( x70 & ~n6032 ) | ( x70 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n7297 = x69 &  n6027 ;
  assign n7298 = n7296 | n7297 ;
  assign n7300 = ( x68 & ~n7299 ) | ( x68 & n7298 ) | ( ~n7299 & n7298 ) ;
  assign n7301 = ( n282 & ~n6035 ) | ( n282 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n7302 = n7300 | n7301 ;
  assign n7303 = ( x50 & ~n7302 ) | ( x50 & 1'b0 ) | ( ~n7302 & 1'b0 ) ;
  assign n7304 = ~x50 & n7302 ;
  assign n7305 = n7303 | n7304 ;
  assign n7306 = ( n7294 & ~n7295 ) | ( n7294 & n7305 ) | ( ~n7295 & n7305 ) ;
  assign n7307 = ( n7295 & ~n7294 ) | ( n7295 & n7305 ) | ( ~n7294 & n7305 ) ;
  assign n7308 = ( n7306 & ~n7305 ) | ( n7306 & n7307 ) | ( ~n7305 & n7307 ) ;
  assign n7309 = ( n7273 & ~n7274 ) | ( n7273 & n7308 ) | ( ~n7274 & n7308 ) ;
  assign n7310 = ( n7273 & ~n7308 ) | ( n7273 & n7274 ) | ( ~n7308 & n7274 ) ;
  assign n7311 = ( n7309 & ~n7273 ) | ( n7309 & n7310 ) | ( ~n7273 & n7310 ) ;
  assign n7312 = ( n7263 & ~n7023 ) | ( n7263 & n7311 ) | ( ~n7023 & n7311 ) ;
  assign n7313 = ( n7023 & ~n7311 ) | ( n7023 & n7263 ) | ( ~n7311 & n7263 ) ;
  assign n7314 = ( n7312 & ~n7263 ) | ( n7312 & n7313 ) | ( ~n7263 & n7313 ) ;
  assign n7315 = ( n7253 & ~n7037 ) | ( n7253 & n7314 ) | ( ~n7037 & n7314 ) ;
  assign n7316 = ( n7037 & ~n7314 ) | ( n7037 & n7253 ) | ( ~n7314 & n7253 ) ;
  assign n7317 = ( n7315 & ~n7253 ) | ( n7315 & n7316 ) | ( ~n7253 & n7316 ) ;
  assign n7318 = ( n7243 & ~n7040 ) | ( n7243 & n7317 ) | ( ~n7040 & n7317 ) ;
  assign n7319 = ( n7040 & ~n7317 ) | ( n7040 & n7243 ) | ( ~n7317 & n7243 ) ;
  assign n7320 = ( n7318 & ~n7243 ) | ( n7318 & n7319 ) | ( ~n7243 & n7319 ) ;
  assign n7321 = ( n7232 & ~n7233 ) | ( n7232 & n7320 ) | ( ~n7233 & n7320 ) ;
  assign n7322 = ( n7232 & ~n7320 ) | ( n7232 & n7233 ) | ( ~n7320 & n7233 ) ;
  assign n7323 = ( n7321 & ~n7232 ) | ( n7321 & n7322 ) | ( ~n7232 & n7322 ) ;
  assign n7324 = ( n7222 & ~n7057 ) | ( n7222 & n7323 ) | ( ~n7057 & n7323 ) ;
  assign n7325 = ( n7057 & ~n7323 ) | ( n7057 & n7222 ) | ( ~n7323 & n7222 ) ;
  assign n7326 = ( n7324 & ~n7222 ) | ( n7324 & n7325 ) | ( ~n7222 & n7325 ) ;
  assign n7327 = ( n7211 & ~n7212 ) | ( n7211 & n7326 ) | ( ~n7212 & n7326 ) ;
  assign n7328 = ( n7211 & ~n7326 ) | ( n7211 & n7212 ) | ( ~n7326 & n7212 ) ;
  assign n7329 = ( n7327 & ~n7211 ) | ( n7327 & n7328 ) | ( ~n7211 & n7328 ) ;
  assign n7330 = ( n7201 & ~n7074 ) | ( n7201 & n7329 ) | ( ~n7074 & n7329 ) ;
  assign n7331 = ( n7074 & ~n7329 ) | ( n7074 & n7201 ) | ( ~n7329 & n7201 ) ;
  assign n7332 = ( n7330 & ~n7201 ) | ( n7330 & n7331 ) | ( ~n7201 & n7331 ) ;
  assign n7336 = x95 &  n1551 ;
  assign n7333 = ( x97 & ~n1451 ) | ( x97 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n7334 = x96 &  n1446 ;
  assign n7335 = n7333 | n7334 ;
  assign n7337 = ( x95 & ~n7336 ) | ( x95 & n7335 ) | ( ~n7336 & n7335 ) ;
  assign n7338 = ~n1454 & n2999 ;
  assign n7339 = n7337 | n7338 ;
  assign n7340 = ( x23 & ~n7339 ) | ( x23 & 1'b0 ) | ( ~n7339 & 1'b0 ) ;
  assign n7341 = ~x23 & n7339 ;
  assign n7342 = n7340 | n7341 ;
  assign n7343 = ( n7332 & ~n7077 ) | ( n7332 & n7342 ) | ( ~n7077 & n7342 ) ;
  assign n7344 = ( n7077 & ~n7342 ) | ( n7077 & n7332 ) | ( ~n7342 & n7332 ) ;
  assign n7345 = ( n7343 & ~n7332 ) | ( n7343 & n7344 ) | ( ~n7332 & n7344 ) ;
  assign n7346 = ( n6840 & ~n7078 ) | ( n6840 & n7088 ) | ( ~n7078 & n7088 ) ;
  assign n7350 = x98 &  n1227 ;
  assign n7347 = ( x100 & ~n1154 ) | ( x100 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n7348 = x99 &  n1149 ;
  assign n7349 = n7347 | n7348 ;
  assign n7351 = ( x98 & ~n7350 ) | ( x98 & n7349 ) | ( ~n7350 & n7349 ) ;
  assign n7352 = n1157 | n3354 ;
  assign n7353 = ~n7351 & n7352 ;
  assign n7354 = x20 &  n7353 ;
  assign n7355 = x20 | n7353 ;
  assign n7356 = ~n7354 & n7355 ;
  assign n7357 = ( n7345 & n7346 ) | ( n7345 & n7356 ) | ( n7346 & n7356 ) ;
  assign n7358 = ( n7346 & ~n7345 ) | ( n7346 & n7356 ) | ( ~n7345 & n7356 ) ;
  assign n7359 = ( n7345 & ~n7357 ) | ( n7345 & n7358 ) | ( ~n7357 & n7358 ) ;
  assign n7360 = ( n7181 & n7191 ) | ( n7181 & n7359 ) | ( n7191 & n7359 ) ;
  assign n7361 = ( n7191 & ~n7181 ) | ( n7191 & n7359 ) | ( ~n7181 & n7359 ) ;
  assign n7362 = ( n7181 & ~n7360 ) | ( n7181 & n7361 ) | ( ~n7360 & n7361 ) ;
  assign n7366 = x104 &  n713 ;
  assign n7363 = ( x106 & ~n641 ) | ( x106 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n7364 = x105 &  n636 ;
  assign n7365 = n7363 | n7364 ;
  assign n7367 = ( x104 & ~n7366 ) | ( x104 & n7365 ) | ( ~n7366 & n7365 ) ;
  assign n7368 = ~n644 & n4458 ;
  assign n7369 = n7367 | n7368 ;
  assign n7370 = ( x14 & ~n7369 ) | ( x14 & 1'b0 ) | ( ~n7369 & 1'b0 ) ;
  assign n7371 = ~x14 & n7369 ;
  assign n7372 = n7370 | n7371 ;
  assign n7374 = ( n7095 & n7362 ) | ( n7095 & n7372 ) | ( n7362 & n7372 ) ;
  assign n7373 = ( n7095 & ~n7362 ) | ( n7095 & n7372 ) | ( ~n7362 & n7372 ) ;
  assign n7375 = ( n7362 & ~n7374 ) | ( n7362 & n7373 ) | ( ~n7374 & n7373 ) ;
  assign n7376 = ( n7179 & ~n7180 ) | ( n7179 & n7375 ) | ( ~n7180 & n7375 ) ;
  assign n7377 = ( n7179 & ~n7375 ) | ( n7179 & n7180 ) | ( ~n7375 & n7180 ) ;
  assign n7378 = ( n7376 & ~n7179 ) | ( n7376 & n7377 ) | ( ~n7179 & n7377 ) ;
  assign n7389 = ( n7122 & ~n7388 ) | ( n7122 & n7378 ) | ( ~n7388 & n7378 ) ;
  assign n7390 = ( n7122 & ~n7378 ) | ( n7122 & n7388 ) | ( ~n7378 & n7388 ) ;
  assign n7391 = ( n7389 & ~n7122 ) | ( n7389 & n7390 ) | ( ~n7122 & n7390 ) ;
  assign n7392 = ( n7159 & ~n7169 ) | ( n7159 & n7391 ) | ( ~n7169 & n7391 ) ;
  assign n7393 = ( n7159 & ~n7391 ) | ( n7159 & n7169 ) | ( ~n7391 & n7169 ) ;
  assign n7394 = ( n7392 & ~n7159 ) | ( n7392 & n7393 ) | ( ~n7159 & n7393 ) ;
  assign n7396 = ( n7157 & n7158 ) | ( n7157 & n7394 ) | ( n7158 & n7394 ) ;
  assign n7395 = ( n7158 & ~n7157 ) | ( n7158 & n7394 ) | ( ~n7157 & n7394 ) ;
  assign n7397 = ( n7157 & ~n7396 ) | ( n7157 & n7395 ) | ( ~n7396 & n7395 ) ;
  assign n7398 = ( n7169 & ~n7159 ) | ( n7169 & n7391 ) | ( ~n7159 & n7391 ) ;
  assign n7402 = x114 &  n225 ;
  assign n7399 = ( x116 & ~n197 ) | ( x116 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n7400 = x115 &  n192 ;
  assign n7401 = n7399 | n7400 ;
  assign n7403 = ( x114 & ~n7402 ) | ( x114 & n7401 ) | ( ~n7402 & n7401 ) ;
  assign n7404 = n200 | n6885 ;
  assign n7405 = ~n7403 & n7404 ;
  assign n7406 = x5 &  n7405 ;
  assign n7407 = x5 | n7405 ;
  assign n7408 = ~n7406 & n7407 ;
  assign n7419 = ( n7181 & ~n7359 ) | ( n7181 & n7191 ) | ( ~n7359 & n7191 ) ;
  assign n7423 = x102 &  n942 ;
  assign n7420 = ( x104 & ~n896 ) | ( x104 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n7421 = x103 &  n891 ;
  assign n7422 = n7420 | n7421 ;
  assign n7424 = ( x102 & ~n7423 ) | ( x102 & n7422 ) | ( ~n7423 & n7422 ) ;
  assign n7425 = n899 | n4249 ;
  assign n7426 = ~n7424 & n7425 ;
  assign n7427 = x17 &  n7426 ;
  assign n7428 = x17 | n7426 ;
  assign n7429 = ~n7427 & n7428 ;
  assign n7433 = x99 &  n1227 ;
  assign n7430 = ( x101 & ~n1154 ) | ( x101 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n7431 = x100 &  n1149 ;
  assign n7432 = n7430 | n7431 ;
  assign n7434 = ( x99 & ~n7433 ) | ( x99 & n7432 ) | ( ~n7433 & n7432 ) ;
  assign n7435 = n1157 | n3694 ;
  assign n7436 = ~n7434 & n7435 ;
  assign n7437 = x20 &  n7436 ;
  assign n7438 = x20 | n7436 ;
  assign n7439 = ~n7437 & n7438 ;
  assign n7443 = x96 &  n1551 ;
  assign n7440 = ( x98 & ~n1451 ) | ( x98 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n7441 = x97 &  n1446 ;
  assign n7442 = n7440 | n7441 ;
  assign n7444 = ( x96 & ~n7443 ) | ( x96 & n7442 ) | ( ~n7443 & n7442 ) ;
  assign n7445 = ~n1454 & n3170 ;
  assign n7446 = n7444 | n7445 ;
  assign n7447 = ( x23 & ~n7446 ) | ( x23 & 1'b0 ) | ( ~n7446 & 1'b0 ) ;
  assign n7448 = ~x23 & n7446 ;
  assign n7449 = n7447 | n7448 ;
  assign n7453 = x93 &  n1894 ;
  assign n7450 = ( x95 & ~n1816 ) | ( x95 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n7451 = x94 &  n1811 ;
  assign n7452 = n7450 | n7451 ;
  assign n7454 = ( x93 & ~n7453 ) | ( x93 & n7452 ) | ( ~n7453 & n7452 ) ;
  assign n7455 = ~n1819 & n2547 ;
  assign n7456 = n7454 | n7455 ;
  assign n7457 = ( x26 & ~n7456 ) | ( x26 & 1'b0 ) | ( ~n7456 & 1'b0 ) ;
  assign n7458 = ~x26 & n7456 ;
  assign n7459 = n7457 | n7458 ;
  assign n7463 = x90 &  n2312 ;
  assign n7460 = ( x92 & ~n2195 ) | ( x92 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n7461 = x91 &  n2190 ;
  assign n7462 = n7460 | n7461 ;
  assign n7464 = ( x90 & ~n7463 ) | ( x90 & n7462 ) | ( ~n7463 & n7462 ) ;
  assign n7465 = ~n2198 & n2248 ;
  assign n7466 = n7464 | n7465 ;
  assign n7467 = ( x29 & ~n7466 ) | ( x29 & 1'b0 ) | ( ~n7466 & 1'b0 ) ;
  assign n7468 = ~x29 & n7466 ;
  assign n7469 = n7467 | n7468 ;
  assign n7473 = x87 &  n2718 ;
  assign n7470 = ( x89 & ~n2642 ) | ( x89 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n7471 = x88 &  n2637 ;
  assign n7472 = n7470 | n7471 ;
  assign n7474 = ( x87 & ~n7473 ) | ( x87 & n7472 ) | ( ~n7473 & n7472 ) ;
  assign n7475 = ( n1741 & ~n2645 ) | ( n1741 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n7476 = n7474 | n7475 ;
  assign n7477 = ( x32 & ~n7476 ) | ( x32 & 1'b0 ) | ( ~n7476 & 1'b0 ) ;
  assign n7478 = ~x32 & n7476 ;
  assign n7479 = n7477 | n7478 ;
  assign n7575 = x81 &  n3756 ;
  assign n7572 = ( x83 & ~n3602 ) | ( x83 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n7573 = x82 &  n3597 ;
  assign n7574 = n7572 | n7573 ;
  assign n7576 = ( x81 & ~n7575 ) | ( x81 & n7574 ) | ( ~n7575 & n7574 ) ;
  assign n7577 = ( n1100 & ~n3605 ) | ( n1100 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n7578 = n7576 | n7577 ;
  assign n7579 = ( x38 & ~n7578 ) | ( x38 & 1'b0 ) | ( ~n7578 & 1'b0 ) ;
  assign n7580 = ~x38 & n7578 ;
  assign n7581 = n7579 | n7580 ;
  assign n7493 = x75 &  n4934 ;
  assign n7490 = ( x77 & ~n4725 ) | ( x77 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n7491 = x76 &  n4720 ;
  assign n7492 = n7490 | n7491 ;
  assign n7494 = ( x75 & ~n7493 ) | ( x75 & n7492 ) | ( ~n7493 & n7492 ) ;
  assign n7495 = ( n677 & ~n4728 ) | ( n677 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n7496 = n7494 | n7495 ;
  assign n7497 = ( x44 & ~n7496 ) | ( x44 & 1'b0 ) | ( ~n7496 & 1'b0 ) ;
  assign n7498 = ~x44 & n7496 ;
  assign n7499 = n7497 | n7498 ;
  assign n7503 = x72 &  n5586 ;
  assign n7500 = ( x74 & ~n5389 ) | ( x74 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n7501 = x73 &  n5384 ;
  assign n7502 = n7500 | n7501 ;
  assign n7504 = ( x72 & ~n7503 ) | ( x72 & n7502 ) | ( ~n7503 & n7502 ) ;
  assign n7505 = ( n482 & ~n5392 ) | ( n482 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n7506 = n7504 | n7505 ;
  assign n7507 = ( x47 & ~n7506 ) | ( x47 & 1'b0 ) | ( ~n7506 & 1'b0 ) ;
  assign n7508 = ~x47 & n7506 ;
  assign n7509 = n7507 | n7508 ;
  assign n7513 = x69 &  n6288 ;
  assign n7510 = ( x71 & ~n6032 ) | ( x71 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n7511 = x70 &  n6027 ;
  assign n7512 = n7510 | n7511 ;
  assign n7514 = ( x69 & ~n7513 ) | ( x69 & n7512 ) | ( ~n7513 & n7512 ) ;
  assign n7515 = ( n298 & ~n6035 ) | ( n298 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n7516 = n7514 | n7515 ;
  assign n7517 = ( x50 & ~n7516 ) | ( x50 & 1'b0 ) | ( ~n7516 & 1'b0 ) ;
  assign n7518 = ~x50 & n7516 ;
  assign n7519 = n7517 | n7518 ;
  assign n7523 = x66 &  n6982 ;
  assign n7520 = ( x68 & ~n6727 ) | ( x68 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n7521 = x67 &  n6722 ;
  assign n7522 = n7520 | n7521 ;
  assign n7524 = ( x66 & ~n7523 ) | ( x66 & n7522 ) | ( ~n7523 & n7522 ) ;
  assign n7525 = ( n213 & ~n6730 ) | ( n213 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n7526 = n7524 | n7525 ;
  assign n7527 = ( x53 & ~n7526 ) | ( x53 & 1'b0 ) | ( ~n7526 & 1'b0 ) ;
  assign n7528 = ~x53 & n7526 ;
  assign n7529 = n7527 | n7528 ;
  assign n7530 = ( x56 & ~n7278 ) | ( x56 & 1'b0 ) | ( ~n7278 & 1'b0 ) ;
  assign n7531 = ( x54 & x55 ) | ( x54 & n7275 ) | ( x55 & n7275 ) ;
  assign n7532 = ( x54 & ~n7276 ) | ( x54 & x55 ) | ( ~n7276 & x55 ) ;
  assign n7533 = ~n7531 &  n7532 ;
  assign n7534 = x64 &  n7533 ;
  assign n7535 = ~x55 & x56 ;
  assign n7536 = ( x55 & ~x56 ) | ( x55 & 1'b0 ) | ( ~x56 & 1'b0 ) ;
  assign n7537 = n7535 | n7536 ;
  assign n7538 = ~n7277 |  n7537 ;
  assign n7539 = ( x65 & ~n7538 ) | ( x65 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n7540 = n7534 | n7539 ;
  assign n7541 = ~n7277 | ~n7537 ;
  assign n7542 = ( n142 & ~n7541 ) | ( n142 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n7543 = n7540 | n7542 ;
  assign n7545 = ( x56 & n7530 ) | ( x56 & n7543 ) | ( n7530 & n7543 ) ;
  assign n7544 = ( x56 & ~n7530 ) | ( x56 & n7543 ) | ( ~n7530 & n7543 ) ;
  assign n7546 = ( n7530 & ~n7545 ) | ( n7530 & n7544 ) | ( ~n7545 & n7544 ) ;
  assign n7548 = ( n7293 & n7529 ) | ( n7293 & n7546 ) | ( n7529 & n7546 ) ;
  assign n7547 = ( n7293 & ~n7529 ) | ( n7293 & n7546 ) | ( ~n7529 & n7546 ) ;
  assign n7549 = ( n7529 & ~n7548 ) | ( n7529 & n7547 ) | ( ~n7548 & n7547 ) ;
  assign n7551 = ( n7307 & n7519 ) | ( n7307 & n7549 ) | ( n7519 & n7549 ) ;
  assign n7550 = ( n7307 & ~n7519 ) | ( n7307 & n7549 ) | ( ~n7519 & n7549 ) ;
  assign n7552 = ( n7519 & ~n7551 ) | ( n7519 & n7550 ) | ( ~n7551 & n7550 ) ;
  assign n7554 = ( n7310 & n7509 ) | ( n7310 & n7552 ) | ( n7509 & n7552 ) ;
  assign n7553 = ( n7310 & ~n7509 ) | ( n7310 & n7552 ) | ( ~n7509 & n7552 ) ;
  assign n7555 = ( n7509 & ~n7554 ) | ( n7509 & n7553 ) | ( ~n7554 & n7553 ) ;
  assign n7557 = ( n7313 & n7499 ) | ( n7313 & n7555 ) | ( n7499 & n7555 ) ;
  assign n7556 = ( n7313 & ~n7499 ) | ( n7313 & n7555 ) | ( ~n7499 & n7555 ) ;
  assign n7558 = ( n7499 & ~n7557 ) | ( n7499 & n7556 ) | ( ~n7557 & n7556 ) ;
  assign n7562 = x78 &  n4344 ;
  assign n7559 = ( x80 & ~n4143 ) | ( x80 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n7560 = x79 &  n4138 ;
  assign n7561 = n7559 | n7560 ;
  assign n7563 = ( x78 & ~n7562 ) | ( x78 & n7561 ) | ( ~n7562 & n7561 ) ;
  assign n7564 = ( n842 & ~n4146 ) | ( n842 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n7565 = n7563 | n7564 ;
  assign n7566 = ( x41 & ~n7565 ) | ( x41 & 1'b0 ) | ( ~n7565 & 1'b0 ) ;
  assign n7567 = ~x41 & n7565 ;
  assign n7568 = n7566 | n7567 ;
  assign n7569 = ( n7558 & ~n7316 ) | ( n7558 & n7568 ) | ( ~n7316 & n7568 ) ;
  assign n7570 = ( n7316 & ~n7568 ) | ( n7316 & n7558 ) | ( ~n7568 & n7558 ) ;
  assign n7571 = ( n7569 & ~n7558 ) | ( n7569 & n7570 ) | ( ~n7558 & n7570 ) ;
  assign n7582 = ( n7319 & ~n7581 ) | ( n7319 & n7571 ) | ( ~n7581 & n7571 ) ;
  assign n7583 = ( n7571 & ~n7319 ) | ( n7571 & n7581 ) | ( ~n7319 & n7581 ) ;
  assign n7584 = ( n7582 & ~n7571 ) | ( n7582 & n7583 ) | ( ~n7571 & n7583 ) ;
  assign n7483 = x84 &  n3214 ;
  assign n7480 = ( x86 & ~n3087 ) | ( x86 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n7481 = x85 &  n3082 ;
  assign n7482 = n7480 | n7481 ;
  assign n7484 = ( x84 & ~n7483 ) | ( x84 & n7482 ) | ( ~n7483 & n7482 ) ;
  assign n7485 = ( n1496 & ~n3090 ) | ( n1496 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n7486 = n7484 | n7485 ;
  assign n7487 = ( x35 & ~n7486 ) | ( x35 & 1'b0 ) | ( ~n7486 & 1'b0 ) ;
  assign n7488 = ~x35 & n7486 ;
  assign n7489 = n7487 | n7488 ;
  assign n7585 = ( n7322 & ~n7584 ) | ( n7322 & n7489 ) | ( ~n7584 & n7489 ) ;
  assign n7586 = ( n7489 & ~n7322 ) | ( n7489 & n7584 ) | ( ~n7322 & n7584 ) ;
  assign n7587 = ( n7585 & ~n7489 ) | ( n7585 & n7586 ) | ( ~n7489 & n7586 ) ;
  assign n7588 = ( n7325 & n7479 ) | ( n7325 & n7587 ) | ( n7479 & n7587 ) ;
  assign n7589 = ( n7325 & ~n7479 ) | ( n7325 & n7587 ) | ( ~n7479 & n7587 ) ;
  assign n7590 = ( n7479 & ~n7588 ) | ( n7479 & n7589 ) | ( ~n7588 & n7589 ) ;
  assign n7591 = ( n7328 & n7469 ) | ( n7328 & n7590 ) | ( n7469 & n7590 ) ;
  assign n7592 = ( n7328 & ~n7469 ) | ( n7328 & n7590 ) | ( ~n7469 & n7590 ) ;
  assign n7593 = ( n7469 & ~n7591 ) | ( n7469 & n7592 ) | ( ~n7591 & n7592 ) ;
  assign n7594 = ( n7331 & n7459 ) | ( n7331 & n7593 ) | ( n7459 & n7593 ) ;
  assign n7595 = ( n7331 & ~n7459 ) | ( n7331 & n7593 ) | ( ~n7459 & n7593 ) ;
  assign n7596 = ( n7459 & ~n7594 ) | ( n7459 & n7595 ) | ( ~n7594 & n7595 ) ;
  assign n7597 = ( n7077 & ~n7332 ) | ( n7077 & n7342 ) | ( ~n7332 & n7342 ) ;
  assign n7598 = ( n7449 & n7596 ) | ( n7449 & n7597 ) | ( n7596 & n7597 ) ;
  assign n7599 = ( n7596 & ~n7449 ) | ( n7596 & n7597 ) | ( ~n7449 & n7597 ) ;
  assign n7600 = ( n7449 & ~n7598 ) | ( n7449 & n7599 ) | ( ~n7598 & n7599 ) ;
  assign n7601 = ( n7345 & ~n7346 ) | ( n7345 & n7356 ) | ( ~n7346 & n7356 ) ;
  assign n7602 = ( n7439 & ~n7600 ) | ( n7439 & n7601 ) | ( ~n7600 & n7601 ) ;
  assign n7603 = ( n7439 & ~n7601 ) | ( n7439 & n7600 ) | ( ~n7601 & n7600 ) ;
  assign n7604 = ( n7602 & ~n7439 ) | ( n7602 & n7603 ) | ( ~n7439 & n7603 ) ;
  assign n7605 = ( n7419 & n7429 ) | ( n7419 & n7604 ) | ( n7429 & n7604 ) ;
  assign n7606 = ( n7429 & ~n7419 ) | ( n7429 & n7604 ) | ( ~n7419 & n7604 ) ;
  assign n7607 = ( n7419 & ~n7605 ) | ( n7419 & n7606 ) | ( ~n7605 & n7606 ) ;
  assign n7612 = x105 &  n713 ;
  assign n7609 = ( x107 & ~n641 ) | ( x107 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n7610 = x106 &  n636 ;
  assign n7611 = n7609 | n7610 ;
  assign n7613 = ( x105 & ~n7612 ) | ( x105 & n7611 ) | ( ~n7612 & n7611 ) ;
  assign n7614 = ~n644 & n4848 ;
  assign n7615 = n7613 | n7614 ;
  assign n7616 = ( x14 & ~n7615 ) | ( x14 & 1'b0 ) | ( ~n7615 & 1'b0 ) ;
  assign n7617 = ~x14 & n7615 ;
  assign n7618 = n7616 | n7617 ;
  assign n7608 = ( n7362 & ~n7095 ) | ( n7362 & n7372 ) | ( ~n7095 & n7372 ) ;
  assign n7619 = ( n7607 & ~n7618 ) | ( n7607 & n7608 ) | ( ~n7618 & n7608 ) ;
  assign n7620 = ( n7607 & ~n7608 ) | ( n7607 & n7618 ) | ( ~n7608 & n7618 ) ;
  assign n7621 = ( n7619 & ~n7607 ) | ( n7619 & n7620 ) | ( ~n7607 & n7620 ) ;
  assign n7625 = x108 &  n503 ;
  assign n7622 = ( x110 & ~n450 ) | ( x110 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n7623 = x109 &  n445 ;
  assign n7624 = n7622 | n7623 ;
  assign n7626 = ( x108 & ~n7625 ) | ( x108 & n7624 ) | ( ~n7625 & n7624 ) ;
  assign n7627 = n453 | n5283 ;
  assign n7628 = ~n7626 & n7627 ;
  assign n7629 = x11 &  n7628 ;
  assign n7630 = x11 | n7628 ;
  assign n7631 = ~n7629 & n7630 ;
  assign n7633 = ( n7377 & n7621 ) | ( n7377 & n7631 ) | ( n7621 & n7631 ) ;
  assign n7632 = ( n7377 & ~n7621 ) | ( n7377 & n7631 ) | ( ~n7621 & n7631 ) ;
  assign n7634 = ( n7621 & ~n7633 ) | ( n7621 & n7632 ) | ( ~n7633 & n7632 ) ;
  assign n7412 = x111 &  n353 ;
  assign n7409 = ( x113 & ~n313 ) | ( x113 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n7410 = x112 &  n308 ;
  assign n7411 = n7409 | n7410 ;
  assign n7413 = ( x111 & ~n7412 ) | ( x111 & n7411 ) | ( ~n7412 & n7411 ) ;
  assign n7414 = n316 | n6169 ;
  assign n7415 = ~n7413 & n7414 ;
  assign n7416 = x8 &  n7415 ;
  assign n7417 = x8 | n7415 ;
  assign n7418 = ~n7416 & n7417 ;
  assign n7635 = ( n7389 & n7418 ) | ( n7389 & n7634 ) | ( n7418 & n7634 ) ;
  assign n7636 = ( n7389 & ~n7634 ) | ( n7389 & n7418 ) | ( ~n7634 & n7418 ) ;
  assign n7637 = ( n7634 & ~n7635 ) | ( n7634 & n7636 ) | ( ~n7635 & n7636 ) ;
  assign n7638 = ( n7398 & ~n7408 ) | ( n7398 & n7637 ) | ( ~n7408 & n7637 ) ;
  assign n7639 = ( n7408 & ~n7398 ) | ( n7408 & n7637 ) | ( ~n7398 & n7637 ) ;
  assign n7640 = ( n7638 & ~n7637 ) | ( n7638 & n7639 ) | ( ~n7637 & n7639 ) ;
  assign n7644 = ~n136 & x119 ;
  assign n7641 = ( x117 & ~n150 ) | ( x117 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n7642 = ( x118 & ~n131 ) | ( x118 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n7643 = n7641 | n7642 ;
  assign n7645 = ( x119 & ~n7644 ) | ( x119 & n7643 ) | ( ~n7644 & n7643 ) ;
  assign n7647 = ( x118 & x119 ) | ( x118 & n7151 ) | ( x119 & n7151 ) ;
  assign n7646 = ( x118 & ~x119 ) | ( x118 & n7151 ) | ( ~x119 & n7151 ) ;
  assign n7648 = ( x119 & ~n7647 ) | ( x119 & n7646 ) | ( ~n7647 & n7646 ) ;
  assign n7649 = ( n139 & ~n7645 ) | ( n139 & n7648 ) | ( ~n7645 & n7648 ) ;
  assign n7650 = ~n139 & n7649 ;
  assign n7651 = ( x2 & n7645 ) | ( x2 & n7650 ) | ( n7645 & n7650 ) ;
  assign n7652 = ( x2 & ~n7650 ) | ( x2 & n7645 ) | ( ~n7650 & n7645 ) ;
  assign n7653 = ( n7650 & ~n7651 ) | ( n7650 & n7652 ) | ( ~n7651 & n7652 ) ;
  assign n7654 = ( n7396 & n7640 ) | ( n7396 & n7653 ) | ( n7640 & n7653 ) ;
  assign n7655 = ( n7396 & ~n7640 ) | ( n7396 & n7653 ) | ( ~n7640 & n7653 ) ;
  assign n7656 = ( n7640 & ~n7654 ) | ( n7640 & n7655 ) | ( ~n7654 & n7655 ) ;
  assign n7677 = ( n7419 & ~n7604 ) | ( n7419 & n7429 ) | ( ~n7604 & n7429 ) ;
  assign n7681 = x103 &  n942 ;
  assign n7678 = ( x105 & ~n896 ) | ( x105 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n7679 = x104 &  n891 ;
  assign n7680 = n7678 | n7679 ;
  assign n7682 = ( x103 & ~n7681 ) | ( x103 & n7680 ) | ( ~n7681 & n7680 ) ;
  assign n7683 = ~n899 & n4442 ;
  assign n7684 = n7682 | n7683 ;
  assign n7685 = ( x17 & ~n7684 ) | ( x17 & 1'b0 ) | ( ~n7684 & 1'b0 ) ;
  assign n7686 = ~x17 & n7684 ;
  assign n7687 = n7685 | n7686 ;
  assign n7691 = x100 &  n1227 ;
  assign n7688 = ( x102 & ~n1154 ) | ( x102 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n7689 = x101 &  n1149 ;
  assign n7690 = n7688 | n7689 ;
  assign n7692 = ( x100 & ~n7691 ) | ( x100 & n7690 ) | ( ~n7691 & n7690 ) ;
  assign n7693 = n1157 | n3872 ;
  assign n7694 = ~n7692 & n7693 ;
  assign n7695 = x20 &  n7694 ;
  assign n7696 = x20 | n7694 ;
  assign n7697 = ~n7695 & n7696 ;
  assign n7849 = x97 &  n1551 ;
  assign n7846 = ( x99 & ~n1451 ) | ( x99 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n7847 = x98 &  n1446 ;
  assign n7848 = n7846 | n7847 ;
  assign n7850 = ( x97 & ~n7849 ) | ( x97 & n7848 ) | ( ~n7849 & n7848 ) ;
  assign n7851 = ~n1454 & n3338 ;
  assign n7852 = n7850 | n7851 ;
  assign n7853 = ( x23 & ~n7852 ) | ( x23 & 1'b0 ) | ( ~n7852 & 1'b0 ) ;
  assign n7854 = ~x23 & n7852 ;
  assign n7855 = n7853 | n7854 ;
  assign n7701 = x94 &  n1894 ;
  assign n7698 = ( x96 & ~n1816 ) | ( x96 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n7699 = x95 &  n1811 ;
  assign n7700 = n7698 | n7699 ;
  assign n7702 = ( x94 & ~n7701 ) | ( x94 & n7700 ) | ( ~n7701 & n7700 ) ;
  assign n7703 = ~n1819 & n2836 ;
  assign n7704 = n7702 | n7703 ;
  assign n7705 = ( x26 & ~n7704 ) | ( x26 & 1'b0 ) | ( ~n7704 & 1'b0 ) ;
  assign n7706 = ~x26 & n7704 ;
  assign n7707 = n7705 | n7706 ;
  assign n7820 = x88 &  n2718 ;
  assign n7817 = ( x90 & ~n2642 ) | ( x90 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n7818 = x89 &  n2637 ;
  assign n7819 = n7817 | n7818 ;
  assign n7821 = ( x88 & ~n7820 ) | ( x88 & n7819 ) | ( ~n7820 & n7819 ) ;
  assign n7822 = ( n1976 & ~n2645 ) | ( n1976 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n7823 = n7821 | n7822 ;
  assign n7824 = ( x32 & ~n7823 ) | ( x32 & 1'b0 ) | ( ~n7823 & 1'b0 ) ;
  assign n7825 = ~x32 & n7823 ;
  assign n7826 = n7824 | n7825 ;
  assign n7711 = x79 &  n4344 ;
  assign n7708 = ( x81 & ~n4143 ) | ( x81 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n7709 = x80 &  n4138 ;
  assign n7710 = n7708 | n7709 ;
  assign n7712 = ( x79 & ~n7711 ) | ( x79 & n7710 ) | ( ~n7711 & n7710 ) ;
  assign n7713 = ( n994 & ~n4146 ) | ( n994 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n7714 = n7712 | n7713 ;
  assign n7715 = ( x41 & ~n7714 ) | ( x41 & 1'b0 ) | ( ~n7714 & 1'b0 ) ;
  assign n7716 = ~x41 & n7714 ;
  assign n7717 = n7715 | n7716 ;
  assign n7718 = ( n7316 & n7558 ) | ( n7316 & n7568 ) | ( n7558 & n7568 ) ;
  assign n7776 = x76 &  n4934 ;
  assign n7773 = ( x78 & ~n4725 ) | ( x78 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n7774 = x77 &  n4720 ;
  assign n7775 = n7773 | n7774 ;
  assign n7777 = ( x76 & ~n7776 ) | ( x76 & n7775 ) | ( ~n7776 & n7775 ) ;
  assign n7778 = ( n693 & ~n4728 ) | ( n693 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n7779 = n7777 | n7778 ;
  assign n7780 = ( x44 & ~n7779 ) | ( x44 & 1'b0 ) | ( ~n7779 & 1'b0 ) ;
  assign n7781 = ~x44 & n7779 ;
  assign n7782 = n7780 | n7781 ;
  assign n7722 = x73 &  n5586 ;
  assign n7719 = ( x75 & ~n5389 ) | ( x75 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n7720 = x74 &  n5384 ;
  assign n7721 = n7719 | n7720 ;
  assign n7723 = ( x73 & ~n7722 ) | ( x73 & n7721 ) | ( ~n7722 & n7721 ) ;
  assign n7724 = ( n540 & ~n5392 ) | ( n540 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n7725 = n7723 | n7724 ;
  assign n7726 = ( x47 & ~n7725 ) | ( x47 & 1'b0 ) | ( ~n7725 & 1'b0 ) ;
  assign n7727 = ~x47 & n7725 ;
  assign n7728 = n7726 | n7727 ;
  assign n7747 = x67 &  n6982 ;
  assign n7744 = ( x69 & ~n6727 ) | ( x69 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n7745 = x68 &  n6722 ;
  assign n7746 = n7744 | n7745 ;
  assign n7748 = ( x67 & ~n7747 ) | ( x67 & n7746 ) | ( ~n7747 & n7746 ) ;
  assign n7749 = ( n246 & ~n6730 ) | ( n246 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n7750 = n7748 | n7749 ;
  assign n7751 = ( x53 & ~n7750 ) | ( x53 & 1'b0 ) | ( ~n7750 & 1'b0 ) ;
  assign n7752 = ~x53 & n7750 ;
  assign n7753 = n7751 | n7752 ;
  assign n7730 = ( x54 & ~x55 ) | ( x54 & n7537 ) | ( ~x55 & n7537 ) ;
  assign n7729 = ( x54 & ~x55 ) | ( x54 & n7277 ) | ( ~x55 & n7277 ) ;
  assign n7731 = ~n7730 |  n7729 ;
  assign n7735 = x64 &  n7731 ;
  assign n7732 = ( x66 & ~n7538 ) | ( x66 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n7733 = x65 &  n7533 ;
  assign n7734 = n7732 | n7733 ;
  assign n7736 = ( x64 & ~n7735 ) | ( x64 & n7734 ) | ( ~n7735 & n7734 ) ;
  assign n7737 = ( n157 & ~n7541 ) | ( n157 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n7738 = n7736 | n7737 ;
  assign n7739 = ( x56 & ~n7278 ) | ( x56 & n7543 ) | ( ~n7278 & n7543 ) ;
  assign n7740 = ~n7543 & n7739 ;
  assign n7741 = ( n7738 & ~x56 ) | ( n7738 & n7740 ) | ( ~x56 & n7740 ) ;
  assign n7742 = ( x56 & ~n7738 ) | ( x56 & n7740 ) | ( ~n7738 & n7740 ) ;
  assign n7743 = ( n7741 & ~n7740 ) | ( n7741 & n7742 ) | ( ~n7740 & n7742 ) ;
  assign n7754 = ( n7548 & ~n7753 ) | ( n7548 & n7743 ) | ( ~n7753 & n7743 ) ;
  assign n7755 = ( n7743 & ~n7548 ) | ( n7743 & n7753 ) | ( ~n7548 & n7753 ) ;
  assign n7756 = ( n7754 & ~n7743 ) | ( n7754 & n7755 ) | ( ~n7743 & n7755 ) ;
  assign n7760 = x70 &  n6288 ;
  assign n7757 = ( x72 & ~n6032 ) | ( x72 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n7758 = x71 &  n6027 ;
  assign n7759 = n7757 | n7758 ;
  assign n7761 = ( x70 & ~n7760 ) | ( x70 & n7759 ) | ( ~n7760 & n7759 ) ;
  assign n7762 = ( n345 & ~n6035 ) | ( n345 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n7763 = n7761 | n7762 ;
  assign n7764 = ( x50 & ~n7763 ) | ( x50 & 1'b0 ) | ( ~n7763 & 1'b0 ) ;
  assign n7765 = ~x50 & n7763 ;
  assign n7766 = n7764 | n7765 ;
  assign n7767 = ( n7756 & ~n7551 ) | ( n7756 & n7766 ) | ( ~n7551 & n7766 ) ;
  assign n7768 = ( n7551 & ~n7766 ) | ( n7551 & n7756 ) | ( ~n7766 & n7756 ) ;
  assign n7769 = ( n7767 & ~n7756 ) | ( n7767 & n7768 ) | ( ~n7756 & n7768 ) ;
  assign n7771 = ( n7554 & n7728 ) | ( n7554 & n7769 ) | ( n7728 & n7769 ) ;
  assign n7770 = ( n7554 & ~n7728 ) | ( n7554 & n7769 ) | ( ~n7728 & n7769 ) ;
  assign n7772 = ( n7728 & ~n7771 ) | ( n7728 & n7770 ) | ( ~n7771 & n7770 ) ;
  assign n7784 = ( n7557 & n7772 ) | ( n7557 & n7782 ) | ( n7772 & n7782 ) ;
  assign n7783 = ( n7557 & ~n7782 ) | ( n7557 & n7772 ) | ( ~n7782 & n7772 ) ;
  assign n7785 = ( n7782 & ~n7784 ) | ( n7782 & n7783 ) | ( ~n7784 & n7783 ) ;
  assign n7787 = ( n7717 & n7718 ) | ( n7717 & n7785 ) | ( n7718 & n7785 ) ;
  assign n7786 = ( n7718 & ~n7717 ) | ( n7718 & n7785 ) | ( ~n7717 & n7785 ) ;
  assign n7788 = ( n7717 & ~n7787 ) | ( n7717 & n7786 ) | ( ~n7787 & n7786 ) ;
  assign n7789 = ( n7319 & n7571 ) | ( n7319 & n7581 ) | ( n7571 & n7581 ) ;
  assign n7793 = x82 &  n3756 ;
  assign n7790 = ( x84 & ~n3602 ) | ( x84 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n7791 = x83 &  n3597 ;
  assign n7792 = n7790 | n7791 ;
  assign n7794 = ( x82 & ~n7793 ) | ( x82 & n7792 ) | ( ~n7793 & n7792 ) ;
  assign n7795 = ( n1199 & ~n3605 ) | ( n1199 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n7796 = n7794 | n7795 ;
  assign n7797 = ( x38 & ~n7796 ) | ( x38 & 1'b0 ) | ( ~n7796 & 1'b0 ) ;
  assign n7798 = ~x38 & n7796 ;
  assign n7799 = n7797 | n7798 ;
  assign n7800 = ( n7788 & ~n7789 ) | ( n7788 & n7799 ) | ( ~n7789 & n7799 ) ;
  assign n7801 = ( n7788 & ~n7799 ) | ( n7788 & n7789 ) | ( ~n7799 & n7789 ) ;
  assign n7802 = ( n7800 & ~n7788 ) | ( n7800 & n7801 ) | ( ~n7788 & n7801 ) ;
  assign n7803 = ( n7322 & n7489 ) | ( n7322 & n7584 ) | ( n7489 & n7584 ) ;
  assign n7807 = x85 &  n3214 ;
  assign n7804 = ( x87 & ~n3087 ) | ( x87 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n7805 = x86 &  n3082 ;
  assign n7806 = n7804 | n7805 ;
  assign n7808 = ( x85 & ~n7807 ) | ( x85 & n7806 ) | ( ~n7807 & n7806 ) ;
  assign n7809 = ( n1512 & ~n3090 ) | ( n1512 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n7810 = n7808 | n7809 ;
  assign n7811 = ( x35 & ~n7810 ) | ( x35 & 1'b0 ) | ( ~n7810 & 1'b0 ) ;
  assign n7812 = ~x35 & n7810 ;
  assign n7813 = n7811 | n7812 ;
  assign n7814 = ( n7802 & ~n7803 ) | ( n7802 & n7813 ) | ( ~n7803 & n7813 ) ;
  assign n7815 = ( n7802 & ~n7813 ) | ( n7802 & n7803 ) | ( ~n7813 & n7803 ) ;
  assign n7816 = ( n7814 & ~n7802 ) | ( n7814 & n7815 ) | ( ~n7802 & n7815 ) ;
  assign n7827 = ( n7588 & ~n7826 ) | ( n7588 & n7816 ) | ( ~n7826 & n7816 ) ;
  assign n7828 = ( n7816 & ~n7588 ) | ( n7816 & n7826 ) | ( ~n7588 & n7826 ) ;
  assign n7829 = ( n7827 & ~n7816 ) | ( n7827 & n7828 ) | ( ~n7816 & n7828 ) ;
  assign n7833 = x91 &  n2312 ;
  assign n7830 = ( x93 & ~n2195 ) | ( x93 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n7831 = x92 &  n2190 ;
  assign n7832 = n7830 | n7831 ;
  assign n7834 = ( x91 & ~n7833 ) | ( x91 & n7832 ) | ( ~n7833 & n7832 ) ;
  assign n7835 = n2198 | n2264 ;
  assign n7836 = ~n7834 & n7835 ;
  assign n7837 = x29 &  n7836 ;
  assign n7838 = x29 | n7836 ;
  assign n7839 = ~n7837 & n7838 ;
  assign n7841 = ( n7591 & n7829 ) | ( n7591 & n7839 ) | ( n7829 & n7839 ) ;
  assign n7840 = ( n7591 & ~n7829 ) | ( n7591 & n7839 ) | ( ~n7829 & n7839 ) ;
  assign n7842 = ( n7829 & ~n7841 ) | ( n7829 & n7840 ) | ( ~n7841 & n7840 ) ;
  assign n7843 = ( n7707 & ~n7594 ) | ( n7707 & n7842 ) | ( ~n7594 & n7842 ) ;
  assign n7844 = ( n7594 & ~n7842 ) | ( n7594 & n7707 ) | ( ~n7842 & n7707 ) ;
  assign n7845 = ( n7843 & ~n7707 ) | ( n7843 & n7844 ) | ( ~n7707 & n7844 ) ;
  assign n7856 = ( n7598 & ~n7855 ) | ( n7598 & n7845 ) | ( ~n7855 & n7845 ) ;
  assign n7857 = ( n7845 & ~n7598 ) | ( n7845 & n7855 ) | ( ~n7598 & n7855 ) ;
  assign n7858 = ( n7856 & ~n7845 ) | ( n7856 & n7857 ) | ( ~n7845 & n7857 ) ;
  assign n7859 = ( n7602 & n7697 ) | ( n7602 & n7858 ) | ( n7697 & n7858 ) ;
  assign n7860 = ( n7602 & ~n7697 ) | ( n7602 & n7858 ) | ( ~n7697 & n7858 ) ;
  assign n7861 = ( n7697 & ~n7859 ) | ( n7697 & n7860 ) | ( ~n7859 & n7860 ) ;
  assign n7863 = ( n7677 & n7687 ) | ( n7677 & n7861 ) | ( n7687 & n7861 ) ;
  assign n7862 = ( n7687 & ~n7677 ) | ( n7687 & n7861 ) | ( ~n7677 & n7861 ) ;
  assign n7864 = ( n7677 & ~n7863 ) | ( n7677 & n7862 ) | ( ~n7863 & n7862 ) ;
  assign n7865 = ( n7607 & n7608 ) | ( n7607 & n7618 ) | ( n7608 & n7618 ) ;
  assign n7869 = x106 &  n713 ;
  assign n7866 = ( x108 & ~n641 ) | ( x108 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n7867 = x107 &  n636 ;
  assign n7868 = n7866 | n7867 ;
  assign n7870 = ( x106 & ~n7869 ) | ( x106 & n7868 ) | ( ~n7869 & n7868 ) ;
  assign n7871 = n644 | n5055 ;
  assign n7872 = ~n7870 & n7871 ;
  assign n7873 = x14 &  n7872 ;
  assign n7874 = x14 | n7872 ;
  assign n7875 = ~n7873 & n7874 ;
  assign n7876 = ( n7864 & n7865 ) | ( n7864 & n7875 ) | ( n7865 & n7875 ) ;
  assign n7877 = ( n7865 & ~n7864 ) | ( n7865 & n7875 ) | ( ~n7864 & n7875 ) ;
  assign n7878 = ( n7864 & ~n7876 ) | ( n7864 & n7877 ) | ( ~n7876 & n7877 ) ;
  assign n7879 = ( n7377 & ~n7631 ) | ( n7377 & n7621 ) | ( ~n7631 & n7621 ) ;
  assign n7883 = x109 &  n503 ;
  assign n7880 = ( x111 & ~n450 ) | ( x111 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n7881 = x110 &  n445 ;
  assign n7882 = n7880 | n7881 ;
  assign n7884 = ( x109 & ~n7883 ) | ( x109 & n7882 ) | ( ~n7883 & n7882 ) ;
  assign n7885 = n453 | n5711 ;
  assign n7886 = ~n7884 & n7885 ;
  assign n7887 = x11 &  n7886 ;
  assign n7888 = x11 | n7886 ;
  assign n7889 = ~n7887 & n7888 ;
  assign n7890 = ( n7878 & n7879 ) | ( n7878 & n7889 ) | ( n7879 & n7889 ) ;
  assign n7891 = ( n7879 & ~n7878 ) | ( n7879 & n7889 ) | ( ~n7878 & n7889 ) ;
  assign n7892 = ( n7878 & ~n7890 ) | ( n7878 & n7891 ) | ( ~n7890 & n7891 ) ;
  assign n7670 = x112 &  n353 ;
  assign n7667 = ( x114 & ~n313 ) | ( x114 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n7668 = x113 &  n308 ;
  assign n7669 = n7667 | n7668 ;
  assign n7671 = ( x112 & ~n7670 ) | ( x112 & n7669 ) | ( ~n7670 & n7669 ) ;
  assign n7672 = n316 | n6185 ;
  assign n7673 = ~n7671 & n7672 ;
  assign n7674 = x8 &  n7673 ;
  assign n7675 = x8 | n7673 ;
  assign n7676 = ~n7674 & n7675 ;
  assign n7894 = ( n7635 & n7676 ) | ( n7635 & n7892 ) | ( n7676 & n7892 ) ;
  assign n7893 = ( n7635 & ~n7892 ) | ( n7635 & n7676 ) | ( ~n7892 & n7676 ) ;
  assign n7895 = ( n7892 & ~n7894 ) | ( n7892 & n7893 ) | ( ~n7894 & n7893 ) ;
  assign n7660 = x115 &  n225 ;
  assign n7657 = ( x117 & ~n197 ) | ( x117 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n7658 = x116 &  n192 ;
  assign n7659 = n7657 | n7658 ;
  assign n7661 = ( x115 & ~n7660 ) | ( x115 & n7659 ) | ( ~n7660 & n7659 ) ;
  assign n7662 = n200 | n7136 ;
  assign n7663 = ~n7661 & n7662 ;
  assign n7664 = x5 &  n7663 ;
  assign n7665 = x5 | n7663 ;
  assign n7666 = ~n7664 & n7665 ;
  assign n7896 = ( n7639 & ~n7895 ) | ( n7639 & n7666 ) | ( ~n7895 & n7666 ) ;
  assign n7897 = ( n7639 & ~n7666 ) | ( n7639 & n7895 ) | ( ~n7666 & n7895 ) ;
  assign n7898 = ( n7896 & ~n7639 ) | ( n7896 & n7897 ) | ( ~n7639 & n7897 ) ;
  assign n7899 = ( n7640 & ~n7396 ) | ( n7640 & n7653 ) | ( ~n7396 & n7653 ) ;
  assign n7903 = ~n136 & x120 ;
  assign n7900 = ( x118 & ~n150 ) | ( x118 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n7901 = ( x119 & ~n131 ) | ( x119 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n7902 = n7900 | n7901 ;
  assign n7904 = ( x120 & ~n7903 ) | ( x120 & n7902 ) | ( ~n7903 & n7902 ) ;
  assign n7905 = x119 | x120 ;
  assign n7906 = x119 &  x120 ;
  assign n7907 = ( n7905 & ~n7906 ) | ( n7905 & 1'b0 ) | ( ~n7906 & 1'b0 ) ;
  assign n7908 = n7647 &  n7907 ;
  assign n7909 = ( n7647 & ~n139 ) | ( n7647 & n7907 ) | ( ~n139 & n7907 ) ;
  assign n7910 = ( n7904 & ~n7908 ) | ( n7904 & n7909 ) | ( ~n7908 & n7909 ) ;
  assign n7911 = ( x2 & ~n7910 ) | ( x2 & 1'b0 ) | ( ~n7910 & 1'b0 ) ;
  assign n7912 = ~x2 & n7910 ;
  assign n7913 = n7911 | n7912 ;
  assign n7914 = ( n7898 & n7899 ) | ( n7898 & n7913 ) | ( n7899 & n7913 ) ;
  assign n7915 = ( n7899 & ~n7898 ) | ( n7899 & n7913 ) | ( ~n7898 & n7913 ) ;
  assign n7916 = ( n7898 & ~n7914 ) | ( n7898 & n7915 ) | ( ~n7914 & n7915 ) ;
  assign n8171 = ~n136 & x121 ;
  assign n8168 = ( x119 & ~n150 ) | ( x119 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n8169 = ( x120 & ~n131 ) | ( x120 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n8170 = n8168 | n8169 ;
  assign n8172 = ( x121 & ~n8171 ) | ( x121 & n8170 ) | ( ~n8171 & n8170 ) ;
  assign n8173 = ( x119 & ~x121 ) | ( x119 & x120 ) | ( ~x121 & x120 ) ;
  assign n8175 = ( x120 & ~n8173 ) | ( x120 & n7647 ) | ( ~n8173 & n7647 ) ;
  assign n8174 = ( n7647 & ~x119 ) | ( n7647 & n8173 ) | ( ~x119 & n8173 ) ;
  assign n8176 = ( x121 & ~n8175 ) | ( x121 & n8174 ) | ( ~n8175 & n8174 ) ;
  assign n8177 = ( n139 & ~n8172 ) | ( n139 & n8176 ) | ( ~n8172 & n8176 ) ;
  assign n8178 = ~n139 & n8177 ;
  assign n8179 = ( x2 & n8172 ) | ( x2 & n8178 ) | ( n8172 & n8178 ) ;
  assign n8180 = ( x2 & ~n8178 ) | ( x2 & n8172 ) | ( ~n8178 & n8172 ) ;
  assign n8181 = ( n8178 & ~n8179 ) | ( n8178 & n8180 ) | ( ~n8179 & n8180 ) ;
  assign n7930 = x113 &  n353 ;
  assign n7927 = ( x115 & ~n313 ) | ( x115 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n7928 = x114 &  n308 ;
  assign n7929 = n7927 | n7928 ;
  assign n7931 = ( x113 & ~n7930 ) | ( x113 & n7929 ) | ( ~n7930 & n7929 ) ;
  assign n7932 = ~n316 & n6420 ;
  assign n7933 = n7931 | n7932 ;
  assign n7934 = ( x8 & ~n7933 ) | ( x8 & 1'b0 ) | ( ~n7933 & 1'b0 ) ;
  assign n7935 = ~x8 & n7933 ;
  assign n7936 = n7934 | n7935 ;
  assign n7940 = x110 &  n503 ;
  assign n7937 = ( x112 & ~n450 ) | ( x112 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n7938 = x111 &  n445 ;
  assign n7939 = n7937 | n7938 ;
  assign n7941 = ( x110 & ~n7940 ) | ( x110 & n7939 ) | ( ~n7940 & n7939 ) ;
  assign n7942 = ~n453 & n5727 ;
  assign n7943 = n7941 | n7942 ;
  assign n7944 = ( x11 & ~n7943 ) | ( x11 & 1'b0 ) | ( ~n7943 & 1'b0 ) ;
  assign n7945 = ~x11 & n7943 ;
  assign n7946 = n7944 | n7945 ;
  assign n7947 = ( n7878 & ~n7879 ) | ( n7878 & n7889 ) | ( ~n7879 & n7889 ) ;
  assign n7951 = x107 &  n713 ;
  assign n7948 = ( x109 & ~n641 ) | ( x109 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n7949 = x108 &  n636 ;
  assign n7950 = n7948 | n7949 ;
  assign n7952 = ( x107 & ~n7951 ) | ( x107 & n7950 ) | ( ~n7951 & n7950 ) ;
  assign n7953 = ~n644 & n5267 ;
  assign n7954 = n7952 | n7953 ;
  assign n7955 = ( x14 & ~n7954 ) | ( x14 & 1'b0 ) | ( ~n7954 & 1'b0 ) ;
  assign n7956 = ~x14 & n7954 ;
  assign n7957 = n7955 | n7956 ;
  assign n7958 = ( n7864 & ~n7875 ) | ( n7864 & n7865 ) | ( ~n7875 & n7865 ) ;
  assign n7959 = ( n7677 & ~n7687 ) | ( n7677 & n7861 ) | ( ~n7687 & n7861 ) ;
  assign n7963 = x104 &  n942 ;
  assign n7960 = ( x106 & ~n896 ) | ( x106 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n7961 = x105 &  n891 ;
  assign n7962 = n7960 | n7961 ;
  assign n7964 = ( x104 & ~n7963 ) | ( x104 & n7962 ) | ( ~n7963 & n7962 ) ;
  assign n7965 = ~n899 & n4458 ;
  assign n7966 = n7964 | n7965 ;
  assign n7967 = ( x17 & ~n7966 ) | ( x17 & 1'b0 ) | ( ~n7966 & 1'b0 ) ;
  assign n7968 = ~x17 & n7966 ;
  assign n7969 = n7967 | n7968 ;
  assign n7983 = x92 &  n2312 ;
  assign n7980 = ( x94 & ~n2195 ) | ( x94 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n7981 = x93 &  n2190 ;
  assign n7982 = n7980 | n7981 ;
  assign n7984 = ( x92 & ~n7983 ) | ( x92 & n7982 ) | ( ~n7983 & n7982 ) ;
  assign n7985 = ~n2198 & n2401 ;
  assign n7986 = n7984 | n7985 ;
  assign n7987 = ( x29 & ~n7986 ) | ( x29 & 1'b0 ) | ( ~n7986 & 1'b0 ) ;
  assign n7988 = ~x29 & n7986 ;
  assign n7989 = n7987 | n7988 ;
  assign n7990 = ( n7591 & ~n7839 ) | ( n7591 & n7829 ) | ( ~n7839 & n7829 ) ;
  assign n7994 = x86 &  n3214 ;
  assign n7991 = ( x88 & ~n3087 ) | ( x88 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n7992 = x87 &  n3082 ;
  assign n7993 = n7991 | n7992 ;
  assign n7995 = ( x86 & ~n7994 ) | ( x86 & n7993 ) | ( ~n7994 & n7993 ) ;
  assign n7996 = ( n1624 & ~n3090 ) | ( n1624 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n7997 = n7995 | n7996 ;
  assign n7998 = ( x35 & ~n7997 ) | ( x35 & 1'b0 ) | ( ~n7997 & 1'b0 ) ;
  assign n7999 = ~x35 & n7997 ;
  assign n8000 = n7998 | n7999 ;
  assign n8004 = x83 &  n3756 ;
  assign n8001 = ( x85 & ~n3602 ) | ( x85 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n8002 = x84 &  n3597 ;
  assign n8003 = n8001 | n8002 ;
  assign n8005 = ( x83 & ~n8004 ) | ( x83 & n8003 ) | ( ~n8004 & n8003 ) ;
  assign n8006 = ( n1295 & ~n3605 ) | ( n1295 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n8007 = n8005 | n8006 ;
  assign n8008 = ( x38 & ~n8007 ) | ( x38 & 1'b0 ) | ( ~n8007 & 1'b0 ) ;
  assign n8009 = ~x38 & n8007 ;
  assign n8010 = n8008 | n8009 ;
  assign n8011 = ( n7788 & n7789 ) | ( n7788 & n7799 ) | ( n7789 & n7799 ) ;
  assign n8015 = x80 &  n4344 ;
  assign n8012 = ( x82 & ~n4143 ) | ( x82 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n8013 = x81 &  n4138 ;
  assign n8014 = n8012 | n8013 ;
  assign n8016 = ( x80 & ~n8015 ) | ( x80 & n8014 ) | ( ~n8015 & n8014 ) ;
  assign n8017 = ( n1084 & ~n4146 ) | ( n1084 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n8018 = n8016 | n8017 ;
  assign n8019 = ( x41 & ~n8018 ) | ( x41 & 1'b0 ) | ( ~n8018 & 1'b0 ) ;
  assign n8020 = ~x41 & n8018 ;
  assign n8021 = n8019 | n8020 ;
  assign n8025 = x77 &  n4934 ;
  assign n8022 = ( x79 & ~n4725 ) | ( x79 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n8023 = x78 &  n4720 ;
  assign n8024 = n8022 | n8023 ;
  assign n8026 = ( x77 & ~n8025 ) | ( x77 & n8024 ) | ( ~n8025 & n8024 ) ;
  assign n8027 = ( n766 & ~n4728 ) | ( n766 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n8028 = n8026 | n8027 ;
  assign n8029 = ( x44 & ~n8028 ) | ( x44 & 1'b0 ) | ( ~n8028 & 1'b0 ) ;
  assign n8030 = ~x44 & n8028 ;
  assign n8031 = n8029 | n8030 ;
  assign n8035 = x74 &  n5586 ;
  assign n8032 = ( x76 & ~n5389 ) | ( x76 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n8033 = x75 &  n5384 ;
  assign n8034 = n8032 | n8033 ;
  assign n8036 = ( x74 & ~n8035 ) | ( x74 & n8034 ) | ( ~n8035 & n8034 ) ;
  assign n8037 = ( n603 & ~n5392 ) | ( n603 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n8038 = n8036 | n8037 ;
  assign n8039 = ( x47 & ~n8038 ) | ( x47 & 1'b0 ) | ( ~n8038 & 1'b0 ) ;
  assign n8040 = ~x47 & n8038 ;
  assign n8041 = n8039 | n8040 ;
  assign n8042 = ( x56 & ~x57 ) | ( x56 & 1'b0 ) | ( ~x57 & 1'b0 ) ;
  assign n8043 = ~x56 & x57 ;
  assign n8044 = n8042 | n8043 ;
  assign n8045 = x64 &  n8044 ;
  assign n8046 = ( n7278 & ~n7543 ) | ( n7278 & n7738 ) | ( ~n7543 & n7738 ) ;
  assign n8047 = ( x56 & n7543 ) | ( x56 & n8046 ) | ( n7543 & n8046 ) ;
  assign n8048 = ( x56 & ~n8047 ) | ( x56 & 1'b0 ) | ( ~n8047 & 1'b0 ) ;
  assign n8052 = x65 &  n7731 ;
  assign n8049 = ( x67 & ~n7538 ) | ( x67 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n8050 = x66 &  n7533 ;
  assign n8051 = n8049 | n8050 ;
  assign n8053 = ( x65 & ~n8052 ) | ( x65 & n8051 ) | ( ~n8052 & n8051 ) ;
  assign n8054 = n173 | n7541 ;
  assign n8055 = ~n8053 & n8054 ;
  assign n8056 = x56 &  n8055 ;
  assign n8057 = x56 | n8055 ;
  assign n8058 = ~n8056 & n8057 ;
  assign n8059 = ( n8045 & ~n8048 ) | ( n8045 & n8058 ) | ( ~n8048 & n8058 ) ;
  assign n8060 = ( n8045 & ~n8058 ) | ( n8045 & n8048 ) | ( ~n8058 & n8048 ) ;
  assign n8061 = ( n8059 & ~n8045 ) | ( n8059 & n8060 ) | ( ~n8045 & n8060 ) ;
  assign n8062 = ( n7548 & n7743 ) | ( n7548 & n7753 ) | ( n7743 & n7753 ) ;
  assign n8066 = x68 &  n6982 ;
  assign n8063 = ( x70 & ~n6727 ) | ( x70 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n8064 = x69 &  n6722 ;
  assign n8065 = n8063 | n8064 ;
  assign n8067 = ( x68 & ~n8066 ) | ( x68 & n8065 ) | ( ~n8066 & n8065 ) ;
  assign n8068 = ( n282 & ~n6730 ) | ( n282 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n8069 = n8067 | n8068 ;
  assign n8070 = ( x53 & ~n8069 ) | ( x53 & 1'b0 ) | ( ~n8069 & 1'b0 ) ;
  assign n8071 = ~x53 & n8069 ;
  assign n8072 = n8070 | n8071 ;
  assign n8073 = ( n8061 & ~n8062 ) | ( n8061 & n8072 ) | ( ~n8062 & n8072 ) ;
  assign n8074 = ( n8062 & ~n8061 ) | ( n8062 & n8072 ) | ( ~n8061 & n8072 ) ;
  assign n8075 = ( n8073 & ~n8072 ) | ( n8073 & n8074 ) | ( ~n8072 & n8074 ) ;
  assign n8080 = x71 &  n6288 ;
  assign n8077 = ( x73 & ~n6032 ) | ( x73 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n8078 = x72 &  n6027 ;
  assign n8079 = n8077 | n8078 ;
  assign n8081 = ( x71 & ~n8080 ) | ( x71 & n8079 ) | ( ~n8080 & n8079 ) ;
  assign n8082 = ( n389 & ~n6035 ) | ( n389 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n8083 = n8081 | n8082 ;
  assign n8084 = ( x50 & ~n8083 ) | ( x50 & 1'b0 ) | ( ~n8083 & 1'b0 ) ;
  assign n8085 = ~x50 & n8083 ;
  assign n8086 = n8084 | n8085 ;
  assign n8076 = ( n7551 & n7756 ) | ( n7551 & n7766 ) | ( n7756 & n7766 ) ;
  assign n8087 = ( n8075 & ~n8086 ) | ( n8075 & n8076 ) | ( ~n8086 & n8076 ) ;
  assign n8088 = ( n8075 & ~n8076 ) | ( n8075 & n8086 ) | ( ~n8076 & n8086 ) ;
  assign n8089 = ( n8087 & ~n8075 ) | ( n8087 & n8088 ) | ( ~n8075 & n8088 ) ;
  assign n8090 = ( n8041 & ~n7771 ) | ( n8041 & n8089 ) | ( ~n7771 & n8089 ) ;
  assign n8091 = ( n7771 & ~n8089 ) | ( n7771 & n8041 ) | ( ~n8089 & n8041 ) ;
  assign n8092 = ( n8090 & ~n8041 ) | ( n8090 & n8091 ) | ( ~n8041 & n8091 ) ;
  assign n8093 = ( n8031 & ~n7784 ) | ( n8031 & n8092 ) | ( ~n7784 & n8092 ) ;
  assign n8094 = ( n7784 & ~n8092 ) | ( n7784 & n8031 ) | ( ~n8092 & n8031 ) ;
  assign n8095 = ( n8093 & ~n8031 ) | ( n8093 & n8094 ) | ( ~n8031 & n8094 ) ;
  assign n8096 = ( n8021 & ~n7787 ) | ( n8021 & n8095 ) | ( ~n7787 & n8095 ) ;
  assign n8097 = ( n7787 & ~n8095 ) | ( n7787 & n8021 ) | ( ~n8095 & n8021 ) ;
  assign n8098 = ( n8096 & ~n8021 ) | ( n8096 & n8097 ) | ( ~n8021 & n8097 ) ;
  assign n8099 = ( n8010 & ~n8011 ) | ( n8010 & n8098 ) | ( ~n8011 & n8098 ) ;
  assign n8100 = ( n8010 & ~n8098 ) | ( n8010 & n8011 ) | ( ~n8098 & n8011 ) ;
  assign n8101 = ( n8099 & ~n8010 ) | ( n8099 & n8100 ) | ( ~n8010 & n8100 ) ;
  assign n8102 = ( n7802 & n7803 ) | ( n7802 & n7813 ) | ( n7803 & n7813 ) ;
  assign n8103 = ( n8000 & ~n8101 ) | ( n8000 & n8102 ) | ( ~n8101 & n8102 ) ;
  assign n8104 = ( n8000 & ~n8102 ) | ( n8000 & n8101 ) | ( ~n8102 & n8101 ) ;
  assign n8105 = ( n8103 & ~n8000 ) | ( n8103 & n8104 ) | ( ~n8000 & n8104 ) ;
  assign n8106 = ( n7588 & n7816 ) | ( n7588 & n7826 ) | ( n7816 & n7826 ) ;
  assign n8110 = x89 &  n2718 ;
  assign n8107 = ( x91 & ~n2642 ) | ( x91 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n8108 = x90 &  n2637 ;
  assign n8109 = n8107 | n8108 ;
  assign n8111 = ( x89 & ~n8110 ) | ( x89 & n8109 ) | ( ~n8110 & n8109 ) ;
  assign n8112 = ( n2108 & ~n2645 ) | ( n2108 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n8113 = n8111 | n8112 ;
  assign n8114 = ( x32 & ~n8113 ) | ( x32 & 1'b0 ) | ( ~n8113 & 1'b0 ) ;
  assign n8115 = ~x32 & n8113 ;
  assign n8116 = n8114 | n8115 ;
  assign n8117 = ( n8105 & ~n8106 ) | ( n8105 & n8116 ) | ( ~n8106 & n8116 ) ;
  assign n8118 = ( n8105 & ~n8116 ) | ( n8105 & n8106 ) | ( ~n8116 & n8106 ) ;
  assign n8119 = ( n8117 & ~n8105 ) | ( n8117 & n8118 ) | ( ~n8105 & n8118 ) ;
  assign n8120 = ( n7989 & ~n7990 ) | ( n7989 & n8119 ) | ( ~n7990 & n8119 ) ;
  assign n8121 = ( n7989 & ~n8119 ) | ( n7989 & n7990 ) | ( ~n8119 & n7990 ) ;
  assign n8122 = ( n8120 & ~n7989 ) | ( n8120 & n8121 ) | ( ~n7989 & n8121 ) ;
  assign n8126 = x95 &  n1894 ;
  assign n8123 = ( x97 & ~n1816 ) | ( x97 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n8124 = x96 &  n1811 ;
  assign n8125 = n8123 | n8124 ;
  assign n8127 = ( x95 & ~n8126 ) | ( x95 & n8125 ) | ( ~n8126 & n8125 ) ;
  assign n8128 = ~n1819 & n2999 ;
  assign n8129 = n8127 | n8128 ;
  assign n8130 = ( x26 & ~n8129 ) | ( x26 & 1'b0 ) | ( ~n8129 & 1'b0 ) ;
  assign n8131 = ~x26 & n8129 ;
  assign n8132 = n8130 | n8131 ;
  assign n8133 = ( n8122 & ~n7844 ) | ( n8122 & n8132 ) | ( ~n7844 & n8132 ) ;
  assign n8134 = ( n7844 & ~n8132 ) | ( n7844 & n8122 ) | ( ~n8132 & n8122 ) ;
  assign n8135 = ( n8133 & ~n8122 ) | ( n8133 & n8134 ) | ( ~n8122 & n8134 ) ;
  assign n8136 = ( n7598 & ~n7845 ) | ( n7598 & n7855 ) | ( ~n7845 & n7855 ) ;
  assign n8140 = x98 &  n1551 ;
  assign n8137 = ( x100 & ~n1451 ) | ( x100 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n8138 = x99 &  n1446 ;
  assign n8139 = n8137 | n8138 ;
  assign n8141 = ( x98 & ~n8140 ) | ( x98 & n8139 ) | ( ~n8140 & n8139 ) ;
  assign n8142 = n1454 | n3354 ;
  assign n8143 = ~n8141 & n8142 ;
  assign n8144 = x23 &  n8143 ;
  assign n8145 = x23 | n8143 ;
  assign n8146 = ~n8144 & n8145 ;
  assign n8147 = ( n8135 & n8136 ) | ( n8135 & n8146 ) | ( n8136 & n8146 ) ;
  assign n8148 = ( n8136 & ~n8135 ) | ( n8136 & n8146 ) | ( ~n8135 & n8146 ) ;
  assign n8149 = ( n8135 & ~n8147 ) | ( n8135 & n8148 ) | ( ~n8147 & n8148 ) ;
  assign n7973 = x101 &  n1227 ;
  assign n7970 = ( x103 & ~n1154 ) | ( x103 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n7971 = x102 &  n1149 ;
  assign n7972 = n7970 | n7971 ;
  assign n7974 = ( x101 & ~n7973 ) | ( x101 & n7972 ) | ( ~n7973 & n7972 ) ;
  assign n7975 = n1157 | n4056 ;
  assign n7976 = ~n7974 & n7975 ;
  assign n7977 = x20 &  n7976 ;
  assign n7978 = x20 | n7976 ;
  assign n7979 = ~n7977 & n7978 ;
  assign n8150 = ( n7859 & ~n8149 ) | ( n7859 & n7979 ) | ( ~n8149 & n7979 ) ;
  assign n8151 = ( n7979 & ~n7859 ) | ( n7979 & n8149 ) | ( ~n7859 & n8149 ) ;
  assign n8152 = ( n8150 & ~n7979 ) | ( n8150 & n8151 ) | ( ~n7979 & n8151 ) ;
  assign n8153 = ( n7959 & ~n7969 ) | ( n7959 & n8152 ) | ( ~n7969 & n8152 ) ;
  assign n8154 = ( n7959 & ~n8152 ) | ( n7959 & n7969 ) | ( ~n8152 & n7969 ) ;
  assign n8155 = ( n8153 & ~n7959 ) | ( n8153 & n8154 ) | ( ~n7959 & n8154 ) ;
  assign n8156 = ( n7957 & ~n7958 ) | ( n7957 & n8155 ) | ( ~n7958 & n8155 ) ;
  assign n8157 = ( n7957 & ~n8155 ) | ( n7957 & n7958 ) | ( ~n8155 & n7958 ) ;
  assign n8158 = ( n8156 & ~n7957 ) | ( n8156 & n8157 ) | ( ~n7957 & n8157 ) ;
  assign n8159 = ( n7946 & n7947 ) | ( n7946 & n8158 ) | ( n7947 & n8158 ) ;
  assign n8160 = ( n7947 & ~n7946 ) | ( n7947 & n8158 ) | ( ~n7946 & n8158 ) ;
  assign n8161 = ( n7946 & ~n8159 ) | ( n7946 & n8160 ) | ( ~n8159 & n8160 ) ;
  assign n8162 = ( n7936 & ~n7893 ) | ( n7936 & n8161 ) | ( ~n7893 & n8161 ) ;
  assign n8163 = ( n7893 & ~n7936 ) | ( n7893 & n8161 ) | ( ~n7936 & n8161 ) ;
  assign n8164 = ( n8162 & ~n8161 ) | ( n8162 & n8163 ) | ( ~n8161 & n8163 ) ;
  assign n7920 = x116 &  n225 ;
  assign n7917 = ( x118 & ~n197 ) | ( x118 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n7918 = x117 &  n192 ;
  assign n7919 = n7917 | n7918 ;
  assign n7921 = ( x116 & ~n7920 ) | ( x116 & n7919 ) | ( ~n7920 & n7919 ) ;
  assign n7922 = n200 | n7152 ;
  assign n7923 = ~n7921 & n7922 ;
  assign n7924 = x5 &  n7923 ;
  assign n7925 = x5 | n7923 ;
  assign n7926 = ~n7924 & n7925 ;
  assign n8165 = ( n7896 & n7926 ) | ( n7896 & n8164 ) | ( n7926 & n8164 ) ;
  assign n8166 = ( n7896 & ~n8164 ) | ( n7896 & n7926 ) | ( ~n8164 & n7926 ) ;
  assign n8167 = ( n8164 & ~n8165 ) | ( n8164 & n8166 ) | ( ~n8165 & n8166 ) ;
  assign n8182 = ( n7914 & n8167 ) | ( n7914 & n8181 ) | ( n8167 & n8181 ) ;
  assign n8183 = ( n7914 & ~n8181 ) | ( n7914 & n8167 ) | ( ~n8181 & n8167 ) ;
  assign n8184 = ( n8181 & ~n8182 ) | ( n8181 & n8183 ) | ( ~n8182 & n8183 ) ;
  assign n8188 = x117 &  n225 ;
  assign n8185 = ( x119 & ~n197 ) | ( x119 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n8186 = x118 &  n192 ;
  assign n8187 = n8185 | n8186 ;
  assign n8189 = ( x117 & ~n8188 ) | ( x117 & n8187 ) | ( ~n8188 & n8187 ) ;
  assign n8190 = ~n200 & n7648 ;
  assign n8191 = n8189 | n8190 ;
  assign n8192 = ( x5 & ~n8191 ) | ( x5 & 1'b0 ) | ( ~n8191 & 1'b0 ) ;
  assign n8193 = ~x5 & n8191 ;
  assign n8194 = n8192 | n8193 ;
  assign n8198 = x114 &  n353 ;
  assign n8195 = ( x116 & ~n313 ) | ( x116 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n8196 = x115 &  n308 ;
  assign n8197 = n8195 | n8196 ;
  assign n8199 = ( x114 & ~n8198 ) | ( x114 & n8197 ) | ( ~n8198 & n8197 ) ;
  assign n8200 = n316 | n6885 ;
  assign n8201 = ~n8199 & n8200 ;
  assign n8202 = x8 &  n8201 ;
  assign n8203 = x8 | n8201 ;
  assign n8204 = ~n8202 & n8203 ;
  assign n8208 = x111 &  n503 ;
  assign n8205 = ( x113 & ~n450 ) | ( x113 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n8206 = x112 &  n445 ;
  assign n8207 = n8205 | n8206 ;
  assign n8209 = ( x111 & ~n8208 ) | ( x111 & n8207 ) | ( ~n8208 & n8207 ) ;
  assign n8210 = n453 | n6169 ;
  assign n8211 = ~n8209 & n8210 ;
  assign n8212 = x11 &  n8211 ;
  assign n8213 = x11 | n8211 ;
  assign n8214 = ~n8212 & n8213 ;
  assign n8215 = ( n7969 & ~n7959 ) | ( n7969 & n8152 ) | ( ~n7959 & n8152 ) ;
  assign n8239 = x99 &  n1551 ;
  assign n8236 = ( x101 & ~n1451 ) | ( x101 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n8237 = x100 &  n1446 ;
  assign n8238 = n8236 | n8237 ;
  assign n8240 = ( x99 & ~n8239 ) | ( x99 & n8238 ) | ( ~n8239 & n8238 ) ;
  assign n8241 = n1454 | n3694 ;
  assign n8242 = ~n8240 & n8241 ;
  assign n8243 = x23 &  n8242 ;
  assign n8244 = x23 | n8242 ;
  assign n8245 = ~n8243 & n8244 ;
  assign n8249 = x96 &  n1894 ;
  assign n8246 = ( x98 & ~n1816 ) | ( x98 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n8247 = x97 &  n1811 ;
  assign n8248 = n8246 | n8247 ;
  assign n8250 = ( x96 & ~n8249 ) | ( x96 & n8248 ) | ( ~n8249 & n8248 ) ;
  assign n8251 = ~n1819 & n3170 ;
  assign n8252 = n8250 | n8251 ;
  assign n8253 = ( x26 & ~n8252 ) | ( x26 & 1'b0 ) | ( ~n8252 & 1'b0 ) ;
  assign n8254 = ~x26 & n8252 ;
  assign n8255 = n8253 | n8254 ;
  assign n8259 = x87 &  n3214 ;
  assign n8256 = ( x89 & ~n3087 ) | ( x89 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n8257 = x88 &  n3082 ;
  assign n8258 = n8256 | n8257 ;
  assign n8260 = ( x87 & ~n8259 ) | ( x87 & n8258 ) | ( ~n8259 & n8258 ) ;
  assign n8261 = ( n1741 & ~n3090 ) | ( n1741 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n8262 = n8260 | n8261 ;
  assign n8263 = ( x35 & ~n8262 ) | ( x35 & 1'b0 ) | ( ~n8262 & 1'b0 ) ;
  assign n8264 = ~x35 & n8262 ;
  assign n8265 = n8263 | n8264 ;
  assign n8362 = x81 &  n4344 ;
  assign n8359 = ( x83 & ~n4143 ) | ( x83 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n8360 = x82 &  n4138 ;
  assign n8361 = n8359 | n8360 ;
  assign n8363 = ( x81 & ~n8362 ) | ( x81 & n8361 ) | ( ~n8362 & n8361 ) ;
  assign n8364 = ( n1100 & ~n4146 ) | ( n1100 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n8365 = n8363 | n8364 ;
  assign n8366 = ( x41 & ~n8365 ) | ( x41 & 1'b0 ) | ( ~n8365 & 1'b0 ) ;
  assign n8367 = ~x41 & n8365 ;
  assign n8368 = n8366 | n8367 ;
  assign n8346 = x75 &  n5586 ;
  assign n8343 = ( x77 & ~n5389 ) | ( x77 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n8344 = x76 &  n5384 ;
  assign n8345 = n8343 | n8344 ;
  assign n8347 = ( x75 & ~n8346 ) | ( x75 & n8345 ) | ( ~n8346 & n8345 ) ;
  assign n8348 = ( n677 & ~n5392 ) | ( n677 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n8349 = n8347 | n8348 ;
  assign n8350 = ( x47 & ~n8349 ) | ( x47 & 1'b0 ) | ( ~n8349 & 1'b0 ) ;
  assign n8351 = ~x47 & n8349 ;
  assign n8352 = n8350 | n8351 ;
  assign n8289 = x69 &  n6982 ;
  assign n8286 = ( x71 & ~n6727 ) | ( x71 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n8287 = x70 &  n6722 ;
  assign n8288 = n8286 | n8287 ;
  assign n8290 = ( x69 & ~n8289 ) | ( x69 & n8288 ) | ( ~n8289 & n8288 ) ;
  assign n8291 = ( n298 & ~n6730 ) | ( n298 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n8292 = n8290 | n8291 ;
  assign n8293 = ( x53 & ~n8292 ) | ( x53 & 1'b0 ) | ( ~n8292 & 1'b0 ) ;
  assign n8294 = ~x53 & n8292 ;
  assign n8295 = n8293 | n8294 ;
  assign n8299 = x66 &  n7731 ;
  assign n8296 = ( x68 & ~n7538 ) | ( x68 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n8297 = x67 &  n7533 ;
  assign n8298 = n8296 | n8297 ;
  assign n8300 = ( x66 & ~n8299 ) | ( x66 & n8298 ) | ( ~n8299 & n8298 ) ;
  assign n8301 = ( n213 & ~n7541 ) | ( n213 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n8302 = n8300 | n8301 ;
  assign n8303 = ( x56 & ~n8302 ) | ( x56 & 1'b0 ) | ( ~n8302 & 1'b0 ) ;
  assign n8304 = ~x56 & n8302 ;
  assign n8305 = n8303 | n8304 ;
  assign n8306 = ( x59 & ~n8045 ) | ( x59 & 1'b0 ) | ( ~n8045 & 1'b0 ) ;
  assign n8307 = ( x57 & x58 ) | ( x57 & n8042 ) | ( x58 & n8042 ) ;
  assign n8308 = ( x57 & ~n8043 ) | ( x57 & x58 ) | ( ~n8043 & x58 ) ;
  assign n8309 = ~n8307 &  n8308 ;
  assign n8310 = x64 &  n8309 ;
  assign n8311 = ~x58 & x59 ;
  assign n8312 = ( x58 & ~x59 ) | ( x58 & 1'b0 ) | ( ~x59 & 1'b0 ) ;
  assign n8313 = n8311 | n8312 ;
  assign n8314 = ~n8044 |  n8313 ;
  assign n8315 = ( x65 & ~n8314 ) | ( x65 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n8316 = n8310 | n8315 ;
  assign n8317 = ~n8044 | ~n8313 ;
  assign n8318 = ( n142 & ~n8317 ) | ( n142 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n8319 = n8316 | n8318 ;
  assign n8321 = ( x59 & n8306 ) | ( x59 & n8319 ) | ( n8306 & n8319 ) ;
  assign n8320 = ( x59 & ~n8306 ) | ( x59 & n8319 ) | ( ~n8306 & n8319 ) ;
  assign n8322 = ( n8306 & ~n8321 ) | ( n8306 & n8320 ) | ( ~n8321 & n8320 ) ;
  assign n8324 = ( n8060 & n8305 ) | ( n8060 & n8322 ) | ( n8305 & n8322 ) ;
  assign n8323 = ( n8060 & ~n8305 ) | ( n8060 & n8322 ) | ( ~n8305 & n8322 ) ;
  assign n8325 = ( n8305 & ~n8324 ) | ( n8305 & n8323 ) | ( ~n8324 & n8323 ) ;
  assign n8327 = ( n8074 & n8295 ) | ( n8074 & n8325 ) | ( n8295 & n8325 ) ;
  assign n8326 = ( n8074 & ~n8295 ) | ( n8074 & n8325 ) | ( ~n8295 & n8325 ) ;
  assign n8328 = ( n8295 & ~n8327 ) | ( n8295 & n8326 ) | ( ~n8327 & n8326 ) ;
  assign n8339 = ( n8076 & ~n8075 ) | ( n8076 & n8086 ) | ( ~n8075 & n8086 ) ;
  assign n8332 = x72 &  n6288 ;
  assign n8329 = ( x74 & ~n6032 ) | ( x74 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n8330 = x73 &  n6027 ;
  assign n8331 = n8329 | n8330 ;
  assign n8333 = ( x72 & ~n8332 ) | ( x72 & n8331 ) | ( ~n8332 & n8331 ) ;
  assign n8334 = ( n482 & ~n6035 ) | ( n482 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n8335 = n8333 | n8334 ;
  assign n8336 = ( x50 & ~n8335 ) | ( x50 & 1'b0 ) | ( ~n8335 & 1'b0 ) ;
  assign n8337 = ~x50 & n8335 ;
  assign n8338 = n8336 | n8337 ;
  assign n8340 = ( n8328 & ~n8339 ) | ( n8328 & n8338 ) | ( ~n8339 & n8338 ) ;
  assign n8341 = ( n8328 & ~n8338 ) | ( n8328 & n8339 ) | ( ~n8338 & n8339 ) ;
  assign n8342 = ( n8340 & ~n8328 ) | ( n8340 & n8341 ) | ( ~n8328 & n8341 ) ;
  assign n8353 = ( n8091 & ~n8352 ) | ( n8091 & n8342 ) | ( ~n8352 & n8342 ) ;
  assign n8354 = ( n8342 & ~n8091 ) | ( n8342 & n8352 ) | ( ~n8091 & n8352 ) ;
  assign n8355 = ( n8353 & ~n8342 ) | ( n8353 & n8354 ) | ( ~n8342 & n8354 ) ;
  assign n8279 = x78 &  n4934 ;
  assign n8276 = ( x80 & ~n4725 ) | ( x80 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n8277 = x79 &  n4720 ;
  assign n8278 = n8276 | n8277 ;
  assign n8280 = ( x78 & ~n8279 ) | ( x78 & n8278 ) | ( ~n8279 & n8278 ) ;
  assign n8281 = ( n842 & ~n4728 ) | ( n842 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n8282 = n8280 | n8281 ;
  assign n8283 = ( x44 & ~n8282 ) | ( x44 & 1'b0 ) | ( ~n8282 & 1'b0 ) ;
  assign n8284 = ~x44 & n8282 ;
  assign n8285 = n8283 | n8284 ;
  assign n8356 = ( n8094 & ~n8355 ) | ( n8094 & n8285 ) | ( ~n8355 & n8285 ) ;
  assign n8357 = ( n8285 & ~n8094 ) | ( n8285 & n8355 ) | ( ~n8094 & n8355 ) ;
  assign n8358 = ( n8356 & ~n8285 ) | ( n8356 & n8357 ) | ( ~n8285 & n8357 ) ;
  assign n8369 = ( n8097 & ~n8368 ) | ( n8097 & n8358 ) | ( ~n8368 & n8358 ) ;
  assign n8370 = ( n8358 & ~n8097 ) | ( n8358 & n8368 ) | ( ~n8097 & n8368 ) ;
  assign n8371 = ( n8369 & ~n8358 ) | ( n8369 & n8370 ) | ( ~n8358 & n8370 ) ;
  assign n8269 = x84 &  n3756 ;
  assign n8266 = ( x86 & ~n3602 ) | ( x86 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n8267 = x85 &  n3597 ;
  assign n8268 = n8266 | n8267 ;
  assign n8270 = ( x84 & ~n8269 ) | ( x84 & n8268 ) | ( ~n8269 & n8268 ) ;
  assign n8271 = ( n1496 & ~n3605 ) | ( n1496 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n8272 = n8270 | n8271 ;
  assign n8273 = ( x38 & ~n8272 ) | ( x38 & 1'b0 ) | ( ~n8272 & 1'b0 ) ;
  assign n8274 = ~x38 & n8272 ;
  assign n8275 = n8273 | n8274 ;
  assign n8372 = ( n8100 & ~n8371 ) | ( n8100 & n8275 ) | ( ~n8371 & n8275 ) ;
  assign n8373 = ( n8275 & ~n8100 ) | ( n8275 & n8371 ) | ( ~n8100 & n8371 ) ;
  assign n8374 = ( n8372 & ~n8275 ) | ( n8372 & n8373 ) | ( ~n8275 & n8373 ) ;
  assign n8375 = ( n8103 & n8265 ) | ( n8103 & n8374 ) | ( n8265 & n8374 ) ;
  assign n8376 = ( n8103 & ~n8265 ) | ( n8103 & n8374 ) | ( ~n8265 & n8374 ) ;
  assign n8377 = ( n8265 & ~n8375 ) | ( n8265 & n8376 ) | ( ~n8375 & n8376 ) ;
  assign n8382 = x90 &  n2718 ;
  assign n8379 = ( x92 & ~n2642 ) | ( x92 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n8380 = x91 &  n2637 ;
  assign n8381 = n8379 | n8380 ;
  assign n8383 = ( x90 & ~n8382 ) | ( x90 & n8381 ) | ( ~n8382 & n8381 ) ;
  assign n8384 = ( n2248 & ~n2645 ) | ( n2248 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n8385 = n8383 | n8384 ;
  assign n8386 = ( x32 & ~n8385 ) | ( x32 & 1'b0 ) | ( ~n8385 & 1'b0 ) ;
  assign n8387 = ~x32 & n8385 ;
  assign n8388 = n8386 | n8387 ;
  assign n8378 = ( n8106 & ~n8105 ) | ( n8106 & n8116 ) | ( ~n8105 & n8116 ) ;
  assign n8389 = ( n8377 & ~n8388 ) | ( n8377 & n8378 ) | ( ~n8388 & n8378 ) ;
  assign n8390 = ( n8377 & ~n8378 ) | ( n8377 & n8388 ) | ( ~n8378 & n8388 ) ;
  assign n8391 = ( n8389 & ~n8377 ) | ( n8389 & n8390 ) | ( ~n8377 & n8390 ) ;
  assign n8395 = x93 &  n2312 ;
  assign n8392 = ( x95 & ~n2195 ) | ( x95 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n8393 = x94 &  n2190 ;
  assign n8394 = n8392 | n8393 ;
  assign n8396 = ( x93 & ~n8395 ) | ( x93 & n8394 ) | ( ~n8395 & n8394 ) ;
  assign n8397 = ~n2198 & n2547 ;
  assign n8398 = n8396 | n8397 ;
  assign n8399 = ( x29 & ~n8398 ) | ( x29 & 1'b0 ) | ( ~n8398 & 1'b0 ) ;
  assign n8400 = ~x29 & n8398 ;
  assign n8401 = n8399 | n8400 ;
  assign n8402 = ( n8391 & ~n8121 ) | ( n8391 & n8401 ) | ( ~n8121 & n8401 ) ;
  assign n8403 = ( n8121 & ~n8401 ) | ( n8121 & n8391 ) | ( ~n8401 & n8391 ) ;
  assign n8404 = ( n8402 & ~n8391 ) | ( n8402 & n8403 ) | ( ~n8391 & n8403 ) ;
  assign n8405 = ( n7844 & ~n8122 ) | ( n7844 & n8132 ) | ( ~n8122 & n8132 ) ;
  assign n8406 = ( n8255 & n8404 ) | ( n8255 & n8405 ) | ( n8404 & n8405 ) ;
  assign n8407 = ( n8404 & ~n8255 ) | ( n8404 & n8405 ) | ( ~n8255 & n8405 ) ;
  assign n8408 = ( n8255 & ~n8406 ) | ( n8255 & n8407 ) | ( ~n8406 & n8407 ) ;
  assign n8409 = ( n8135 & ~n8136 ) | ( n8135 & n8146 ) | ( ~n8136 & n8146 ) ;
  assign n8410 = ( n8245 & ~n8408 ) | ( n8245 & n8409 ) | ( ~n8408 & n8409 ) ;
  assign n8411 = ( n8245 & ~n8409 ) | ( n8245 & n8408 ) | ( ~n8409 & n8408 ) ;
  assign n8412 = ( n8410 & ~n8245 ) | ( n8410 & n8411 ) | ( ~n8245 & n8411 ) ;
  assign n8229 = x102 &  n1227 ;
  assign n8226 = ( x104 & ~n1154 ) | ( x104 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n8227 = x103 &  n1149 ;
  assign n8228 = n8226 | n8227 ;
  assign n8230 = ( x102 & ~n8229 ) | ( x102 & n8228 ) | ( ~n8229 & n8228 ) ;
  assign n8231 = n1157 | n4249 ;
  assign n8232 = ~n8230 & n8231 ;
  assign n8233 = x20 &  n8232 ;
  assign n8234 = x20 | n8232 ;
  assign n8235 = ~n8233 & n8234 ;
  assign n8413 = ( n8150 & ~n8412 ) | ( n8150 & n8235 ) | ( ~n8412 & n8235 ) ;
  assign n8414 = ( n8235 & ~n8150 ) | ( n8235 & n8412 ) | ( ~n8150 & n8412 ) ;
  assign n8415 = ( n8413 & ~n8235 ) | ( n8413 & n8414 ) | ( ~n8235 & n8414 ) ;
  assign n8219 = x105 &  n942 ;
  assign n8216 = ( x107 & ~n896 ) | ( x107 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n8217 = x106 &  n891 ;
  assign n8218 = n8216 | n8217 ;
  assign n8220 = ( x105 & ~n8219 ) | ( x105 & n8218 ) | ( ~n8219 & n8218 ) ;
  assign n8221 = ~n899 & n4848 ;
  assign n8222 = n8220 | n8221 ;
  assign n8223 = ( x17 & ~n8222 ) | ( x17 & 1'b0 ) | ( ~n8222 & 1'b0 ) ;
  assign n8224 = ~x17 & n8222 ;
  assign n8225 = n8223 | n8224 ;
  assign n8416 = ( n8215 & ~n8415 ) | ( n8215 & n8225 ) | ( ~n8415 & n8225 ) ;
  assign n8417 = ( n8215 & ~n8225 ) | ( n8215 & n8415 ) | ( ~n8225 & n8415 ) ;
  assign n8418 = ( n8416 & ~n8215 ) | ( n8416 & n8417 ) | ( ~n8215 & n8417 ) ;
  assign n8422 = x108 &  n713 ;
  assign n8419 = ( x110 & ~n641 ) | ( x110 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n8420 = x109 &  n636 ;
  assign n8421 = n8419 | n8420 ;
  assign n8423 = ( x108 & ~n8422 ) | ( x108 & n8421 ) | ( ~n8422 & n8421 ) ;
  assign n8424 = n644 | n5283 ;
  assign n8425 = ~n8423 & n8424 ;
  assign n8426 = x14 &  n8425 ;
  assign n8427 = x14 | n8425 ;
  assign n8428 = ~n8426 & n8427 ;
  assign n8430 = ( n8157 & n8418 ) | ( n8157 & n8428 ) | ( n8418 & n8428 ) ;
  assign n8429 = ( n8157 & ~n8418 ) | ( n8157 & n8428 ) | ( ~n8418 & n8428 ) ;
  assign n8431 = ( n8418 & ~n8430 ) | ( n8418 & n8429 ) | ( ~n8430 & n8429 ) ;
  assign n8433 = ( n8160 & n8214 ) | ( n8160 & n8431 ) | ( n8214 & n8431 ) ;
  assign n8432 = ( n8160 & ~n8214 ) | ( n8160 & n8431 ) | ( ~n8214 & n8431 ) ;
  assign n8434 = ( n8214 & ~n8433 ) | ( n8214 & n8432 ) | ( ~n8433 & n8432 ) ;
  assign n8435 = ( n8204 & ~n8162 ) | ( n8204 & n8434 ) | ( ~n8162 & n8434 ) ;
  assign n8436 = ( n8162 & ~n8204 ) | ( n8162 & n8434 ) | ( ~n8204 & n8434 ) ;
  assign n8437 = ( n8435 & ~n8434 ) | ( n8435 & n8436 ) | ( ~n8434 & n8436 ) ;
  assign n8438 = ( n8194 & ~n8165 ) | ( n8194 & n8437 ) | ( ~n8165 & n8437 ) ;
  assign n8439 = ( n8165 & ~n8194 ) | ( n8165 & n8437 ) | ( ~n8194 & n8437 ) ;
  assign n8440 = ( n8438 & ~n8437 ) | ( n8438 & n8439 ) | ( ~n8437 & n8439 ) ;
  assign n8441 = ( n7914 & ~n8167 ) | ( n7914 & n8181 ) | ( ~n8167 & n8181 ) ;
  assign n8445 = ~n136 & x122 ;
  assign n8442 = ( x120 & ~n150 ) | ( x120 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n8443 = ( x121 & ~n131 ) | ( x121 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n8444 = n8442 | n8443 ;
  assign n8446 = ( x122 & ~n8445 ) | ( x122 & n8444 ) | ( ~n8445 & n8444 ) ;
  assign n8447 = ( x119 & x120 ) | ( x119 & n7647 ) | ( x120 & n7647 ) ;
  assign n8448 = ( x120 & x121 ) | ( x120 & n8447 ) | ( x121 & n8447 ) ;
  assign n8449 = x121 | x122 ;
  assign n8450 = x121 &  x122 ;
  assign n8451 = ( n8449 & ~n8450 ) | ( n8449 & 1'b0 ) | ( ~n8450 & 1'b0 ) ;
  assign n8452 = n8448 &  n8451 ;
  assign n8453 = ( n8448 & ~n139 ) | ( n8448 & n8451 ) | ( ~n139 & n8451 ) ;
  assign n8454 = ( n8446 & ~n8452 ) | ( n8446 & n8453 ) | ( ~n8452 & n8453 ) ;
  assign n8455 = ( x2 & ~n8454 ) | ( x2 & 1'b0 ) | ( ~n8454 & 1'b0 ) ;
  assign n8456 = ~x2 & n8454 ;
  assign n8457 = n8455 | n8456 ;
  assign n8459 = ( n8440 & n8441 ) | ( n8440 & n8457 ) | ( n8441 & n8457 ) ;
  assign n8458 = ( n8441 & ~n8440 ) | ( n8441 & n8457 ) | ( ~n8440 & n8457 ) ;
  assign n8460 = ( n8440 & ~n8459 ) | ( n8440 & n8458 ) | ( ~n8459 & n8458 ) ;
  assign n8464 = ~n136 & x123 ;
  assign n8461 = ( x121 & ~n150 ) | ( x121 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n8462 = ( x122 & ~n131 ) | ( x122 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n8463 = n8461 | n8462 ;
  assign n8465 = ( x123 & ~n8464 ) | ( x123 & n8463 ) | ( ~n8464 & n8463 ) ;
  assign n8466 = ( x121 & x122 ) | ( x121 & n8448 ) | ( x122 & n8448 ) ;
  assign n8467 = x122 | x123 ;
  assign n8468 = x122 &  x123 ;
  assign n8469 = ( n8467 & ~n8468 ) | ( n8467 & 1'b0 ) | ( ~n8468 & 1'b0 ) ;
  assign n8470 = n8466 &  n8469 ;
  assign n8471 = n8466 | n8469 ;
  assign n8472 = ~n8470 & n8471 ;
  assign n8473 = ~n139 & n8472 ;
  assign n8474 = n8465 | n8473 ;
  assign n8478 = x118 &  n225 ;
  assign n8475 = ( x120 & ~n197 ) | ( x120 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n8476 = x119 &  n192 ;
  assign n8477 = n8475 | n8476 ;
  assign n8479 = ( x118 & ~n8478 ) | ( x118 & n8477 ) | ( ~n8478 & n8477 ) ;
  assign n8480 = ( n7647 & ~n200 ) | ( n7647 & n7907 ) | ( ~n200 & n7907 ) ;
  assign n8481 = ( n8479 & ~n7908 ) | ( n8479 & n8480 ) | ( ~n7908 & n8480 ) ;
  assign n8482 = ( x5 & ~n8481 ) | ( x5 & 1'b0 ) | ( ~n8481 & 1'b0 ) ;
  assign n8483 = ~x5 & n8481 ;
  assign n8484 = n8482 | n8483 ;
  assign n8488 = x112 &  n503 ;
  assign n8485 = ( x114 & ~n450 ) | ( x114 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n8486 = x113 &  n445 ;
  assign n8487 = n8485 | n8486 ;
  assign n8489 = ( x112 & ~n8488 ) | ( x112 & n8487 ) | ( ~n8488 & n8487 ) ;
  assign n8490 = n453 | n6185 ;
  assign n8491 = ~n8489 & n8490 ;
  assign n8492 = ( n8157 & ~n8428 ) | ( n8157 & n8418 ) | ( ~n8428 & n8418 ) ;
  assign n8496 = x109 &  n713 ;
  assign n8493 = ( x111 & ~n641 ) | ( x111 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n8494 = x110 &  n636 ;
  assign n8495 = n8493 | n8494 ;
  assign n8497 = ( x109 & ~n8496 ) | ( x109 & n8495 ) | ( ~n8496 & n8495 ) ;
  assign n8498 = n644 | n5711 ;
  assign n8499 = ~n8497 & n8498 ;
  assign n8500 = x14 &  n8499 ;
  assign n8501 = x14 | n8499 ;
  assign n8502 = ~n8500 & n8501 ;
  assign n8503 = ( n8215 & n8225 ) | ( n8215 & n8415 ) | ( n8225 & n8415 ) ;
  assign n8507 = x106 &  n942 ;
  assign n8504 = ( x108 & ~n896 ) | ( x108 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n8505 = x107 &  n891 ;
  assign n8506 = n8504 | n8505 ;
  assign n8508 = ( x106 & ~n8507 ) | ( x106 & n8506 ) | ( ~n8507 & n8506 ) ;
  assign n8509 = n899 | n5055 ;
  assign n8510 = ~n8508 & n8509 ;
  assign n8511 = x17 &  n8510 ;
  assign n8512 = x17 | n8510 ;
  assign n8513 = ~n8511 & n8512 ;
  assign n8517 = x100 &  n1551 ;
  assign n8514 = ( x102 & ~n1451 ) | ( x102 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n8515 = x101 &  n1446 ;
  assign n8516 = n8514 | n8515 ;
  assign n8518 = ( x100 & ~n8517 ) | ( x100 & n8516 ) | ( ~n8517 & n8516 ) ;
  assign n8519 = n1454 | n3872 ;
  assign n8520 = ~n8518 & n8519 ;
  assign n8521 = x23 &  n8520 ;
  assign n8522 = x23 | n8520 ;
  assign n8523 = ~n8521 & n8522 ;
  assign n8679 = x97 &  n1894 ;
  assign n8676 = ( x99 & ~n1816 ) | ( x99 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n8677 = x98 &  n1811 ;
  assign n8678 = n8676 | n8677 ;
  assign n8680 = ( x97 & ~n8679 ) | ( x97 & n8678 ) | ( ~n8679 & n8678 ) ;
  assign n8681 = ~n1819 & n3338 ;
  assign n8682 = n8680 | n8681 ;
  assign n8683 = ( x26 & ~n8682 ) | ( x26 & 1'b0 ) | ( ~n8682 & 1'b0 ) ;
  assign n8684 = ~x26 & n8682 ;
  assign n8685 = n8683 | n8684 ;
  assign n8527 = x88 &  n3214 ;
  assign n8524 = ( x90 & ~n3087 ) | ( x90 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n8525 = x89 &  n3082 ;
  assign n8526 = n8524 | n8525 ;
  assign n8528 = ( x88 & ~n8527 ) | ( x88 & n8526 ) | ( ~n8527 & n8526 ) ;
  assign n8529 = ( n1976 & ~n3090 ) | ( n1976 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n8530 = n8528 | n8529 ;
  assign n8531 = ( x35 & ~n8530 ) | ( x35 & 1'b0 ) | ( ~n8530 & 1'b0 ) ;
  assign n8532 = ~x35 & n8530 ;
  assign n8533 = n8531 | n8532 ;
  assign n8537 = x79 &  n4934 ;
  assign n8534 = ( x81 & ~n4725 ) | ( x81 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n8535 = x80 &  n4720 ;
  assign n8536 = n8534 | n8535 ;
  assign n8538 = ( x79 & ~n8537 ) | ( x79 & n8536 ) | ( ~n8537 & n8536 ) ;
  assign n8539 = ( n994 & ~n4728 ) | ( n994 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n8540 = n8538 | n8539 ;
  assign n8541 = ( x44 & ~n8540 ) | ( x44 & 1'b0 ) | ( ~n8540 & 1'b0 ) ;
  assign n8542 = ~x44 & n8540 ;
  assign n8543 = n8541 | n8542 ;
  assign n8544 = ( n8094 & n8285 ) | ( n8094 & n8355 ) | ( n8285 & n8355 ) ;
  assign n8604 = x76 &  n5586 ;
  assign n8601 = ( x78 & ~n5389 ) | ( x78 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n8602 = x77 &  n5384 ;
  assign n8603 = n8601 | n8602 ;
  assign n8605 = ( x76 & ~n8604 ) | ( x76 & n8603 ) | ( ~n8604 & n8603 ) ;
  assign n8606 = ( n693 & ~n5392 ) | ( n693 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n8607 = n8605 | n8606 ;
  assign n8608 = ( x47 & ~n8607 ) | ( x47 & 1'b0 ) | ( ~n8607 & 1'b0 ) ;
  assign n8609 = ~x47 & n8607 ;
  assign n8610 = n8608 | n8609 ;
  assign n8548 = x73 &  n6288 ;
  assign n8545 = ( x75 & ~n6032 ) | ( x75 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n8546 = x74 &  n6027 ;
  assign n8547 = n8545 | n8546 ;
  assign n8549 = ( x73 & ~n8548 ) | ( x73 & n8547 ) | ( ~n8548 & n8547 ) ;
  assign n8550 = ( n540 & ~n6035 ) | ( n540 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n8551 = n8549 | n8550 ;
  assign n8552 = ( x50 & ~n8551 ) | ( x50 & 1'b0 ) | ( ~n8551 & 1'b0 ) ;
  assign n8553 = ~x50 & n8551 ;
  assign n8554 = n8552 | n8553 ;
  assign n8555 = ( n8328 & n8338 ) | ( n8328 & n8339 ) | ( n8338 & n8339 ) ;
  assign n8574 = x67 &  n7731 ;
  assign n8571 = ( x69 & ~n7538 ) | ( x69 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n8572 = x68 &  n7533 ;
  assign n8573 = n8571 | n8572 ;
  assign n8575 = ( x67 & ~n8574 ) | ( x67 & n8573 ) | ( ~n8574 & n8573 ) ;
  assign n8576 = ( n246 & ~n7541 ) | ( n246 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n8577 = n8575 | n8576 ;
  assign n8578 = ( x56 & ~n8577 ) | ( x56 & 1'b0 ) | ( ~n8577 & 1'b0 ) ;
  assign n8579 = ~x56 & n8577 ;
  assign n8580 = n8578 | n8579 ;
  assign n8557 = ( x57 & ~x58 ) | ( x57 & n8313 ) | ( ~x58 & n8313 ) ;
  assign n8556 = ( x57 & ~x58 ) | ( x57 & n8044 ) | ( ~x58 & n8044 ) ;
  assign n8558 = ~n8557 |  n8556 ;
  assign n8562 = x64 &  n8558 ;
  assign n8559 = ( x66 & ~n8314 ) | ( x66 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n8560 = x65 &  n8309 ;
  assign n8561 = n8559 | n8560 ;
  assign n8563 = ( x64 & ~n8562 ) | ( x64 & n8561 ) | ( ~n8562 & n8561 ) ;
  assign n8564 = ( n157 & ~n8317 ) | ( n157 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n8565 = n8563 | n8564 ;
  assign n8566 = ( x59 & ~n8045 ) | ( x59 & n8319 ) | ( ~n8045 & n8319 ) ;
  assign n8567 = ~n8319 & n8566 ;
  assign n8568 = ( n8565 & ~x59 ) | ( n8565 & n8567 ) | ( ~x59 & n8567 ) ;
  assign n8569 = ( x59 & ~n8565 ) | ( x59 & n8567 ) | ( ~n8565 & n8567 ) ;
  assign n8570 = ( n8568 & ~n8567 ) | ( n8568 & n8569 ) | ( ~n8567 & n8569 ) ;
  assign n8581 = ( n8324 & ~n8580 ) | ( n8324 & n8570 ) | ( ~n8580 & n8570 ) ;
  assign n8582 = ( n8570 & ~n8324 ) | ( n8570 & n8580 ) | ( ~n8324 & n8580 ) ;
  assign n8583 = ( n8581 & ~n8570 ) | ( n8581 & n8582 ) | ( ~n8570 & n8582 ) ;
  assign n8587 = x70 &  n6982 ;
  assign n8584 = ( x72 & ~n6727 ) | ( x72 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n8585 = x71 &  n6722 ;
  assign n8586 = n8584 | n8585 ;
  assign n8588 = ( x70 & ~n8587 ) | ( x70 & n8586 ) | ( ~n8587 & n8586 ) ;
  assign n8589 = ( n345 & ~n6730 ) | ( n345 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n8590 = n8588 | n8589 ;
  assign n8591 = ( x53 & ~n8590 ) | ( x53 & 1'b0 ) | ( ~n8590 & 1'b0 ) ;
  assign n8592 = ~x53 & n8590 ;
  assign n8593 = n8591 | n8592 ;
  assign n8594 = ( n8583 & ~n8327 ) | ( n8583 & n8593 ) | ( ~n8327 & n8593 ) ;
  assign n8595 = ( n8327 & ~n8593 ) | ( n8327 & n8583 ) | ( ~n8593 & n8583 ) ;
  assign n8596 = ( n8594 & ~n8583 ) | ( n8594 & n8595 ) | ( ~n8583 & n8595 ) ;
  assign n8598 = ( n8554 & n8555 ) | ( n8554 & n8596 ) | ( n8555 & n8596 ) ;
  assign n8597 = ( n8555 & ~n8554 ) | ( n8555 & n8596 ) | ( ~n8554 & n8596 ) ;
  assign n8599 = ( n8554 & ~n8598 ) | ( n8554 & n8597 ) | ( ~n8598 & n8597 ) ;
  assign n8600 = ( n8091 & n8342 ) | ( n8091 & n8352 ) | ( n8342 & n8352 ) ;
  assign n8612 = ( n8599 & n8600 ) | ( n8599 & n8610 ) | ( n8600 & n8610 ) ;
  assign n8611 = ( n8599 & ~n8610 ) | ( n8599 & n8600 ) | ( ~n8610 & n8600 ) ;
  assign n8613 = ( n8610 & ~n8612 ) | ( n8610 & n8611 ) | ( ~n8612 & n8611 ) ;
  assign n8615 = ( n8543 & n8544 ) | ( n8543 & n8613 ) | ( n8544 & n8613 ) ;
  assign n8614 = ( n8544 & ~n8543 ) | ( n8544 & n8613 ) | ( ~n8543 & n8613 ) ;
  assign n8616 = ( n8543 & ~n8615 ) | ( n8543 & n8614 ) | ( ~n8615 & n8614 ) ;
  assign n8617 = ( n8097 & n8358 ) | ( n8097 & n8368 ) | ( n8358 & n8368 ) ;
  assign n8621 = x82 &  n4344 ;
  assign n8618 = ( x84 & ~n4143 ) | ( x84 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n8619 = x83 &  n4138 ;
  assign n8620 = n8618 | n8619 ;
  assign n8622 = ( x82 & ~n8621 ) | ( x82 & n8620 ) | ( ~n8621 & n8620 ) ;
  assign n8623 = ( n1199 & ~n4146 ) | ( n1199 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n8624 = n8622 | n8623 ;
  assign n8625 = ( x41 & ~n8624 ) | ( x41 & 1'b0 ) | ( ~n8624 & 1'b0 ) ;
  assign n8626 = ~x41 & n8624 ;
  assign n8627 = n8625 | n8626 ;
  assign n8628 = ( n8616 & ~n8617 ) | ( n8616 & n8627 ) | ( ~n8617 & n8627 ) ;
  assign n8629 = ( n8616 & ~n8627 ) | ( n8616 & n8617 ) | ( ~n8627 & n8617 ) ;
  assign n8630 = ( n8628 & ~n8616 ) | ( n8628 & n8629 ) | ( ~n8616 & n8629 ) ;
  assign n8631 = ( n8100 & n8275 ) | ( n8100 & n8371 ) | ( n8275 & n8371 ) ;
  assign n8635 = x85 &  n3756 ;
  assign n8632 = ( x87 & ~n3602 ) | ( x87 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n8633 = x86 &  n3597 ;
  assign n8634 = n8632 | n8633 ;
  assign n8636 = ( x85 & ~n8635 ) | ( x85 & n8634 ) | ( ~n8635 & n8634 ) ;
  assign n8637 = ( n1512 & ~n3605 ) | ( n1512 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n8638 = n8636 | n8637 ;
  assign n8639 = ( x38 & ~n8638 ) | ( x38 & 1'b0 ) | ( ~n8638 & 1'b0 ) ;
  assign n8640 = ~x38 & n8638 ;
  assign n8641 = n8639 | n8640 ;
  assign n8642 = ( n8630 & ~n8631 ) | ( n8630 & n8641 ) | ( ~n8631 & n8641 ) ;
  assign n8643 = ( n8630 & ~n8641 ) | ( n8630 & n8631 ) | ( ~n8641 & n8631 ) ;
  assign n8644 = ( n8642 & ~n8630 ) | ( n8642 & n8643 ) | ( ~n8630 & n8643 ) ;
  assign n8645 = ( n8375 & n8533 ) | ( n8375 & n8644 ) | ( n8533 & n8644 ) ;
  assign n8646 = ( n8375 & ~n8533 ) | ( n8375 & n8644 ) | ( ~n8533 & n8644 ) ;
  assign n8647 = ( n8533 & ~n8645 ) | ( n8533 & n8646 ) | ( ~n8645 & n8646 ) ;
  assign n8648 = ( n8377 & n8378 ) | ( n8377 & n8388 ) | ( n8378 & n8388 ) ;
  assign n8652 = x91 &  n2718 ;
  assign n8649 = ( x93 & ~n2642 ) | ( x93 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n8650 = x92 &  n2637 ;
  assign n8651 = n8649 | n8650 ;
  assign n8653 = ( x91 & ~n8652 ) | ( x91 & n8651 ) | ( ~n8652 & n8651 ) ;
  assign n8654 = n2264 | n2645 ;
  assign n8655 = ~n8653 & n8654 ;
  assign n8656 = x32 &  n8655 ;
  assign n8657 = x32 | n8655 ;
  assign n8658 = ~n8656 & n8657 ;
  assign n8659 = ( n8647 & n8648 ) | ( n8647 & n8658 ) | ( n8648 & n8658 ) ;
  assign n8660 = ( n8648 & ~n8647 ) | ( n8648 & n8658 ) | ( ~n8647 & n8658 ) ;
  assign n8661 = ( n8647 & ~n8659 ) | ( n8647 & n8660 ) | ( ~n8659 & n8660 ) ;
  assign n8666 = x94 &  n2312 ;
  assign n8663 = ( x96 & ~n2195 ) | ( x96 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n8664 = x95 &  n2190 ;
  assign n8665 = n8663 | n8664 ;
  assign n8667 = ( x94 & ~n8666 ) | ( x94 & n8665 ) | ( ~n8666 & n8665 ) ;
  assign n8668 = ~n2198 & n2836 ;
  assign n8669 = n8667 | n8668 ;
  assign n8670 = ( x29 & ~n8669 ) | ( x29 & 1'b0 ) | ( ~n8669 & 1'b0 ) ;
  assign n8671 = ~x29 & n8669 ;
  assign n8672 = n8670 | n8671 ;
  assign n8662 = ( n8121 & n8391 ) | ( n8121 & n8401 ) | ( n8391 & n8401 ) ;
  assign n8673 = ( n8661 & ~n8672 ) | ( n8661 & n8662 ) | ( ~n8672 & n8662 ) ;
  assign n8674 = ( n8661 & ~n8662 ) | ( n8661 & n8672 ) | ( ~n8662 & n8672 ) ;
  assign n8675 = ( n8673 & ~n8661 ) | ( n8673 & n8674 ) | ( ~n8661 & n8674 ) ;
  assign n8686 = ( n8406 & ~n8685 ) | ( n8406 & n8675 ) | ( ~n8685 & n8675 ) ;
  assign n8687 = ( n8675 & ~n8406 ) | ( n8675 & n8685 ) | ( ~n8406 & n8685 ) ;
  assign n8688 = ( n8686 & ~n8675 ) | ( n8686 & n8687 ) | ( ~n8675 & n8687 ) ;
  assign n8689 = ( n8410 & n8523 ) | ( n8410 & n8688 ) | ( n8523 & n8688 ) ;
  assign n8690 = ( n8410 & ~n8523 ) | ( n8410 & n8688 ) | ( ~n8523 & n8688 ) ;
  assign n8691 = ( n8523 & ~n8689 ) | ( n8523 & n8690 ) | ( ~n8689 & n8690 ) ;
  assign n8695 = x103 &  n1227 ;
  assign n8692 = ( x105 & ~n1154 ) | ( x105 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n8693 = x104 &  n1149 ;
  assign n8694 = n8692 | n8693 ;
  assign n8696 = ( x103 & ~n8695 ) | ( x103 & n8694 ) | ( ~n8695 & n8694 ) ;
  assign n8697 = ~n1157 & n4442 ;
  assign n8698 = n8696 | n8697 ;
  assign n8699 = ( x20 & ~n8698 ) | ( x20 & 1'b0 ) | ( ~n8698 & 1'b0 ) ;
  assign n8700 = ~x20 & n8698 ;
  assign n8701 = n8699 | n8700 ;
  assign n8702 = ( n8413 & n8691 ) | ( n8413 & n8701 ) | ( n8691 & n8701 ) ;
  assign n8703 = ( n8413 & ~n8691 ) | ( n8413 & n8701 ) | ( ~n8691 & n8701 ) ;
  assign n8704 = ( n8691 & ~n8702 ) | ( n8691 & n8703 ) | ( ~n8702 & n8703 ) ;
  assign n8705 = ( n8503 & ~n8513 ) | ( n8503 & n8704 ) | ( ~n8513 & n8704 ) ;
  assign n8706 = ( n8503 & ~n8704 ) | ( n8503 & n8513 ) | ( ~n8704 & n8513 ) ;
  assign n8707 = ( n8705 & ~n8503 ) | ( n8705 & n8706 ) | ( ~n8503 & n8706 ) ;
  assign n8709 = ( n8492 & n8502 ) | ( n8492 & n8707 ) | ( n8502 & n8707 ) ;
  assign n8708 = ( n8502 & ~n8492 ) | ( n8502 & n8707 ) | ( ~n8492 & n8707 ) ;
  assign n8710 = ( n8492 & ~n8709 ) | ( n8492 & n8708 ) | ( ~n8709 & n8708 ) ;
  assign n8711 = ( n8491 & ~x11 ) | ( n8491 & n8710 ) | ( ~x11 & n8710 ) ;
  assign n8712 = ( x11 & ~n8491 ) | ( x11 & n8710 ) | ( ~n8491 & n8710 ) ;
  assign n8713 = ( n8711 & ~n8710 ) | ( n8711 & n8712 ) | ( ~n8710 & n8712 ) ;
  assign n8717 = x115 &  n353 ;
  assign n8714 = ( x117 & ~n313 ) | ( x117 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n8715 = x116 &  n308 ;
  assign n8716 = n8714 | n8715 ;
  assign n8718 = ( x115 & ~n8717 ) | ( x115 & n8716 ) | ( ~n8717 & n8716 ) ;
  assign n8719 = n316 | n7136 ;
  assign n8720 = ~n8718 & n8719 ;
  assign n8721 = x8 | n8720 ;
  assign n8722 = ~x8 & n8720 ;
  assign n8723 = ( n8721 & ~n8720 ) | ( n8721 & n8722 ) | ( ~n8720 & n8722 ) ;
  assign n8724 = ( n8433 & ~n8713 ) | ( n8433 & n8723 ) | ( ~n8713 & n8723 ) ;
  assign n8725 = ( n8713 & ~n8433 ) | ( n8713 & n8723 ) | ( ~n8433 & n8723 ) ;
  assign n8726 = ( n8724 & ~n8723 ) | ( n8724 & n8725 ) | ( ~n8723 & n8725 ) ;
  assign n8727 = ( n8435 & ~n8484 ) | ( n8435 & n8726 ) | ( ~n8484 & n8726 ) ;
  assign n8728 = ( n8435 & ~n8726 ) | ( n8435 & n8484 ) | ( ~n8726 & n8484 ) ;
  assign n8729 = ( n8727 & ~n8435 ) | ( n8727 & n8728 ) | ( ~n8435 & n8728 ) ;
  assign n8730 = ( x2 & ~n8474 ) | ( x2 & n8729 ) | ( ~n8474 & n8729 ) ;
  assign n8731 = ( x2 & ~n8729 ) | ( x2 & n8474 ) | ( ~n8729 & n8474 ) ;
  assign n8732 = ( n8730 & ~x2 ) | ( n8730 & n8731 ) | ( ~x2 & n8731 ) ;
  assign n8733 = ( n8438 & ~n8458 ) | ( n8438 & n8732 ) | ( ~n8458 & n8732 ) ;
  assign n8734 = ( n8438 & ~n8732 ) | ( n8438 & n8458 ) | ( ~n8732 & n8458 ) ;
  assign n8735 = ( n8733 & ~n8438 ) | ( n8733 & n8734 ) | ( ~n8438 & n8734 ) ;
  assign n8736 = n8435 &  n8726 ;
  assign n8737 = n8435 | n8726 ;
  assign n8738 = ~n8736 & n8737 ;
  assign n8739 = ( x2 & ~n8474 ) | ( x2 & 1'b0 ) | ( ~n8474 & 1'b0 ) ;
  assign n8740 = ~x2 & n8474 ;
  assign n8741 = n8739 | n8740 ;
  assign n8742 = ( n8484 & n8738 ) | ( n8484 & n8741 ) | ( n8738 & n8741 ) ;
  assign n8743 = ( n8438 & n8458 ) | ( n8438 & n8732 ) | ( n8458 & n8732 ) ;
  assign n8760 = x11 &  n8491 ;
  assign n8761 = x11 | n8491 ;
  assign n8762 = ~n8760 & n8761 ;
  assign n8764 = ( n8433 & ~n8710 ) | ( n8433 & n8762 ) | ( ~n8710 & n8762 ) ;
  assign n8780 = x113 &  n503 ;
  assign n8777 = ( x115 & ~n450 ) | ( x115 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n8778 = x114 &  n445 ;
  assign n8779 = n8777 | n8778 ;
  assign n8781 = ( x113 & ~n8780 ) | ( x113 & n8779 ) | ( ~n8780 & n8779 ) ;
  assign n8782 = ~n453 & n6420 ;
  assign n8783 = n8781 | n8782 ;
  assign n8784 = ( x11 & ~n8783 ) | ( x11 & 1'b0 ) | ( ~n8783 & 1'b0 ) ;
  assign n8785 = ~x11 & n8783 ;
  assign n8786 = n8784 | n8785 ;
  assign n8790 = x110 &  n713 ;
  assign n8787 = ( x112 & ~n641 ) | ( x112 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n8788 = x111 &  n636 ;
  assign n8789 = n8787 | n8788 ;
  assign n8791 = ( x110 & ~n8790 ) | ( x110 & n8789 ) | ( ~n8790 & n8789 ) ;
  assign n8792 = ~n644 & n5727 ;
  assign n8793 = n8791 | n8792 ;
  assign n8794 = ( x14 & ~n8793 ) | ( x14 & 1'b0 ) | ( ~n8793 & 1'b0 ) ;
  assign n8795 = ~x14 & n8793 ;
  assign n8796 = n8794 | n8795 ;
  assign n8830 = x86 &  n3756 ;
  assign n8827 = ( x88 & ~n3602 ) | ( x88 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n8828 = x87 &  n3597 ;
  assign n8829 = n8827 | n8828 ;
  assign n8831 = ( x86 & ~n8830 ) | ( x86 & n8829 ) | ( ~n8830 & n8829 ) ;
  assign n8832 = ( n1624 & ~n3605 ) | ( n1624 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n8833 = n8831 | n8832 ;
  assign n8834 = ( x38 & ~n8833 ) | ( x38 & 1'b0 ) | ( ~n8833 & 1'b0 ) ;
  assign n8835 = ~x38 & n8833 ;
  assign n8836 = n8834 | n8835 ;
  assign n8840 = x83 &  n4344 ;
  assign n8837 = ( x85 & ~n4143 ) | ( x85 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n8838 = x84 &  n4138 ;
  assign n8839 = n8837 | n8838 ;
  assign n8841 = ( x83 & ~n8840 ) | ( x83 & n8839 ) | ( ~n8840 & n8839 ) ;
  assign n8842 = ( n1295 & ~n4146 ) | ( n1295 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n8843 = n8841 | n8842 ;
  assign n8844 = ( x41 & ~n8843 ) | ( x41 & 1'b0 ) | ( ~n8843 & 1'b0 ) ;
  assign n8845 = ~x41 & n8843 ;
  assign n8846 = n8844 | n8845 ;
  assign n8847 = ( n8616 & n8617 ) | ( n8616 & n8627 ) | ( n8617 & n8627 ) ;
  assign n8851 = x80 &  n4934 ;
  assign n8848 = ( x82 & ~n4725 ) | ( x82 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n8849 = x81 &  n4720 ;
  assign n8850 = n8848 | n8849 ;
  assign n8852 = ( x80 & ~n8851 ) | ( x80 & n8850 ) | ( ~n8851 & n8850 ) ;
  assign n8853 = ( n1084 & ~n4728 ) | ( n1084 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n8854 = n8852 | n8853 ;
  assign n8855 = ( x44 & ~n8854 ) | ( x44 & 1'b0 ) | ( ~n8854 & 1'b0 ) ;
  assign n8856 = ~x44 & n8854 ;
  assign n8857 = n8855 | n8856 ;
  assign n8861 = x77 &  n5586 ;
  assign n8858 = ( x79 & ~n5389 ) | ( x79 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n8859 = x78 &  n5384 ;
  assign n8860 = n8858 | n8859 ;
  assign n8862 = ( x77 & ~n8861 ) | ( x77 & n8860 ) | ( ~n8861 & n8860 ) ;
  assign n8863 = ( n766 & ~n5392 ) | ( n766 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n8864 = n8862 | n8863 ;
  assign n8865 = ( x47 & ~n8864 ) | ( x47 & 1'b0 ) | ( ~n8864 & 1'b0 ) ;
  assign n8866 = ~x47 & n8864 ;
  assign n8867 = n8865 | n8866 ;
  assign n8871 = x74 &  n6288 ;
  assign n8868 = ( x76 & ~n6032 ) | ( x76 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n8869 = x75 &  n6027 ;
  assign n8870 = n8868 | n8869 ;
  assign n8872 = ( x74 & ~n8871 ) | ( x74 & n8870 ) | ( ~n8871 & n8870 ) ;
  assign n8873 = ( n603 & ~n6035 ) | ( n603 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n8874 = n8872 | n8873 ;
  assign n8875 = ( x50 & ~n8874 ) | ( x50 & 1'b0 ) | ( ~n8874 & 1'b0 ) ;
  assign n8876 = ~x50 & n8874 ;
  assign n8877 = n8875 | n8876 ;
  assign n8878 = ( x59 & ~x60 ) | ( x59 & 1'b0 ) | ( ~x60 & 1'b0 ) ;
  assign n8879 = ~x59 & x60 ;
  assign n8880 = n8878 | n8879 ;
  assign n8881 = x64 &  n8880 ;
  assign n8882 = ( n8045 & ~n8319 ) | ( n8045 & n8565 ) | ( ~n8319 & n8565 ) ;
  assign n8883 = ( x59 & n8319 ) | ( x59 & n8882 ) | ( n8319 & n8882 ) ;
  assign n8884 = ( x59 & ~n8883 ) | ( x59 & 1'b0 ) | ( ~n8883 & 1'b0 ) ;
  assign n8888 = x65 &  n8558 ;
  assign n8885 = ( x67 & ~n8314 ) | ( x67 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n8886 = x66 &  n8309 ;
  assign n8887 = n8885 | n8886 ;
  assign n8889 = ( x65 & ~n8888 ) | ( x65 & n8887 ) | ( ~n8888 & n8887 ) ;
  assign n8890 = n173 | n8317 ;
  assign n8891 = ~n8889 & n8890 ;
  assign n8892 = x59 &  n8891 ;
  assign n8893 = x59 | n8891 ;
  assign n8894 = ~n8892 & n8893 ;
  assign n8895 = ( n8881 & ~n8884 ) | ( n8881 & n8894 ) | ( ~n8884 & n8894 ) ;
  assign n8896 = ( n8881 & ~n8894 ) | ( n8881 & n8884 ) | ( ~n8894 & n8884 ) ;
  assign n8897 = ( n8895 & ~n8881 ) | ( n8895 & n8896 ) | ( ~n8881 & n8896 ) ;
  assign n8898 = ( n8324 & n8570 ) | ( n8324 & n8580 ) | ( n8570 & n8580 ) ;
  assign n8902 = x68 &  n7731 ;
  assign n8899 = ( x70 & ~n7538 ) | ( x70 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n8900 = x69 &  n7533 ;
  assign n8901 = n8899 | n8900 ;
  assign n8903 = ( x68 & ~n8902 ) | ( x68 & n8901 ) | ( ~n8902 & n8901 ) ;
  assign n8904 = ( n282 & ~n7541 ) | ( n282 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n8905 = n8903 | n8904 ;
  assign n8906 = ( x56 & ~n8905 ) | ( x56 & 1'b0 ) | ( ~n8905 & 1'b0 ) ;
  assign n8907 = ~x56 & n8905 ;
  assign n8908 = n8906 | n8907 ;
  assign n8909 = ( n8897 & ~n8898 ) | ( n8897 & n8908 ) | ( ~n8898 & n8908 ) ;
  assign n8910 = ( n8898 & ~n8897 ) | ( n8898 & n8908 ) | ( ~n8897 & n8908 ) ;
  assign n8911 = ( n8909 & ~n8908 ) | ( n8909 & n8910 ) | ( ~n8908 & n8910 ) ;
  assign n8916 = x71 &  n6982 ;
  assign n8913 = ( x73 & ~n6727 ) | ( x73 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n8914 = x72 &  n6722 ;
  assign n8915 = n8913 | n8914 ;
  assign n8917 = ( x71 & ~n8916 ) | ( x71 & n8915 ) | ( ~n8916 & n8915 ) ;
  assign n8918 = ( n389 & ~n6730 ) | ( n389 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n8919 = n8917 | n8918 ;
  assign n8920 = ( x53 & ~n8919 ) | ( x53 & 1'b0 ) | ( ~n8919 & 1'b0 ) ;
  assign n8921 = ~x53 & n8919 ;
  assign n8922 = n8920 | n8921 ;
  assign n8912 = ( n8327 & n8583 ) | ( n8327 & n8593 ) | ( n8583 & n8593 ) ;
  assign n8923 = ( n8911 & ~n8922 ) | ( n8911 & n8912 ) | ( ~n8922 & n8912 ) ;
  assign n8924 = ( n8911 & ~n8912 ) | ( n8911 & n8922 ) | ( ~n8912 & n8922 ) ;
  assign n8925 = ( n8923 & ~n8911 ) | ( n8923 & n8924 ) | ( ~n8911 & n8924 ) ;
  assign n8926 = ( n8877 & ~n8598 ) | ( n8877 & n8925 ) | ( ~n8598 & n8925 ) ;
  assign n8927 = ( n8598 & ~n8925 ) | ( n8598 & n8877 ) | ( ~n8925 & n8877 ) ;
  assign n8928 = ( n8926 & ~n8877 ) | ( n8926 & n8927 ) | ( ~n8877 & n8927 ) ;
  assign n8929 = ( n8867 & ~n8612 ) | ( n8867 & n8928 ) | ( ~n8612 & n8928 ) ;
  assign n8930 = ( n8612 & ~n8928 ) | ( n8612 & n8867 ) | ( ~n8928 & n8867 ) ;
  assign n8931 = ( n8929 & ~n8867 ) | ( n8929 & n8930 ) | ( ~n8867 & n8930 ) ;
  assign n8932 = ( n8857 & ~n8615 ) | ( n8857 & n8931 ) | ( ~n8615 & n8931 ) ;
  assign n8933 = ( n8615 & ~n8931 ) | ( n8615 & n8857 ) | ( ~n8931 & n8857 ) ;
  assign n8934 = ( n8932 & ~n8857 ) | ( n8932 & n8933 ) | ( ~n8857 & n8933 ) ;
  assign n8935 = ( n8846 & ~n8847 ) | ( n8846 & n8934 ) | ( ~n8847 & n8934 ) ;
  assign n8936 = ( n8846 & ~n8934 ) | ( n8846 & n8847 ) | ( ~n8934 & n8847 ) ;
  assign n8937 = ( n8935 & ~n8846 ) | ( n8935 & n8936 ) | ( ~n8846 & n8936 ) ;
  assign n8938 = ( n8630 & n8631 ) | ( n8630 & n8641 ) | ( n8631 & n8641 ) ;
  assign n8939 = ( n8836 & ~n8937 ) | ( n8836 & n8938 ) | ( ~n8937 & n8938 ) ;
  assign n8940 = ( n8836 & ~n8938 ) | ( n8836 & n8937 ) | ( ~n8938 & n8937 ) ;
  assign n8941 = ( n8939 & ~n8836 ) | ( n8939 & n8940 ) | ( ~n8836 & n8940 ) ;
  assign n8820 = x89 &  n3214 ;
  assign n8817 = ( x91 & ~n3087 ) | ( x91 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n8818 = x90 &  n3082 ;
  assign n8819 = n8817 | n8818 ;
  assign n8821 = ( x89 & ~n8820 ) | ( x89 & n8819 ) | ( ~n8820 & n8819 ) ;
  assign n8822 = ( n2108 & ~n3090 ) | ( n2108 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n8823 = n8821 | n8822 ;
  assign n8824 = ( x35 & ~n8823 ) | ( x35 & 1'b0 ) | ( ~n8823 & 1'b0 ) ;
  assign n8825 = ~x35 & n8823 ;
  assign n8826 = n8824 | n8825 ;
  assign n8942 = ( n8645 & ~n8941 ) | ( n8645 & n8826 ) | ( ~n8941 & n8826 ) ;
  assign n8943 = ( n8826 & ~n8645 ) | ( n8826 & n8941 ) | ( ~n8645 & n8941 ) ;
  assign n8944 = ( n8942 & ~n8826 ) | ( n8942 & n8943 ) | ( ~n8826 & n8943 ) ;
  assign n8945 = ( n8647 & ~n8658 ) | ( n8647 & n8648 ) | ( ~n8658 & n8648 ) ;
  assign n8949 = x92 &  n2718 ;
  assign n8946 = ( x94 & ~n2642 ) | ( x94 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n8947 = x93 &  n2637 ;
  assign n8948 = n8946 | n8947 ;
  assign n8950 = ( x92 & ~n8949 ) | ( x92 & n8948 ) | ( ~n8949 & n8948 ) ;
  assign n8951 = ( n2401 & ~n2645 ) | ( n2401 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n8952 = n8950 | n8951 ;
  assign n8953 = ( x32 & ~n8952 ) | ( x32 & 1'b0 ) | ( ~n8952 & 1'b0 ) ;
  assign n8954 = ~x32 & n8952 ;
  assign n8955 = n8953 | n8954 ;
  assign n8956 = ( n8944 & ~n8945 ) | ( n8944 & n8955 ) | ( ~n8945 & n8955 ) ;
  assign n8957 = ( n8944 & ~n8955 ) | ( n8944 & n8945 ) | ( ~n8955 & n8945 ) ;
  assign n8958 = ( n8956 & ~n8944 ) | ( n8956 & n8957 ) | ( ~n8944 & n8957 ) ;
  assign n8959 = ( n8662 & ~n8661 ) | ( n8662 & n8672 ) | ( ~n8661 & n8672 ) ;
  assign n8963 = x95 &  n2312 ;
  assign n8960 = ( x97 & ~n2195 ) | ( x97 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n8961 = x96 &  n2190 ;
  assign n8962 = n8960 | n8961 ;
  assign n8964 = ( x95 & ~n8963 ) | ( x95 & n8962 ) | ( ~n8963 & n8962 ) ;
  assign n8965 = ~n2198 & n2999 ;
  assign n8966 = n8964 | n8965 ;
  assign n8967 = ( x29 & ~n8966 ) | ( x29 & 1'b0 ) | ( ~n8966 & 1'b0 ) ;
  assign n8968 = ~x29 & n8966 ;
  assign n8969 = n8967 | n8968 ;
  assign n8970 = ( n8958 & ~n8959 ) | ( n8958 & n8969 ) | ( ~n8959 & n8969 ) ;
  assign n8971 = ( n8959 & ~n8958 ) | ( n8959 & n8969 ) | ( ~n8958 & n8969 ) ;
  assign n8972 = ( n8970 & ~n8969 ) | ( n8970 & n8971 ) | ( ~n8969 & n8971 ) ;
  assign n8973 = ( n8406 & ~n8675 ) | ( n8406 & n8685 ) | ( ~n8675 & n8685 ) ;
  assign n8977 = x98 &  n1894 ;
  assign n8974 = ( x100 & ~n1816 ) | ( x100 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n8975 = x99 &  n1811 ;
  assign n8976 = n8974 | n8975 ;
  assign n8978 = ( x98 & ~n8977 ) | ( x98 & n8976 ) | ( ~n8977 & n8976 ) ;
  assign n8979 = n1819 | n3354 ;
  assign n8980 = ~n8978 & n8979 ;
  assign n8981 = x26 &  n8980 ;
  assign n8982 = x26 | n8980 ;
  assign n8983 = ~n8981 & n8982 ;
  assign n8984 = ( n8972 & n8973 ) | ( n8972 & n8983 ) | ( n8973 & n8983 ) ;
  assign n8985 = ( n8973 & ~n8972 ) | ( n8973 & n8983 ) | ( ~n8972 & n8983 ) ;
  assign n8986 = ( n8972 & ~n8984 ) | ( n8972 & n8985 ) | ( ~n8984 & n8985 ) ;
  assign n8810 = x101 &  n1551 ;
  assign n8807 = ( x103 & ~n1451 ) | ( x103 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n8808 = x102 &  n1446 ;
  assign n8809 = n8807 | n8808 ;
  assign n8811 = ( x101 & ~n8810 ) | ( x101 & n8809 ) | ( ~n8810 & n8809 ) ;
  assign n8812 = n1454 | n4056 ;
  assign n8813 = ~n8811 & n8812 ;
  assign n8814 = x23 &  n8813 ;
  assign n8815 = x23 | n8813 ;
  assign n8816 = ~n8814 & n8815 ;
  assign n8987 = ( n8689 & ~n8986 ) | ( n8689 & n8816 ) | ( ~n8986 & n8816 ) ;
  assign n8988 = ( n8816 & ~n8689 ) | ( n8816 & n8986 ) | ( ~n8689 & n8986 ) ;
  assign n8989 = ( n8987 & ~n8816 ) | ( n8987 & n8988 ) | ( ~n8816 & n8988 ) ;
  assign n8990 = ( n8413 & ~n8701 ) | ( n8413 & n8691 ) | ( ~n8701 & n8691 ) ;
  assign n8994 = x104 &  n1227 ;
  assign n8991 = ( x106 & ~n1154 ) | ( x106 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n8992 = x105 &  n1149 ;
  assign n8993 = n8991 | n8992 ;
  assign n8995 = ( x104 & ~n8994 ) | ( x104 & n8993 ) | ( ~n8994 & n8993 ) ;
  assign n8996 = ~n1157 & n4458 ;
  assign n8997 = n8995 | n8996 ;
  assign n8998 = ( x20 & ~n8997 ) | ( x20 & 1'b0 ) | ( ~n8997 & 1'b0 ) ;
  assign n8999 = ~x20 & n8997 ;
  assign n9000 = n8998 | n8999 ;
  assign n9002 = ( n8989 & n8990 ) | ( n8989 & n9000 ) | ( n8990 & n9000 ) ;
  assign n9001 = ( n8990 & ~n8989 ) | ( n8990 & n9000 ) | ( ~n8989 & n9000 ) ;
  assign n9003 = ( n8989 & ~n9002 ) | ( n8989 & n9001 ) | ( ~n9002 & n9001 ) ;
  assign n8800 = x107 &  n942 ;
  assign n8797 = ( x109 & ~n896 ) | ( x109 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n8798 = x108 &  n891 ;
  assign n8799 = n8797 | n8798 ;
  assign n8801 = ( x107 & ~n8800 ) | ( x107 & n8799 ) | ( ~n8800 & n8799 ) ;
  assign n8802 = ~n899 & n5267 ;
  assign n8803 = n8801 | n8802 ;
  assign n8804 = ( x17 & ~n8803 ) | ( x17 & 1'b0 ) | ( ~n8803 & 1'b0 ) ;
  assign n8805 = ~x17 & n8803 ;
  assign n8806 = n8804 | n8805 ;
  assign n9005 = ( n8705 & n8806 ) | ( n8705 & n9003 ) | ( n8806 & n9003 ) ;
  assign n9004 = ( n8705 & ~n9003 ) | ( n8705 & n8806 ) | ( ~n9003 & n8806 ) ;
  assign n9006 = ( n9003 & ~n9005 ) | ( n9003 & n9004 ) | ( ~n9005 & n9004 ) ;
  assign n9007 = ( n8708 & ~n8796 ) | ( n8708 & n9006 ) | ( ~n8796 & n9006 ) ;
  assign n9008 = ( n8796 & ~n8708 ) | ( n8796 & n9006 ) | ( ~n8708 & n9006 ) ;
  assign n9009 = ( n9007 & ~n9006 ) | ( n9007 & n9008 ) | ( ~n9006 & n9008 ) ;
  assign n9010 = ( n8786 & ~n9009 ) | ( n8786 & 1'b0 ) | ( ~n9009 & 1'b0 ) ;
  assign n9011 = ~n8786 & n9009 ;
  assign n9012 = n9010 | n9011 ;
  assign n8770 = x116 &  n353 ;
  assign n8767 = ( x118 & ~n313 ) | ( x118 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n8768 = x117 &  n308 ;
  assign n8769 = n8767 | n8768 ;
  assign n8771 = ( x116 & ~n8770 ) | ( x116 & n8769 ) | ( ~n8770 & n8769 ) ;
  assign n8772 = ( n316 & ~n7152 ) | ( n316 & n8771 ) | ( ~n7152 & n8771 ) ;
  assign n8773 = n7152 | n8772 ;
  assign n8775 = ( x8 & n8771 ) | ( x8 & n8773 ) | ( n8771 & n8773 ) ;
  assign n8774 = ( x8 & ~n8773 ) | ( x8 & n8771 ) | ( ~n8773 & n8771 ) ;
  assign n8776 = ( n8773 & ~n8775 ) | ( n8773 & n8774 ) | ( ~n8775 & n8774 ) ;
  assign n9013 = ( n8764 & ~n9012 ) | ( n8764 & n8776 ) | ( ~n9012 & n8776 ) ;
  assign n9014 = ( n8776 & ~n8764 ) | ( n8776 & n9012 ) | ( ~n8764 & n9012 ) ;
  assign n9015 = ( n9013 & ~n8776 ) | ( n9013 & n9014 ) | ( ~n8776 & n9014 ) ;
  assign n8763 = ( n8710 & ~n8433 ) | ( n8710 & n8762 ) | ( ~n8433 & n8762 ) ;
  assign n8765 = ( n8763 & ~n8762 ) | ( n8763 & n8764 ) | ( ~n8762 & n8764 ) ;
  assign n8758 = ( x8 & ~n8720 ) | ( x8 & 1'b0 ) | ( ~n8720 & 1'b0 ) ;
  assign n8759 = ( n8721 & ~x8 ) | ( n8721 & n8758 ) | ( ~x8 & n8758 ) ;
  assign n8766 = ( n8435 & ~n8765 ) | ( n8435 & n8759 ) | ( ~n8765 & n8759 ) ;
  assign n9019 = x119 &  n225 ;
  assign n9016 = ( x121 & ~n197 ) | ( x121 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n9017 = x120 &  n192 ;
  assign n9018 = n9016 | n9017 ;
  assign n9020 = ( x119 & ~n9019 ) | ( x119 & n9018 ) | ( ~n9019 & n9018 ) ;
  assign n9021 = ~n200 & n8176 ;
  assign n9022 = n9020 | n9021 ;
  assign n9023 = ~x5 & n9022 ;
  assign n9024 = x5 | n9022 ;
  assign n9025 = ( n9023 & ~n9022 ) | ( n9023 & n9024 ) | ( ~n9022 & n9024 ) ;
  assign n9026 = ( n9015 & ~n8766 ) | ( n9015 & n9025 ) | ( ~n8766 & n9025 ) ;
  assign n9027 = ( n8766 & ~n9015 ) | ( n8766 & n9025 ) | ( ~n9015 & n9025 ) ;
  assign n9028 = ( n9026 & ~n9025 ) | ( n9026 & n9027 ) | ( ~n9025 & n9027 ) ;
  assign n8747 = ~n136 & x124 ;
  assign n8744 = ( x122 & ~n150 ) | ( x122 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n8745 = ( x123 & ~n131 ) | ( x123 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n8746 = n8744 | n8745 ;
  assign n8748 = ( x124 & ~n8747 ) | ( x124 & n8746 ) | ( ~n8747 & n8746 ) ;
  assign n8749 = ( x122 & x123 ) | ( x122 & n8466 ) | ( x123 & n8466 ) ;
  assign n8750 = x123 | x124 ;
  assign n8751 = x123 &  x124 ;
  assign n8752 = ( n8750 & ~n8751 ) | ( n8750 & 1'b0 ) | ( ~n8751 & 1'b0 ) ;
  assign n8753 = n8749 &  n8752 ;
  assign n8754 = n8749 | n8752 ;
  assign n8755 = ~n8753 & n8754 ;
  assign n8756 = ~n139 & n8755 ;
  assign n8757 = n8748 | n8756 ;
  assign n9029 = ( x2 & n8757 ) | ( x2 & n9028 ) | ( n8757 & n9028 ) ;
  assign n9030 = ( x2 & ~n9028 ) | ( x2 & n8757 ) | ( ~n9028 & n8757 ) ;
  assign n9031 = ( n9028 & ~n9029 ) | ( n9028 & n9030 ) | ( ~n9029 & n9030 ) ;
  assign n9032 = ( n8742 & ~n8743 ) | ( n8742 & n9031 ) | ( ~n8743 & n9031 ) ;
  assign n9033 = ( n8742 & ~n9031 ) | ( n8742 & n8743 ) | ( ~n9031 & n8743 ) ;
  assign n9034 = ( n9032 & ~n8742 ) | ( n9032 & n9033 ) | ( ~n8742 & n9033 ) ;
  assign n9035 = ( x2 & ~n8757 ) | ( x2 & 1'b0 ) | ( ~n8757 & 1'b0 ) ;
  assign n9036 = ~x2 & n8757 ;
  assign n9037 = n9035 | n9036 ;
  assign n9040 = n8766 &  n9015 ;
  assign n9041 = n8766 | n9015 ;
  assign n9042 = ~n9040 & n9041 ;
  assign n9038 = x5 &  n9022 ;
  assign n9039 = ( x5 & ~n9038 ) | ( x5 & n9023 ) | ( ~n9038 & n9023 ) ;
  assign n9043 = ( n9037 & ~n9042 ) | ( n9037 & n9039 ) | ( ~n9042 & n9039 ) ;
  assign n9044 = ( n8786 & ~n8764 ) | ( n8786 & n9009 ) | ( ~n8764 & n9009 ) ;
  assign n9058 = x111 &  n713 ;
  assign n9055 = ( x113 & ~n641 ) | ( x113 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n9056 = x112 &  n636 ;
  assign n9057 = n9055 | n9056 ;
  assign n9059 = ( x111 & ~n9058 ) | ( x111 & n9057 ) | ( ~n9058 & n9057 ) ;
  assign n9060 = n644 | n6169 ;
  assign n9061 = ~n9059 & n9060 ;
  assign n9075 = x99 &  n1894 ;
  assign n9072 = ( x101 & ~n1816 ) | ( x101 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n9073 = x100 &  n1811 ;
  assign n9074 = n9072 | n9073 ;
  assign n9076 = ( x99 & ~n9075 ) | ( x99 & n9074 ) | ( ~n9075 & n9074 ) ;
  assign n9077 = n1819 | n3694 ;
  assign n9078 = ~n9076 & n9077 ;
  assign n9079 = x26 &  n9078 ;
  assign n9080 = x26 | n9078 ;
  assign n9081 = ~n9079 & n9080 ;
  assign n9085 = x90 &  n3214 ;
  assign n9082 = ( x92 & ~n3087 ) | ( x92 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n9083 = x91 &  n3082 ;
  assign n9084 = n9082 | n9083 ;
  assign n9086 = ( x90 & ~n9085 ) | ( x90 & n9084 ) | ( ~n9085 & n9084 ) ;
  assign n9087 = ( n2248 & ~n3090 ) | ( n2248 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n9088 = n9086 | n9087 ;
  assign n9089 = ( x35 & ~n9088 ) | ( x35 & 1'b0 ) | ( ~n9088 & 1'b0 ) ;
  assign n9090 = ~x35 & n9088 ;
  assign n9091 = n9089 | n9090 ;
  assign n9095 = x87 &  n3756 ;
  assign n9092 = ( x89 & ~n3602 ) | ( x89 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n9093 = x88 &  n3597 ;
  assign n9094 = n9092 | n9093 ;
  assign n9096 = ( x87 & ~n9095 ) | ( x87 & n9094 ) | ( ~n9095 & n9094 ) ;
  assign n9097 = ( n1741 & ~n3605 ) | ( n1741 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n9098 = n9096 | n9097 ;
  assign n9099 = ( x38 & ~n9098 ) | ( x38 & 1'b0 ) | ( ~n9098 & 1'b0 ) ;
  assign n9100 = ~x38 & n9098 ;
  assign n9101 = n9099 | n9100 ;
  assign n9198 = x81 &  n4934 ;
  assign n9195 = ( x83 & ~n4725 ) | ( x83 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n9196 = x82 &  n4720 ;
  assign n9197 = n9195 | n9196 ;
  assign n9199 = ( x81 & ~n9198 ) | ( x81 & n9197 ) | ( ~n9198 & n9197 ) ;
  assign n9200 = ( n1100 & ~n4728 ) | ( n1100 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n9201 = n9199 | n9200 ;
  assign n9202 = ( x44 & ~n9201 ) | ( x44 & 1'b0 ) | ( ~n9201 & 1'b0 ) ;
  assign n9203 = ~x44 & n9201 ;
  assign n9204 = n9202 | n9203 ;
  assign n9182 = x75 &  n6288 ;
  assign n9179 = ( x77 & ~n6032 ) | ( x77 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n9180 = x76 &  n6027 ;
  assign n9181 = n9179 | n9180 ;
  assign n9183 = ( x75 & ~n9182 ) | ( x75 & n9181 ) | ( ~n9182 & n9181 ) ;
  assign n9184 = ( n677 & ~n6035 ) | ( n677 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n9185 = n9183 | n9184 ;
  assign n9186 = ( x50 & ~n9185 ) | ( x50 & 1'b0 ) | ( ~n9185 & 1'b0 ) ;
  assign n9187 = ~x50 & n9185 ;
  assign n9188 = n9186 | n9187 ;
  assign n9125 = x69 &  n7731 ;
  assign n9122 = ( x71 & ~n7538 ) | ( x71 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n9123 = x70 &  n7533 ;
  assign n9124 = n9122 | n9123 ;
  assign n9126 = ( x69 & ~n9125 ) | ( x69 & n9124 ) | ( ~n9125 & n9124 ) ;
  assign n9127 = ( n298 & ~n7541 ) | ( n298 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n9128 = n9126 | n9127 ;
  assign n9129 = ( x56 & ~n9128 ) | ( x56 & 1'b0 ) | ( ~n9128 & 1'b0 ) ;
  assign n9130 = ~x56 & n9128 ;
  assign n9131 = n9129 | n9130 ;
  assign n9135 = x66 &  n8558 ;
  assign n9132 = ( x68 & ~n8314 ) | ( x68 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n9133 = x67 &  n8309 ;
  assign n9134 = n9132 | n9133 ;
  assign n9136 = ( x66 & ~n9135 ) | ( x66 & n9134 ) | ( ~n9135 & n9134 ) ;
  assign n9137 = ( n213 & ~n8317 ) | ( n213 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n9138 = n9136 | n9137 ;
  assign n9139 = ( x59 & ~n9138 ) | ( x59 & 1'b0 ) | ( ~n9138 & 1'b0 ) ;
  assign n9140 = ~x59 & n9138 ;
  assign n9141 = n9139 | n9140 ;
  assign n9142 = ( x62 & ~n8881 ) | ( x62 & 1'b0 ) | ( ~n8881 & 1'b0 ) ;
  assign n9143 = ( x60 & x61 ) | ( x60 & n8878 ) | ( x61 & n8878 ) ;
  assign n9144 = ( x60 & ~n8879 ) | ( x60 & x61 ) | ( ~n8879 & x61 ) ;
  assign n9145 = ~n9143 &  n9144 ;
  assign n9146 = x64 &  n9145 ;
  assign n9147 = ~x61 & x62 ;
  assign n9148 = ( x61 & ~x62 ) | ( x61 & 1'b0 ) | ( ~x62 & 1'b0 ) ;
  assign n9149 = n9147 | n9148 ;
  assign n9150 = ~n8880 |  n9149 ;
  assign n9151 = ( x65 & ~n9150 ) | ( x65 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n9152 = n9146 | n9151 ;
  assign n9153 = ~n8880 | ~n9149 ;
  assign n9154 = ( n142 & ~n9153 ) | ( n142 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n9155 = n9152 | n9154 ;
  assign n9157 = ( x62 & n9142 ) | ( x62 & n9155 ) | ( n9142 & n9155 ) ;
  assign n9156 = ( x62 & ~n9142 ) | ( x62 & n9155 ) | ( ~n9142 & n9155 ) ;
  assign n9158 = ( n9142 & ~n9157 ) | ( n9142 & n9156 ) | ( ~n9157 & n9156 ) ;
  assign n9160 = ( n8896 & n9141 ) | ( n8896 & n9158 ) | ( n9141 & n9158 ) ;
  assign n9159 = ( n8896 & ~n9141 ) | ( n8896 & n9158 ) | ( ~n9141 & n9158 ) ;
  assign n9161 = ( n9141 & ~n9160 ) | ( n9141 & n9159 ) | ( ~n9160 & n9159 ) ;
  assign n9163 = ( n8910 & n9131 ) | ( n8910 & n9161 ) | ( n9131 & n9161 ) ;
  assign n9162 = ( n8910 & ~n9131 ) | ( n8910 & n9161 ) | ( ~n9131 & n9161 ) ;
  assign n9164 = ( n9131 & ~n9163 ) | ( n9131 & n9162 ) | ( ~n9163 & n9162 ) ;
  assign n9175 = ( n8912 & ~n8911 ) | ( n8912 & n8922 ) | ( ~n8911 & n8922 ) ;
  assign n9168 = x72 &  n6982 ;
  assign n9165 = ( x74 & ~n6727 ) | ( x74 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n9166 = x73 &  n6722 ;
  assign n9167 = n9165 | n9166 ;
  assign n9169 = ( x72 & ~n9168 ) | ( x72 & n9167 ) | ( ~n9168 & n9167 ) ;
  assign n9170 = ( n482 & ~n6730 ) | ( n482 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n9171 = n9169 | n9170 ;
  assign n9172 = ( x53 & ~n9171 ) | ( x53 & 1'b0 ) | ( ~n9171 & 1'b0 ) ;
  assign n9173 = ~x53 & n9171 ;
  assign n9174 = n9172 | n9173 ;
  assign n9176 = ( n9164 & ~n9175 ) | ( n9164 & n9174 ) | ( ~n9175 & n9174 ) ;
  assign n9177 = ( n9164 & ~n9174 ) | ( n9164 & n9175 ) | ( ~n9174 & n9175 ) ;
  assign n9178 = ( n9176 & ~n9164 ) | ( n9176 & n9177 ) | ( ~n9164 & n9177 ) ;
  assign n9189 = ( n8927 & ~n9188 ) | ( n8927 & n9178 ) | ( ~n9188 & n9178 ) ;
  assign n9190 = ( n9178 & ~n8927 ) | ( n9178 & n9188 ) | ( ~n8927 & n9188 ) ;
  assign n9191 = ( n9189 & ~n9178 ) | ( n9189 & n9190 ) | ( ~n9178 & n9190 ) ;
  assign n9115 = x78 &  n5586 ;
  assign n9112 = ( x80 & ~n5389 ) | ( x80 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n9113 = x79 &  n5384 ;
  assign n9114 = n9112 | n9113 ;
  assign n9116 = ( x78 & ~n9115 ) | ( x78 & n9114 ) | ( ~n9115 & n9114 ) ;
  assign n9117 = ( n842 & ~n5392 ) | ( n842 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n9118 = n9116 | n9117 ;
  assign n9119 = ( x47 & ~n9118 ) | ( x47 & 1'b0 ) | ( ~n9118 & 1'b0 ) ;
  assign n9120 = ~x47 & n9118 ;
  assign n9121 = n9119 | n9120 ;
  assign n9192 = ( n8930 & ~n9191 ) | ( n8930 & n9121 ) | ( ~n9191 & n9121 ) ;
  assign n9193 = ( n9121 & ~n8930 ) | ( n9121 & n9191 ) | ( ~n8930 & n9191 ) ;
  assign n9194 = ( n9192 & ~n9121 ) | ( n9192 & n9193 ) | ( ~n9121 & n9193 ) ;
  assign n9205 = ( n8933 & ~n9204 ) | ( n8933 & n9194 ) | ( ~n9204 & n9194 ) ;
  assign n9206 = ( n9194 & ~n8933 ) | ( n9194 & n9204 ) | ( ~n8933 & n9204 ) ;
  assign n9207 = ( n9205 & ~n9194 ) | ( n9205 & n9206 ) | ( ~n9194 & n9206 ) ;
  assign n9105 = x84 &  n4344 ;
  assign n9102 = ( x86 & ~n4143 ) | ( x86 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n9103 = x85 &  n4138 ;
  assign n9104 = n9102 | n9103 ;
  assign n9106 = ( x84 & ~n9105 ) | ( x84 & n9104 ) | ( ~n9105 & n9104 ) ;
  assign n9107 = ( n1496 & ~n4146 ) | ( n1496 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n9108 = n9106 | n9107 ;
  assign n9109 = ( x41 & ~n9108 ) | ( x41 & 1'b0 ) | ( ~n9108 & 1'b0 ) ;
  assign n9110 = ~x41 & n9108 ;
  assign n9111 = n9109 | n9110 ;
  assign n9208 = ( n8936 & ~n9207 ) | ( n8936 & n9111 ) | ( ~n9207 & n9111 ) ;
  assign n9209 = ( n9111 & ~n8936 ) | ( n9111 & n9207 ) | ( ~n8936 & n9207 ) ;
  assign n9210 = ( n9208 & ~n9111 ) | ( n9208 & n9209 ) | ( ~n9111 & n9209 ) ;
  assign n9211 = ( n8939 & n9101 ) | ( n8939 & n9210 ) | ( n9101 & n9210 ) ;
  assign n9212 = ( n8939 & ~n9101 ) | ( n8939 & n9210 ) | ( ~n9101 & n9210 ) ;
  assign n9213 = ( n9101 & ~n9211 ) | ( n9101 & n9212 ) | ( ~n9211 & n9212 ) ;
  assign n9214 = ( n8942 & n9091 ) | ( n8942 & n9213 ) | ( n9091 & n9213 ) ;
  assign n9215 = ( n8942 & ~n9091 ) | ( n8942 & n9213 ) | ( ~n9091 & n9213 ) ;
  assign n9216 = ( n9091 & ~n9214 ) | ( n9091 & n9215 ) | ( ~n9214 & n9215 ) ;
  assign n9221 = x93 &  n2718 ;
  assign n9218 = ( x95 & ~n2642 ) | ( x95 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n9219 = x94 &  n2637 ;
  assign n9220 = n9218 | n9219 ;
  assign n9222 = ( x93 & ~n9221 ) | ( x93 & n9220 ) | ( ~n9221 & n9220 ) ;
  assign n9223 = ( n2547 & ~n2645 ) | ( n2547 & 1'b0 ) | ( ~n2645 & 1'b0 ) ;
  assign n9224 = n9222 | n9223 ;
  assign n9225 = ( x32 & ~n9224 ) | ( x32 & 1'b0 ) | ( ~n9224 & 1'b0 ) ;
  assign n9226 = ~x32 & n9224 ;
  assign n9227 = n9225 | n9226 ;
  assign n9217 = ( n8945 & ~n8944 ) | ( n8945 & n8955 ) | ( ~n8944 & n8955 ) ;
  assign n9228 = ( n9216 & ~n9227 ) | ( n9216 & n9217 ) | ( ~n9227 & n9217 ) ;
  assign n9229 = ( n9216 & ~n9217 ) | ( n9216 & n9227 ) | ( ~n9217 & n9227 ) ;
  assign n9230 = ( n9228 & ~n9216 ) | ( n9228 & n9229 ) | ( ~n9216 & n9229 ) ;
  assign n9234 = x96 &  n2312 ;
  assign n9231 = ( x98 & ~n2195 ) | ( x98 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n9232 = x97 &  n2190 ;
  assign n9233 = n9231 | n9232 ;
  assign n9235 = ( x96 & ~n9234 ) | ( x96 & n9233 ) | ( ~n9234 & n9233 ) ;
  assign n9236 = ~n2198 & n3170 ;
  assign n9237 = n9235 | n9236 ;
  assign n9238 = ( x29 & ~n9237 ) | ( x29 & 1'b0 ) | ( ~n9237 & 1'b0 ) ;
  assign n9239 = ~x29 & n9237 ;
  assign n9240 = n9238 | n9239 ;
  assign n9241 = ( n9230 & ~n8971 ) | ( n9230 & n9240 ) | ( ~n8971 & n9240 ) ;
  assign n9242 = ( n8971 & ~n9240 ) | ( n8971 & n9230 ) | ( ~n9240 & n9230 ) ;
  assign n9243 = ( n9241 & ~n9230 ) | ( n9241 & n9242 ) | ( ~n9230 & n9242 ) ;
  assign n9244 = ( n8972 & ~n8973 ) | ( n8972 & n8983 ) | ( ~n8973 & n8983 ) ;
  assign n9245 = ( n9081 & ~n9243 ) | ( n9081 & n9244 ) | ( ~n9243 & n9244 ) ;
  assign n9246 = ( n9081 & ~n9244 ) | ( n9081 & n9243 ) | ( ~n9244 & n9243 ) ;
  assign n9247 = ( n9245 & ~n9081 ) | ( n9245 & n9246 ) | ( ~n9081 & n9246 ) ;
  assign n9065 = x102 &  n1551 ;
  assign n9062 = ( x104 & ~n1451 ) | ( x104 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n9063 = x103 &  n1446 ;
  assign n9064 = n9062 | n9063 ;
  assign n9066 = ( x102 & ~n9065 ) | ( x102 & n9064 ) | ( ~n9065 & n9064 ) ;
  assign n9067 = n1454 | n4249 ;
  assign n9068 = ~n9066 & n9067 ;
  assign n9069 = x23 &  n9068 ;
  assign n9070 = x23 | n9068 ;
  assign n9071 = ~n9069 & n9070 ;
  assign n9248 = ( n8987 & ~n9247 ) | ( n8987 & n9071 ) | ( ~n9247 & n9071 ) ;
  assign n9249 = ( n9071 & ~n8987 ) | ( n9071 & n9247 ) | ( ~n8987 & n9247 ) ;
  assign n9250 = ( n9248 & ~n9071 ) | ( n9248 & n9249 ) | ( ~n9071 & n9249 ) ;
  assign n9255 = x105 &  n1227 ;
  assign n9252 = ( x107 & ~n1154 ) | ( x107 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n9253 = x106 &  n1149 ;
  assign n9254 = n9252 | n9253 ;
  assign n9256 = ( x105 & ~n9255 ) | ( x105 & n9254 ) | ( ~n9255 & n9254 ) ;
  assign n9257 = ~n1157 & n4848 ;
  assign n9258 = n9256 | n9257 ;
  assign n9259 = ( x20 & ~n9258 ) | ( x20 & 1'b0 ) | ( ~n9258 & 1'b0 ) ;
  assign n9260 = ~x20 & n9258 ;
  assign n9261 = n9259 | n9260 ;
  assign n9251 = ( n8989 & ~n8990 ) | ( n8989 & n9000 ) | ( ~n8990 & n9000 ) ;
  assign n9262 = ( n9250 & ~n9261 ) | ( n9250 & n9251 ) | ( ~n9261 & n9251 ) ;
  assign n9263 = ( n9250 & ~n9251 ) | ( n9250 & n9261 ) | ( ~n9251 & n9261 ) ;
  assign n9264 = ( n9262 & ~n9250 ) | ( n9262 & n9263 ) | ( ~n9250 & n9263 ) ;
  assign n9268 = x108 &  n942 ;
  assign n9265 = ( x110 & ~n896 ) | ( x110 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n9266 = x109 &  n891 ;
  assign n9267 = n9265 | n9266 ;
  assign n9269 = ( x108 & ~n9268 ) | ( x108 & n9267 ) | ( ~n9268 & n9267 ) ;
  assign n9270 = n899 | n5283 ;
  assign n9271 = ~n9269 & n9270 ;
  assign n9272 = x17 &  n9271 ;
  assign n9273 = x17 | n9271 ;
  assign n9274 = ~n9272 & n9273 ;
  assign n9276 = ( n9004 & n9264 ) | ( n9004 & n9274 ) | ( n9264 & n9274 ) ;
  assign n9275 = ( n9004 & ~n9264 ) | ( n9004 & n9274 ) | ( ~n9264 & n9274 ) ;
  assign n9277 = ( n9264 & ~n9276 ) | ( n9264 & n9275 ) | ( ~n9276 & n9275 ) ;
  assign n9278 = ( x14 & ~n9061 ) | ( x14 & n9277 ) | ( ~n9061 & n9277 ) ;
  assign n9279 = ( n9061 & ~x14 ) | ( n9061 & n9277 ) | ( ~x14 & n9277 ) ;
  assign n9280 = ( n9278 & ~n9277 ) | ( n9278 & n9279 ) | ( ~n9277 & n9279 ) ;
  assign n9284 = x114 &  n503 ;
  assign n9281 = ( x116 & ~n450 ) | ( x116 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n9282 = x115 &  n445 ;
  assign n9283 = n9281 | n9282 ;
  assign n9285 = ( x114 & ~n9284 ) | ( x114 & n9283 ) | ( ~n9284 & n9283 ) ;
  assign n9286 = n453 | n6885 ;
  assign n9287 = ~n9285 & n9286 ;
  assign n9288 = x11 | n9287 ;
  assign n9289 = ~x11 & n9287 ;
  assign n9290 = ( n9288 & ~n9287 ) | ( n9288 & n9289 ) | ( ~n9287 & n9289 ) ;
  assign n9291 = ( n9007 & ~n9280 ) | ( n9007 & n9290 ) | ( ~n9280 & n9290 ) ;
  assign n9292 = ( n9280 & ~n9007 ) | ( n9280 & n9290 ) | ( ~n9007 & n9290 ) ;
  assign n9293 = ( n9291 & ~n9290 ) | ( n9291 & n9292 ) | ( ~n9290 & n9292 ) ;
  assign n9048 = x117 &  n353 ;
  assign n9045 = ( x119 & ~n313 ) | ( x119 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n9046 = x118 &  n308 ;
  assign n9047 = n9045 | n9046 ;
  assign n9049 = ( x117 & ~n9048 ) | ( x117 & n9047 ) | ( ~n9048 & n9047 ) ;
  assign n9050 = ~n316 & n7648 ;
  assign n9051 = n9049 | n9050 ;
  assign n9052 = ( x8 & ~n9051 ) | ( x8 & 1'b0 ) | ( ~n9051 & 1'b0 ) ;
  assign n9053 = ~x8 & n9051 ;
  assign n9054 = n9052 | n9053 ;
  assign n9294 = ( n9044 & ~n9293 ) | ( n9044 & n9054 ) | ( ~n9293 & n9054 ) ;
  assign n9295 = ( n9044 & ~n9054 ) | ( n9044 & n9293 ) | ( ~n9054 & n9293 ) ;
  assign n9296 = ( n9294 & ~n9044 ) | ( n9294 & n9295 ) | ( ~n9044 & n9295 ) ;
  assign n9307 = ( n8764 & ~n9009 ) | ( n8764 & n8786 ) | ( ~n9009 & n8786 ) ;
  assign n9308 = ( n9044 & ~n8786 ) | ( n9044 & n9307 ) | ( ~n8786 & n9307 ) ;
  assign n9309 = ( n8766 & n8776 ) | ( n8766 & n9308 ) | ( n8776 & n9308 ) ;
  assign n9300 = x120 &  n225 ;
  assign n9297 = ( x122 & ~n197 ) | ( x122 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n9298 = x121 &  n192 ;
  assign n9299 = n9297 | n9298 ;
  assign n9301 = ( x120 & ~n9300 ) | ( x120 & n9299 ) | ( ~n9300 & n9299 ) ;
  assign n9302 = ( n8448 & ~n200 ) | ( n8448 & n8451 ) | ( ~n200 & n8451 ) ;
  assign n9303 = ( n9301 & ~n8452 ) | ( n9301 & n9302 ) | ( ~n8452 & n9302 ) ;
  assign n9304 = ( x5 & ~n9303 ) | ( x5 & 1'b0 ) | ( ~n9303 & 1'b0 ) ;
  assign n9305 = ~x5 & n9303 ;
  assign n9306 = n9304 | n9305 ;
  assign n9310 = ( n9296 & ~n9309 ) | ( n9296 & n9306 ) | ( ~n9309 & n9306 ) ;
  assign n9311 = ( n9296 & ~n9306 ) | ( n9296 & n9309 ) | ( ~n9306 & n9309 ) ;
  assign n9312 = ( n9310 & ~n9296 ) | ( n9310 & n9311 ) | ( ~n9296 & n9311 ) ;
  assign n9316 = ~n136 & x125 ;
  assign n9313 = ( x123 & ~n150 ) | ( x123 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n9314 = ( x124 & ~n131 ) | ( x124 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n9315 = n9313 | n9314 ;
  assign n9317 = ( x125 & ~n9316 ) | ( x125 & n9315 ) | ( ~n9316 & n9315 ) ;
  assign n9318 = ( x123 & x124 ) | ( x123 & n8749 ) | ( x124 & n8749 ) ;
  assign n9319 = x124 | x125 ;
  assign n9320 = x124 &  x125 ;
  assign n9321 = ( n9319 & ~n9320 ) | ( n9319 & 1'b0 ) | ( ~n9320 & 1'b0 ) ;
  assign n9322 = n9318 &  n9321 ;
  assign n9323 = n9318 | n9321 ;
  assign n9324 = ~n9322 & n9323 ;
  assign n9325 = ~n139 & n9324 ;
  assign n9326 = n9317 | n9325 ;
  assign n9327 = ( x2 & ~n9312 ) | ( x2 & n9326 ) | ( ~n9312 & n9326 ) ;
  assign n9328 = ( x2 & ~n9326 ) | ( x2 & n9312 ) | ( ~n9326 & n9312 ) ;
  assign n9329 = ( n9327 & ~x2 ) | ( n9327 & n9328 ) | ( ~x2 & n9328 ) ;
  assign n9330 = ( n9033 & n9043 ) | ( n9033 & n9329 ) | ( n9043 & n9329 ) ;
  assign n9331 = ( n9033 & ~n9043 ) | ( n9033 & n9329 ) | ( ~n9043 & n9329 ) ;
  assign n9332 = ( n9043 & ~n9330 ) | ( n9043 & n9331 ) | ( ~n9330 & n9331 ) ;
  assign n9333 = ~n9296 & n9309 ;
  assign n9334 = ( n9296 & ~n9309 ) | ( n9296 & 1'b0 ) | ( ~n9309 & 1'b0 ) ;
  assign n9335 = n9333 | n9334 ;
  assign n9336 = ( x2 & ~n9326 ) | ( x2 & 1'b0 ) | ( ~n9326 & 1'b0 ) ;
  assign n9337 = ~x2 & n9326 ;
  assign n9338 = n9336 | n9337 ;
  assign n9339 = ( n9306 & ~n9335 ) | ( n9306 & n9338 ) | ( ~n9335 & n9338 ) ;
  assign n9340 = ( n9033 & ~n9329 ) | ( n9033 & n9043 ) | ( ~n9329 & n9043 ) ;
  assign n9624 = x121 &  n225 ;
  assign n9621 = ( x123 & ~n197 ) | ( x123 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n9622 = x122 &  n192 ;
  assign n9623 = n9621 | n9622 ;
  assign n9625 = ( x121 & ~n9624 ) | ( x121 & n9623 ) | ( ~n9624 & n9623 ) ;
  assign n9626 = ( n8466 & ~n200 ) | ( n8466 & n8469 ) | ( ~n200 & n8469 ) ;
  assign n9627 = ( n9625 & ~n8470 ) | ( n9625 & n9626 ) | ( ~n8470 & n9626 ) ;
  assign n9628 = ( x5 & ~n9627 ) | ( x5 & 1'b0 ) | ( ~n9627 & 1'b0 ) ;
  assign n9629 = ~x5 & n9627 ;
  assign n9630 = n9628 | n9629 ;
  assign n9352 = ( x11 & ~n9287 ) | ( x11 & 1'b0 ) | ( ~n9287 & 1'b0 ) ;
  assign n9353 = ( n9288 & ~x11 ) | ( n9288 & n9352 ) | ( ~x11 & n9352 ) ;
  assign n9354 = n9007 &  n9280 ;
  assign n9355 = n9007 | n9280 ;
  assign n9356 = ~n9354 & n9355 ;
  assign n9357 = ( n9353 & ~n9044 ) | ( n9353 & n9356 ) | ( ~n9044 & n9356 ) ;
  assign n9361 = x118 &  n353 ;
  assign n9358 = ( x120 & ~n313 ) | ( x120 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n9359 = x119 &  n308 ;
  assign n9360 = n9358 | n9359 ;
  assign n9362 = ( x118 & ~n9361 ) | ( x118 & n9360 ) | ( ~n9361 & n9360 ) ;
  assign n9363 = n7647 | n7907 ;
  assign n9364 = ~n7908 & n9363 ;
  assign n9365 = ~n316 & n9364 ;
  assign n9366 = n9362 | n9365 ;
  assign n9367 = ( x8 & ~n9366 ) | ( x8 & 1'b0 ) | ( ~n9366 & 1'b0 ) ;
  assign n9368 = ~x8 & n9366 ;
  assign n9369 = n9367 | n9368 ;
  assign n9370 = ( n644 & ~n6169 ) | ( n644 & n9059 ) | ( ~n6169 & n9059 ) ;
  assign n9371 = n6169 | n9370 ;
  assign n9373 = ( x14 & n9059 ) | ( x14 & n9371 ) | ( n9059 & n9371 ) ;
  assign n9372 = ( x14 & ~n9371 ) | ( x14 & n9059 ) | ( ~n9371 & n9059 ) ;
  assign n9374 = ( n9371 & ~n9373 ) | ( n9371 & n9372 ) | ( ~n9373 & n9372 ) ;
  assign n9375 = ( n9007 & n9277 ) | ( n9007 & n9374 ) | ( n9277 & n9374 ) ;
  assign n9379 = x115 &  n503 ;
  assign n9376 = ( x117 & ~n450 ) | ( x117 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n9377 = x116 &  n445 ;
  assign n9378 = n9376 | n9377 ;
  assign n9380 = ( x115 & ~n9379 ) | ( x115 & n9378 ) | ( ~n9379 & n9378 ) ;
  assign n9381 = n453 | n7136 ;
  assign n9382 = ~n9380 & n9381 ;
  assign n9383 = x11 &  n9382 ;
  assign n9384 = x11 | n9382 ;
  assign n9385 = ~n9383 & n9384 ;
  assign n9389 = x112 &  n713 ;
  assign n9386 = ( x114 & ~n641 ) | ( x114 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n9387 = x113 &  n636 ;
  assign n9388 = n9386 | n9387 ;
  assign n9390 = ( x112 & ~n9389 ) | ( x112 & n9388 ) | ( ~n9389 & n9388 ) ;
  assign n9391 = n644 | n6185 ;
  assign n9392 = ~n9390 & n9391 ;
  assign n9396 = x100 &  n1894 ;
  assign n9393 = ( x102 & ~n1816 ) | ( x102 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n9394 = x101 &  n1811 ;
  assign n9395 = n9393 | n9394 ;
  assign n9397 = ( x100 & ~n9396 ) | ( x100 & n9395 ) | ( ~n9396 & n9395 ) ;
  assign n9398 = n1819 | n3872 ;
  assign n9399 = ~n9397 & n9398 ;
  assign n9400 = x26 &  n9399 ;
  assign n9401 = x26 | n9399 ;
  assign n9402 = ~n9400 & n9401 ;
  assign n9406 = x97 &  n2312 ;
  assign n9403 = ( x99 & ~n2195 ) | ( x99 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n9404 = x98 &  n2190 ;
  assign n9405 = n9403 | n9404 ;
  assign n9407 = ( x97 & ~n9406 ) | ( x97 & n9405 ) | ( ~n9406 & n9405 ) ;
  assign n9408 = ~n2198 & n3338 ;
  assign n9409 = n9407 | n9408 ;
  assign n9410 = ( x29 & ~n9409 ) | ( x29 & 1'b0 ) | ( ~n9409 & 1'b0 ) ;
  assign n9411 = ~x29 & n9409 ;
  assign n9412 = n9410 | n9411 ;
  assign n9416 = x91 &  n3214 ;
  assign n9413 = ( x93 & ~n3087 ) | ( x93 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n9414 = x92 &  n3082 ;
  assign n9415 = n9413 | n9414 ;
  assign n9417 = ( x91 & ~n9416 ) | ( x91 & n9415 ) | ( ~n9416 & n9415 ) ;
  assign n9418 = n2264 | n3090 ;
  assign n9419 = ~n9417 & n9418 ;
  assign n9420 = x35 &  n9419 ;
  assign n9421 = x35 | n9419 ;
  assign n9422 = ~n9420 & n9421 ;
  assign n9426 = x88 &  n3756 ;
  assign n9423 = ( x90 & ~n3602 ) | ( x90 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n9424 = x89 &  n3597 ;
  assign n9425 = n9423 | n9424 ;
  assign n9427 = ( x88 & ~n9426 ) | ( x88 & n9425 ) | ( ~n9426 & n9425 ) ;
  assign n9428 = ( n1976 & ~n3605 ) | ( n1976 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n9429 = n9427 | n9428 ;
  assign n9430 = ( x38 & ~n9429 ) | ( x38 & 1'b0 ) | ( ~n9429 & 1'b0 ) ;
  assign n9431 = ~x38 & n9429 ;
  assign n9432 = n9430 | n9431 ;
  assign n9436 = x79 &  n5586 ;
  assign n9433 = ( x81 & ~n5389 ) | ( x81 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n9434 = x80 &  n5384 ;
  assign n9435 = n9433 | n9434 ;
  assign n9437 = ( x79 & ~n9436 ) | ( x79 & n9435 ) | ( ~n9436 & n9435 ) ;
  assign n9438 = ( n994 & ~n5392 ) | ( n994 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n9439 = n9437 | n9438 ;
  assign n9440 = ( x47 & ~n9439 ) | ( x47 & 1'b0 ) | ( ~n9439 & 1'b0 ) ;
  assign n9441 = ~x47 & n9439 ;
  assign n9442 = n9440 | n9441 ;
  assign n9443 = ( n8930 & n9121 ) | ( n8930 & n9191 ) | ( n9121 & n9191 ) ;
  assign n9503 = x76 &  n6288 ;
  assign n9500 = ( x78 & ~n6032 ) | ( x78 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n9501 = x77 &  n6027 ;
  assign n9502 = n9500 | n9501 ;
  assign n9504 = ( x76 & ~n9503 ) | ( x76 & n9502 ) | ( ~n9503 & n9502 ) ;
  assign n9505 = ( n693 & ~n6035 ) | ( n693 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n9506 = n9504 | n9505 ;
  assign n9507 = ( x50 & ~n9506 ) | ( x50 & 1'b0 ) | ( ~n9506 & 1'b0 ) ;
  assign n9508 = ~x50 & n9506 ;
  assign n9509 = n9507 | n9508 ;
  assign n9447 = x73 &  n6982 ;
  assign n9444 = ( x75 & ~n6727 ) | ( x75 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n9445 = x74 &  n6722 ;
  assign n9446 = n9444 | n9445 ;
  assign n9448 = ( x73 & ~n9447 ) | ( x73 & n9446 ) | ( ~n9447 & n9446 ) ;
  assign n9449 = ( n540 & ~n6730 ) | ( n540 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n9450 = n9448 | n9449 ;
  assign n9451 = ( x53 & ~n9450 ) | ( x53 & 1'b0 ) | ( ~n9450 & 1'b0 ) ;
  assign n9452 = ~x53 & n9450 ;
  assign n9453 = n9451 | n9452 ;
  assign n9454 = ( n9164 & n9174 ) | ( n9164 & n9175 ) | ( n9174 & n9175 ) ;
  assign n9473 = x67 &  n8558 ;
  assign n9470 = ( x69 & ~n8314 ) | ( x69 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n9471 = x68 &  n8309 ;
  assign n9472 = n9470 | n9471 ;
  assign n9474 = ( x67 & ~n9473 ) | ( x67 & n9472 ) | ( ~n9473 & n9472 ) ;
  assign n9475 = ( n246 & ~n8317 ) | ( n246 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n9476 = n9474 | n9475 ;
  assign n9477 = ( x59 & ~n9476 ) | ( x59 & 1'b0 ) | ( ~n9476 & 1'b0 ) ;
  assign n9478 = ~x59 & n9476 ;
  assign n9479 = n9477 | n9478 ;
  assign n9456 = ( x60 & ~x61 ) | ( x60 & n9149 ) | ( ~x61 & n9149 ) ;
  assign n9455 = ( x60 & ~x61 ) | ( x60 & n8880 ) | ( ~x61 & n8880 ) ;
  assign n9457 = ~n9456 |  n9455 ;
  assign n9461 = x64 &  n9457 ;
  assign n9458 = ( x66 & ~n9150 ) | ( x66 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n9459 = x65 &  n9145 ;
  assign n9460 = n9458 | n9459 ;
  assign n9462 = ( x64 & ~n9461 ) | ( x64 & n9460 ) | ( ~n9461 & n9460 ) ;
  assign n9463 = ( n157 & ~n9153 ) | ( n157 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n9464 = n9462 | n9463 ;
  assign n9465 = ( x62 & ~n8881 ) | ( x62 & n9155 ) | ( ~n8881 & n9155 ) ;
  assign n9466 = ~n9155 & n9465 ;
  assign n9467 = ( n9464 & ~x62 ) | ( n9464 & n9466 ) | ( ~x62 & n9466 ) ;
  assign n9468 = ( x62 & ~n9464 ) | ( x62 & n9466 ) | ( ~n9464 & n9466 ) ;
  assign n9469 = ( n9467 & ~n9466 ) | ( n9467 & n9468 ) | ( ~n9466 & n9468 ) ;
  assign n9480 = ( n9160 & ~n9479 ) | ( n9160 & n9469 ) | ( ~n9479 & n9469 ) ;
  assign n9481 = ( n9469 & ~n9160 ) | ( n9469 & n9479 ) | ( ~n9160 & n9479 ) ;
  assign n9482 = ( n9480 & ~n9469 ) | ( n9480 & n9481 ) | ( ~n9469 & n9481 ) ;
  assign n9486 = x70 &  n7731 ;
  assign n9483 = ( x72 & ~n7538 ) | ( x72 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n9484 = x71 &  n7533 ;
  assign n9485 = n9483 | n9484 ;
  assign n9487 = ( x70 & ~n9486 ) | ( x70 & n9485 ) | ( ~n9486 & n9485 ) ;
  assign n9488 = ( n345 & ~n7541 ) | ( n345 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n9489 = n9487 | n9488 ;
  assign n9490 = ( x56 & ~n9489 ) | ( x56 & 1'b0 ) | ( ~n9489 & 1'b0 ) ;
  assign n9491 = ~x56 & n9489 ;
  assign n9492 = n9490 | n9491 ;
  assign n9493 = ( n9482 & ~n9163 ) | ( n9482 & n9492 ) | ( ~n9163 & n9492 ) ;
  assign n9494 = ( n9163 & ~n9492 ) | ( n9163 & n9482 ) | ( ~n9492 & n9482 ) ;
  assign n9495 = ( n9493 & ~n9482 ) | ( n9493 & n9494 ) | ( ~n9482 & n9494 ) ;
  assign n9497 = ( n9453 & n9454 ) | ( n9453 & n9495 ) | ( n9454 & n9495 ) ;
  assign n9496 = ( n9454 & ~n9453 ) | ( n9454 & n9495 ) | ( ~n9453 & n9495 ) ;
  assign n9498 = ( n9453 & ~n9497 ) | ( n9453 & n9496 ) | ( ~n9497 & n9496 ) ;
  assign n9499 = ( n8927 & n9178 ) | ( n8927 & n9188 ) | ( n9178 & n9188 ) ;
  assign n9511 = ( n9498 & n9499 ) | ( n9498 & n9509 ) | ( n9499 & n9509 ) ;
  assign n9510 = ( n9498 & ~n9509 ) | ( n9498 & n9499 ) | ( ~n9509 & n9499 ) ;
  assign n9512 = ( n9509 & ~n9511 ) | ( n9509 & n9510 ) | ( ~n9511 & n9510 ) ;
  assign n9514 = ( n9442 & n9443 ) | ( n9442 & n9512 ) | ( n9443 & n9512 ) ;
  assign n9513 = ( n9443 & ~n9442 ) | ( n9443 & n9512 ) | ( ~n9442 & n9512 ) ;
  assign n9515 = ( n9442 & ~n9514 ) | ( n9442 & n9513 ) | ( ~n9514 & n9513 ) ;
  assign n9516 = ( n8933 & n9194 ) | ( n8933 & n9204 ) | ( n9194 & n9204 ) ;
  assign n9520 = x82 &  n4934 ;
  assign n9517 = ( x84 & ~n4725 ) | ( x84 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n9518 = x83 &  n4720 ;
  assign n9519 = n9517 | n9518 ;
  assign n9521 = ( x82 & ~n9520 ) | ( x82 & n9519 ) | ( ~n9520 & n9519 ) ;
  assign n9522 = ( n1199 & ~n4728 ) | ( n1199 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n9523 = n9521 | n9522 ;
  assign n9524 = ( x44 & ~n9523 ) | ( x44 & 1'b0 ) | ( ~n9523 & 1'b0 ) ;
  assign n9525 = ~x44 & n9523 ;
  assign n9526 = n9524 | n9525 ;
  assign n9527 = ( n9515 & ~n9516 ) | ( n9515 & n9526 ) | ( ~n9516 & n9526 ) ;
  assign n9528 = ( n9515 & ~n9526 ) | ( n9515 & n9516 ) | ( ~n9526 & n9516 ) ;
  assign n9529 = ( n9527 & ~n9515 ) | ( n9527 & n9528 ) | ( ~n9515 & n9528 ) ;
  assign n9530 = ( n8936 & n9111 ) | ( n8936 & n9207 ) | ( n9111 & n9207 ) ;
  assign n9534 = x85 &  n4344 ;
  assign n9531 = ( x87 & ~n4143 ) | ( x87 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n9532 = x86 &  n4138 ;
  assign n9533 = n9531 | n9532 ;
  assign n9535 = ( x85 & ~n9534 ) | ( x85 & n9533 ) | ( ~n9534 & n9533 ) ;
  assign n9536 = ( n1512 & ~n4146 ) | ( n1512 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n9537 = n9535 | n9536 ;
  assign n9538 = ( x41 & ~n9537 ) | ( x41 & 1'b0 ) | ( ~n9537 & 1'b0 ) ;
  assign n9539 = ~x41 & n9537 ;
  assign n9540 = n9538 | n9539 ;
  assign n9541 = ( n9529 & ~n9530 ) | ( n9529 & n9540 ) | ( ~n9530 & n9540 ) ;
  assign n9542 = ( n9529 & ~n9540 ) | ( n9529 & n9530 ) | ( ~n9540 & n9530 ) ;
  assign n9543 = ( n9541 & ~n9529 ) | ( n9541 & n9542 ) | ( ~n9529 & n9542 ) ;
  assign n9544 = ( n9211 & n9432 ) | ( n9211 & n9543 ) | ( n9432 & n9543 ) ;
  assign n9545 = ( n9211 & ~n9432 ) | ( n9211 & n9543 ) | ( ~n9432 & n9543 ) ;
  assign n9546 = ( n9432 & ~n9544 ) | ( n9432 & n9545 ) | ( ~n9544 & n9545 ) ;
  assign n9548 = ( n9214 & n9422 ) | ( n9214 & n9546 ) | ( n9422 & n9546 ) ;
  assign n9547 = ( n9214 & ~n9422 ) | ( n9214 & n9546 ) | ( ~n9422 & n9546 ) ;
  assign n9549 = ( n9422 & ~n9548 ) | ( n9422 & n9547 ) | ( ~n9548 & n9547 ) ;
  assign n9550 = ( n9216 & n9217 ) | ( n9216 & n9227 ) | ( n9217 & n9227 ) ;
  assign n9554 = x94 &  n2718 ;
  assign n9551 = ( x96 & ~n2642 ) | ( x96 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n9552 = x95 &  n2637 ;
  assign n9553 = n9551 | n9552 ;
  assign n9555 = ( x94 & ~n9554 ) | ( x94 & n9553 ) | ( ~n9554 & n9553 ) ;
  assign n9556 = ~n2645 & n2836 ;
  assign n9557 = n9555 | n9556 ;
  assign n9558 = ( x32 & ~n9557 ) | ( x32 & 1'b0 ) | ( ~n9557 & 1'b0 ) ;
  assign n9559 = ~x32 & n9557 ;
  assign n9560 = n9558 | n9559 ;
  assign n9561 = ( n9549 & ~n9550 ) | ( n9549 & n9560 ) | ( ~n9550 & n9560 ) ;
  assign n9562 = ( n9549 & ~n9560 ) | ( n9549 & n9550 ) | ( ~n9560 & n9550 ) ;
  assign n9563 = ( n9561 & ~n9549 ) | ( n9561 & n9562 ) | ( ~n9549 & n9562 ) ;
  assign n9564 = ( n8971 & n9230 ) | ( n8971 & n9240 ) | ( n9230 & n9240 ) ;
  assign n9565 = ( n9412 & n9563 ) | ( n9412 & n9564 ) | ( n9563 & n9564 ) ;
  assign n9566 = ( n9563 & ~n9412 ) | ( n9563 & n9564 ) | ( ~n9412 & n9564 ) ;
  assign n9567 = ( n9412 & ~n9565 ) | ( n9412 & n9566 ) | ( ~n9565 & n9566 ) ;
  assign n9568 = ( n9245 & n9402 ) | ( n9245 & n9567 ) | ( n9402 & n9567 ) ;
  assign n9569 = ( n9245 & ~n9402 ) | ( n9245 & n9567 ) | ( ~n9402 & n9567 ) ;
  assign n9570 = ( n9402 & ~n9568 ) | ( n9402 & n9569 ) | ( ~n9568 & n9569 ) ;
  assign n9574 = x103 &  n1551 ;
  assign n9571 = ( x105 & ~n1451 ) | ( x105 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n9572 = x104 &  n1446 ;
  assign n9573 = n9571 | n9572 ;
  assign n9575 = ( x103 & ~n9574 ) | ( x103 & n9573 ) | ( ~n9574 & n9573 ) ;
  assign n9576 = ~n1454 & n4442 ;
  assign n9577 = n9575 | n9576 ;
  assign n9578 = ( x23 & ~n9577 ) | ( x23 & 1'b0 ) | ( ~n9577 & 1'b0 ) ;
  assign n9579 = ~x23 & n9577 ;
  assign n9580 = n9578 | n9579 ;
  assign n9581 = ( n9248 & n9570 ) | ( n9248 & n9580 ) | ( n9570 & n9580 ) ;
  assign n9582 = ( n9248 & ~n9570 ) | ( n9248 & n9580 ) | ( ~n9570 & n9580 ) ;
  assign n9583 = ( n9570 & ~n9581 ) | ( n9570 & n9582 ) | ( ~n9581 & n9582 ) ;
  assign n9584 = ( n9250 & n9251 ) | ( n9250 & n9261 ) | ( n9251 & n9261 ) ;
  assign n9588 = x106 &  n1227 ;
  assign n9585 = ( x108 & ~n1154 ) | ( x108 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n9586 = x107 &  n1149 ;
  assign n9587 = n9585 | n9586 ;
  assign n9589 = ( x106 & ~n9588 ) | ( x106 & n9587 ) | ( ~n9588 & n9587 ) ;
  assign n9590 = n1157 | n5055 ;
  assign n9591 = ~n9589 & n9590 ;
  assign n9592 = x20 &  n9591 ;
  assign n9593 = x20 | n9591 ;
  assign n9594 = ~n9592 & n9593 ;
  assign n9596 = ( n9583 & n9584 ) | ( n9583 & n9594 ) | ( n9584 & n9594 ) ;
  assign n9595 = ( n9584 & ~n9583 ) | ( n9584 & n9594 ) | ( ~n9583 & n9594 ) ;
  assign n9597 = ( n9583 & ~n9596 ) | ( n9583 & n9595 ) | ( ~n9596 & n9595 ) ;
  assign n9598 = ( n9004 & ~n9274 ) | ( n9004 & n9264 ) | ( ~n9274 & n9264 ) ;
  assign n9602 = x109 &  n942 ;
  assign n9599 = ( x111 & ~n896 ) | ( x111 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n9600 = x110 &  n891 ;
  assign n9601 = n9599 | n9600 ;
  assign n9603 = ( x109 & ~n9602 ) | ( x109 & n9601 ) | ( ~n9602 & n9601 ) ;
  assign n9604 = n899 | n5711 ;
  assign n9605 = ~n9603 & n9604 ;
  assign n9606 = x17 &  n9605 ;
  assign n9607 = x17 | n9605 ;
  assign n9608 = ~n9606 & n9607 ;
  assign n9609 = ( n9597 & n9598 ) | ( n9597 & n9608 ) | ( n9598 & n9608 ) ;
  assign n9610 = ( n9598 & ~n9597 ) | ( n9598 & n9608 ) | ( ~n9597 & n9608 ) ;
  assign n9611 = ( n9597 & ~n9609 ) | ( n9597 & n9610 ) | ( ~n9609 & n9610 ) ;
  assign n9612 = ( n9392 & ~x14 ) | ( n9392 & n9611 ) | ( ~x14 & n9611 ) ;
  assign n9613 = ( x14 & ~n9392 ) | ( x14 & n9611 ) | ( ~n9392 & n9611 ) ;
  assign n9614 = ( n9612 & ~n9611 ) | ( n9612 & n9613 ) | ( ~n9611 & n9613 ) ;
  assign n9615 = ( n9375 & n9385 ) | ( n9375 & n9614 ) | ( n9385 & n9614 ) ;
  assign n9616 = ( n9385 & ~n9375 ) | ( n9385 & n9614 ) | ( ~n9375 & n9614 ) ;
  assign n9617 = ( n9375 & ~n9615 ) | ( n9375 & n9616 ) | ( ~n9615 & n9616 ) ;
  assign n9619 = ( n9357 & n9369 ) | ( n9357 & n9617 ) | ( n9369 & n9617 ) ;
  assign n9618 = ( n9369 & ~n9357 ) | ( n9369 & n9617 ) | ( ~n9357 & n9617 ) ;
  assign n9620 = ( n9357 & ~n9619 ) | ( n9357 & n9618 ) | ( ~n9619 & n9618 ) ;
  assign n9631 = ~n9044 & n9293 ;
  assign n9632 = ( n9044 & ~n9293 ) | ( n9044 & 1'b0 ) | ( ~n9293 & 1'b0 ) ;
  assign n9633 = n9631 | n9632 ;
  assign n9634 = ( n9054 & ~n9309 ) | ( n9054 & n9633 ) | ( ~n9309 & n9633 ) ;
  assign n9635 = ( n9630 & ~n9620 ) | ( n9630 & n9634 ) | ( ~n9620 & n9634 ) ;
  assign n9636 = ( n9620 & ~n9630 ) | ( n9620 & n9634 ) | ( ~n9630 & n9634 ) ;
  assign n9637 = ( n9635 & ~n9634 ) | ( n9635 & n9636 ) | ( ~n9634 & n9636 ) ;
  assign n9344 = ~n136 & x126 ;
  assign n9341 = ( x124 & ~n150 ) | ( x124 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n9342 = ( x125 & ~n131 ) | ( x125 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n9343 = n9341 | n9342 ;
  assign n9345 = ( x126 & ~n9344 ) | ( x126 & n9343 ) | ( ~n9344 & n9343 ) ;
  assign n9346 = ( x124 & x125 ) | ( x124 & n9318 ) | ( x125 & n9318 ) ;
  assign n9347 = ( x125 & ~x126 ) | ( x125 & n9346 ) | ( ~x126 & n9346 ) ;
  assign n9348 = ( x125 & x126 ) | ( x125 & n9346 ) | ( x126 & n9346 ) ;
  assign n9349 = ( ~x126 & ~n9347 ) | ( ~x126 & n9348 ) | ( ~n9347 & n9348 ) ;
  assign n9350 = n139 | n9349 ;
  assign n9351 = ~n9345 & n9350 ;
  assign n9638 = ( x2 & ~n9637 ) | ( x2 & n9351 ) | ( ~n9637 & n9351 ) ;
  assign n9639 = ( x2 & ~n9351 ) | ( x2 & n9637 ) | ( ~n9351 & n9637 ) ;
  assign n9640 = ( n9638 & ~x2 ) | ( n9638 & n9639 ) | ( ~x2 & n9639 ) ;
  assign n9641 = ( n9339 & ~n9340 ) | ( n9339 & n9640 ) | ( ~n9340 & n9640 ) ;
  assign n9642 = ( n9339 & ~n9640 ) | ( n9339 & n9340 ) | ( ~n9640 & n9340 ) ;
  assign n9643 = ( n9641 & ~n9339 ) | ( n9641 & n9642 ) | ( ~n9339 & n9642 ) ;
  assign n9649 = ( n9357 & ~n9617 ) | ( n9357 & 1'b0 ) | ( ~n9617 & 1'b0 ) ;
  assign n9650 = ~n9357 & n9617 ;
  assign n9651 = n9649 | n9650 ;
  assign n9652 = ( n9369 & n9630 ) | ( n9369 & n9651 ) | ( n9630 & n9651 ) ;
  assign n9663 = x14 &  n9392 ;
  assign n9664 = x14 | n9392 ;
  assign n9665 = ~n9663 & n9664 ;
  assign n9666 = ( n9375 & ~n9611 ) | ( n9375 & n9665 ) | ( ~n9611 & n9665 ) ;
  assign n9670 = x116 &  n503 ;
  assign n9667 = ( x118 & ~n450 ) | ( x118 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n9668 = x117 &  n445 ;
  assign n9669 = n9667 | n9668 ;
  assign n9671 = ( x116 & ~n9670 ) | ( x116 & n9669 ) | ( ~n9670 & n9669 ) ;
  assign n9672 = n453 | n7152 ;
  assign n9673 = ~n9671 & n9672 ;
  assign n9674 = x11 &  n9673 ;
  assign n9675 = x11 | n9673 ;
  assign n9676 = ~n9674 & n9675 ;
  assign n9687 = x110 &  n942 ;
  assign n9684 = ( x112 & ~n896 ) | ( x112 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n9685 = x111 &  n891 ;
  assign n9686 = n9684 | n9685 ;
  assign n9688 = ( x110 & ~n9687 ) | ( x110 & n9686 ) | ( ~n9687 & n9686 ) ;
  assign n9689 = ~n899 & n5727 ;
  assign n9690 = n9688 | n9689 ;
  assign n9691 = ( x17 & ~n9690 ) | ( x17 & 1'b0 ) | ( ~n9690 & 1'b0 ) ;
  assign n9692 = ~x17 & n9690 ;
  assign n9693 = n9691 | n9692 ;
  assign n9694 = ( n9597 & ~n9598 ) | ( n9597 & n9608 ) | ( ~n9598 & n9608 ) ;
  assign n9698 = x107 &  n1227 ;
  assign n9695 = ( x109 & ~n1154 ) | ( x109 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n9696 = x108 &  n1149 ;
  assign n9697 = n9695 | n9696 ;
  assign n9699 = ( x107 & ~n9698 ) | ( x107 & n9697 ) | ( ~n9698 & n9697 ) ;
  assign n9700 = ~n1157 & n5267 ;
  assign n9701 = n9699 | n9700 ;
  assign n9702 = ( x20 & ~n9701 ) | ( x20 & 1'b0 ) | ( ~n9701 & 1'b0 ) ;
  assign n9703 = ~x20 & n9701 ;
  assign n9704 = n9702 | n9703 ;
  assign n9705 = ( n9583 & ~n9594 ) | ( n9583 & n9584 ) | ( ~n9594 & n9584 ) ;
  assign n9709 = x104 &  n1551 ;
  assign n9706 = ( x106 & ~n1451 ) | ( x106 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n9707 = x105 &  n1446 ;
  assign n9708 = n9706 | n9707 ;
  assign n9710 = ( x104 & ~n9709 ) | ( x104 & n9708 ) | ( ~n9709 & n9708 ) ;
  assign n9711 = ~n1454 & n4458 ;
  assign n9712 = n9710 | n9711 ;
  assign n9713 = ( x23 & ~n9712 ) | ( x23 & 1'b0 ) | ( ~n9712 & 1'b0 ) ;
  assign n9714 = ~x23 & n9712 ;
  assign n9715 = n9713 | n9714 ;
  assign n9740 = x86 &  n4344 ;
  assign n9737 = ( x88 & ~n4143 ) | ( x88 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n9738 = x87 &  n4138 ;
  assign n9739 = n9737 | n9738 ;
  assign n9741 = ( x86 & ~n9740 ) | ( x86 & n9739 ) | ( ~n9740 & n9739 ) ;
  assign n9742 = ( n1624 & ~n4146 ) | ( n1624 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n9743 = n9741 | n9742 ;
  assign n9744 = ( x41 & ~n9743 ) | ( x41 & 1'b0 ) | ( ~n9743 & 1'b0 ) ;
  assign n9745 = ~x41 & n9743 ;
  assign n9746 = n9744 | n9745 ;
  assign n9750 = x83 &  n4934 ;
  assign n9747 = ( x85 & ~n4725 ) | ( x85 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n9748 = x84 &  n4720 ;
  assign n9749 = n9747 | n9748 ;
  assign n9751 = ( x83 & ~n9750 ) | ( x83 & n9749 ) | ( ~n9750 & n9749 ) ;
  assign n9752 = ( n1295 & ~n4728 ) | ( n1295 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n9753 = n9751 | n9752 ;
  assign n9754 = ( x44 & ~n9753 ) | ( x44 & 1'b0 ) | ( ~n9753 & 1'b0 ) ;
  assign n9755 = ~x44 & n9753 ;
  assign n9756 = n9754 | n9755 ;
  assign n9757 = ( n9515 & n9516 ) | ( n9515 & n9526 ) | ( n9516 & n9526 ) ;
  assign n9822 = x77 &  n6288 ;
  assign n9819 = ( x79 & ~n6032 ) | ( x79 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n9820 = x78 &  n6027 ;
  assign n9821 = n9819 | n9820 ;
  assign n9823 = ( x77 & ~n9822 ) | ( x77 & n9821 ) | ( ~n9822 & n9821 ) ;
  assign n9824 = ( n766 & ~n6035 ) | ( n766 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n9825 = n9823 | n9824 ;
  assign n9826 = ( x50 & ~n9825 ) | ( x50 & 1'b0 ) | ( ~n9825 & 1'b0 ) ;
  assign n9827 = ~x50 & n9825 ;
  assign n9828 = n9826 | n9827 ;
  assign n9809 = x74 &  n6982 ;
  assign n9806 = ( x76 & ~n6727 ) | ( x76 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n9807 = x75 &  n6722 ;
  assign n9808 = n9806 | n9807 ;
  assign n9810 = ( x74 & ~n9809 ) | ( x74 & n9808 ) | ( ~n9809 & n9808 ) ;
  assign n9811 = ( n603 & ~n6730 ) | ( n603 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n9812 = n9810 | n9811 ;
  assign n9813 = ( x53 & ~n9812 ) | ( x53 & 1'b0 ) | ( ~n9812 & 1'b0 ) ;
  assign n9814 = ~x53 & n9812 ;
  assign n9815 = n9813 | n9814 ;
  assign n9758 = ( x62 & ~x63 ) | ( x62 & 1'b0 ) | ( ~x63 & 1'b0 ) ;
  assign n9759 = ~x62 & x63 ;
  assign n9760 = ~n9758 &  ~n9759 ;
  assign n9761 = ( x64 & ~n9760 ) | ( x64 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n9762 = ( n8881 & ~n9155 ) | ( n8881 & n9464 ) | ( ~n9155 & n9464 ) ;
  assign n9763 = ( x62 & n9155 ) | ( x62 & n9762 ) | ( n9155 & n9762 ) ;
  assign n9764 = ( x62 & ~n9763 ) | ( x62 & 1'b0 ) | ( ~n9763 & 1'b0 ) ;
  assign n9768 = x65 &  n9457 ;
  assign n9765 = ( x67 & ~n9150 ) | ( x67 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n9766 = x66 &  n9145 ;
  assign n9767 = n9765 | n9766 ;
  assign n9769 = ( x65 & ~n9768 ) | ( x65 & n9767 ) | ( ~n9768 & n9767 ) ;
  assign n9770 = n173 | n9153 ;
  assign n9771 = ~n9769 & n9770 ;
  assign n9772 = x62 &  n9771 ;
  assign n9773 = x62 | n9771 ;
  assign n9774 = ~n9772 & n9773 ;
  assign n9775 = ( n9761 & ~n9764 ) | ( n9761 & n9774 ) | ( ~n9764 & n9774 ) ;
  assign n9776 = ( n9761 & ~n9774 ) | ( n9761 & n9764 ) | ( ~n9774 & n9764 ) ;
  assign n9777 = ( n9775 & ~n9761 ) | ( n9775 & n9776 ) | ( ~n9761 & n9776 ) ;
  assign n9782 = x68 &  n8558 ;
  assign n9779 = ( x70 & ~n8314 ) | ( x70 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n9780 = x69 &  n8309 ;
  assign n9781 = n9779 | n9780 ;
  assign n9783 = ( x68 & ~n9782 ) | ( x68 & n9781 ) | ( ~n9782 & n9781 ) ;
  assign n9784 = ( n282 & ~n8317 ) | ( n282 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n9785 = n9783 | n9784 ;
  assign n9786 = ( x59 & ~n9785 ) | ( x59 & 1'b0 ) | ( ~n9785 & 1'b0 ) ;
  assign n9787 = ~x59 & n9785 ;
  assign n9788 = n9786 | n9787 ;
  assign n9778 = ( n9160 & n9469 ) | ( n9160 & n9479 ) | ( n9469 & n9479 ) ;
  assign n9789 = ( n9777 & ~n9788 ) | ( n9777 & n9778 ) | ( ~n9788 & n9778 ) ;
  assign n9790 = ( n9777 & ~n9778 ) | ( n9777 & n9788 ) | ( ~n9778 & n9788 ) ;
  assign n9791 = ( n9789 & ~n9777 ) | ( n9789 & n9790 ) | ( ~n9777 & n9790 ) ;
  assign n9792 = ( n9163 & n9482 ) | ( n9163 & n9492 ) | ( n9482 & n9492 ) ;
  assign n9796 = x71 &  n7731 ;
  assign n9793 = ( x73 & ~n7538 ) | ( x73 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n9794 = x72 &  n7533 ;
  assign n9795 = n9793 | n9794 ;
  assign n9797 = ( x71 & ~n9796 ) | ( x71 & n9795 ) | ( ~n9796 & n9795 ) ;
  assign n9798 = ( n389 & ~n7541 ) | ( n389 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n9799 = n9797 | n9798 ;
  assign n9800 = ( x56 & ~n9799 ) | ( x56 & 1'b0 ) | ( ~n9799 & 1'b0 ) ;
  assign n9801 = ~x56 & n9799 ;
  assign n9802 = n9800 | n9801 ;
  assign n9803 = ( n9791 & ~n9792 ) | ( n9791 & n9802 ) | ( ~n9792 & n9802 ) ;
  assign n9804 = ( n9792 & ~n9791 ) | ( n9792 & n9802 ) | ( ~n9791 & n9802 ) ;
  assign n9805 = ( n9803 & ~n9802 ) | ( n9803 & n9804 ) | ( ~n9802 & n9804 ) ;
  assign n9816 = ( n9497 & ~n9815 ) | ( n9497 & n9805 ) | ( ~n9815 & n9805 ) ;
  assign n9817 = ( n9805 & ~n9497 ) | ( n9805 & n9815 ) | ( ~n9497 & n9815 ) ;
  assign n9818 = ( n9816 & ~n9805 ) | ( n9816 & n9817 ) | ( ~n9805 & n9817 ) ;
  assign n9829 = ( n9511 & ~n9828 ) | ( n9511 & n9818 ) | ( ~n9828 & n9818 ) ;
  assign n9830 = ( n9818 & ~n9511 ) | ( n9818 & n9828 ) | ( ~n9511 & n9828 ) ;
  assign n9831 = ( n9829 & ~n9818 ) | ( n9829 & n9830 ) | ( ~n9818 & n9830 ) ;
  assign n9835 = x80 &  n5586 ;
  assign n9832 = ( x82 & ~n5389 ) | ( x82 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n9833 = x81 &  n5384 ;
  assign n9834 = n9832 | n9833 ;
  assign n9836 = ( x80 & ~n9835 ) | ( x80 & n9834 ) | ( ~n9835 & n9834 ) ;
  assign n9837 = ( n1084 & ~n5392 ) | ( n1084 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n9838 = n9836 | n9837 ;
  assign n9839 = ( x47 & ~n9838 ) | ( x47 & 1'b0 ) | ( ~n9838 & 1'b0 ) ;
  assign n9840 = ~x47 & n9838 ;
  assign n9841 = n9839 | n9840 ;
  assign n9842 = ( n9831 & ~n9514 ) | ( n9831 & n9841 ) | ( ~n9514 & n9841 ) ;
  assign n9843 = ( n9514 & ~n9841 ) | ( n9514 & n9831 ) | ( ~n9841 & n9831 ) ;
  assign n9844 = ( n9842 & ~n9831 ) | ( n9842 & n9843 ) | ( ~n9831 & n9843 ) ;
  assign n9845 = ( n9756 & ~n9757 ) | ( n9756 & n9844 ) | ( ~n9757 & n9844 ) ;
  assign n9846 = ( n9756 & ~n9844 ) | ( n9756 & n9757 ) | ( ~n9844 & n9757 ) ;
  assign n9847 = ( n9845 & ~n9756 ) | ( n9845 & n9846 ) | ( ~n9756 & n9846 ) ;
  assign n9848 = ( n9529 & n9530 ) | ( n9529 & n9540 ) | ( n9530 & n9540 ) ;
  assign n9849 = ( n9746 & ~n9847 ) | ( n9746 & n9848 ) | ( ~n9847 & n9848 ) ;
  assign n9850 = ( n9746 & ~n9848 ) | ( n9746 & n9847 ) | ( ~n9848 & n9847 ) ;
  assign n9851 = ( n9849 & ~n9746 ) | ( n9849 & n9850 ) | ( ~n9746 & n9850 ) ;
  assign n9730 = x89 &  n3756 ;
  assign n9727 = ( x91 & ~n3602 ) | ( x91 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n9728 = x90 &  n3597 ;
  assign n9729 = n9727 | n9728 ;
  assign n9731 = ( x89 & ~n9730 ) | ( x89 & n9729 ) | ( ~n9730 & n9729 ) ;
  assign n9732 = ( n2108 & ~n3605 ) | ( n2108 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n9733 = n9731 | n9732 ;
  assign n9734 = ( x38 & ~n9733 ) | ( x38 & 1'b0 ) | ( ~n9733 & 1'b0 ) ;
  assign n9735 = ~x38 & n9733 ;
  assign n9736 = n9734 | n9735 ;
  assign n9852 = ( n9544 & ~n9851 ) | ( n9544 & n9736 ) | ( ~n9851 & n9736 ) ;
  assign n9853 = ( n9736 & ~n9544 ) | ( n9736 & n9851 ) | ( ~n9544 & n9851 ) ;
  assign n9854 = ( n9852 & ~n9736 ) | ( n9852 & n9853 ) | ( ~n9736 & n9853 ) ;
  assign n9720 = x92 &  n3214 ;
  assign n9717 = ( x94 & ~n3087 ) | ( x94 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n9718 = x93 &  n3082 ;
  assign n9719 = n9717 | n9718 ;
  assign n9721 = ( x92 & ~n9720 ) | ( x92 & n9719 ) | ( ~n9720 & n9719 ) ;
  assign n9722 = ( n2401 & ~n3090 ) | ( n2401 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n9723 = n9721 | n9722 ;
  assign n9724 = ( x35 & ~n9723 ) | ( x35 & 1'b0 ) | ( ~n9723 & 1'b0 ) ;
  assign n9725 = ~x35 & n9723 ;
  assign n9726 = n9724 | n9725 ;
  assign n9855 = ( n9547 & ~n9854 ) | ( n9547 & n9726 ) | ( ~n9854 & n9726 ) ;
  assign n9856 = ( n9726 & ~n9547 ) | ( n9726 & n9854 ) | ( ~n9547 & n9854 ) ;
  assign n9857 = ( n9855 & ~n9726 ) | ( n9855 & n9856 ) | ( ~n9726 & n9856 ) ;
  assign n9858 = ( n9550 & ~n9549 ) | ( n9550 & n9560 ) | ( ~n9549 & n9560 ) ;
  assign n9862 = x95 &  n2718 ;
  assign n9859 = ( x97 & ~n2642 ) | ( x97 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n9860 = x96 &  n2637 ;
  assign n9861 = n9859 | n9860 ;
  assign n9863 = ( x95 & ~n9862 ) | ( x95 & n9861 ) | ( ~n9862 & n9861 ) ;
  assign n9864 = ~n2645 & n2999 ;
  assign n9865 = n9863 | n9864 ;
  assign n9866 = ( x32 & ~n9865 ) | ( x32 & 1'b0 ) | ( ~n9865 & 1'b0 ) ;
  assign n9867 = ~x32 & n9865 ;
  assign n9868 = n9866 | n9867 ;
  assign n9869 = ( n9857 & ~n9858 ) | ( n9857 & n9868 ) | ( ~n9858 & n9868 ) ;
  assign n9870 = ( n9858 & ~n9857 ) | ( n9858 & n9868 ) | ( ~n9857 & n9868 ) ;
  assign n9871 = ( n9869 & ~n9868 ) | ( n9869 & n9870 ) | ( ~n9868 & n9870 ) ;
  assign n9872 = ( n9412 & ~n9563 ) | ( n9412 & n9564 ) | ( ~n9563 & n9564 ) ;
  assign n9876 = x98 &  n2312 ;
  assign n9873 = ( x100 & ~n2195 ) | ( x100 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n9874 = x99 &  n2190 ;
  assign n9875 = n9873 | n9874 ;
  assign n9877 = ( x98 & ~n9876 ) | ( x98 & n9875 ) | ( ~n9876 & n9875 ) ;
  assign n9878 = n2198 | n3354 ;
  assign n9879 = ~n9877 & n9878 ;
  assign n9880 = x29 &  n9879 ;
  assign n9881 = x29 | n9879 ;
  assign n9882 = ~n9880 & n9881 ;
  assign n9883 = ( n9871 & n9872 ) | ( n9871 & n9882 ) | ( n9872 & n9882 ) ;
  assign n9884 = ( n9872 & ~n9871 ) | ( n9872 & n9882 ) | ( ~n9871 & n9882 ) ;
  assign n9885 = ( n9871 & ~n9883 ) | ( n9871 & n9884 ) | ( ~n9883 & n9884 ) ;
  assign n9889 = x101 &  n1894 ;
  assign n9886 = ( x103 & ~n1816 ) | ( x103 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n9887 = x102 &  n1811 ;
  assign n9888 = n9886 | n9887 ;
  assign n9890 = ( x101 & ~n9889 ) | ( x101 & n9888 ) | ( ~n9889 & n9888 ) ;
  assign n9891 = n1819 | n4056 ;
  assign n9892 = ~n9890 & n9891 ;
  assign n9893 = x26 &  n9892 ;
  assign n9894 = x26 | n9892 ;
  assign n9895 = ~n9893 & n9894 ;
  assign n9896 = ( n9885 & ~n9568 ) | ( n9885 & n9895 ) | ( ~n9568 & n9895 ) ;
  assign n9897 = ( n9568 & ~n9895 ) | ( n9568 & n9885 ) | ( ~n9895 & n9885 ) ;
  assign n9898 = ( n9896 & ~n9885 ) | ( n9896 & n9897 ) | ( ~n9885 & n9897 ) ;
  assign n9716 = ( n9248 & ~n9580 ) | ( n9248 & n9570 ) | ( ~n9580 & n9570 ) ;
  assign n9899 = ( n9715 & ~n9898 ) | ( n9715 & n9716 ) | ( ~n9898 & n9716 ) ;
  assign n9900 = ( n9715 & ~n9716 ) | ( n9715 & n9898 ) | ( ~n9716 & n9898 ) ;
  assign n9901 = ( n9899 & ~n9715 ) | ( n9899 & n9900 ) | ( ~n9715 & n9900 ) ;
  assign n9902 = ( n9704 & ~n9705 ) | ( n9704 & n9901 ) | ( ~n9705 & n9901 ) ;
  assign n9903 = ( n9704 & ~n9901 ) | ( n9704 & n9705 ) | ( ~n9901 & n9705 ) ;
  assign n9904 = ( n9902 & ~n9704 ) | ( n9902 & n9903 ) | ( ~n9704 & n9903 ) ;
  assign n9905 = ( n9693 & n9694 ) | ( n9693 & n9904 ) | ( n9694 & n9904 ) ;
  assign n9906 = ( n9694 & ~n9693 ) | ( n9694 & n9904 ) | ( ~n9693 & n9904 ) ;
  assign n9907 = ( n9693 & ~n9905 ) | ( n9693 & n9906 ) | ( ~n9905 & n9906 ) ;
  assign n9680 = x113 &  n713 ;
  assign n9677 = ( x115 & ~n641 ) | ( x115 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n9678 = x114 &  n636 ;
  assign n9679 = n9677 | n9678 ;
  assign n9681 = ( x113 & ~n9680 ) | ( x113 & n9679 ) | ( ~n9680 & n9679 ) ;
  assign n9682 = ~n644 & n6420 ;
  assign n9683 = n9681 | n9682 ;
  assign n9909 = ( x14 & n9683 ) | ( x14 & n9907 ) | ( n9683 & n9907 ) ;
  assign n9908 = ( x14 & ~n9907 ) | ( x14 & n9683 ) | ( ~n9907 & n9683 ) ;
  assign n9910 = ( n9907 & ~n9909 ) | ( n9907 & n9908 ) | ( ~n9909 & n9908 ) ;
  assign n9911 = ( n9666 & n9676 ) | ( n9666 & n9910 ) | ( n9676 & n9910 ) ;
  assign n9912 = ( n9676 & ~n9666 ) | ( n9676 & n9910 ) | ( ~n9666 & n9910 ) ;
  assign n9913 = ( n9666 & ~n9911 ) | ( n9666 & n9912 ) | ( ~n9911 & n9912 ) ;
  assign n9924 = n9375 &  n9614 ;
  assign n9925 = n9375 | n9614 ;
  assign n9926 = ~n9924 & n9925 ;
  assign n9927 = ( n9357 & ~n9926 ) | ( n9357 & n9385 ) | ( ~n9926 & n9385 ) ;
  assign n9917 = x119 &  n353 ;
  assign n9914 = ( x121 & ~n313 ) | ( x121 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n9915 = x120 &  n308 ;
  assign n9916 = n9914 | n9915 ;
  assign n9918 = ( x119 & ~n9917 ) | ( x119 & n9916 ) | ( ~n9917 & n9916 ) ;
  assign n9919 = ~n316 & n8176 ;
  assign n9920 = n9918 | n9919 ;
  assign n9921 = ( x8 & ~n9920 ) | ( x8 & 1'b0 ) | ( ~n9920 & 1'b0 ) ;
  assign n9922 = ~x8 & n9920 ;
  assign n9923 = n9921 | n9922 ;
  assign n9928 = ( n9913 & ~n9927 ) | ( n9913 & n9923 ) | ( ~n9927 & n9923 ) ;
  assign n9929 = ( n9913 & ~n9923 ) | ( n9913 & n9927 ) | ( ~n9923 & n9927 ) ;
  assign n9930 = ( n9928 & ~n9913 ) | ( n9928 & n9929 ) | ( ~n9913 & n9929 ) ;
  assign n9656 = x122 &  n225 ;
  assign n9653 = ( x124 & ~n197 ) | ( x124 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n9654 = x123 &  n192 ;
  assign n9655 = n9653 | n9654 ;
  assign n9657 = ( x122 & ~n9656 ) | ( x122 & n9655 ) | ( ~n9656 & n9655 ) ;
  assign n9658 = ( n8749 & ~n200 ) | ( n8749 & n8752 ) | ( ~n200 & n8752 ) ;
  assign n9659 = ( n9657 & ~n8753 ) | ( n9657 & n9658 ) | ( ~n8753 & n9658 ) ;
  assign n9660 = ( x5 & ~n9659 ) | ( x5 & 1'b0 ) | ( ~n9659 & 1'b0 ) ;
  assign n9661 = ~x5 & n9659 ;
  assign n9662 = n9660 | n9661 ;
  assign n9931 = ( n9652 & ~n9930 ) | ( n9652 & n9662 ) | ( ~n9930 & n9662 ) ;
  assign n9932 = ( n9652 & ~n9662 ) | ( n9652 & n9930 ) | ( ~n9662 & n9930 ) ;
  assign n9933 = ( n9931 & ~n9652 ) | ( n9931 & n9932 ) | ( ~n9652 & n9932 ) ;
  assign n9937 = ~n136 & x127 ;
  assign n9934 = ( x125 & ~n150 ) | ( x125 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n9935 = ( x126 & ~n131 ) | ( x126 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n9936 = n9934 | n9935 ;
  assign n9938 = ( x127 & ~n9937 ) | ( x127 & n9936 ) | ( ~n9937 & n9936 ) ;
  assign n9939 = ( x126 & ~x127 ) | ( x126 & n9348 ) | ( ~x127 & n9348 ) ;
  assign n9940 = ( x126 & x127 ) | ( x126 & n9348 ) | ( x127 & n9348 ) ;
  assign n9941 = ( ~x127 & ~n9939 ) | ( ~x127 & n9940 ) | ( ~n9939 & n9940 ) ;
  assign n9942 = n139 | n9941 ;
  assign n9943 = ~n9938 & n9942 ;
  assign n9945 = ( x2 & n9933 ) | ( x2 & n9943 ) | ( n9933 & n9943 ) ;
  assign n9944 = ( n9933 & ~x2 ) | ( n9933 & n9943 ) | ( ~x2 & n9943 ) ;
  assign n9946 = ( x2 & ~n9945 ) | ( x2 & n9944 ) | ( ~n9945 & n9944 ) ;
  assign n9647 = ( x2 & ~n9351 ) | ( x2 & 1'b0 ) | ( ~n9351 & 1'b0 ) ;
  assign n9644 = ( n9620 & ~n9634 ) | ( n9620 & n9630 ) | ( ~n9634 & n9630 ) ;
  assign n9645 = ( n9620 & n9630 ) | ( n9620 & n9634 ) | ( n9630 & n9634 ) ;
  assign n9646 = ~n9644 & n9645 ;
  assign n9648 = ( n9639 & ~n9647 ) | ( n9639 & n9646 ) | ( ~n9647 & n9646 ) ;
  assign n9947 = ( n9642 & ~n9946 ) | ( n9642 & n9648 ) | ( ~n9946 & n9648 ) ;
  assign n9948 = ( n9648 & ~n9642 ) | ( n9648 & n9946 ) | ( ~n9642 & n9946 ) ;
  assign n9949 = ( n9947 & ~n9648 ) | ( n9947 & n9948 ) | ( ~n9648 & n9948 ) ;
  assign n9950 = n9931 &  n9932 ;
  assign n9951 = ( x2 & ~n9943 ) | ( x2 & 1'b0 ) | ( ~n9943 & 1'b0 ) ;
  assign n9952 = ( n9944 & ~n9950 ) | ( n9944 & n9951 ) | ( ~n9950 & n9951 ) ;
  assign n9963 = n9666 &  n9910 ;
  assign n9964 = n9666 | n9910 ;
  assign n9965 = ~n9963 & n9964 ;
  assign n9966 = ( n9676 & ~n9965 ) | ( n9676 & n9927 ) | ( ~n9965 & n9927 ) ;
  assign n9967 = ( n9927 & ~n9676 ) | ( n9927 & n9965 ) | ( ~n9676 & n9965 ) ;
  assign n9968 = ( n9966 & ~n9927 ) | ( n9966 & n9967 ) | ( ~n9927 & n9967 ) ;
  assign n9969 = ( n9662 & ~n9968 ) | ( n9662 & n9923 ) | ( ~n9968 & n9923 ) ;
  assign n9980 = ( n9676 & n9927 ) | ( n9676 & n9965 ) | ( n9927 & n9965 ) ;
  assign n9984 = x120 &  n353 ;
  assign n9981 = ( x122 & ~n313 ) | ( x122 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n9982 = x121 &  n308 ;
  assign n9983 = n9981 | n9982 ;
  assign n9985 = ( x120 & ~n9984 ) | ( x120 & n9983 ) | ( ~n9984 & n9983 ) ;
  assign n9986 = n8448 | n8451 ;
  assign n9987 = ~n8452 & n9986 ;
  assign n9988 = ~n316 & n9987 ;
  assign n9989 = n9985 | n9988 ;
  assign n9990 = ( x8 & ~n9989 ) | ( x8 & 1'b0 ) | ( ~n9989 & 1'b0 ) ;
  assign n9991 = ~x8 & n9989 ;
  assign n9992 = n9990 | n9991 ;
  assign n10228 = x117 &  n503 ;
  assign n10225 = ( x119 & ~n450 ) | ( x119 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n10226 = x118 &  n445 ;
  assign n10227 = n10225 | n10226 ;
  assign n10229 = ( x117 & ~n10228 ) | ( x117 & n10227 ) | ( ~n10228 & n10227 ) ;
  assign n10230 = ~n453 & n7648 ;
  assign n10231 = n10229 | n10230 ;
  assign n10232 = ~x11 & n10231 ;
  assign n10233 = x11 | n10231 ;
  assign n10234 = ( n10232 & ~n10231 ) | ( n10232 & n10233 ) | ( ~n10231 & n10233 ) ;
  assign n9993 = ( x14 & ~n9683 ) | ( x14 & 1'b0 ) | ( ~n9683 & 1'b0 ) ;
  assign n9994 = ~x14 & n9683 ;
  assign n9995 = n9993 | n9994 ;
  assign n9996 = ( n9907 & ~n9666 ) | ( n9907 & n9995 ) | ( ~n9666 & n9995 ) ;
  assign n10000 = x114 &  n713 ;
  assign n9997 = ( x116 & ~n641 ) | ( x116 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n9998 = x115 &  n636 ;
  assign n9999 = n9997 | n9998 ;
  assign n10001 = ( x114 & ~n10000 ) | ( x114 & n9999 ) | ( ~n10000 & n9999 ) ;
  assign n10002 = n644 | n6885 ;
  assign n10003 = ~n10001 & n10002 ;
  assign n10007 = x111 &  n942 ;
  assign n10004 = ( x113 & ~n896 ) | ( x113 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n10005 = x112 &  n891 ;
  assign n10006 = n10004 | n10005 ;
  assign n10008 = ( x111 & ~n10007 ) | ( x111 & n10006 ) | ( ~n10007 & n10006 ) ;
  assign n10009 = n899 | n6169 ;
  assign n10010 = ~n10008 & n10009 ;
  assign n10011 = x17 &  n10010 ;
  assign n10012 = x17 | n10010 ;
  assign n10013 = ~n10011 & n10012 ;
  assign n10017 = x108 &  n1227 ;
  assign n10014 = ( x110 & ~n1154 ) | ( x110 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n10015 = x109 &  n1149 ;
  assign n10016 = n10014 | n10015 ;
  assign n10018 = ( x108 & ~n10017 ) | ( x108 & n10016 ) | ( ~n10017 & n10016 ) ;
  assign n10019 = n1157 | n5283 ;
  assign n10020 = ~n10018 & n10019 ;
  assign n10021 = x20 &  n10020 ;
  assign n10022 = x20 | n10020 ;
  assign n10023 = ~n10021 & n10022 ;
  assign n10027 = x102 &  n1894 ;
  assign n10024 = ( x104 & ~n1816 ) | ( x104 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n10025 = x103 &  n1811 ;
  assign n10026 = n10024 | n10025 ;
  assign n10028 = ( x102 & ~n10027 ) | ( x102 & n10026 ) | ( ~n10027 & n10026 ) ;
  assign n10029 = n1819 | n4249 ;
  assign n10030 = ~n10028 & n10029 ;
  assign n10031 = x26 &  n10030 ;
  assign n10032 = x26 | n10030 ;
  assign n10033 = ~n10031 & n10032 ;
  assign n10037 = x99 &  n2312 ;
  assign n10034 = ( x101 & ~n2195 ) | ( x101 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n10035 = x100 &  n2190 ;
  assign n10036 = n10034 | n10035 ;
  assign n10038 = ( x99 & ~n10037 ) | ( x99 & n10036 ) | ( ~n10037 & n10036 ) ;
  assign n10039 = n2198 | n3694 ;
  assign n10040 = ~n10038 & n10039 ;
  assign n10041 = x29 &  n10040 ;
  assign n10042 = x29 | n10040 ;
  assign n10043 = ~n10041 & n10042 ;
  assign n10047 = x93 &  n3214 ;
  assign n10044 = ( x95 & ~n3087 ) | ( x95 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n10045 = x94 &  n3082 ;
  assign n10046 = n10044 | n10045 ;
  assign n10048 = ( x93 & ~n10047 ) | ( x93 & n10046 ) | ( ~n10047 & n10046 ) ;
  assign n10049 = ( n2547 & ~n3090 ) | ( n2547 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n10050 = n10048 | n10049 ;
  assign n10051 = ( x35 & ~n10050 ) | ( x35 & 1'b0 ) | ( ~n10050 & 1'b0 ) ;
  assign n10052 = ~x35 & n10050 ;
  assign n10053 = n10051 | n10052 ;
  assign n10057 = x90 &  n3756 ;
  assign n10054 = ( x92 & ~n3602 ) | ( x92 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n10055 = x91 &  n3597 ;
  assign n10056 = n10054 | n10055 ;
  assign n10058 = ( x90 & ~n10057 ) | ( x90 & n10056 ) | ( ~n10057 & n10056 ) ;
  assign n10059 = ( n2248 & ~n3605 ) | ( n2248 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n10060 = n10058 | n10059 ;
  assign n10061 = ( x38 & ~n10060 ) | ( x38 & 1'b0 ) | ( ~n10060 & 1'b0 ) ;
  assign n10062 = ~x38 & n10060 ;
  assign n10063 = n10061 | n10062 ;
  assign n10067 = x87 &  n4344 ;
  assign n10064 = ( x89 & ~n4143 ) | ( x89 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n10065 = x88 &  n4138 ;
  assign n10066 = n10064 | n10065 ;
  assign n10068 = ( x87 & ~n10067 ) | ( x87 & n10066 ) | ( ~n10067 & n10066 ) ;
  assign n10069 = ( n1741 & ~n4146 ) | ( n1741 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n10070 = n10068 | n10069 ;
  assign n10071 = ( x41 & ~n10070 ) | ( x41 & 1'b0 ) | ( ~n10070 & 1'b0 ) ;
  assign n10072 = ~x41 & n10070 ;
  assign n10073 = n10071 | n10072 ;
  assign n10077 = x81 &  n5586 ;
  assign n10074 = ( x83 & ~n5389 ) | ( x83 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n10075 = x82 &  n5384 ;
  assign n10076 = n10074 | n10075 ;
  assign n10078 = ( x81 & ~n10077 ) | ( x81 & n10076 ) | ( ~n10077 & n10076 ) ;
  assign n10079 = ( n1100 & ~n5392 ) | ( n1100 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n10080 = n10078 | n10079 ;
  assign n10081 = ( x47 & ~n10080 ) | ( x47 & 1'b0 ) | ( ~n10080 & 1'b0 ) ;
  assign n10082 = ~x47 & n10080 ;
  assign n10083 = n10081 | n10082 ;
  assign n10087 = x75 &  n6982 ;
  assign n10084 = ( x77 & ~n6727 ) | ( x77 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n10085 = x76 &  n6722 ;
  assign n10086 = n10084 | n10085 ;
  assign n10088 = ( x75 & ~n10087 ) | ( x75 & n10086 ) | ( ~n10087 & n10086 ) ;
  assign n10089 = ( n677 & ~n6730 ) | ( n677 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n10090 = n10088 | n10089 ;
  assign n10091 = ( x53 & ~n10090 ) | ( x53 & 1'b0 ) | ( ~n10090 & 1'b0 ) ;
  assign n10092 = ~x53 & n10090 ;
  assign n10093 = n10091 | n10092 ;
  assign n10104 = x62 &  x63 ;
  assign n10105 = x64 &  n10104 ;
  assign n10106 = ( x65 & ~n9760 ) | ( x65 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n10107 = n10105 | n10106 ;
  assign n10097 = x66 &  n9457 ;
  assign n10094 = ( x68 & ~n9150 ) | ( x68 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n10095 = x67 &  n9145 ;
  assign n10096 = n10094 | n10095 ;
  assign n10098 = ( x66 & ~n10097 ) | ( x66 & n10096 ) | ( ~n10097 & n10096 ) ;
  assign n10099 = ( n213 & ~n9153 ) | ( n213 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n10100 = n10098 | n10099 ;
  assign n10101 = ( x62 & ~n10100 ) | ( x62 & 1'b0 ) | ( ~n10100 & 1'b0 ) ;
  assign n10102 = ~x62 & n10100 ;
  assign n10103 = n10101 | n10102 ;
  assign n10108 = ( n9776 & ~n10107 ) | ( n9776 & n10103 ) | ( ~n10107 & n10103 ) ;
  assign n10109 = ( n10103 & ~n9776 ) | ( n10103 & n10107 ) | ( ~n9776 & n10107 ) ;
  assign n10110 = ( n10108 & ~n10103 ) | ( n10108 & n10109 ) | ( ~n10103 & n10109 ) ;
  assign n10115 = x69 &  n8558 ;
  assign n10112 = ( x71 & ~n8314 ) | ( x71 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n10113 = x70 &  n8309 ;
  assign n10114 = n10112 | n10113 ;
  assign n10116 = ( x69 & ~n10115 ) | ( x69 & n10114 ) | ( ~n10115 & n10114 ) ;
  assign n10117 = ( n298 & ~n8317 ) | ( n298 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n10118 = n10116 | n10117 ;
  assign n10119 = ( x59 & ~n10118 ) | ( x59 & 1'b0 ) | ( ~n10118 & 1'b0 ) ;
  assign n10120 = ~x59 & n10118 ;
  assign n10121 = n10119 | n10120 ;
  assign n10111 = ( n9778 & ~n9777 ) | ( n9778 & n9788 ) | ( ~n9777 & n9788 ) ;
  assign n10122 = ( n10110 & ~n10121 ) | ( n10110 & n10111 ) | ( ~n10121 & n10111 ) ;
  assign n10123 = ( n10110 & ~n10111 ) | ( n10110 & n10121 ) | ( ~n10111 & n10121 ) ;
  assign n10124 = ( n10122 & ~n10110 ) | ( n10122 & n10123 ) | ( ~n10110 & n10123 ) ;
  assign n10128 = x72 &  n7731 ;
  assign n10125 = ( x74 & ~n7538 ) | ( x74 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n10126 = x73 &  n7533 ;
  assign n10127 = n10125 | n10126 ;
  assign n10129 = ( x72 & ~n10128 ) | ( x72 & n10127 ) | ( ~n10128 & n10127 ) ;
  assign n10130 = ( n482 & ~n7541 ) | ( n482 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n10131 = n10129 | n10130 ;
  assign n10132 = ( x56 & ~n10131 ) | ( x56 & 1'b0 ) | ( ~n10131 & 1'b0 ) ;
  assign n10133 = ~x56 & n10131 ;
  assign n10134 = n10132 | n10133 ;
  assign n10135 = ( n10124 & ~n9804 ) | ( n10124 & n10134 ) | ( ~n9804 & n10134 ) ;
  assign n10136 = ( n9804 & ~n10134 ) | ( n9804 & n10124 ) | ( ~n10134 & n10124 ) ;
  assign n10137 = ( n10135 & ~n10124 ) | ( n10135 & n10136 ) | ( ~n10124 & n10136 ) ;
  assign n10138 = ( n9497 & ~n9805 ) | ( n9497 & n9815 ) | ( ~n9805 & n9815 ) ;
  assign n10139 = ( n10093 & n10137 ) | ( n10093 & n10138 ) | ( n10137 & n10138 ) ;
  assign n10140 = ( n10137 & ~n10093 ) | ( n10137 & n10138 ) | ( ~n10093 & n10138 ) ;
  assign n10141 = ( n10093 & ~n10139 ) | ( n10093 & n10140 ) | ( ~n10139 & n10140 ) ;
  assign n10152 = ( n9511 & ~n9818 ) | ( n9511 & n9828 ) | ( ~n9818 & n9828 ) ;
  assign n10145 = x78 &  n6288 ;
  assign n10142 = ( x80 & ~n6032 ) | ( x80 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n10143 = x79 &  n6027 ;
  assign n10144 = n10142 | n10143 ;
  assign n10146 = ( x78 & ~n10145 ) | ( x78 & n10144 ) | ( ~n10145 & n10144 ) ;
  assign n10147 = ( n842 & ~n6035 ) | ( n842 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n10148 = n10146 | n10147 ;
  assign n10149 = ( x50 & ~n10148 ) | ( x50 & 1'b0 ) | ( ~n10148 & 1'b0 ) ;
  assign n10150 = ~x50 & n10148 ;
  assign n10151 = n10149 | n10150 ;
  assign n10153 = ( n10141 & ~n10152 ) | ( n10141 & n10151 ) | ( ~n10152 & n10151 ) ;
  assign n10154 = ( n10141 & ~n10151 ) | ( n10141 & n10152 ) | ( ~n10151 & n10152 ) ;
  assign n10155 = ( n10153 & ~n10141 ) | ( n10153 & n10154 ) | ( ~n10141 & n10154 ) ;
  assign n10156 = ( n9514 & ~n9831 ) | ( n9514 & n9841 ) | ( ~n9831 & n9841 ) ;
  assign n10157 = ( n10083 & n10155 ) | ( n10083 & n10156 ) | ( n10155 & n10156 ) ;
  assign n10158 = ( n10155 & ~n10083 ) | ( n10155 & n10156 ) | ( ~n10083 & n10156 ) ;
  assign n10159 = ( n10083 & ~n10157 ) | ( n10083 & n10158 ) | ( ~n10157 & n10158 ) ;
  assign n10163 = x84 &  n4934 ;
  assign n10160 = ( x86 & ~n4725 ) | ( x86 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n10161 = x85 &  n4720 ;
  assign n10162 = n10160 | n10161 ;
  assign n10164 = ( x84 & ~n10163 ) | ( x84 & n10162 ) | ( ~n10163 & n10162 ) ;
  assign n10165 = ( n1496 & ~n4728 ) | ( n1496 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n10166 = n10164 | n10165 ;
  assign n10167 = ( x44 & ~n10166 ) | ( x44 & 1'b0 ) | ( ~n10166 & 1'b0 ) ;
  assign n10168 = ~x44 & n10166 ;
  assign n10169 = n10167 | n10168 ;
  assign n10170 = ( n10159 & ~n9846 ) | ( n10159 & n10169 ) | ( ~n9846 & n10169 ) ;
  assign n10171 = ( n9846 & ~n10169 ) | ( n9846 & n10159 ) | ( ~n10169 & n10159 ) ;
  assign n10172 = ( n10170 & ~n10159 ) | ( n10170 & n10171 ) | ( ~n10159 & n10171 ) ;
  assign n10173 = ( n9849 & n10073 ) | ( n9849 & n10172 ) | ( n10073 & n10172 ) ;
  assign n10174 = ( n9849 & ~n10073 ) | ( n9849 & n10172 ) | ( ~n10073 & n10172 ) ;
  assign n10175 = ( n10073 & ~n10173 ) | ( n10073 & n10174 ) | ( ~n10173 & n10174 ) ;
  assign n10176 = ( n9852 & n10063 ) | ( n9852 & n10175 ) | ( n10063 & n10175 ) ;
  assign n10177 = ( n9852 & ~n10063 ) | ( n9852 & n10175 ) | ( ~n10063 & n10175 ) ;
  assign n10178 = ( n10063 & ~n10176 ) | ( n10063 & n10177 ) | ( ~n10176 & n10177 ) ;
  assign n10179 = ( n9855 & n10053 ) | ( n9855 & n10178 ) | ( n10053 & n10178 ) ;
  assign n10180 = ( n9855 & ~n10053 ) | ( n9855 & n10178 ) | ( ~n10053 & n10178 ) ;
  assign n10181 = ( n10053 & ~n10179 ) | ( n10053 & n10180 ) | ( ~n10179 & n10180 ) ;
  assign n10185 = x96 &  n2718 ;
  assign n10182 = ( x98 & ~n2642 ) | ( x98 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n10183 = x97 &  n2637 ;
  assign n10184 = n10182 | n10183 ;
  assign n10186 = ( x96 & ~n10185 ) | ( x96 & n10184 ) | ( ~n10185 & n10184 ) ;
  assign n10187 = ~n2645 & n3170 ;
  assign n10188 = n10186 | n10187 ;
  assign n10189 = ( x32 & ~n10188 ) | ( x32 & 1'b0 ) | ( ~n10188 & 1'b0 ) ;
  assign n10190 = ~x32 & n10188 ;
  assign n10191 = n10189 | n10190 ;
  assign n10192 = ( n10181 & ~n9870 ) | ( n10181 & n10191 ) | ( ~n9870 & n10191 ) ;
  assign n10193 = ( n9870 & ~n10191 ) | ( n9870 & n10181 ) | ( ~n10191 & n10181 ) ;
  assign n10194 = ( n10192 & ~n10181 ) | ( n10192 & n10193 ) | ( ~n10181 & n10193 ) ;
  assign n10195 = ( n9871 & ~n9872 ) | ( n9871 & n9882 ) | ( ~n9872 & n9882 ) ;
  assign n10196 = ( n10043 & ~n10194 ) | ( n10043 & n10195 ) | ( ~n10194 & n10195 ) ;
  assign n10197 = ( n10043 & ~n10195 ) | ( n10043 & n10194 ) | ( ~n10195 & n10194 ) ;
  assign n10198 = ( n10196 & ~n10043 ) | ( n10196 & n10197 ) | ( ~n10043 & n10197 ) ;
  assign n10199 = ( n9568 & ~n9885 ) | ( n9568 & n9895 ) | ( ~n9885 & n9895 ) ;
  assign n10200 = ( n10033 & ~n10198 ) | ( n10033 & n10199 ) | ( ~n10198 & n10199 ) ;
  assign n10201 = ( n10033 & ~n10199 ) | ( n10033 & n10198 ) | ( ~n10199 & n10198 ) ;
  assign n10202 = ( n10200 & ~n10033 ) | ( n10200 & n10201 ) | ( ~n10033 & n10201 ) ;
  assign n10206 = x105 &  n1551 ;
  assign n10203 = ( x107 & ~n1451 ) | ( x107 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n10204 = x106 &  n1446 ;
  assign n10205 = n10203 | n10204 ;
  assign n10207 = ( x105 & ~n10206 ) | ( x105 & n10205 ) | ( ~n10206 & n10205 ) ;
  assign n10208 = ~n1454 & n4848 ;
  assign n10209 = n10207 | n10208 ;
  assign n10210 = ( x23 & ~n10209 ) | ( x23 & 1'b0 ) | ( ~n10209 & 1'b0 ) ;
  assign n10211 = ~x23 & n10209 ;
  assign n10212 = n10210 | n10211 ;
  assign n10213 = ( n10202 & ~n9900 ) | ( n10202 & n10212 ) | ( ~n9900 & n10212 ) ;
  assign n10214 = ( n9900 & ~n10212 ) | ( n9900 & n10202 ) | ( ~n10212 & n10202 ) ;
  assign n10215 = ( n10213 & ~n10202 ) | ( n10213 & n10214 ) | ( ~n10202 & n10214 ) ;
  assign n10216 = ( n9903 & n10023 ) | ( n9903 & n10215 ) | ( n10023 & n10215 ) ;
  assign n10217 = ( n9903 & ~n10023 ) | ( n9903 & n10215 ) | ( ~n10023 & n10215 ) ;
  assign n10218 = ( n10023 & ~n10216 ) | ( n10023 & n10217 ) | ( ~n10216 & n10217 ) ;
  assign n10220 = ( n9906 & n10013 ) | ( n9906 & n10218 ) | ( n10013 & n10218 ) ;
  assign n10219 = ( n9906 & ~n10013 ) | ( n9906 & n10218 ) | ( ~n10013 & n10218 ) ;
  assign n10221 = ( n10013 & ~n10220 ) | ( n10013 & n10219 ) | ( ~n10220 & n10219 ) ;
  assign n10222 = ( x14 & ~n10003 ) | ( x14 & n10221 ) | ( ~n10003 & n10221 ) ;
  assign n10223 = ( n10003 & ~x14 ) | ( n10003 & n10221 ) | ( ~x14 & n10221 ) ;
  assign n10224 = ( n10222 & ~n10221 ) | ( n10222 & n10223 ) | ( ~n10221 & n10223 ) ;
  assign n10235 = ( n9996 & n10224 ) | ( n9996 & n10234 ) | ( n10224 & n10234 ) ;
  assign n10236 = ( n9996 & ~n10234 ) | ( n9996 & n10224 ) | ( ~n10234 & n10224 ) ;
  assign n10237 = ( n10234 & ~n10235 ) | ( n10234 & n10236 ) | ( ~n10235 & n10236 ) ;
  assign n10238 = ( n9980 & ~n9992 ) | ( n9980 & n10237 ) | ( ~n9992 & n10237 ) ;
  assign n10239 = ( n9980 & ~n10237 ) | ( n9980 & n9992 ) | ( ~n10237 & n9992 ) ;
  assign n10240 = ( n10238 & ~n9980 ) | ( n10238 & n10239 ) | ( ~n9980 & n10239 ) ;
  assign n9973 = x123 &  n225 ;
  assign n9970 = ( x125 & ~n197 ) | ( x125 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n9971 = x124 &  n192 ;
  assign n9972 = n9970 | n9971 ;
  assign n9974 = ( x123 & ~n9973 ) | ( x123 & n9972 ) | ( ~n9973 & n9972 ) ;
  assign n9975 = ( n9318 & ~n200 ) | ( n9318 & n9321 ) | ( ~n200 & n9321 ) ;
  assign n9976 = ( n9974 & ~n9322 ) | ( n9974 & n9975 ) | ( ~n9322 & n9975 ) ;
  assign n9977 = ( x5 & ~n9976 ) | ( x5 & 1'b0 ) | ( ~n9976 & 1'b0 ) ;
  assign n9978 = ~x5 & n9976 ;
  assign n9979 = n9977 | n9978 ;
  assign n10241 = ( n9969 & ~n10240 ) | ( n9969 & n9979 ) | ( ~n10240 & n9979 ) ;
  assign n10242 = ( n9969 & ~n9979 ) | ( n9969 & n10240 ) | ( ~n9979 & n10240 ) ;
  assign n10243 = ( n10241 & ~n9969 ) | ( n10241 & n10242 ) | ( ~n9969 & n10242 ) ;
  assign n9954 = ( x126 & ~n150 ) | ( x126 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n9955 = ( x127 & ~n131 ) | ( x127 & 1'b0 ) | ( ~n131 & 1'b0 ) ;
  assign n9956 = n9954 | n9955 ;
  assign n9957 = ~n9348 & x127 ;
  assign n9958 = ~n9348 & x126 ;
  assign n9959 = ~x127 & x126 ;
  assign n9960 = ( n9957 & ~n9958 ) | ( n9957 & n9959 ) | ( ~n9958 & n9959 ) ;
  assign n9961 = ~n139 & n9960 ;
  assign n9962 = n9956 | n9961 ;
  assign n10244 = ( x2 & n9962 ) | ( x2 & n10243 ) | ( n9962 & n10243 ) ;
  assign n10245 = ( x2 & ~n10243 ) | ( x2 & n9962 ) | ( ~n10243 & n9962 ) ;
  assign n10246 = ( n10243 & ~n10244 ) | ( n10243 & n10245 ) | ( ~n10244 & n10245 ) ;
  assign n9953 = ( n9642 & n9648 ) | ( n9642 & n9946 ) | ( n9648 & n9946 ) ;
  assign n10247 = ( n9952 & ~n10246 ) | ( n9952 & n9953 ) | ( ~n10246 & n9953 ) ;
  assign n10248 = ( n9952 & ~n9953 ) | ( n9952 & n10246 ) | ( ~n9953 & n10246 ) ;
  assign n10249 = ( n10247 & ~n9952 ) | ( n10247 & n10248 ) | ( ~n9952 & n10248 ) ;
  assign n10250 = n10241 &  n10242 ;
  assign n10251 = x2 | n9962 ;
  assign n10252 = ( n10250 & ~n10244 ) | ( n10250 & n10251 ) | ( ~n10244 & n10251 ) ;
  assign n10532 = x124 &  n225 ;
  assign n10529 = ( x126 & ~n197 ) | ( x126 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n10530 = x125 &  n192 ;
  assign n10531 = n10529 | n10530 ;
  assign n10533 = ( x124 & ~n10532 ) | ( x124 & n10531 ) | ( ~n10532 & n10531 ) ;
  assign n10534 = n200 | n9349 ;
  assign n10535 = ~n10533 & n10534 ;
  assign n10513 = x121 &  n353 ;
  assign n10510 = ( x123 & ~n313 ) | ( x123 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n10511 = x122 &  n308 ;
  assign n10512 = n10510 | n10511 ;
  assign n10514 = ( x121 & ~n10513 ) | ( x121 & n10512 ) | ( ~n10513 & n10512 ) ;
  assign n10515 = ~n316 & n8472 ;
  assign n10516 = n10514 | n10515 ;
  assign n10517 = ( x8 & ~n10516 ) | ( x8 & 1'b0 ) | ( ~n10516 & 1'b0 ) ;
  assign n10518 = ~x8 & n10516 ;
  assign n10519 = n10517 | n10518 ;
  assign n10268 = x115 &  n713 ;
  assign n10265 = ( x117 & ~n641 ) | ( x117 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n10266 = x116 &  n636 ;
  assign n10267 = n10265 | n10266 ;
  assign n10269 = ( x115 & ~n10268 ) | ( x115 & n10267 ) | ( ~n10268 & n10267 ) ;
  assign n10270 = n644 | n7136 ;
  assign n10271 = ~n10269 & n10270 ;
  assign n10480 = x112 &  n942 ;
  assign n10477 = ( x114 & ~n896 ) | ( x114 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n10478 = x113 &  n891 ;
  assign n10479 = n10477 | n10478 ;
  assign n10481 = ( x112 & ~n10480 ) | ( x112 & n10479 ) | ( ~n10480 & n10479 ) ;
  assign n10482 = n899 | n6185 ;
  assign n10483 = ~n10481 & n10482 ;
  assign n10484 = x17 &  n10483 ;
  assign n10485 = x17 | n10483 ;
  assign n10486 = ~n10484 & n10485 ;
  assign n10285 = x106 &  n1551 ;
  assign n10282 = ( x108 & ~n1451 ) | ( x108 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n10283 = x107 &  n1446 ;
  assign n10284 = n10282 | n10283 ;
  assign n10286 = ( x106 & ~n10285 ) | ( x106 & n10284 ) | ( ~n10285 & n10284 ) ;
  assign n10287 = n1454 | n5055 ;
  assign n10288 = ~n10286 & n10287 ;
  assign n10289 = x23 &  n10288 ;
  assign n10290 = x23 | n10288 ;
  assign n10291 = ~n10289 & n10290 ;
  assign n10470 = ( n9900 & n10202 ) | ( n9900 & n10212 ) | ( n10202 & n10212 ) ;
  assign n10295 = x100 &  n2312 ;
  assign n10292 = ( x102 & ~n2195 ) | ( x102 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n10293 = x101 &  n2190 ;
  assign n10294 = n10292 | n10293 ;
  assign n10296 = ( x100 & ~n10295 ) | ( x100 & n10294 ) | ( ~n10295 & n10294 ) ;
  assign n10297 = n2198 | n3872 ;
  assign n10298 = ~n10296 & n10297 ;
  assign n10299 = x29 &  n10298 ;
  assign n10300 = x29 | n10298 ;
  assign n10301 = ~n10299 & n10300 ;
  assign n10305 = x97 &  n2718 ;
  assign n10302 = ( x99 & ~n2642 ) | ( x99 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n10303 = x98 &  n2637 ;
  assign n10304 = n10302 | n10303 ;
  assign n10306 = ( x97 & ~n10305 ) | ( x97 & n10304 ) | ( ~n10305 & n10304 ) ;
  assign n10307 = ~n2645 & n3338 ;
  assign n10308 = n10306 | n10307 ;
  assign n10309 = ( x32 & ~n10308 ) | ( x32 & 1'b0 ) | ( ~n10308 & 1'b0 ) ;
  assign n10310 = ~x32 & n10308 ;
  assign n10311 = n10309 | n10310 ;
  assign n10315 = x91 &  n3756 ;
  assign n10312 = ( x93 & ~n3602 ) | ( x93 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n10313 = x92 &  n3597 ;
  assign n10314 = n10312 | n10313 ;
  assign n10316 = ( x91 & ~n10315 ) | ( x91 & n10314 ) | ( ~n10315 & n10314 ) ;
  assign n10317 = n2264 | n3605 ;
  assign n10318 = ~n10316 & n10317 ;
  assign n10319 = x38 &  n10318 ;
  assign n10320 = x38 | n10318 ;
  assign n10321 = ~n10319 & n10320 ;
  assign n10325 = x88 &  n4344 ;
  assign n10322 = ( x90 & ~n4143 ) | ( x90 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n10323 = x89 &  n4138 ;
  assign n10324 = n10322 | n10323 ;
  assign n10326 = ( x88 & ~n10325 ) | ( x88 & n10324 ) | ( ~n10325 & n10324 ) ;
  assign n10327 = ( n1976 & ~n4146 ) | ( n1976 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n10328 = n10326 | n10327 ;
  assign n10329 = ( x41 & ~n10328 ) | ( x41 & 1'b0 ) | ( ~n10328 & 1'b0 ) ;
  assign n10330 = ~x41 & n10328 ;
  assign n10331 = n10329 | n10330 ;
  assign n10407 = x82 &  n5586 ;
  assign n10404 = ( x84 & ~n5389 ) | ( x84 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n10405 = x83 &  n5384 ;
  assign n10406 = n10404 | n10405 ;
  assign n10408 = ( x82 & ~n10407 ) | ( x82 & n10406 ) | ( ~n10407 & n10406 ) ;
  assign n10409 = ( n1199 & ~n5392 ) | ( n1199 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n10410 = n10408 | n10409 ;
  assign n10411 = ( x47 & ~n10410 ) | ( x47 & 1'b0 ) | ( ~n10410 & 1'b0 ) ;
  assign n10412 = ~x47 & n10410 ;
  assign n10413 = n10411 | n10412 ;
  assign n10380 = x76 &  n6982 ;
  assign n10377 = ( x78 & ~n6727 ) | ( x78 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n10378 = x77 &  n6722 ;
  assign n10379 = n10377 | n10378 ;
  assign n10381 = ( x76 & ~n10380 ) | ( x76 & n10379 ) | ( ~n10380 & n10379 ) ;
  assign n10382 = ( n693 & ~n6730 ) | ( n693 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n10383 = n10381 | n10382 ;
  assign n10384 = ( x53 & ~n10383 ) | ( x53 & 1'b0 ) | ( ~n10383 & 1'b0 ) ;
  assign n10385 = ~x53 & n10383 ;
  assign n10386 = n10384 | n10385 ;
  assign n10335 = x67 &  n9457 ;
  assign n10332 = ( x69 & ~n9150 ) | ( x69 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n10333 = x68 &  n9145 ;
  assign n10334 = n10332 | n10333 ;
  assign n10336 = ( x67 & ~n10335 ) | ( x67 & n10334 ) | ( ~n10335 & n10334 ) ;
  assign n10337 = ( n246 & ~n9153 ) | ( n246 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n10338 = n10336 | n10337 ;
  assign n10339 = ( x62 & ~n10338 ) | ( x62 & 1'b0 ) | ( ~n10338 & 1'b0 ) ;
  assign n10340 = ~x62 & n10338 ;
  assign n10341 = n10339 | n10340 ;
  assign n10342 = x65 &  n10104 ;
  assign n10343 = ( x66 & ~n9760 ) | ( x66 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n10344 = n10342 | n10343 ;
  assign n10345 = ( n9776 & n10103 ) | ( n9776 & n10107 ) | ( n10103 & n10107 ) ;
  assign n10346 = ( n10341 & ~n10344 ) | ( n10341 & n10345 ) | ( ~n10344 & n10345 ) ;
  assign n10347 = ( n10341 & ~n10345 ) | ( n10341 & n10344 ) | ( ~n10345 & n10344 ) ;
  assign n10348 = ( n10346 & ~n10341 ) | ( n10346 & n10347 ) | ( ~n10341 & n10347 ) ;
  assign n10353 = x70 &  n8558 ;
  assign n10350 = ( x72 & ~n8314 ) | ( x72 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n10351 = x71 &  n8309 ;
  assign n10352 = n10350 | n10351 ;
  assign n10354 = ( x70 & ~n10353 ) | ( x70 & n10352 ) | ( ~n10353 & n10352 ) ;
  assign n10355 = ( n345 & ~n8317 ) | ( n345 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n10356 = n10354 | n10355 ;
  assign n10357 = ( x59 & ~n10356 ) | ( x59 & 1'b0 ) | ( ~n10356 & 1'b0 ) ;
  assign n10358 = ~x59 & n10356 ;
  assign n10359 = n10357 | n10358 ;
  assign n10349 = ( n10110 & n10111 ) | ( n10110 & n10121 ) | ( n10111 & n10121 ) ;
  assign n10360 = ( n10348 & ~n10359 ) | ( n10348 & n10349 ) | ( ~n10359 & n10349 ) ;
  assign n10361 = ( n10348 & ~n10349 ) | ( n10348 & n10359 ) | ( ~n10349 & n10359 ) ;
  assign n10362 = ( n10360 & ~n10348 ) | ( n10360 & n10361 ) | ( ~n10348 & n10361 ) ;
  assign n10363 = ( n9804 & n10124 ) | ( n9804 & n10134 ) | ( n10124 & n10134 ) ;
  assign n10367 = x73 &  n7731 ;
  assign n10364 = ( x75 & ~n7538 ) | ( x75 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n10365 = x74 &  n7533 ;
  assign n10366 = n10364 | n10365 ;
  assign n10368 = ( x73 & ~n10367 ) | ( x73 & n10366 ) | ( ~n10367 & n10366 ) ;
  assign n10369 = ( n540 & ~n7541 ) | ( n540 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n10370 = n10368 | n10369 ;
  assign n10371 = ( x56 & ~n10370 ) | ( x56 & 1'b0 ) | ( ~n10370 & 1'b0 ) ;
  assign n10372 = ~x56 & n10370 ;
  assign n10373 = n10371 | n10372 ;
  assign n10374 = ( n10362 & ~n10363 ) | ( n10362 & n10373 ) | ( ~n10363 & n10373 ) ;
  assign n10375 = ( n10362 & ~n10373 ) | ( n10362 & n10363 ) | ( ~n10373 & n10363 ) ;
  assign n10376 = ( n10374 & ~n10362 ) | ( n10374 & n10375 ) | ( ~n10362 & n10375 ) ;
  assign n10388 = ( n10139 & n10376 ) | ( n10139 & n10386 ) | ( n10376 & n10386 ) ;
  assign n10387 = ( n10139 & ~n10386 ) | ( n10139 & n10376 ) | ( ~n10386 & n10376 ) ;
  assign n10389 = ( n10386 & ~n10388 ) | ( n10386 & n10387 ) | ( ~n10388 & n10387 ) ;
  assign n10390 = ( n10141 & n10151 ) | ( n10141 & n10152 ) | ( n10151 & n10152 ) ;
  assign n10394 = x79 &  n6288 ;
  assign n10391 = ( x81 & ~n6032 ) | ( x81 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n10392 = x80 &  n6027 ;
  assign n10393 = n10391 | n10392 ;
  assign n10395 = ( x79 & ~n10394 ) | ( x79 & n10393 ) | ( ~n10394 & n10393 ) ;
  assign n10396 = ( n994 & ~n6035 ) | ( n994 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n10397 = n10395 | n10396 ;
  assign n10398 = ( x50 & ~n10397 ) | ( x50 & 1'b0 ) | ( ~n10397 & 1'b0 ) ;
  assign n10399 = ~x50 & n10397 ;
  assign n10400 = n10398 | n10399 ;
  assign n10401 = ( n10389 & ~n10390 ) | ( n10389 & n10400 ) | ( ~n10390 & n10400 ) ;
  assign n10402 = ( n10389 & ~n10400 ) | ( n10389 & n10390 ) | ( ~n10400 & n10390 ) ;
  assign n10403 = ( n10401 & ~n10389 ) | ( n10401 & n10402 ) | ( ~n10389 & n10402 ) ;
  assign n10414 = ( n10157 & ~n10413 ) | ( n10157 & n10403 ) | ( ~n10413 & n10403 ) ;
  assign n10415 = ( n10403 & ~n10157 ) | ( n10403 & n10413 ) | ( ~n10157 & n10413 ) ;
  assign n10416 = ( n10414 & ~n10403 ) | ( n10414 & n10415 ) | ( ~n10403 & n10415 ) ;
  assign n10417 = ( n9846 & n10159 ) | ( n9846 & n10169 ) | ( n10159 & n10169 ) ;
  assign n10421 = x85 &  n4934 ;
  assign n10418 = ( x87 & ~n4725 ) | ( x87 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n10419 = x86 &  n4720 ;
  assign n10420 = n10418 | n10419 ;
  assign n10422 = ( x85 & ~n10421 ) | ( x85 & n10420 ) | ( ~n10421 & n10420 ) ;
  assign n10423 = ( n1512 & ~n4728 ) | ( n1512 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n10424 = n10422 | n10423 ;
  assign n10425 = ( x44 & ~n10424 ) | ( x44 & 1'b0 ) | ( ~n10424 & 1'b0 ) ;
  assign n10426 = ~x44 & n10424 ;
  assign n10427 = n10425 | n10426 ;
  assign n10428 = ( n10416 & ~n10417 ) | ( n10416 & n10427 ) | ( ~n10417 & n10427 ) ;
  assign n10429 = ( n10416 & ~n10427 ) | ( n10416 & n10417 ) | ( ~n10427 & n10417 ) ;
  assign n10430 = ( n10428 & ~n10416 ) | ( n10428 & n10429 ) | ( ~n10416 & n10429 ) ;
  assign n10431 = ( n10173 & n10331 ) | ( n10173 & n10430 ) | ( n10331 & n10430 ) ;
  assign n10432 = ( n10173 & ~n10331 ) | ( n10173 & n10430 ) | ( ~n10331 & n10430 ) ;
  assign n10433 = ( n10331 & ~n10431 ) | ( n10331 & n10432 ) | ( ~n10431 & n10432 ) ;
  assign n10435 = ( n10176 & n10321 ) | ( n10176 & n10433 ) | ( n10321 & n10433 ) ;
  assign n10434 = ( n10176 & ~n10321 ) | ( n10176 & n10433 ) | ( ~n10321 & n10433 ) ;
  assign n10436 = ( n10321 & ~n10435 ) | ( n10321 & n10434 ) | ( ~n10435 & n10434 ) ;
  assign n10440 = x94 &  n3214 ;
  assign n10437 = ( x96 & ~n3087 ) | ( x96 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n10438 = x95 &  n3082 ;
  assign n10439 = n10437 | n10438 ;
  assign n10441 = ( x94 & ~n10440 ) | ( x94 & n10439 ) | ( ~n10440 & n10439 ) ;
  assign n10442 = ( n2836 & ~n3090 ) | ( n2836 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n10443 = n10441 | n10442 ;
  assign n10444 = ( x35 & ~n10443 ) | ( x35 & 1'b0 ) | ( ~n10443 & 1'b0 ) ;
  assign n10445 = ~x35 & n10443 ;
  assign n10446 = n10444 | n10445 ;
  assign n10447 = ( n10436 & ~n10179 ) | ( n10436 & n10446 ) | ( ~n10179 & n10446 ) ;
  assign n10448 = ( n10179 & ~n10446 ) | ( n10179 & n10436 ) | ( ~n10446 & n10436 ) ;
  assign n10449 = ( n10447 & ~n10436 ) | ( n10447 & n10448 ) | ( ~n10436 & n10448 ) ;
  assign n10450 = ( n9870 & n10181 ) | ( n9870 & n10191 ) | ( n10181 & n10191 ) ;
  assign n10451 = ( n10311 & n10449 ) | ( n10311 & n10450 ) | ( n10449 & n10450 ) ;
  assign n10452 = ( n10449 & ~n10311 ) | ( n10449 & n10450 ) | ( ~n10311 & n10450 ) ;
  assign n10453 = ( n10311 & ~n10451 ) | ( n10311 & n10452 ) | ( ~n10451 & n10452 ) ;
  assign n10454 = ( n10196 & n10301 ) | ( n10196 & n10453 ) | ( n10301 & n10453 ) ;
  assign n10455 = ( n10196 & ~n10301 ) | ( n10196 & n10453 ) | ( ~n10301 & n10453 ) ;
  assign n10456 = ( n10301 & ~n10454 ) | ( n10301 & n10455 ) | ( ~n10454 & n10455 ) ;
  assign n10460 = x103 &  n1894 ;
  assign n10457 = ( x105 & ~n1816 ) | ( x105 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n10458 = x104 &  n1811 ;
  assign n10459 = n10457 | n10458 ;
  assign n10461 = ( x103 & ~n10460 ) | ( x103 & n10459 ) | ( ~n10460 & n10459 ) ;
  assign n10462 = ~n1819 & n4442 ;
  assign n10463 = n10461 | n10462 ;
  assign n10464 = ( x26 & ~n10463 ) | ( x26 & 1'b0 ) | ( ~n10463 & 1'b0 ) ;
  assign n10465 = ~x26 & n10463 ;
  assign n10466 = n10464 | n10465 ;
  assign n10467 = ( n10200 & n10456 ) | ( n10200 & n10466 ) | ( n10456 & n10466 ) ;
  assign n10468 = ( n10200 & ~n10456 ) | ( n10200 & n10466 ) | ( ~n10456 & n10466 ) ;
  assign n10469 = ( n10456 & ~n10467 ) | ( n10456 & n10468 ) | ( ~n10467 & n10468 ) ;
  assign n10471 = ( n10291 & ~n10470 ) | ( n10291 & n10469 ) | ( ~n10470 & n10469 ) ;
  assign n10472 = ( n10291 & ~n10469 ) | ( n10291 & n10470 ) | ( ~n10469 & n10470 ) ;
  assign n10473 = ( n10471 & ~n10291 ) | ( n10471 & n10472 ) | ( ~n10291 & n10472 ) ;
  assign n10275 = x109 &  n1227 ;
  assign n10272 = ( x111 & ~n1154 ) | ( x111 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n10273 = x110 &  n1149 ;
  assign n10274 = n10272 | n10273 ;
  assign n10276 = ( x109 & ~n10275 ) | ( x109 & n10274 ) | ( ~n10275 & n10274 ) ;
  assign n10277 = n1157 | n5711 ;
  assign n10278 = ~n10276 & n10277 ;
  assign n10279 = x20 &  n10278 ;
  assign n10280 = x20 | n10278 ;
  assign n10281 = ~n10279 & n10280 ;
  assign n10474 = ( n10217 & ~n10473 ) | ( n10217 & n10281 ) | ( ~n10473 & n10281 ) ;
  assign n10475 = ( n10281 & ~n10217 ) | ( n10281 & n10473 ) | ( ~n10217 & n10473 ) ;
  assign n10476 = ( n10474 & ~n10281 ) | ( n10474 & n10475 ) | ( ~n10281 & n10475 ) ;
  assign n10487 = ( n10220 & ~n10486 ) | ( n10220 & n10476 ) | ( ~n10486 & n10476 ) ;
  assign n10488 = ( n10476 & ~n10220 ) | ( n10476 & n10486 ) | ( ~n10220 & n10486 ) ;
  assign n10489 = ( n10487 & ~n10476 ) | ( n10487 & n10488 ) | ( ~n10476 & n10488 ) ;
  assign n10490 = ( n10271 & ~x14 ) | ( n10271 & n10489 ) | ( ~x14 & n10489 ) ;
  assign n10491 = ( x14 & ~n10271 ) | ( x14 & n10489 ) | ( ~n10271 & n10489 ) ;
  assign n10492 = ( n10490 & ~n10489 ) | ( n10490 & n10491 ) | ( ~n10489 & n10491 ) ;
  assign n10496 = x118 &  n503 ;
  assign n10493 = ( x120 & ~n450 ) | ( x120 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n10494 = x119 &  n445 ;
  assign n10495 = n10493 | n10494 ;
  assign n10497 = ( x118 & ~n10496 ) | ( x118 & n10495 ) | ( ~n10496 & n10495 ) ;
  assign n10498 = ~n453 & n9364 ;
  assign n10499 = n10497 | n10498 ;
  assign n10500 = ( x11 & ~n10499 ) | ( x11 & 1'b0 ) | ( ~n10499 & 1'b0 ) ;
  assign n10501 = ~x11 & n10499 ;
  assign n10502 = n10500 | n10501 ;
  assign n10503 = x14 &  n10003 ;
  assign n10504 = x14 | n10003 ;
  assign n10505 = ~n10503 & n10504 ;
  assign n10506 = ( n10221 & ~n9996 ) | ( n10221 & n10505 ) | ( ~n9996 & n10505 ) ;
  assign n10507 = ( n10492 & ~n10502 ) | ( n10492 & n10506 ) | ( ~n10502 & n10506 ) ;
  assign n10508 = ( n10492 & ~n10506 ) | ( n10492 & n10502 ) | ( ~n10506 & n10502 ) ;
  assign n10509 = ( n10507 & ~n10492 ) | ( n10507 & n10508 ) | ( ~n10492 & n10508 ) ;
  assign n10520 = x11 &  n10231 ;
  assign n10521 = ( x11 & ~n10520 ) | ( x11 & n10232 ) | ( ~n10520 & n10232 ) ;
  assign n10522 = ~n9996 & n10224 ;
  assign n10523 = ( n9996 & ~n10224 ) | ( n9996 & 1'b0 ) | ( ~n10224 & 1'b0 ) ;
  assign n10524 = n10522 | n10523 ;
  assign n10525 = ( n10521 & ~n9980 ) | ( n10521 & n10524 ) | ( ~n9980 & n10524 ) ;
  assign n10526 = ( n10519 & ~n10509 ) | ( n10519 & n10525 ) | ( ~n10509 & n10525 ) ;
  assign n10527 = ( n10509 & ~n10519 ) | ( n10509 & n10525 ) | ( ~n10519 & n10525 ) ;
  assign n10528 = ( n10526 & ~n10525 ) | ( n10526 & n10527 ) | ( ~n10525 & n10527 ) ;
  assign n10536 = ( x5 & ~n10535 ) | ( x5 & n10528 ) | ( ~n10535 & n10528 ) ;
  assign n10537 = ( x5 & ~n10528 ) | ( x5 & n10535 ) | ( ~n10528 & n10535 ) ;
  assign n10538 = ( n10536 & ~x5 ) | ( n10536 & n10537 ) | ( ~x5 & n10537 ) ;
  assign n10253 = n9980 | n10237 ;
  assign n10254 = ( n9980 & ~n10237 ) | ( n9980 & 1'b0 ) | ( ~n10237 & 1'b0 ) ;
  assign n10255 = ( n10253 & ~n9980 ) | ( n10253 & n10254 ) | ( ~n9980 & n10254 ) ;
  assign n10256 = ( n9979 & ~n10255 ) | ( n9979 & n9992 ) | ( ~n10255 & n9992 ) ;
  assign n10257 = ~x126 & n9348 ;
  assign n10258 = ( ~x126 & ~x127 ) | ( ~x126 & ~n10257 ) | ( ~x127 & ~n10257 ) ;
  assign n10260 = n139 | n10258 ;
  assign n10261 = ~x2 & n10260 ;
  assign n10259 = ( x127 & ~n150 ) | ( x127 & 1'b0 ) | ( ~n150 & 1'b0 ) ;
  assign n10262 = ~n10259 & n10260 ;
  assign n10263 = x2 | n10260 ;
  assign n10264 = ( n10261 & ~n10262 ) | ( n10261 & n10263 ) | ( ~n10262 & n10263 ) ;
  assign n10540 = ( n10256 & n10264 ) | ( n10256 & n10538 ) | ( n10264 & n10538 ) ;
  assign n10539 = ( n10256 & ~n10538 ) | ( n10256 & n10264 ) | ( ~n10538 & n10264 ) ;
  assign n10541 = ( n10538 & ~n10540 ) | ( n10538 & n10539 ) | ( ~n10540 & n10539 ) ;
  assign n10543 = ( n10248 & n10252 ) | ( n10248 & n10541 ) | ( n10252 & n10541 ) ;
  assign n10542 = ( n10248 & ~n10252 ) | ( n10248 & n10541 ) | ( ~n10252 & n10541 ) ;
  assign n10544 = ( n10252 & ~n10543 ) | ( n10252 & n10542 ) | ( ~n10543 & n10542 ) ;
  assign n10545 = ( n10264 & ~n10256 ) | ( n10264 & n10538 ) | ( ~n10256 & n10538 ) ;
  assign n10549 = x5 &  n10535 ;
  assign n10550 = x5 | n10535 ;
  assign n10551 = ~n10549 & n10550 ;
  assign n10546 = ( x8 & n10509 ) | ( x8 & n10516 ) | ( n10509 & n10516 ) ;
  assign n10547 = ( n10509 & ~x8 ) | ( n10509 & n10516 ) | ( ~x8 & n10516 ) ;
  assign n10548 = ( x8 & ~n10546 ) | ( x8 & n10547 ) | ( ~n10546 & n10547 ) ;
  assign n10552 = ( n10525 & ~n10551 ) | ( n10525 & n10548 ) | ( ~n10551 & n10548 ) ;
  assign n10556 = x125 &  n225 ;
  assign n10553 = ( x127 & ~n197 ) | ( x127 & 1'b0 ) | ( ~n197 & 1'b0 ) ;
  assign n10554 = x126 &  n192 ;
  assign n10555 = n10553 | n10554 ;
  assign n10557 = ( x125 & ~n10556 ) | ( x125 & n10555 ) | ( ~n10556 & n10555 ) ;
  assign n10558 = n200 | n9941 ;
  assign n10559 = ~n10557 & n10558 ;
  assign n10560 = x5 &  n10559 ;
  assign n10561 = x5 | n10559 ;
  assign n10562 = ~n10560 & n10561 ;
  assign n10563 = n10492 &  n10506 ;
  assign n10564 = n10492 | n10506 ;
  assign n10565 = ~n10563 & n10564 ;
  assign n10566 = ( n10502 & n10519 ) | ( n10502 & n10565 ) | ( n10519 & n10565 ) ;
  assign n10567 = ( n644 & ~n7136 ) | ( n644 & n10269 ) | ( ~n7136 & n10269 ) ;
  assign n10568 = n7136 | n10567 ;
  assign n10570 = ( x14 & n10269 ) | ( x14 & n10568 ) | ( n10269 & n10568 ) ;
  assign n10569 = ( x14 & ~n10568 ) | ( x14 & n10269 ) | ( ~n10568 & n10269 ) ;
  assign n10571 = ( n10568 & ~n10570 ) | ( n10568 & n10569 ) | ( ~n10570 & n10569 ) ;
  assign n10572 = ( n10506 & ~n10489 ) | ( n10506 & n10571 ) | ( ~n10489 & n10571 ) ;
  assign n10576 = x119 &  n503 ;
  assign n10573 = ( x121 & ~n450 ) | ( x121 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n10574 = x120 &  n445 ;
  assign n10575 = n10573 | n10574 ;
  assign n10577 = ( x119 & ~n10576 ) | ( x119 & n10575 ) | ( ~n10576 & n10575 ) ;
  assign n10578 = ~n453 & n8176 ;
  assign n10579 = n10577 | n10578 ;
  assign n10580 = ( x11 & ~n10579 ) | ( x11 & 1'b0 ) | ( ~n10579 & 1'b0 ) ;
  assign n10581 = ~x11 & n10579 ;
  assign n10582 = n10580 | n10581 ;
  assign n10583 = ( n10220 & ~n10476 ) | ( n10220 & n10486 ) | ( ~n10476 & n10486 ) ;
  assign n10587 = x113 &  n942 ;
  assign n10584 = ( x115 & ~n896 ) | ( x115 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n10585 = x114 &  n891 ;
  assign n10586 = n10584 | n10585 ;
  assign n10588 = ( x113 & ~n10587 ) | ( x113 & n10586 ) | ( ~n10587 & n10586 ) ;
  assign n10589 = ~n899 & n6420 ;
  assign n10590 = n10588 | n10589 ;
  assign n10591 = ( x17 & ~n10590 ) | ( x17 & 1'b0 ) | ( ~n10590 & 1'b0 ) ;
  assign n10592 = ~x17 & n10590 ;
  assign n10593 = n10591 | n10592 ;
  assign n10597 = x110 &  n1227 ;
  assign n10594 = ( x112 & ~n1154 ) | ( x112 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n10595 = x111 &  n1149 ;
  assign n10596 = n10594 | n10595 ;
  assign n10598 = ( x110 & ~n10597 ) | ( x110 & n10596 ) | ( ~n10597 & n10596 ) ;
  assign n10599 = ~n1157 & n5727 ;
  assign n10600 = n10598 | n10599 ;
  assign n10796 = x20 | n10600 ;
  assign n10797 = ~x20 & n10600 ;
  assign n10798 = ( n10796 & ~n10600 ) | ( n10796 & n10797 ) | ( ~n10600 & n10797 ) ;
  assign n10601 = ( n10469 & ~n10291 ) | ( n10469 & n10470 ) | ( ~n10291 & n10470 ) ;
  assign n10602 = ( n10200 & ~n10466 ) | ( n10200 & n10456 ) | ( ~n10466 & n10456 ) ;
  assign n10606 = x104 &  n1894 ;
  assign n10603 = ( x106 & ~n1816 ) | ( x106 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n10604 = x105 &  n1811 ;
  assign n10605 = n10603 | n10604 ;
  assign n10607 = ( x104 & ~n10606 ) | ( x104 & n10605 ) | ( ~n10606 & n10605 ) ;
  assign n10608 = ~n1819 & n4458 ;
  assign n10609 = n10607 | n10608 ;
  assign n10777 = x26 | n10609 ;
  assign n10778 = ~x26 & n10609 ;
  assign n10779 = ( n10777 & ~n10609 ) | ( n10777 & n10778 ) | ( ~n10609 & n10778 ) ;
  assign n10613 = x101 &  n2312 ;
  assign n10610 = ( x103 & ~n2195 ) | ( x103 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n10611 = x102 &  n2190 ;
  assign n10612 = n10610 | n10611 ;
  assign n10614 = ( x101 & ~n10613 ) | ( x101 & n10612 ) | ( ~n10613 & n10612 ) ;
  assign n10615 = ( n2198 & ~n4056 ) | ( n2198 & n10614 ) | ( ~n4056 & n10614 ) ;
  assign n10616 = n4056 | n10615 ;
  assign n10618 = ( x29 & n10614 ) | ( x29 & n10616 ) | ( n10614 & n10616 ) ;
  assign n10617 = ( x29 & ~n10616 ) | ( x29 & n10614 ) | ( ~n10616 & n10614 ) ;
  assign n10619 = ( n10616 & ~n10618 ) | ( n10616 & n10617 ) | ( ~n10618 & n10617 ) ;
  assign n10620 = ( n10311 & ~n10449 ) | ( n10311 & n10450 ) | ( ~n10449 & n10450 ) ;
  assign n10621 = ( n10416 & n10417 ) | ( n10416 & n10427 ) | ( n10417 & n10427 ) ;
  assign n10622 = ( n10389 & n10390 ) | ( n10389 & n10400 ) | ( n10390 & n10400 ) ;
  assign n10623 = ( n10362 & n10363 ) | ( n10362 & n10373 ) | ( n10363 & n10373 ) ;
  assign n10627 = x77 &  n6982 ;
  assign n10624 = ( x79 & ~n6727 ) | ( x79 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n10625 = x78 &  n6722 ;
  assign n10626 = n10624 | n10625 ;
  assign n10628 = ( x77 & ~n10627 ) | ( x77 & n10626 ) | ( ~n10627 & n10626 ) ;
  assign n10629 = ( n766 & ~n6730 ) | ( n766 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n10630 = n10628 | n10629 ;
  assign n10631 = ( x53 & ~n10630 ) | ( x53 & 1'b0 ) | ( ~n10630 & 1'b0 ) ;
  assign n10632 = ~x53 & n10630 ;
  assign n10633 = n10631 | n10632 ;
  assign n10634 = x66 &  n10104 ;
  assign n10635 = ( x67 & ~n9760 ) | ( x67 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n10636 = n10634 | n10635 ;
  assign n10640 = x68 &  n9457 ;
  assign n10637 = ( x70 & ~n9150 ) | ( x70 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n10638 = x69 &  n9145 ;
  assign n10639 = n10637 | n10638 ;
  assign n10641 = ( x68 & ~n10640 ) | ( x68 & n10639 ) | ( ~n10640 & n10639 ) ;
  assign n10642 = ( n282 & ~n10641 ) | ( n282 & n9153 ) | ( ~n10641 & n9153 ) ;
  assign n10643 = ~n9153 & n10642 ;
  assign n10644 = ( x62 & n10641 ) | ( x62 & n10643 ) | ( n10641 & n10643 ) ;
  assign n10645 = ( x62 & ~n10643 ) | ( x62 & n10641 ) | ( ~n10643 & n10641 ) ;
  assign n10646 = ( n10643 & ~n10644 ) | ( n10643 & n10645 ) | ( ~n10644 & n10645 ) ;
  assign n10647 = ( x2 & n10636 ) | ( x2 & n10646 ) | ( n10636 & n10646 ) ;
  assign n10648 = ( x2 & ~n10636 ) | ( x2 & n10646 ) | ( ~n10636 & n10646 ) ;
  assign n10649 = ( n10636 & ~n10647 ) | ( n10636 & n10648 ) | ( ~n10647 & n10648 ) ;
  assign n10654 = x71 &  n8558 ;
  assign n10651 = ( x73 & ~n8314 ) | ( x73 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n10652 = x72 &  n8309 ;
  assign n10653 = n10651 | n10652 ;
  assign n10655 = ( x71 & ~n10654 ) | ( x71 & n10653 ) | ( ~n10654 & n10653 ) ;
  assign n10656 = ( n389 & ~n8317 ) | ( n389 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n10657 = n10655 | n10656 ;
  assign n10658 = ( x59 & ~n10657 ) | ( x59 & 1'b0 ) | ( ~n10657 & 1'b0 ) ;
  assign n10659 = ~x59 & n10657 ;
  assign n10660 = n10658 | n10659 ;
  assign n10650 = ( n10341 & n10344 ) | ( n10341 & n10345 ) | ( n10344 & n10345 ) ;
  assign n10661 = ( n10649 & ~n10660 ) | ( n10649 & n10650 ) | ( ~n10660 & n10650 ) ;
  assign n10662 = ( n10649 & ~n10650 ) | ( n10649 & n10660 ) | ( ~n10650 & n10660 ) ;
  assign n10663 = ( n10661 & ~n10649 ) | ( n10661 & n10662 ) | ( ~n10649 & n10662 ) ;
  assign n10664 = ( n10348 & n10349 ) | ( n10348 & n10359 ) | ( n10349 & n10359 ) ;
  assign n10668 = x74 &  n7731 ;
  assign n10665 = ( x76 & ~n7538 ) | ( x76 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n10666 = x75 &  n7533 ;
  assign n10667 = n10665 | n10666 ;
  assign n10669 = ( x74 & ~n10668 ) | ( x74 & n10667 ) | ( ~n10668 & n10667 ) ;
  assign n10670 = ( n603 & ~n7541 ) | ( n603 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n10671 = n10669 | n10670 ;
  assign n10672 = ( x56 & ~n10671 ) | ( x56 & 1'b0 ) | ( ~n10671 & 1'b0 ) ;
  assign n10673 = ~x56 & n10671 ;
  assign n10674 = n10672 | n10673 ;
  assign n10675 = ( n10663 & ~n10664 ) | ( n10663 & n10674 ) | ( ~n10664 & n10674 ) ;
  assign n10676 = ( n10663 & ~n10674 ) | ( n10663 & n10664 ) | ( ~n10674 & n10664 ) ;
  assign n10677 = ( n10675 & ~n10663 ) | ( n10675 & n10676 ) | ( ~n10663 & n10676 ) ;
  assign n10679 = ( n10623 & n10633 ) | ( n10623 & n10677 ) | ( n10633 & n10677 ) ;
  assign n10678 = ( n10633 & ~n10623 ) | ( n10633 & n10677 ) | ( ~n10623 & n10677 ) ;
  assign n10680 = ( n10623 & ~n10679 ) | ( n10623 & n10678 ) | ( ~n10679 & n10678 ) ;
  assign n10684 = x80 &  n6288 ;
  assign n10681 = ( x82 & ~n6032 ) | ( x82 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n10682 = x81 &  n6027 ;
  assign n10683 = n10681 | n10682 ;
  assign n10685 = ( x80 & ~n10684 ) | ( x80 & n10683 ) | ( ~n10684 & n10683 ) ;
  assign n10686 = ( n1084 & ~n6035 ) | ( n1084 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n10687 = n10685 | n10686 ;
  assign n10688 = ( x50 & ~n10687 ) | ( x50 & 1'b0 ) | ( ~n10687 & 1'b0 ) ;
  assign n10689 = ~x50 & n10687 ;
  assign n10690 = n10688 | n10689 ;
  assign n10691 = ( n10388 & ~n10680 ) | ( n10388 & n10690 ) | ( ~n10680 & n10690 ) ;
  assign n10692 = ( n10388 & ~n10690 ) | ( n10388 & n10680 ) | ( ~n10690 & n10680 ) ;
  assign n10693 = ( n10691 & ~n10388 ) | ( n10691 & n10692 ) | ( ~n10388 & n10692 ) ;
  assign n10697 = x83 &  n5586 ;
  assign n10694 = ( x85 & ~n5389 ) | ( x85 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n10695 = x84 &  n5384 ;
  assign n10696 = n10694 | n10695 ;
  assign n10698 = ( x83 & ~n10697 ) | ( x83 & n10696 ) | ( ~n10697 & n10696 ) ;
  assign n10699 = ( n1295 & ~n5392 ) | ( n1295 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n10700 = n10698 | n10699 ;
  assign n10701 = ( x47 & ~n10700 ) | ( x47 & 1'b0 ) | ( ~n10700 & 1'b0 ) ;
  assign n10702 = ~x47 & n10700 ;
  assign n10703 = n10701 | n10702 ;
  assign n10704 = ( n10622 & ~n10693 ) | ( n10622 & n10703 ) | ( ~n10693 & n10703 ) ;
  assign n10705 = ( n10622 & ~n10703 ) | ( n10622 & n10693 ) | ( ~n10703 & n10693 ) ;
  assign n10706 = ( n10704 & ~n10622 ) | ( n10704 & n10705 ) | ( ~n10622 & n10705 ) ;
  assign n10717 = ( n10157 & n10403 ) | ( n10157 & n10413 ) | ( n10403 & n10413 ) ;
  assign n10710 = x86 &  n4934 ;
  assign n10707 = ( x88 & ~n4725 ) | ( x88 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n10708 = x87 &  n4720 ;
  assign n10709 = n10707 | n10708 ;
  assign n10711 = ( x86 & ~n10710 ) | ( x86 & n10709 ) | ( ~n10710 & n10709 ) ;
  assign n10712 = ( n1624 & ~n4728 ) | ( n1624 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n10713 = n10711 | n10712 ;
  assign n10714 = ( x44 & ~n10713 ) | ( x44 & 1'b0 ) | ( ~n10713 & 1'b0 ) ;
  assign n10715 = ~x44 & n10713 ;
  assign n10716 = n10714 | n10715 ;
  assign n10718 = ( n10706 & ~n10717 ) | ( n10706 & n10716 ) | ( ~n10717 & n10716 ) ;
  assign n10719 = ( n10706 & ~n10716 ) | ( n10706 & n10717 ) | ( ~n10716 & n10717 ) ;
  assign n10720 = ( n10718 & ~n10706 ) | ( n10718 & n10719 ) | ( ~n10706 & n10719 ) ;
  assign n10724 = x89 &  n4344 ;
  assign n10721 = ( x91 & ~n4143 ) | ( x91 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n10722 = x90 &  n4138 ;
  assign n10723 = n10721 | n10722 ;
  assign n10725 = ( x89 & ~n10724 ) | ( x89 & n10723 ) | ( ~n10724 & n10723 ) ;
  assign n10726 = ( n2108 & ~n4146 ) | ( n2108 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n10727 = n10725 | n10726 ;
  assign n10728 = ( x41 & ~n10727 ) | ( x41 & 1'b0 ) | ( ~n10727 & 1'b0 ) ;
  assign n10729 = ~x41 & n10727 ;
  assign n10730 = n10728 | n10729 ;
  assign n10731 = ( n10621 & ~n10720 ) | ( n10621 & n10730 ) | ( ~n10720 & n10730 ) ;
  assign n10732 = ( n10621 & ~n10730 ) | ( n10621 & n10720 ) | ( ~n10730 & n10720 ) ;
  assign n10733 = ( n10731 & ~n10621 ) | ( n10731 & n10732 ) | ( ~n10621 & n10732 ) ;
  assign n10737 = x92 &  n3756 ;
  assign n10734 = ( x94 & ~n3602 ) | ( x94 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n10735 = x93 &  n3597 ;
  assign n10736 = n10734 | n10735 ;
  assign n10738 = ( x92 & ~n10737 ) | ( x92 & n10736 ) | ( ~n10737 & n10736 ) ;
  assign n10739 = ( n2401 & ~n3605 ) | ( n2401 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n10740 = n10738 | n10739 ;
  assign n10741 = ( x38 & ~n10740 ) | ( x38 & 1'b0 ) | ( ~n10740 & 1'b0 ) ;
  assign n10742 = ~x38 & n10740 ;
  assign n10743 = n10741 | n10742 ;
  assign n10744 = ( n10431 & ~n10733 ) | ( n10431 & n10743 ) | ( ~n10733 & n10743 ) ;
  assign n10745 = ( n10431 & ~n10743 ) | ( n10431 & n10733 ) | ( ~n10743 & n10733 ) ;
  assign n10746 = ( n10744 & ~n10431 ) | ( n10744 & n10745 ) | ( ~n10431 & n10745 ) ;
  assign n10750 = x95 &  n3214 ;
  assign n10747 = ( x97 & ~n3087 ) | ( x97 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n10748 = x96 &  n3082 ;
  assign n10749 = n10747 | n10748 ;
  assign n10751 = ( x95 & ~n10750 ) | ( x95 & n10749 ) | ( ~n10750 & n10749 ) ;
  assign n10752 = ( n2999 & ~n3090 ) | ( n2999 & 1'b0 ) | ( ~n3090 & 1'b0 ) ;
  assign n10753 = n10751 | n10752 ;
  assign n10754 = ( x35 & ~n10753 ) | ( x35 & 1'b0 ) | ( ~n10753 & 1'b0 ) ;
  assign n10755 = ~x35 & n10753 ;
  assign n10756 = n10754 | n10755 ;
  assign n10757 = ( n10746 & ~n10434 ) | ( n10746 & n10756 ) | ( ~n10434 & n10756 ) ;
  assign n10758 = ( n10434 & ~n10756 ) | ( n10434 & n10746 ) | ( ~n10756 & n10746 ) ;
  assign n10759 = ( n10757 & ~n10746 ) | ( n10757 & n10758 ) | ( ~n10746 & n10758 ) ;
  assign n10760 = ( n10179 & ~n10436 ) | ( n10179 & n10446 ) | ( ~n10436 & n10446 ) ;
  assign n10764 = x98 &  n2718 ;
  assign n10761 = ( x100 & ~n2642 ) | ( x100 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n10762 = x99 &  n2637 ;
  assign n10763 = n10761 | n10762 ;
  assign n10765 = ( x98 & ~n10764 ) | ( x98 & n10763 ) | ( ~n10764 & n10763 ) ;
  assign n10766 = ( n2645 & ~n3354 ) | ( n2645 & n10765 ) | ( ~n3354 & n10765 ) ;
  assign n10767 = n3354 | n10766 ;
  assign n10769 = ( x32 & n10765 ) | ( x32 & n10767 ) | ( n10765 & n10767 ) ;
  assign n10768 = ( x32 & ~n10767 ) | ( x32 & n10765 ) | ( ~n10767 & n10765 ) ;
  assign n10770 = ( n10767 & ~n10769 ) | ( n10767 & n10768 ) | ( ~n10769 & n10768 ) ;
  assign n10772 = ( n10759 & n10760 ) | ( n10759 & n10770 ) | ( n10760 & n10770 ) ;
  assign n10771 = ( n10760 & ~n10759 ) | ( n10760 & n10770 ) | ( ~n10759 & n10770 ) ;
  assign n10773 = ( n10759 & ~n10772 ) | ( n10759 & n10771 ) | ( ~n10772 & n10771 ) ;
  assign n10774 = ( n10619 & n10620 ) | ( n10619 & n10773 ) | ( n10620 & n10773 ) ;
  assign n10775 = ( n10620 & ~n10619 ) | ( n10620 & n10773 ) | ( ~n10619 & n10773 ) ;
  assign n10776 = ( n10619 & ~n10774 ) | ( n10619 & n10775 ) | ( ~n10774 & n10775 ) ;
  assign n10781 = ( n10454 & n10776 ) | ( n10454 & n10779 ) | ( n10776 & n10779 ) ;
  assign n10780 = ( n10454 & ~n10779 ) | ( n10454 & n10776 ) | ( ~n10779 & n10776 ) ;
  assign n10782 = ( n10779 & ~n10781 ) | ( n10779 & n10780 ) | ( ~n10781 & n10780 ) ;
  assign n10786 = x107 &  n1551 ;
  assign n10783 = ( x109 & ~n1451 ) | ( x109 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n10784 = x108 &  n1446 ;
  assign n10785 = n10783 | n10784 ;
  assign n10787 = ( x107 & ~n10786 ) | ( x107 & n10785 ) | ( ~n10786 & n10785 ) ;
  assign n10788 = ~n1454 & n5267 ;
  assign n10789 = n10787 | n10788 ;
  assign n10790 = ( x23 & ~n10789 ) | ( x23 & 1'b0 ) | ( ~n10789 & 1'b0 ) ;
  assign n10791 = ~x23 & n10789 ;
  assign n10792 = n10790 | n10791 ;
  assign n10794 = ( n10602 & n10782 ) | ( n10602 & n10792 ) | ( n10782 & n10792 ) ;
  assign n10793 = ( n10782 & ~n10602 ) | ( n10782 & n10792 ) | ( ~n10602 & n10792 ) ;
  assign n10795 = ( n10602 & ~n10794 ) | ( n10602 & n10793 ) | ( ~n10794 & n10793 ) ;
  assign n10800 = ( n10601 & n10795 ) | ( n10601 & n10798 ) | ( n10795 & n10798 ) ;
  assign n10799 = ( n10601 & ~n10798 ) | ( n10601 & n10795 ) | ( ~n10798 & n10795 ) ;
  assign n10801 = ( n10798 & ~n10800 ) | ( n10798 & n10799 ) | ( ~n10800 & n10799 ) ;
  assign n10803 = ( n10475 & n10593 ) | ( n10475 & n10801 ) | ( n10593 & n10801 ) ;
  assign n10802 = ( n10475 & ~n10593 ) | ( n10475 & n10801 ) | ( ~n10593 & n10801 ) ;
  assign n10804 = ( n10593 & ~n10803 ) | ( n10593 & n10802 ) | ( ~n10803 & n10802 ) ;
  assign n10808 = x116 &  n713 ;
  assign n10805 = ( x118 & ~n641 ) | ( x118 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n10806 = x117 &  n636 ;
  assign n10807 = n10805 | n10806 ;
  assign n10809 = ( x116 & ~n10808 ) | ( x116 & n10807 ) | ( ~n10808 & n10807 ) ;
  assign n10810 = ( n644 & ~n7152 ) | ( n644 & n10809 ) | ( ~n7152 & n10809 ) ;
  assign n10811 = n7152 | n10810 ;
  assign n10813 = ( x14 & n10809 ) | ( x14 & n10811 ) | ( n10809 & n10811 ) ;
  assign n10812 = ( x14 & ~n10811 ) | ( x14 & n10809 ) | ( ~n10811 & n10809 ) ;
  assign n10814 = ( n10811 & ~n10813 ) | ( n10811 & n10812 ) | ( ~n10813 & n10812 ) ;
  assign n10815 = ( n10583 & ~n10804 ) | ( n10583 & n10814 ) | ( ~n10804 & n10814 ) ;
  assign n10816 = ( n10583 & ~n10814 ) | ( n10583 & n10804 ) | ( ~n10814 & n10804 ) ;
  assign n10817 = ( n10815 & ~n10583 ) | ( n10815 & n10816 ) | ( ~n10583 & n10816 ) ;
  assign n10818 = ( n10572 & n10582 ) | ( n10572 & n10817 ) | ( n10582 & n10817 ) ;
  assign n10819 = ( n10582 & ~n10572 ) | ( n10582 & n10817 ) | ( ~n10572 & n10817 ) ;
  assign n10820 = ( n10572 & ~n10818 ) | ( n10572 & n10819 ) | ( ~n10818 & n10819 ) ;
  assign n10824 = x122 &  n353 ;
  assign n10821 = ( x124 & ~n313 ) | ( x124 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n10822 = x123 &  n308 ;
  assign n10823 = n10821 | n10822 ;
  assign n10825 = ( x122 & ~n10824 ) | ( x122 & n10823 ) | ( ~n10824 & n10823 ) ;
  assign n10826 = ~n316 & n8755 ;
  assign n10827 = n10825 | n10826 ;
  assign n10828 = ( x8 & ~n10827 ) | ( x8 & 1'b0 ) | ( ~n10827 & 1'b0 ) ;
  assign n10829 = ~x8 & n10827 ;
  assign n10830 = n10828 | n10829 ;
  assign n10831 = ( n10566 & ~n10820 ) | ( n10566 & n10830 ) | ( ~n10820 & n10830 ) ;
  assign n10832 = ( n10820 & ~n10566 ) | ( n10820 & n10830 ) | ( ~n10566 & n10830 ) ;
  assign n10833 = ( n10831 & ~n10830 ) | ( n10831 & n10832 ) | ( ~n10830 & n10832 ) ;
  assign n10834 = ( n10552 & ~n10562 ) | ( n10552 & n10833 ) | ( ~n10562 & n10833 ) ;
  assign n10835 = ( n10562 & ~n10552 ) | ( n10562 & n10833 ) | ( ~n10552 & n10833 ) ;
  assign n10836 = ( n10834 & ~n10833 ) | ( n10834 & n10835 ) | ( ~n10833 & n10835 ) ;
  assign n10837 = ( n10252 & ~n10248 ) | ( n10252 & n10541 ) | ( ~n10248 & n10541 ) ;
  assign n10839 = ( n10545 & n10836 ) | ( n10545 & n10837 ) | ( n10836 & n10837 ) ;
  assign n10838 = ( n10836 & ~n10545 ) | ( n10836 & n10837 ) | ( ~n10545 & n10837 ) ;
  assign n10840 = ( n10545 & ~n10839 ) | ( n10545 & n10838 ) | ( ~n10839 & n10838 ) ;
  assign n10841 = ( n10545 & ~n10837 ) | ( n10545 & n10836 ) | ( ~n10837 & n10836 ) ;
  assign n10842 = ( n10572 & ~n10582 ) | ( n10572 & n10817 ) | ( ~n10582 & n10817 ) ;
  assign n11102 = x123 &  n353 ;
  assign n11099 = ( x125 & ~n313 ) | ( x125 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n11100 = x124 &  n308 ;
  assign n11101 = n11099 | n11100 ;
  assign n11103 = ( x123 & ~n11102 ) | ( x123 & n11101 ) | ( ~n11102 & n11101 ) ;
  assign n11104 = ( n316 & n9324 ) | ( n316 & n11103 ) | ( n9324 & n11103 ) ;
  assign n11105 = ( n9324 & ~n11104 ) | ( n9324 & 1'b0 ) | ( ~n11104 & 1'b0 ) ;
  assign n11106 = ( x8 & n11103 ) | ( x8 & n11105 ) | ( n11103 & n11105 ) ;
  assign n11107 = ( x8 & ~n11105 ) | ( x8 & n11103 ) | ( ~n11105 & n11103 ) ;
  assign n11108 = ( n11105 & ~n11106 ) | ( n11105 & n11107 ) | ( ~n11106 & n11107 ) ;
  assign n10843 = ( n10583 & n10804 ) | ( n10583 & n10814 ) | ( n10804 & n10814 ) ;
  assign n11076 = x117 &  n713 ;
  assign n11073 = ( x119 & ~n641 ) | ( x119 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n11074 = x118 &  n636 ;
  assign n11075 = n11073 | n11074 ;
  assign n11077 = ( x117 & ~n11076 ) | ( x117 & n11075 ) | ( ~n11076 & n11075 ) ;
  assign n11078 = ~n644 & n7648 ;
  assign n11079 = n11077 | n11078 ;
  assign n11080 = ~x14 & n11079 ;
  assign n11081 = x14 | n11079 ;
  assign n11082 = ( n11080 & ~n11079 ) | ( n11080 & n11081 ) | ( ~n11079 & n11081 ) ;
  assign n10844 = ( n10593 & ~n10475 ) | ( n10593 & n10801 ) | ( ~n10475 & n10801 ) ;
  assign n10848 = x114 &  n942 ;
  assign n10845 = ( x116 & ~n896 ) | ( x116 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n10846 = x115 &  n891 ;
  assign n10847 = n10845 | n10846 ;
  assign n10849 = ( x114 & ~n10848 ) | ( x114 & n10847 ) | ( ~n10848 & n10847 ) ;
  assign n10850 = n899 | n6885 ;
  assign n10851 = ~n10849 & n10850 ;
  assign n10852 = x17 &  n10851 ;
  assign n10853 = x17 | n10851 ;
  assign n10854 = ~n10852 & n10853 ;
  assign n11067 = x20 &  n10600 ;
  assign n11068 = ( n10796 & ~n11067 ) | ( n10796 & 1'b0 ) | ( ~n11067 & 1'b0 ) ;
  assign n11069 = ( n10601 & n10795 ) | ( n10601 & n11068 ) | ( n10795 & n11068 ) ;
  assign n10855 = ( n10602 & ~n10792 ) | ( n10602 & n10782 ) | ( ~n10792 & n10782 ) ;
  assign n10859 = x111 &  n1227 ;
  assign n10856 = ( x113 & ~n1154 ) | ( x113 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n10857 = x112 &  n1149 ;
  assign n10858 = n10856 | n10857 ;
  assign n10860 = ( x111 & ~n10859 ) | ( x111 & n10858 ) | ( ~n10859 & n10858 ) ;
  assign n10861 = n1157 | n6169 ;
  assign n10862 = ~n10860 & n10861 ;
  assign n10863 = x20 &  n10862 ;
  assign n10864 = x20 | n10862 ;
  assign n10865 = ~n10863 & n10864 ;
  assign n10869 = x108 &  n1551 ;
  assign n10866 = ( x110 & ~n1451 ) | ( x110 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n10867 = x109 &  n1446 ;
  assign n10868 = n10866 | n10867 ;
  assign n10870 = ( x108 & ~n10869 ) | ( x108 & n10868 ) | ( ~n10869 & n10868 ) ;
  assign n10871 = n1454 | n5283 ;
  assign n10872 = ~n10870 & n10871 ;
  assign n10873 = x23 &  n10872 ;
  assign n10874 = x23 | n10872 ;
  assign n10875 = ~n10873 & n10874 ;
  assign n10876 = ( n10619 & ~n10620 ) | ( n10619 & n10773 ) | ( ~n10620 & n10773 ) ;
  assign n10887 = ( n10759 & ~n10770 ) | ( n10759 & n10760 ) | ( ~n10770 & n10760 ) ;
  assign n10891 = x99 &  n2718 ;
  assign n10888 = ( x101 & ~n2642 ) | ( x101 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n10889 = x100 &  n2637 ;
  assign n10890 = n10888 | n10889 ;
  assign n10892 = ( x99 & ~n10891 ) | ( x99 & n10890 ) | ( ~n10891 & n10890 ) ;
  assign n10893 = ( n2645 & ~n3694 ) | ( n2645 & n10892 ) | ( ~n3694 & n10892 ) ;
  assign n10894 = n3694 | n10893 ;
  assign n10896 = ( x32 & n10892 ) | ( x32 & n10894 ) | ( n10892 & n10894 ) ;
  assign n10895 = ( x32 & ~n10894 ) | ( x32 & n10892 ) | ( ~n10894 & n10892 ) ;
  assign n10897 = ( n10894 & ~n10896 ) | ( n10894 & n10895 ) | ( ~n10896 & n10895 ) ;
  assign n10899 = ( n10431 & n10733 ) | ( n10431 & n10743 ) | ( n10733 & n10743 ) ;
  assign n10903 = x96 &  n3214 ;
  assign n10900 = ( x98 & ~n3087 ) | ( x98 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n10901 = x97 &  n3082 ;
  assign n10902 = n10900 | n10901 ;
  assign n10904 = ( x96 & ~n10903 ) | ( x96 & n10902 ) | ( ~n10903 & n10902 ) ;
  assign n10905 = ~n3090 & n3170 ;
  assign n10906 = n10904 | n10905 ;
  assign n10907 = ( x35 & ~n10906 ) | ( x35 & 1'b0 ) | ( ~n10906 & 1'b0 ) ;
  assign n10908 = ~x35 & n10906 ;
  assign n10909 = n10907 | n10908 ;
  assign n10910 = ( n10621 & n10720 ) | ( n10621 & n10730 ) | ( n10720 & n10730 ) ;
  assign n10911 = ( n10706 & n10716 ) | ( n10706 & n10717 ) | ( n10716 & n10717 ) ;
  assign n10912 = ( n10622 & n10693 ) | ( n10622 & n10703 ) | ( n10693 & n10703 ) ;
  assign n10913 = ( n10388 & n10680 ) | ( n10388 & n10690 ) | ( n10680 & n10690 ) ;
  assign n10914 = ( n10649 & n10650 ) | ( n10649 & n10660 ) | ( n10650 & n10660 ) ;
  assign n10934 = x72 &  n8558 ;
  assign n10931 = ( x74 & ~n8314 ) | ( x74 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n10932 = x73 &  n8309 ;
  assign n10933 = n10931 | n10932 ;
  assign n10935 = ( x72 & ~n10934 ) | ( x72 & n10933 ) | ( ~n10934 & n10933 ) ;
  assign n10936 = ( n482 & ~n8317 ) | ( n482 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n10937 = n10935 | n10936 ;
  assign n10918 = x69 &  n9457 ;
  assign n10915 = ( x71 & ~n9150 ) | ( x71 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n10916 = x70 &  n9145 ;
  assign n10917 = n10915 | n10916 ;
  assign n10919 = ( x69 & ~n10918 ) | ( x69 & n10917 ) | ( ~n10918 & n10917 ) ;
  assign n10920 = ( n298 & ~n9153 ) | ( n298 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n10921 = n10919 | n10920 ;
  assign n10922 = ( x62 & ~n10921 ) | ( x62 & 1'b0 ) | ( ~n10921 & 1'b0 ) ;
  assign n10923 = ~x62 & n10921 ;
  assign n10924 = n10922 | n10923 ;
  assign n10925 = x67 &  n10104 ;
  assign n10926 = ( x68 & ~n9760 ) | ( x68 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n10927 = n10925 | n10926 ;
  assign n10928 = ( x2 & n10924 ) | ( x2 & n10927 ) | ( n10924 & n10927 ) ;
  assign n10929 = ( x2 & ~n10924 ) | ( x2 & n10927 ) | ( ~n10924 & n10927 ) ;
  assign n10930 = ( n10924 & ~n10928 ) | ( n10924 & n10929 ) | ( ~n10928 & n10929 ) ;
  assign n10938 = ~x59 & n10647 ;
  assign n10939 = x59 | n10647 ;
  assign n10940 = ( n10938 & ~n10647 ) | ( n10938 & n10939 ) | ( ~n10647 & n10939 ) ;
  assign n10941 = ( n10937 & ~n10930 ) | ( n10937 & n10940 ) | ( ~n10930 & n10940 ) ;
  assign n10942 = ( n10930 & ~n10937 ) | ( n10930 & n10940 ) | ( ~n10937 & n10940 ) ;
  assign n10943 = ( n10941 & ~n10940 ) | ( n10941 & n10942 ) | ( ~n10940 & n10942 ) ;
  assign n10947 = x75 &  n7731 ;
  assign n10944 = ( x77 & ~n7538 ) | ( x77 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n10945 = x76 &  n7533 ;
  assign n10946 = n10944 | n10945 ;
  assign n10948 = ( x75 & ~n10947 ) | ( x75 & n10946 ) | ( ~n10947 & n10946 ) ;
  assign n10949 = ( n677 & ~n7541 ) | ( n677 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n10950 = n10948 | n10949 ;
  assign n10951 = ( x56 & ~n10950 ) | ( x56 & 1'b0 ) | ( ~n10950 & 1'b0 ) ;
  assign n10952 = ~x56 & n10950 ;
  assign n10953 = n10951 | n10952 ;
  assign n10954 = ( n10914 & ~n10943 ) | ( n10914 & n10953 ) | ( ~n10943 & n10953 ) ;
  assign n10955 = ( n10914 & ~n10953 ) | ( n10914 & n10943 ) | ( ~n10953 & n10943 ) ;
  assign n10956 = ( n10954 & ~n10914 ) | ( n10954 & n10955 ) | ( ~n10914 & n10955 ) ;
  assign n10967 = ( n10663 & n10664 ) | ( n10663 & n10674 ) | ( n10664 & n10674 ) ;
  assign n10960 = x78 &  n6982 ;
  assign n10957 = ( x80 & ~n6727 ) | ( x80 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n10958 = x79 &  n6722 ;
  assign n10959 = n10957 | n10958 ;
  assign n10961 = ( x78 & ~n10960 ) | ( x78 & n10959 ) | ( ~n10960 & n10959 ) ;
  assign n10962 = ( n842 & ~n6730 ) | ( n842 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n10963 = n10961 | n10962 ;
  assign n10964 = ( x53 & ~n10963 ) | ( x53 & 1'b0 ) | ( ~n10963 & 1'b0 ) ;
  assign n10965 = ~x53 & n10963 ;
  assign n10966 = n10964 | n10965 ;
  assign n10968 = ( n10956 & ~n10967 ) | ( n10956 & n10966 ) | ( ~n10967 & n10966 ) ;
  assign n10969 = ( n10956 & ~n10966 ) | ( n10956 & n10967 ) | ( ~n10966 & n10967 ) ;
  assign n10970 = ( n10968 & ~n10956 ) | ( n10968 & n10969 ) | ( ~n10956 & n10969 ) ;
  assign n10974 = x81 &  n6288 ;
  assign n10971 = ( x83 & ~n6032 ) | ( x83 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n10972 = x82 &  n6027 ;
  assign n10973 = n10971 | n10972 ;
  assign n10975 = ( x81 & ~n10974 ) | ( x81 & n10973 ) | ( ~n10974 & n10973 ) ;
  assign n10976 = ( n1100 & ~n6035 ) | ( n1100 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n10977 = n10975 | n10976 ;
  assign n10978 = ( x50 & ~n10977 ) | ( x50 & 1'b0 ) | ( ~n10977 & 1'b0 ) ;
  assign n10979 = ~x50 & n10977 ;
  assign n10980 = n10978 | n10979 ;
  assign n10981 = ( n10679 & ~n10970 ) | ( n10679 & n10980 ) | ( ~n10970 & n10980 ) ;
  assign n10982 = ( n10679 & ~n10980 ) | ( n10679 & n10970 ) | ( ~n10980 & n10970 ) ;
  assign n10983 = ( n10981 & ~n10679 ) | ( n10981 & n10982 ) | ( ~n10679 & n10982 ) ;
  assign n10987 = x84 &  n5586 ;
  assign n10984 = ( x86 & ~n5389 ) | ( x86 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n10985 = x85 &  n5384 ;
  assign n10986 = n10984 | n10985 ;
  assign n10988 = ( x84 & ~n10987 ) | ( x84 & n10986 ) | ( ~n10987 & n10986 ) ;
  assign n10989 = ( n1496 & ~n5392 ) | ( n1496 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n10990 = n10988 | n10989 ;
  assign n10991 = ( x47 & ~n10990 ) | ( x47 & 1'b0 ) | ( ~n10990 & 1'b0 ) ;
  assign n10992 = ~x47 & n10990 ;
  assign n10993 = n10991 | n10992 ;
  assign n10994 = ( n10913 & ~n10983 ) | ( n10913 & n10993 ) | ( ~n10983 & n10993 ) ;
  assign n10995 = ( n10913 & ~n10993 ) | ( n10913 & n10983 ) | ( ~n10993 & n10983 ) ;
  assign n10996 = ( n10994 & ~n10913 ) | ( n10994 & n10995 ) | ( ~n10913 & n10995 ) ;
  assign n11000 = x87 &  n4934 ;
  assign n10997 = ( x89 & ~n4725 ) | ( x89 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n10998 = x88 &  n4720 ;
  assign n10999 = n10997 | n10998 ;
  assign n11001 = ( x87 & ~n11000 ) | ( x87 & n10999 ) | ( ~n11000 & n10999 ) ;
  assign n11002 = ( n1741 & ~n4728 ) | ( n1741 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n11003 = n11001 | n11002 ;
  assign n11004 = ( x44 & ~n11003 ) | ( x44 & 1'b0 ) | ( ~n11003 & 1'b0 ) ;
  assign n11005 = ~x44 & n11003 ;
  assign n11006 = n11004 | n11005 ;
  assign n11007 = ( n10912 & ~n10996 ) | ( n10912 & n11006 ) | ( ~n10996 & n11006 ) ;
  assign n11008 = ( n10912 & ~n11006 ) | ( n10912 & n10996 ) | ( ~n11006 & n10996 ) ;
  assign n11009 = ( n11007 & ~n10912 ) | ( n11007 & n11008 ) | ( ~n10912 & n11008 ) ;
  assign n11013 = x90 &  n4344 ;
  assign n11010 = ( x92 & ~n4143 ) | ( x92 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n11011 = x91 &  n4138 ;
  assign n11012 = n11010 | n11011 ;
  assign n11014 = ( x90 & ~n11013 ) | ( x90 & n11012 ) | ( ~n11013 & n11012 ) ;
  assign n11015 = ( n2248 & ~n4146 ) | ( n2248 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n11016 = n11014 | n11015 ;
  assign n11017 = ( x41 & ~n11016 ) | ( x41 & 1'b0 ) | ( ~n11016 & 1'b0 ) ;
  assign n11018 = ~x41 & n11016 ;
  assign n11019 = n11017 | n11018 ;
  assign n11020 = ( n10911 & ~n11009 ) | ( n10911 & n11019 ) | ( ~n11009 & n11019 ) ;
  assign n11021 = ( n10911 & ~n11019 ) | ( n10911 & n11009 ) | ( ~n11019 & n11009 ) ;
  assign n11022 = ( n11020 & ~n10911 ) | ( n11020 & n11021 ) | ( ~n10911 & n11021 ) ;
  assign n11026 = x93 &  n3756 ;
  assign n11023 = ( x95 & ~n3602 ) | ( x95 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n11024 = x94 &  n3597 ;
  assign n11025 = n11023 | n11024 ;
  assign n11027 = ( x93 & ~n11026 ) | ( x93 & n11025 ) | ( ~n11026 & n11025 ) ;
  assign n11028 = ( n2547 & ~n3605 ) | ( n2547 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n11029 = n11027 | n11028 ;
  assign n11030 = ( x38 & ~n11029 ) | ( x38 & 1'b0 ) | ( ~n11029 & 1'b0 ) ;
  assign n11031 = ~x38 & n11029 ;
  assign n11032 = n11030 | n11031 ;
  assign n11033 = ( n10910 & ~n11022 ) | ( n10910 & n11032 ) | ( ~n11022 & n11032 ) ;
  assign n11034 = ( n10910 & ~n11032 ) | ( n10910 & n11022 ) | ( ~n11032 & n11022 ) ;
  assign n11035 = ( n11033 & ~n10910 ) | ( n11033 & n11034 ) | ( ~n10910 & n11034 ) ;
  assign n11037 = ( n10899 & n10909 ) | ( n10899 & n11035 ) | ( n10909 & n11035 ) ;
  assign n11036 = ( n10909 & ~n10899 ) | ( n10909 & n11035 ) | ( ~n10899 & n11035 ) ;
  assign n11038 = ( n10899 & ~n11037 ) | ( n10899 & n11036 ) | ( ~n11037 & n11036 ) ;
  assign n10898 = ( n10434 & n10746 ) | ( n10434 & n10756 ) | ( n10746 & n10756 ) ;
  assign n11039 = ( n10897 & ~n11038 ) | ( n10897 & n10898 ) | ( ~n11038 & n10898 ) ;
  assign n11040 = ( n10897 & ~n10898 ) | ( n10897 & n11038 ) | ( ~n10898 & n11038 ) ;
  assign n11041 = ( n11039 & ~n10897 ) | ( n11039 & n11040 ) | ( ~n10897 & n11040 ) ;
  assign n11045 = x102 &  n2312 ;
  assign n11042 = ( x104 & ~n2195 ) | ( x104 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n11043 = x103 &  n2190 ;
  assign n11044 = n11042 | n11043 ;
  assign n11046 = ( x102 & ~n11045 ) | ( x102 & n11044 ) | ( ~n11045 & n11044 ) ;
  assign n11047 = ( n2198 & ~n4249 ) | ( n2198 & n11046 ) | ( ~n4249 & n11046 ) ;
  assign n11048 = n4249 | n11047 ;
  assign n11050 = ( x29 & n11046 ) | ( x29 & n11048 ) | ( n11046 & n11048 ) ;
  assign n11049 = ( x29 & ~n11048 ) | ( x29 & n11046 ) | ( ~n11048 & n11046 ) ;
  assign n11051 = ( n11048 & ~n11050 ) | ( n11048 & n11049 ) | ( ~n11050 & n11049 ) ;
  assign n11053 = ( n10887 & n11041 ) | ( n10887 & n11051 ) | ( n11041 & n11051 ) ;
  assign n11052 = ( n11041 & ~n10887 ) | ( n11041 & n11051 ) | ( ~n10887 & n11051 ) ;
  assign n11054 = ( n10887 & ~n11053 ) | ( n10887 & n11052 ) | ( ~n11053 & n11052 ) ;
  assign n10880 = x105 &  n1894 ;
  assign n10877 = ( x107 & ~n1816 ) | ( x107 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n10878 = x106 &  n1811 ;
  assign n10879 = n10877 | n10878 ;
  assign n10881 = ( x105 & ~n10880 ) | ( x105 & n10879 ) | ( ~n10880 & n10879 ) ;
  assign n10882 = ~n1819 & n4848 ;
  assign n10883 = n10881 | n10882 ;
  assign n10885 = x26 &  n10883 ;
  assign n10884 = ~x26 & n10883 ;
  assign n10886 = ( x26 & ~n10885 ) | ( x26 & n10884 ) | ( ~n10885 & n10884 ) ;
  assign n11055 = ( n10876 & ~n11054 ) | ( n10876 & n10886 ) | ( ~n11054 & n10886 ) ;
  assign n11056 = ( n10876 & ~n10886 ) | ( n10876 & n11054 ) | ( ~n10886 & n11054 ) ;
  assign n11057 = ( n11055 & ~n10876 ) | ( n11055 & n11056 ) | ( ~n10876 & n11056 ) ;
  assign n11058 = x26 &  n10609 ;
  assign n11059 = ( n10777 & ~n11058 ) | ( n10777 & 1'b0 ) | ( ~n11058 & 1'b0 ) ;
  assign n11060 = ( n10776 & ~n10454 ) | ( n10776 & n11059 ) | ( ~n10454 & n11059 ) ;
  assign n11062 = ( n10875 & n11057 ) | ( n10875 & n11060 ) | ( n11057 & n11060 ) ;
  assign n11061 = ( n11057 & ~n10875 ) | ( n11057 & n11060 ) | ( ~n10875 & n11060 ) ;
  assign n11063 = ( n10875 & ~n11062 ) | ( n10875 & n11061 ) | ( ~n11062 & n11061 ) ;
  assign n11065 = ( n10855 & n10865 ) | ( n10855 & n11063 ) | ( n10865 & n11063 ) ;
  assign n11064 = ( n10865 & ~n10855 ) | ( n10865 & n11063 ) | ( ~n10855 & n11063 ) ;
  assign n11066 = ( n10855 & ~n11065 ) | ( n10855 & n11064 ) | ( ~n11065 & n11064 ) ;
  assign n11070 = ( n10854 & ~n11069 ) | ( n10854 & n11066 ) | ( ~n11069 & n11066 ) ;
  assign n11071 = ( n10854 & ~n11066 ) | ( n10854 & n11069 ) | ( ~n11066 & n11069 ) ;
  assign n11072 = ( n11070 & ~n10854 ) | ( n11070 & n11071 ) | ( ~n10854 & n11071 ) ;
  assign n11083 = ( n10844 & n11072 ) | ( n10844 & n11082 ) | ( n11072 & n11082 ) ;
  assign n11084 = ( n10844 & ~n11082 ) | ( n10844 & n11072 ) | ( ~n11082 & n11072 ) ;
  assign n11085 = ( n11082 & ~n11083 ) | ( n11082 & n11084 ) | ( ~n11083 & n11084 ) ;
  assign n11089 = x120 &  n503 ;
  assign n11086 = ( x122 & ~n450 ) | ( x122 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n11087 = x121 &  n445 ;
  assign n11088 = n11086 | n11087 ;
  assign n11090 = ( x120 & ~n11089 ) | ( x120 & n11088 ) | ( ~n11089 & n11088 ) ;
  assign n11091 = ( n453 & n9987 ) | ( n453 & n11090 ) | ( n9987 & n11090 ) ;
  assign n11092 = ( n9987 & ~n11091 ) | ( n9987 & 1'b0 ) | ( ~n11091 & 1'b0 ) ;
  assign n11093 = ( x11 & n11090 ) | ( x11 & n11092 ) | ( n11090 & n11092 ) ;
  assign n11094 = ( x11 & ~n11092 ) | ( x11 & n11090 ) | ( ~n11092 & n11090 ) ;
  assign n11095 = ( n11092 & ~n11093 ) | ( n11092 & n11094 ) | ( ~n11093 & n11094 ) ;
  assign n11097 = ( n10843 & n11085 ) | ( n10843 & n11095 ) | ( n11085 & n11095 ) ;
  assign n11096 = ( n11085 & ~n10843 ) | ( n11085 & n11095 ) | ( ~n10843 & n11095 ) ;
  assign n11098 = ( n10843 & ~n11097 ) | ( n10843 & n11096 ) | ( ~n11097 & n11096 ) ;
  assign n11109 = ( n10842 & ~n11108 ) | ( n10842 & n11098 ) | ( ~n11108 & n11098 ) ;
  assign n11110 = ( n10842 & ~n11098 ) | ( n10842 & n11108 ) | ( ~n11098 & n11108 ) ;
  assign n11111 = ( n11109 & ~n10842 ) | ( n11109 & n11110 ) | ( ~n10842 & n11110 ) ;
  assign n11112 = ( x126 & ~n225 ) | ( x126 & 1'b0 ) | ( ~n225 & 1'b0 ) ;
  assign n11113 = x127 &  n192 ;
  assign n11114 = n11112 | n11113 ;
  assign n11115 = n200 | n9960 ;
  assign n11116 = ( n11114 & ~n200 ) | ( n11114 & n11115 ) | ( ~n200 & n11115 ) ;
  assign n11117 = ( x5 & ~n11116 ) | ( x5 & 1'b0 ) | ( ~n11116 & 1'b0 ) ;
  assign n11118 = ~x5 & n11116 ;
  assign n11119 = n11117 | n11118 ;
  assign n11120 = ( n10566 & n10820 ) | ( n10566 & n10830 ) | ( n10820 & n10830 ) ;
  assign n11122 = ( n11111 & n11119 ) | ( n11111 & n11120 ) | ( n11119 & n11120 ) ;
  assign n11121 = ( n11119 & ~n11111 ) | ( n11119 & n11120 ) | ( ~n11111 & n11120 ) ;
  assign n11123 = ( n11111 & ~n11122 ) | ( n11111 & n11121 ) | ( ~n11122 & n11121 ) ;
  assign n11124 = ( n10834 & n10841 ) | ( n10834 & n11123 ) | ( n10841 & n11123 ) ;
  assign n11125 = ( n10841 & ~n10834 ) | ( n10841 & n11123 ) | ( ~n10834 & n11123 ) ;
  assign n11126 = ( n10834 & ~n11124 ) | ( n10834 & n11125 ) | ( ~n11124 & n11125 ) ;
  assign n11127 = ( n11098 & ~n10842 ) | ( n11098 & n11108 ) | ( ~n10842 & n11108 ) ;
  assign n11128 = ( x127 & ~n225 ) | ( x127 & 1'b0 ) | ( ~n225 & 1'b0 ) ;
  assign n11129 = n200 | n10258 ;
  assign n11130 = ~n11128 & n11129 ;
  assign n11131 = x5 &  n11130 ;
  assign n11132 = x5 | n11130 ;
  assign n11133 = ~n11131 & n11132 ;
  assign n11134 = x14 &  n11079 ;
  assign n11135 = ( x14 & ~n11134 ) | ( x14 & n11080 ) | ( ~n11134 & n11080 ) ;
  assign n11136 = ( n10844 & ~n11072 ) | ( n10844 & n11135 ) | ( ~n11072 & n11135 ) ;
  assign n11140 = x121 &  n503 ;
  assign n11137 = ( x123 & ~n450 ) | ( x123 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n11138 = x122 &  n445 ;
  assign n11139 = n11137 | n11138 ;
  assign n11141 = ( x121 & ~n11140 ) | ( x121 & n11139 ) | ( ~n11140 & n11139 ) ;
  assign n11142 = ~n453 & n8472 ;
  assign n11143 = n11141 | n11142 ;
  assign n11144 = ( x11 & ~n11143 ) | ( x11 & 1'b0 ) | ( ~n11143 & 1'b0 ) ;
  assign n11145 = ~x11 & n11143 ;
  assign n11146 = n11144 | n11145 ;
  assign n11147 = ( n11066 & ~n10854 ) | ( n11066 & n11069 ) | ( ~n10854 & n11069 ) ;
  assign n11151 = x118 &  n713 ;
  assign n11148 = ( x120 & ~n641 ) | ( x120 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n11149 = x119 &  n636 ;
  assign n11150 = n11148 | n11149 ;
  assign n11152 = ( x118 & ~n11151 ) | ( x118 & n11150 ) | ( ~n11151 & n11150 ) ;
  assign n11153 = ~n644 & n9364 ;
  assign n11154 = n11152 | n11153 ;
  assign n11155 = ( x14 & ~n11154 ) | ( x14 & 1'b0 ) | ( ~n11154 & 1'b0 ) ;
  assign n11156 = ~x14 & n11154 ;
  assign n11157 = n11155 | n11156 ;
  assign n11161 = x115 &  n942 ;
  assign n11158 = ( x117 & ~n896 ) | ( x117 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n11159 = x116 &  n891 ;
  assign n11160 = n11158 | n11159 ;
  assign n11162 = ( x115 & ~n11161 ) | ( x115 & n11160 ) | ( ~n11161 & n11160 ) ;
  assign n11163 = ( n899 & ~n7136 ) | ( n899 & n11162 ) | ( ~n7136 & n11162 ) ;
  assign n11164 = n7136 | n11163 ;
  assign n11166 = ( x17 & n11162 ) | ( x17 & n11164 ) | ( n11162 & n11164 ) ;
  assign n11165 = ( x17 & ~n11164 ) | ( x17 & n11162 ) | ( ~n11164 & n11162 ) ;
  assign n11167 = ( n11164 & ~n11166 ) | ( n11164 & n11165 ) | ( ~n11166 & n11165 ) ;
  assign n11168 = ( n10855 & ~n11063 ) | ( n10855 & n10865 ) | ( ~n11063 & n10865 ) ;
  assign n11169 = ( n10875 & ~n11060 ) | ( n10875 & n11057 ) | ( ~n11060 & n11057 ) ;
  assign n11173 = x112 &  n1227 ;
  assign n11170 = ( x114 & ~n1154 ) | ( x114 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n11171 = x113 &  n1149 ;
  assign n11172 = n11170 | n11171 ;
  assign n11174 = ( x112 & ~n11173 ) | ( x112 & n11172 ) | ( ~n11173 & n11172 ) ;
  assign n11175 = n1157 | n6185 ;
  assign n11176 = ~n11174 & n11175 ;
  assign n11177 = x20 &  n11176 ;
  assign n11178 = x20 | n11176 ;
  assign n11179 = ~n11177 & n11178 ;
  assign n11180 = ( n10886 & ~n10876 ) | ( n10886 & n11054 ) | ( ~n10876 & n11054 ) ;
  assign n11184 = x109 &  n1551 ;
  assign n11181 = ( x111 & ~n1451 ) | ( x111 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n11182 = x110 &  n1446 ;
  assign n11183 = n11181 | n11182 ;
  assign n11185 = ( x109 & ~n11184 ) | ( x109 & n11183 ) | ( ~n11184 & n11183 ) ;
  assign n11186 = n1454 | n5711 ;
  assign n11187 = ~n11185 & n11186 ;
  assign n11188 = x23 &  n11187 ;
  assign n11189 = x23 | n11187 ;
  assign n11190 = ~n11188 & n11189 ;
  assign n11191 = ( n10898 & ~n10897 ) | ( n10898 & n11038 ) | ( ~n10897 & n11038 ) ;
  assign n11195 = x103 &  n2312 ;
  assign n11192 = ( x105 & ~n2195 ) | ( x105 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n11193 = x104 &  n2190 ;
  assign n11194 = n11192 | n11193 ;
  assign n11196 = ( x103 & ~n11195 ) | ( x103 & n11194 ) | ( ~n11195 & n11194 ) ;
  assign n11197 = ~n2198 & n4442 ;
  assign n11198 = n11196 | n11197 ;
  assign n11199 = ( x29 & ~n11198 ) | ( x29 & 1'b0 ) | ( ~n11198 & 1'b0 ) ;
  assign n11200 = ~x29 & n11198 ;
  assign n11201 = n11199 | n11200 ;
  assign n11349 = x100 &  n2718 ;
  assign n11346 = ( x102 & ~n2642 ) | ( x102 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n11347 = x101 &  n2637 ;
  assign n11348 = n11346 | n11347 ;
  assign n11350 = ( x100 & ~n11349 ) | ( x100 & n11348 ) | ( ~n11349 & n11348 ) ;
  assign n11351 = ( n2645 & ~n3872 ) | ( n2645 & n11350 ) | ( ~n3872 & n11350 ) ;
  assign n11352 = n3872 | n11351 ;
  assign n11354 = ( x32 & n11350 ) | ( x32 & n11352 ) | ( n11350 & n11352 ) ;
  assign n11353 = ( x32 & ~n11352 ) | ( x32 & n11350 ) | ( ~n11352 & n11350 ) ;
  assign n11355 = ( n11352 & ~n11354 ) | ( n11352 & n11353 ) | ( ~n11354 & n11353 ) ;
  assign n11202 = ( n10911 & n11009 ) | ( n10911 & n11019 ) | ( n11009 & n11019 ) ;
  assign n11203 = ( n10912 & n10996 ) | ( n10912 & n11006 ) | ( n10996 & n11006 ) ;
  assign n11204 = ( n10913 & n10983 ) | ( n10913 & n10993 ) | ( n10983 & n10993 ) ;
  assign n11205 = ( n10956 & n10966 ) | ( n10956 & n10967 ) | ( n10966 & n10967 ) ;
  assign n11206 = ( n10914 & n10943 ) | ( n10914 & n10953 ) | ( n10943 & n10953 ) ;
  assign n11210 = x70 &  n9457 ;
  assign n11207 = ( x72 & ~n9150 ) | ( x72 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n11208 = x71 &  n9145 ;
  assign n11209 = n11207 | n11208 ;
  assign n11211 = ( x70 & ~n11210 ) | ( x70 & n11209 ) | ( ~n11210 & n11209 ) ;
  assign n11212 = ( n345 & ~n11211 ) | ( n345 & n9153 ) | ( ~n11211 & n9153 ) ;
  assign n11213 = ~n9153 & n11212 ;
  assign n11214 = ( x62 & n11211 ) | ( x62 & n11213 ) | ( n11211 & n11213 ) ;
  assign n11215 = ( x62 & ~n11213 ) | ( x62 & n11211 ) | ( ~n11213 & n11211 ) ;
  assign n11216 = ( n11213 & ~n11214 ) | ( n11213 & n11215 ) | ( ~n11214 & n11215 ) ;
  assign n11217 = x68 &  n10104 ;
  assign n11218 = ( x69 & ~n9760 ) | ( x69 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n11219 = n11217 | n11218 ;
  assign n11220 = ( x2 & n11216 ) | ( x2 & n11219 ) | ( n11216 & n11219 ) ;
  assign n11221 = ( x2 & ~n11216 ) | ( x2 & n11219 ) | ( ~n11216 & n11219 ) ;
  assign n11222 = ( n11216 & ~n11220 ) | ( n11216 & n11221 ) | ( ~n11220 & n11221 ) ;
  assign n11226 = x73 &  n8558 ;
  assign n11223 = ( x75 & ~n8314 ) | ( x75 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n11224 = x74 &  n8309 ;
  assign n11225 = n11223 | n11224 ;
  assign n11227 = ( x73 & ~n11226 ) | ( x73 & n11225 ) | ( ~n11226 & n11225 ) ;
  assign n11228 = ( n540 & ~n11227 ) | ( n540 & n8317 ) | ( ~n11227 & n8317 ) ;
  assign n11229 = ~n8317 & n11228 ;
  assign n11230 = ( x59 & n11227 ) | ( x59 & n11229 ) | ( n11227 & n11229 ) ;
  assign n11231 = ( x59 & ~n11229 ) | ( x59 & n11227 ) | ( ~n11229 & n11227 ) ;
  assign n11232 = ( n11229 & ~n11230 ) | ( n11229 & n11231 ) | ( ~n11230 & n11231 ) ;
  assign n11233 = ( n10928 & ~n11222 ) | ( n10928 & n11232 ) | ( ~n11222 & n11232 ) ;
  assign n11234 = ( n10928 & ~n11232 ) | ( n10928 & n11222 ) | ( ~n11232 & n11222 ) ;
  assign n11235 = ( n11233 & ~n10928 ) | ( n11233 & n11234 ) | ( ~n10928 & n11234 ) ;
  assign n11246 = x59 | n10937 ;
  assign n11247 = x59 &  n10937 ;
  assign n11248 = ( n11246 & ~n11247 ) | ( n11246 & 1'b0 ) | ( ~n11247 & 1'b0 ) ;
  assign n11249 = ( n10647 & n10930 ) | ( n10647 & n11248 ) | ( n10930 & n11248 ) ;
  assign n11239 = x76 &  n7731 ;
  assign n11236 = ( x78 & ~n7538 ) | ( x78 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n11237 = x77 &  n7533 ;
  assign n11238 = n11236 | n11237 ;
  assign n11240 = ( x76 & ~n11239 ) | ( x76 & n11238 ) | ( ~n11239 & n11238 ) ;
  assign n11241 = ( n693 & ~n11240 ) | ( n693 & n7541 ) | ( ~n11240 & n7541 ) ;
  assign n11242 = ~n7541 & n11241 ;
  assign n11243 = ( x56 & n11240 ) | ( x56 & n11242 ) | ( n11240 & n11242 ) ;
  assign n11244 = ( x56 & ~n11242 ) | ( x56 & n11240 ) | ( ~n11242 & n11240 ) ;
  assign n11245 = ( n11242 & ~n11243 ) | ( n11242 & n11244 ) | ( ~n11243 & n11244 ) ;
  assign n11250 = ( n11235 & ~n11249 ) | ( n11235 & n11245 ) | ( ~n11249 & n11245 ) ;
  assign n11251 = ( n11235 & ~n11245 ) | ( n11235 & n11249 ) | ( ~n11245 & n11249 ) ;
  assign n11252 = ( n11250 & ~n11235 ) | ( n11250 & n11251 ) | ( ~n11235 & n11251 ) ;
  assign n11256 = x79 &  n6982 ;
  assign n11253 = ( x81 & ~n6727 ) | ( x81 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n11254 = x80 &  n6722 ;
  assign n11255 = n11253 | n11254 ;
  assign n11257 = ( x79 & ~n11256 ) | ( x79 & n11255 ) | ( ~n11256 & n11255 ) ;
  assign n11258 = ( n994 & ~n6730 ) | ( n994 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n11259 = n11257 | n11258 ;
  assign n11261 = x53 &  n11259 ;
  assign n11260 = ~x53 & n11259 ;
  assign n11262 = ( x53 & ~n11261 ) | ( x53 & n11260 ) | ( ~n11261 & n11260 ) ;
  assign n11263 = ( n11206 & ~n11252 ) | ( n11206 & n11262 ) | ( ~n11252 & n11262 ) ;
  assign n11264 = ( n11206 & ~n11262 ) | ( n11206 & n11252 ) | ( ~n11262 & n11252 ) ;
  assign n11265 = ( n11263 & ~n11206 ) | ( n11263 & n11264 ) | ( ~n11206 & n11264 ) ;
  assign n11269 = x82 &  n6288 ;
  assign n11266 = ( x84 & ~n6032 ) | ( x84 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n11267 = x83 &  n6027 ;
  assign n11268 = n11266 | n11267 ;
  assign n11270 = ( x82 & ~n11269 ) | ( x82 & n11268 ) | ( ~n11269 & n11268 ) ;
  assign n11271 = ( n1199 & ~n6035 ) | ( n1199 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n11272 = n11270 | n11271 ;
  assign n11273 = ( x50 & ~n11272 ) | ( x50 & 1'b0 ) | ( ~n11272 & 1'b0 ) ;
  assign n11274 = ~x50 & n11272 ;
  assign n11275 = n11273 | n11274 ;
  assign n11276 = ( n11205 & ~n11265 ) | ( n11205 & n11275 ) | ( ~n11265 & n11275 ) ;
  assign n11277 = ( n11205 & ~n11275 ) | ( n11205 & n11265 ) | ( ~n11275 & n11265 ) ;
  assign n11278 = ( n11276 & ~n11205 ) | ( n11276 & n11277 ) | ( ~n11205 & n11277 ) ;
  assign n11289 = ( n10679 & n10970 ) | ( n10679 & n10980 ) | ( n10970 & n10980 ) ;
  assign n11282 = x85 &  n5586 ;
  assign n11279 = ( x87 & ~n5389 ) | ( x87 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n11280 = x86 &  n5384 ;
  assign n11281 = n11279 | n11280 ;
  assign n11283 = ( x85 & ~n11282 ) | ( x85 & n11281 ) | ( ~n11282 & n11281 ) ;
  assign n11284 = ( n1512 & ~n5392 ) | ( n1512 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n11285 = n11283 | n11284 ;
  assign n11286 = ( x47 & ~n11285 ) | ( x47 & 1'b0 ) | ( ~n11285 & 1'b0 ) ;
  assign n11287 = ~x47 & n11285 ;
  assign n11288 = n11286 | n11287 ;
  assign n11290 = ( n11278 & ~n11289 ) | ( n11278 & n11288 ) | ( ~n11289 & n11288 ) ;
  assign n11291 = ( n11278 & ~n11288 ) | ( n11278 & n11289 ) | ( ~n11288 & n11289 ) ;
  assign n11292 = ( n11290 & ~n11278 ) | ( n11290 & n11291 ) | ( ~n11278 & n11291 ) ;
  assign n11296 = x88 &  n4934 ;
  assign n11293 = ( x90 & ~n4725 ) | ( x90 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n11294 = x89 &  n4720 ;
  assign n11295 = n11293 | n11294 ;
  assign n11297 = ( x88 & ~n11296 ) | ( x88 & n11295 ) | ( ~n11296 & n11295 ) ;
  assign n11298 = ( n1976 & ~n4728 ) | ( n1976 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n11299 = n11297 | n11298 ;
  assign n11300 = ( x44 & ~n11299 ) | ( x44 & 1'b0 ) | ( ~n11299 & 1'b0 ) ;
  assign n11301 = ~x44 & n11299 ;
  assign n11302 = n11300 | n11301 ;
  assign n11303 = ( n11204 & ~n11292 ) | ( n11204 & n11302 ) | ( ~n11292 & n11302 ) ;
  assign n11304 = ( n11204 & ~n11302 ) | ( n11204 & n11292 ) | ( ~n11302 & n11292 ) ;
  assign n11305 = ( n11303 & ~n11204 ) | ( n11303 & n11304 ) | ( ~n11204 & n11304 ) ;
  assign n11309 = x91 &  n4344 ;
  assign n11306 = ( x93 & ~n4143 ) | ( x93 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n11307 = x92 &  n4138 ;
  assign n11308 = n11306 | n11307 ;
  assign n11310 = ( x91 & ~n11309 ) | ( x91 & n11308 ) | ( ~n11309 & n11308 ) ;
  assign n11311 = n2264 | n4146 ;
  assign n11312 = ~n11310 & n11311 ;
  assign n11313 = x41 &  n11312 ;
  assign n11314 = x41 | n11312 ;
  assign n11315 = ~n11313 & n11314 ;
  assign n11317 = ( n11203 & n11305 ) | ( n11203 & n11315 ) | ( n11305 & n11315 ) ;
  assign n11316 = ( n11305 & ~n11203 ) | ( n11305 & n11315 ) | ( ~n11203 & n11315 ) ;
  assign n11318 = ( n11203 & ~n11317 ) | ( n11203 & n11316 ) | ( ~n11317 & n11316 ) ;
  assign n11322 = x94 &  n3756 ;
  assign n11319 = ( x96 & ~n3602 ) | ( x96 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n11320 = x95 &  n3597 ;
  assign n11321 = n11319 | n11320 ;
  assign n11323 = ( x94 & ~n11322 ) | ( x94 & n11321 ) | ( ~n11322 & n11321 ) ;
  assign n11324 = ( n2836 & ~n3605 ) | ( n2836 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n11325 = n11323 | n11324 ;
  assign n11326 = ( x38 & ~n11325 ) | ( x38 & 1'b0 ) | ( ~n11325 & 1'b0 ) ;
  assign n11327 = ~x38 & n11325 ;
  assign n11328 = n11326 | n11327 ;
  assign n11329 = ( n11202 & n11318 ) | ( n11202 & n11328 ) | ( n11318 & n11328 ) ;
  assign n11330 = ( n11318 & ~n11202 ) | ( n11318 & n11328 ) | ( ~n11202 & n11328 ) ;
  assign n11331 = ( n11202 & ~n11329 ) | ( n11202 & n11330 ) | ( ~n11329 & n11330 ) ;
  assign n11335 = x97 &  n3214 ;
  assign n11332 = ( x99 & ~n3087 ) | ( x99 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n11333 = x98 &  n3082 ;
  assign n11334 = n11332 | n11333 ;
  assign n11336 = ( x97 & ~n11335 ) | ( x97 & n11334 ) | ( ~n11335 & n11334 ) ;
  assign n11337 = ~n3090 & n3338 ;
  assign n11338 = n11336 | n11337 ;
  assign n11339 = ( x35 & ~n11338 ) | ( x35 & 1'b0 ) | ( ~n11338 & 1'b0 ) ;
  assign n11340 = ~x35 & n11338 ;
  assign n11341 = n11339 | n11340 ;
  assign n11342 = ( n10910 & n11022 ) | ( n10910 & n11032 ) | ( n11022 & n11032 ) ;
  assign n11343 = ( n11331 & ~n11341 ) | ( n11331 & n11342 ) | ( ~n11341 & n11342 ) ;
  assign n11344 = ( n11331 & ~n11342 ) | ( n11331 & n11341 ) | ( ~n11342 & n11341 ) ;
  assign n11345 = ( n11343 & ~n11331 ) | ( n11343 & n11344 ) | ( ~n11331 & n11344 ) ;
  assign n11356 = ( n11037 & ~n11355 ) | ( n11037 & n11345 ) | ( ~n11355 & n11345 ) ;
  assign n11357 = ( n11037 & ~n11345 ) | ( n11037 & n11355 ) | ( ~n11345 & n11355 ) ;
  assign n11358 = ( n11356 & ~n11037 ) | ( n11356 & n11357 ) | ( ~n11037 & n11357 ) ;
  assign n11359 = ( n11191 & ~n11201 ) | ( n11191 & n11358 ) | ( ~n11201 & n11358 ) ;
  assign n11360 = ( n11191 & ~n11358 ) | ( n11191 & n11201 ) | ( ~n11358 & n11201 ) ;
  assign n11361 = ( n11359 & ~n11191 ) | ( n11359 & n11360 ) | ( ~n11191 & n11360 ) ;
  assign n11365 = x106 &  n1894 ;
  assign n11362 = ( x108 & ~n1816 ) | ( x108 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n11363 = x107 &  n1811 ;
  assign n11364 = n11362 | n11363 ;
  assign n11366 = ( x106 & ~n11365 ) | ( x106 & n11364 ) | ( ~n11365 & n11364 ) ;
  assign n11367 = ( n1819 & ~n5055 ) | ( n1819 & n11366 ) | ( ~n5055 & n11366 ) ;
  assign n11368 = n5055 | n11367 ;
  assign n11370 = ( x26 & n11366 ) | ( x26 & n11368 ) | ( n11366 & n11368 ) ;
  assign n11369 = ( x26 & ~n11368 ) | ( x26 & n11366 ) | ( ~n11368 & n11366 ) ;
  assign n11371 = ( n11368 & ~n11370 ) | ( n11368 & n11369 ) | ( ~n11370 & n11369 ) ;
  assign n11372 = ( n11052 & n11361 ) | ( n11052 & n11371 ) | ( n11361 & n11371 ) ;
  assign n11373 = ( n11361 & ~n11052 ) | ( n11361 & n11371 ) | ( ~n11052 & n11371 ) ;
  assign n11374 = ( n11052 & ~n11372 ) | ( n11052 & n11373 ) | ( ~n11372 & n11373 ) ;
  assign n11375 = ( n11180 & n11190 ) | ( n11180 & n11374 ) | ( n11190 & n11374 ) ;
  assign n11376 = ( n11190 & ~n11180 ) | ( n11190 & n11374 ) | ( ~n11180 & n11374 ) ;
  assign n11377 = ( n11180 & ~n11375 ) | ( n11180 & n11376 ) | ( ~n11375 & n11376 ) ;
  assign n11378 = ( n11169 & ~n11179 ) | ( n11169 & n11377 ) | ( ~n11179 & n11377 ) ;
  assign n11379 = ( n11169 & ~n11377 ) | ( n11169 & n11179 ) | ( ~n11377 & n11179 ) ;
  assign n11380 = ( n11378 & ~n11169 ) | ( n11378 & n11379 ) | ( ~n11169 & n11379 ) ;
  assign n11381 = ( n11167 & ~n11168 ) | ( n11167 & n11380 ) | ( ~n11168 & n11380 ) ;
  assign n11382 = ( n11167 & ~n11380 ) | ( n11167 & n11168 ) | ( ~n11380 & n11168 ) ;
  assign n11383 = ( n11381 & ~n11167 ) | ( n11381 & n11382 ) | ( ~n11167 & n11382 ) ;
  assign n11385 = ( n11147 & n11157 ) | ( n11147 & n11383 ) | ( n11157 & n11383 ) ;
  assign n11384 = ( n11157 & ~n11147 ) | ( n11157 & n11383 ) | ( ~n11147 & n11383 ) ;
  assign n11386 = ( n11147 & ~n11385 ) | ( n11147 & n11384 ) | ( ~n11385 & n11384 ) ;
  assign n11388 = ( n11136 & n11146 ) | ( n11136 & n11386 ) | ( n11146 & n11386 ) ;
  assign n11387 = ( n11146 & ~n11136 ) | ( n11146 & n11386 ) | ( ~n11136 & n11386 ) ;
  assign n11389 = ( n11136 & ~n11388 ) | ( n11136 & n11387 ) | ( ~n11388 & n11387 ) ;
  assign n11393 = x124 &  n353 ;
  assign n11390 = ( x126 & ~n313 ) | ( x126 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n11391 = x125 &  n308 ;
  assign n11392 = n11390 | n11391 ;
  assign n11394 = ( x124 & ~n11393 ) | ( x124 & n11392 ) | ( ~n11393 & n11392 ) ;
  assign n11395 = ~n316 & n9349 ;
  assign n11396 = ( n316 & ~n11394 ) | ( n316 & n11395 ) | ( ~n11394 & n11395 ) ;
  assign n11397 = x8 &  n11396 ;
  assign n11398 = x8 | n11396 ;
  assign n11399 = ~n11397 & n11398 ;
  assign n11400 = ( n10843 & ~n11095 ) | ( n10843 & n11085 ) | ( ~n11095 & n11085 ) ;
  assign n11401 = ( n11389 & n11399 ) | ( n11389 & n11400 ) | ( n11399 & n11400 ) ;
  assign n11402 = ( n11399 & ~n11389 ) | ( n11399 & n11400 ) | ( ~n11389 & n11400 ) ;
  assign n11403 = ( n11389 & ~n11401 ) | ( n11389 & n11402 ) | ( ~n11401 & n11402 ) ;
  assign n11404 = ( n11127 & ~n11133 ) | ( n11127 & n11403 ) | ( ~n11133 & n11403 ) ;
  assign n11405 = ( n11133 & ~n11127 ) | ( n11133 & n11403 ) | ( ~n11127 & n11403 ) ;
  assign n11406 = ( n11404 & ~n11403 ) | ( n11404 & n11405 ) | ( ~n11403 & n11405 ) ;
  assign n11407 = ( n11121 & ~n11406 ) | ( n11121 & n11125 ) | ( ~n11406 & n11125 ) ;
  assign n11408 = ( n11121 & ~n11125 ) | ( n11121 & n11406 ) | ( ~n11125 & n11406 ) ;
  assign n11409 = ( n11407 & ~n11121 ) | ( n11407 & n11408 ) | ( ~n11121 & n11408 ) ;
  assign n11420 = ( n11136 & ~n11386 ) | ( n11136 & n11146 ) | ( ~n11386 & n11146 ) ;
  assign n11424 = x122 &  n503 ;
  assign n11421 = ( x124 & ~n450 ) | ( x124 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n11422 = x123 &  n445 ;
  assign n11423 = n11421 | n11422 ;
  assign n11425 = ( x122 & ~n11424 ) | ( x122 & n11423 ) | ( ~n11424 & n11423 ) ;
  assign n11426 = ~n453 & n8755 ;
  assign n11427 = n11425 | n11426 ;
  assign n11429 = x11 &  n11427 ;
  assign n11428 = ~x11 & n11427 ;
  assign n11430 = ( x11 & ~n11429 ) | ( x11 & n11428 ) | ( ~n11429 & n11428 ) ;
  assign n11434 = x119 &  n713 ;
  assign n11431 = ( x121 & ~n641 ) | ( x121 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n11432 = x120 &  n636 ;
  assign n11433 = n11431 | n11432 ;
  assign n11435 = ( x119 & ~n11434 ) | ( x119 & n11433 ) | ( ~n11434 & n11433 ) ;
  assign n11436 = ~n644 & n8176 ;
  assign n11437 = n11435 | n11436 ;
  assign n11438 = ( x14 & ~n11437 ) | ( x14 & 1'b0 ) | ( ~n11437 & 1'b0 ) ;
  assign n11439 = ~x14 & n11437 ;
  assign n11440 = n11438 | n11439 ;
  assign n11444 = x116 &  n942 ;
  assign n11441 = ( x118 & ~n896 ) | ( x118 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n11442 = x117 &  n891 ;
  assign n11443 = n11441 | n11442 ;
  assign n11445 = ( x116 & ~n11444 ) | ( x116 & n11443 ) | ( ~n11444 & n11443 ) ;
  assign n11446 = n899 | n7152 ;
  assign n11447 = ~n11445 & n11446 ;
  assign n11448 = x17 &  n11447 ;
  assign n11449 = x17 | n11447 ;
  assign n11450 = ~n11448 & n11449 ;
  assign n11451 = ( n11167 & n11168 ) | ( n11167 & n11380 ) | ( n11168 & n11380 ) ;
  assign n11455 = x113 &  n1227 ;
  assign n11452 = ( x115 & ~n1154 ) | ( x115 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n11453 = x114 &  n1149 ;
  assign n11454 = n11452 | n11453 ;
  assign n11456 = ( x113 & ~n11455 ) | ( x113 & n11454 ) | ( ~n11455 & n11454 ) ;
  assign n11457 = ~n1157 & n6420 ;
  assign n11458 = n11456 | n11457 ;
  assign n11459 = ( x20 & ~n11458 ) | ( x20 & 1'b0 ) | ( ~n11458 & 1'b0 ) ;
  assign n11460 = ~x20 & n11458 ;
  assign n11461 = n11459 | n11460 ;
  assign n11462 = ( n11180 & ~n11190 ) | ( n11180 & n11374 ) | ( ~n11190 & n11374 ) ;
  assign n11466 = x110 &  n1551 ;
  assign n11463 = ( x112 & ~n1451 ) | ( x112 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n11464 = x111 &  n1446 ;
  assign n11465 = n11463 | n11464 ;
  assign n11467 = ( x110 & ~n11466 ) | ( x110 & n11465 ) | ( ~n11466 & n11465 ) ;
  assign n11468 = ~n1454 & n5727 ;
  assign n11469 = n11467 | n11468 ;
  assign n11471 = x23 &  n11469 ;
  assign n11470 = ~x23 & n11469 ;
  assign n11472 = ( x23 & ~n11471 ) | ( x23 & n11470 ) | ( ~n11471 & n11470 ) ;
  assign n11476 = x107 &  n1894 ;
  assign n11473 = ( x109 & ~n1816 ) | ( x109 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n11474 = x108 &  n1811 ;
  assign n11475 = n11473 | n11474 ;
  assign n11477 = ( x107 & ~n11476 ) | ( x107 & n11475 ) | ( ~n11476 & n11475 ) ;
  assign n11478 = ~n1819 & n5267 ;
  assign n11479 = n11477 | n11478 ;
  assign n11480 = ( x26 & ~n11479 ) | ( x26 & 1'b0 ) | ( ~n11479 & 1'b0 ) ;
  assign n11481 = ~x26 & n11479 ;
  assign n11482 = n11480 | n11481 ;
  assign n11483 = ( n11052 & ~n11361 ) | ( n11052 & n11371 ) | ( ~n11361 & n11371 ) ;
  assign n11484 = ( n11191 & n11201 ) | ( n11191 & n11358 ) | ( n11201 & n11358 ) ;
  assign n11488 = x104 &  n2312 ;
  assign n11485 = ( x106 & ~n2195 ) | ( x106 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n11486 = x105 &  n2190 ;
  assign n11487 = n11485 | n11486 ;
  assign n11489 = ( x104 & ~n11488 ) | ( x104 & n11487 ) | ( ~n11488 & n11487 ) ;
  assign n11490 = ~n2198 & n4458 ;
  assign n11491 = n11489 | n11490 ;
  assign n11492 = ( x29 & ~n11491 ) | ( x29 & 1'b0 ) | ( ~n11491 & 1'b0 ) ;
  assign n11493 = ~x29 & n11491 ;
  assign n11494 = n11492 | n11493 ;
  assign n11498 = x101 &  n2718 ;
  assign n11495 = ( x103 & ~n2642 ) | ( x103 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n11496 = x102 &  n2637 ;
  assign n11497 = n11495 | n11496 ;
  assign n11499 = ( x101 & ~n11498 ) | ( x101 & n11497 ) | ( ~n11498 & n11497 ) ;
  assign n11500 = n2645 | n4056 ;
  assign n11501 = ~n11499 & n11500 ;
  assign n11502 = x32 &  n11501 ;
  assign n11503 = x32 | n11501 ;
  assign n11504 = ~n11502 & n11503 ;
  assign n11508 = x89 &  n4934 ;
  assign n11505 = ( x91 & ~n4725 ) | ( x91 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n11506 = x90 &  n4720 ;
  assign n11507 = n11505 | n11506 ;
  assign n11509 = ( x89 & ~n11508 ) | ( x89 & n11507 ) | ( ~n11508 & n11507 ) ;
  assign n11510 = ( n2108 & ~n4728 ) | ( n2108 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n11511 = n11509 | n11510 ;
  assign n11512 = ( x44 & ~n11511 ) | ( x44 & 1'b0 ) | ( ~n11511 & 1'b0 ) ;
  assign n11513 = ~x44 & n11511 ;
  assign n11514 = n11512 | n11513 ;
  assign n11518 = x80 &  n6982 ;
  assign n11515 = ( x82 & ~n6727 ) | ( x82 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n11516 = x81 &  n6722 ;
  assign n11517 = n11515 | n11516 ;
  assign n11519 = ( x80 & ~n11518 ) | ( x80 & n11517 ) | ( ~n11518 & n11517 ) ;
  assign n11520 = ( n1084 & ~n6730 ) | ( n1084 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n11521 = n11519 | n11520 ;
  assign n11522 = ( x53 & ~n11521 ) | ( x53 & 1'b0 ) | ( ~n11521 & 1'b0 ) ;
  assign n11523 = ~x53 & n11521 ;
  assign n11524 = n11522 | n11523 ;
  assign n11528 = x77 &  n7731 ;
  assign n11525 = ( x79 & ~n7538 ) | ( x79 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n11526 = x78 &  n7533 ;
  assign n11527 = n11525 | n11526 ;
  assign n11529 = ( x77 & ~n11528 ) | ( x77 & n11527 ) | ( ~n11528 & n11527 ) ;
  assign n11530 = ( n766 & ~n7541 ) | ( n766 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n11531 = n11529 | n11530 ;
  assign n11532 = ( x56 & ~n11531 ) | ( x56 & 1'b0 ) | ( ~n11531 & 1'b0 ) ;
  assign n11533 = ~x56 & n11531 ;
  assign n11534 = n11532 | n11533 ;
  assign n11538 = x74 &  n8558 ;
  assign n11535 = ( x76 & ~n8314 ) | ( x76 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n11536 = x75 &  n8309 ;
  assign n11537 = n11535 | n11536 ;
  assign n11539 = ( x74 & ~n11538 ) | ( x74 & n11537 ) | ( ~n11538 & n11537 ) ;
  assign n11540 = ( n603 & ~n8317 ) | ( n603 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n11541 = n11539 | n11540 ;
  assign n11542 = ( x59 & ~n11541 ) | ( x59 & 1'b0 ) | ( ~n11541 & 1'b0 ) ;
  assign n11543 = ~x59 & n11541 ;
  assign n11544 = n11542 | n11543 ;
  assign n11545 = ( n10928 & n11222 ) | ( n10928 & n11232 ) | ( n11222 & n11232 ) ;
  assign n11555 = x71 &  n9457 ;
  assign n11552 = ( x73 & ~n9150 ) | ( x73 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n11553 = x72 &  n9145 ;
  assign n11554 = n11552 | n11553 ;
  assign n11556 = ( x71 & ~n11555 ) | ( x71 & n11554 ) | ( ~n11555 & n11554 ) ;
  assign n11557 = ( n389 & ~n9153 ) | ( n389 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n11558 = n11556 | n11557 ;
  assign n11559 = ( x62 & ~n11558 ) | ( x62 & 1'b0 ) | ( ~n11558 & 1'b0 ) ;
  assign n11560 = ~x62 & n11558 ;
  assign n11561 = n11559 | n11560 ;
  assign n11546 = x69 &  n10104 ;
  assign n11547 = ( x70 & ~n9760 ) | ( x70 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n11548 = n11546 | n11547 ;
  assign n11550 = ( x2 & x5 ) | ( x2 & n11548 ) | ( x5 & n11548 ) ;
  assign n11549 = ( x2 & ~x5 ) | ( x2 & n11548 ) | ( ~x5 & n11548 ) ;
  assign n11551 = ( x5 & ~n11550 ) | ( x5 & n11549 ) | ( ~n11550 & n11549 ) ;
  assign n11562 = ( n11220 & ~n11561 ) | ( n11220 & n11551 ) | ( ~n11561 & n11551 ) ;
  assign n11563 = ( n11551 & ~n11220 ) | ( n11551 & n11561 ) | ( ~n11220 & n11561 ) ;
  assign n11564 = ( n11562 & ~n11551 ) | ( n11562 & n11563 ) | ( ~n11551 & n11563 ) ;
  assign n11566 = ( n11544 & n11545 ) | ( n11544 & n11564 ) | ( n11545 & n11564 ) ;
  assign n11565 = ( n11545 & ~n11544 ) | ( n11545 & n11564 ) | ( ~n11544 & n11564 ) ;
  assign n11567 = ( n11544 & ~n11566 ) | ( n11544 & n11565 ) | ( ~n11566 & n11565 ) ;
  assign n11568 = ( n11235 & n11245 ) | ( n11235 & n11249 ) | ( n11245 & n11249 ) ;
  assign n11569 = ( n11534 & ~n11567 ) | ( n11534 & n11568 ) | ( ~n11567 & n11568 ) ;
  assign n11570 = ( n11534 & ~n11568 ) | ( n11534 & n11567 ) | ( ~n11568 & n11567 ) ;
  assign n11571 = ( n11569 & ~n11534 ) | ( n11569 & n11570 ) | ( ~n11534 & n11570 ) ;
  assign n11572 = ( n11206 & n11252 ) | ( n11206 & n11262 ) | ( n11252 & n11262 ) ;
  assign n11573 = ( n11524 & n11571 ) | ( n11524 & n11572 ) | ( n11571 & n11572 ) ;
  assign n11574 = ( n11571 & ~n11524 ) | ( n11571 & n11572 ) | ( ~n11524 & n11572 ) ;
  assign n11575 = ( n11524 & ~n11573 ) | ( n11524 & n11574 ) | ( ~n11573 & n11574 ) ;
  assign n11580 = x83 &  n6288 ;
  assign n11577 = ( x85 & ~n6032 ) | ( x85 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n11578 = x84 &  n6027 ;
  assign n11579 = n11577 | n11578 ;
  assign n11581 = ( x83 & ~n11580 ) | ( x83 & n11579 ) | ( ~n11580 & n11579 ) ;
  assign n11582 = ( n1295 & ~n6035 ) | ( n1295 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n11583 = n11581 | n11582 ;
  assign n11584 = ( x50 & ~n11583 ) | ( x50 & 1'b0 ) | ( ~n11583 & 1'b0 ) ;
  assign n11585 = ~x50 & n11583 ;
  assign n11586 = n11584 | n11585 ;
  assign n11576 = ( n11205 & n11265 ) | ( n11205 & n11275 ) | ( n11265 & n11275 ) ;
  assign n11587 = ( n11575 & ~n11586 ) | ( n11575 & n11576 ) | ( ~n11586 & n11576 ) ;
  assign n11588 = ( n11575 & ~n11576 ) | ( n11575 & n11586 ) | ( ~n11576 & n11586 ) ;
  assign n11589 = ( n11587 & ~n11575 ) | ( n11587 & n11588 ) | ( ~n11575 & n11588 ) ;
  assign n11590 = ( n11278 & n11288 ) | ( n11278 & n11289 ) | ( n11288 & n11289 ) ;
  assign n11594 = x86 &  n5586 ;
  assign n11591 = ( x88 & ~n5389 ) | ( x88 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n11592 = x87 &  n5384 ;
  assign n11593 = n11591 | n11592 ;
  assign n11595 = ( x86 & ~n11594 ) | ( x86 & n11593 ) | ( ~n11594 & n11593 ) ;
  assign n11596 = ( n1624 & ~n5392 ) | ( n1624 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n11597 = n11595 | n11596 ;
  assign n11598 = ( x47 & ~n11597 ) | ( x47 & 1'b0 ) | ( ~n11597 & 1'b0 ) ;
  assign n11599 = ~x47 & n11597 ;
  assign n11600 = n11598 | n11599 ;
  assign n11601 = ( n11589 & ~n11590 ) | ( n11589 & n11600 ) | ( ~n11590 & n11600 ) ;
  assign n11602 = ( n11589 & ~n11600 ) | ( n11589 & n11590 ) | ( ~n11600 & n11590 ) ;
  assign n11603 = ( n11601 & ~n11589 ) | ( n11601 & n11602 ) | ( ~n11589 & n11602 ) ;
  assign n11604 = ( n11204 & n11292 ) | ( n11204 & n11302 ) | ( n11292 & n11302 ) ;
  assign n11605 = ( n11514 & n11603 ) | ( n11514 & n11604 ) | ( n11603 & n11604 ) ;
  assign n11606 = ( n11603 & ~n11514 ) | ( n11603 & n11604 ) | ( ~n11514 & n11604 ) ;
  assign n11607 = ( n11514 & ~n11605 ) | ( n11514 & n11606 ) | ( ~n11605 & n11606 ) ;
  assign n11612 = x92 &  n4344 ;
  assign n11609 = ( x94 & ~n4143 ) | ( x94 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n11610 = x93 &  n4138 ;
  assign n11611 = n11609 | n11610 ;
  assign n11613 = ( x92 & ~n11612 ) | ( x92 & n11611 ) | ( ~n11612 & n11611 ) ;
  assign n11614 = ( n2401 & ~n4146 ) | ( n2401 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n11615 = n11613 | n11614 ;
  assign n11616 = ( x41 & ~n11615 ) | ( x41 & 1'b0 ) | ( ~n11615 & 1'b0 ) ;
  assign n11617 = ~x41 & n11615 ;
  assign n11618 = n11616 | n11617 ;
  assign n11608 = ( n11203 & ~n11315 ) | ( n11203 & n11305 ) | ( ~n11315 & n11305 ) ;
  assign n11619 = ( n11607 & ~n11618 ) | ( n11607 & n11608 ) | ( ~n11618 & n11608 ) ;
  assign n11620 = ( n11607 & ~n11608 ) | ( n11607 & n11618 ) | ( ~n11608 & n11618 ) ;
  assign n11621 = ( n11619 & ~n11607 ) | ( n11619 & n11620 ) | ( ~n11607 & n11620 ) ;
  assign n11622 = ( n11202 & ~n11318 ) | ( n11202 & n11328 ) | ( ~n11318 & n11328 ) ;
  assign n11626 = x95 &  n3756 ;
  assign n11623 = ( x97 & ~n3602 ) | ( x97 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n11624 = x96 &  n3597 ;
  assign n11625 = n11623 | n11624 ;
  assign n11627 = ( x95 & ~n11626 ) | ( x95 & n11625 ) | ( ~n11626 & n11625 ) ;
  assign n11628 = ( n2999 & ~n3605 ) | ( n2999 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n11629 = n11627 | n11628 ;
  assign n11630 = ( x38 & ~n11629 ) | ( x38 & 1'b0 ) | ( ~n11629 & 1'b0 ) ;
  assign n11631 = ~x38 & n11629 ;
  assign n11632 = n11630 | n11631 ;
  assign n11633 = ( n11621 & ~n11622 ) | ( n11621 & n11632 ) | ( ~n11622 & n11632 ) ;
  assign n11634 = ( n11621 & ~n11632 ) | ( n11621 & n11622 ) | ( ~n11632 & n11622 ) ;
  assign n11635 = ( n11633 & ~n11621 ) | ( n11633 & n11634 ) | ( ~n11621 & n11634 ) ;
  assign n11636 = ( n11341 & ~n11331 ) | ( n11341 & n11342 ) | ( ~n11331 & n11342 ) ;
  assign n11640 = x98 &  n3214 ;
  assign n11637 = ( x100 & ~n3087 ) | ( x100 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n11638 = x99 &  n3082 ;
  assign n11639 = n11637 | n11638 ;
  assign n11641 = ( x98 & ~n11640 ) | ( x98 & n11639 ) | ( ~n11640 & n11639 ) ;
  assign n11642 = n3090 | n3354 ;
  assign n11643 = ~n11641 & n11642 ;
  assign n11644 = x35 &  n11643 ;
  assign n11645 = x35 | n11643 ;
  assign n11646 = ~n11644 & n11645 ;
  assign n11648 = ( n11635 & n11636 ) | ( n11635 & n11646 ) | ( n11636 & n11646 ) ;
  assign n11647 = ( n11636 & ~n11635 ) | ( n11636 & n11646 ) | ( ~n11635 & n11646 ) ;
  assign n11649 = ( n11635 & ~n11648 ) | ( n11635 & n11647 ) | ( ~n11648 & n11647 ) ;
  assign n11650 = ( n11345 & ~n11037 ) | ( n11345 & n11355 ) | ( ~n11037 & n11355 ) ;
  assign n11651 = ( n11504 & n11649 ) | ( n11504 & n11650 ) | ( n11649 & n11650 ) ;
  assign n11652 = ( n11649 & ~n11504 ) | ( n11649 & n11650 ) | ( ~n11504 & n11650 ) ;
  assign n11653 = ( n11504 & ~n11651 ) | ( n11504 & n11652 ) | ( ~n11651 & n11652 ) ;
  assign n11654 = ( n11484 & ~n11494 ) | ( n11484 & n11653 ) | ( ~n11494 & n11653 ) ;
  assign n11655 = ( n11484 & ~n11653 ) | ( n11484 & n11494 ) | ( ~n11653 & n11494 ) ;
  assign n11656 = ( n11654 & ~n11484 ) | ( n11654 & n11655 ) | ( ~n11484 & n11655 ) ;
  assign n11657 = ( n11482 & n11483 ) | ( n11482 & n11656 ) | ( n11483 & n11656 ) ;
  assign n11658 = ( n11483 & ~n11482 ) | ( n11483 & n11656 ) | ( ~n11482 & n11656 ) ;
  assign n11659 = ( n11482 & ~n11657 ) | ( n11482 & n11658 ) | ( ~n11657 & n11658 ) ;
  assign n11660 = ( n11462 & ~n11472 ) | ( n11462 & n11659 ) | ( ~n11472 & n11659 ) ;
  assign n11661 = ( n11462 & ~n11659 ) | ( n11462 & n11472 ) | ( ~n11659 & n11472 ) ;
  assign n11662 = ( n11660 & ~n11462 ) | ( n11660 & n11661 ) | ( ~n11462 & n11661 ) ;
  assign n11663 = ( n11169 & n11179 ) | ( n11169 & n11377 ) | ( n11179 & n11377 ) ;
  assign n11665 = ( n11461 & n11662 ) | ( n11461 & n11663 ) | ( n11662 & n11663 ) ;
  assign n11664 = ( n11662 & ~n11461 ) | ( n11662 & n11663 ) | ( ~n11461 & n11663 ) ;
  assign n11666 = ( n11461 & ~n11665 ) | ( n11461 & n11664 ) | ( ~n11665 & n11664 ) ;
  assign n11667 = ( n11450 & ~n11451 ) | ( n11450 & n11666 ) | ( ~n11451 & n11666 ) ;
  assign n11668 = ( n11450 & ~n11666 ) | ( n11450 & n11451 ) | ( ~n11666 & n11451 ) ;
  assign n11669 = ( n11667 & ~n11450 ) | ( n11667 & n11668 ) | ( ~n11450 & n11668 ) ;
  assign n11670 = ( n11147 & ~n11383 ) | ( n11147 & n11157 ) | ( ~n11383 & n11157 ) ;
  assign n11671 = ( n11440 & n11669 ) | ( n11440 & n11670 ) | ( n11669 & n11670 ) ;
  assign n11672 = ( n11669 & ~n11440 ) | ( n11669 & n11670 ) | ( ~n11440 & n11670 ) ;
  assign n11673 = ( n11440 & ~n11671 ) | ( n11440 & n11672 ) | ( ~n11671 & n11672 ) ;
  assign n11675 = ( n11420 & n11430 ) | ( n11420 & n11673 ) | ( n11430 & n11673 ) ;
  assign n11674 = ( n11430 & ~n11420 ) | ( n11430 & n11673 ) | ( ~n11420 & n11673 ) ;
  assign n11676 = ( n11420 & ~n11675 ) | ( n11420 & n11674 ) | ( ~n11675 & n11674 ) ;
  assign n11413 = x125 &  n353 ;
  assign n11410 = ( x127 & ~n313 ) | ( x127 & 1'b0 ) | ( ~n313 & 1'b0 ) ;
  assign n11411 = x126 &  n308 ;
  assign n11412 = n11410 | n11411 ;
  assign n11414 = ( x125 & ~n11413 ) | ( x125 & n11412 ) | ( ~n11413 & n11412 ) ;
  assign n11415 = n316 | n9941 ;
  assign n11416 = ~n11414 & n11415 ;
  assign n11417 = x8 &  n11416 ;
  assign n11418 = x8 | n11416 ;
  assign n11419 = ~n11417 & n11418 ;
  assign n11677 = ( n11401 & n11419 ) | ( n11401 & n11676 ) | ( n11419 & n11676 ) ;
  assign n11678 = ( n11401 & ~n11676 ) | ( n11401 & n11419 ) | ( ~n11676 & n11419 ) ;
  assign n11679 = ( n11676 & ~n11677 ) | ( n11676 & n11678 ) | ( ~n11677 & n11678 ) ;
  assign n11680 = ( n11405 & n11408 ) | ( n11405 & n11679 ) | ( n11408 & n11679 ) ;
  assign n11681 = ( n11408 & ~n11405 ) | ( n11408 & n11679 ) | ( ~n11405 & n11679 ) ;
  assign n11682 = ( n11405 & ~n11680 ) | ( n11405 & n11681 ) | ( ~n11680 & n11681 ) ;
  assign n11683 = ( n11420 & ~n11673 ) | ( n11420 & n11430 ) | ( ~n11673 & n11430 ) ;
  assign n11691 = ( n11440 & ~n11669 ) | ( n11440 & n11670 ) | ( ~n11669 & n11670 ) ;
  assign n11687 = x123 &  n503 ;
  assign n11684 = ( x125 & ~n450 ) | ( x125 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n11685 = x124 &  n445 ;
  assign n11686 = n11684 | n11685 ;
  assign n11688 = ( x123 & ~n11687 ) | ( x123 & n11686 ) | ( ~n11687 & n11686 ) ;
  assign n11689 = ~n453 & n9324 ;
  assign n11690 = n11688 | n11689 ;
  assign n11692 = ( x11 & n11690 ) | ( x11 & n11691 ) | ( n11690 & n11691 ) ;
  assign n11693 = ( x11 & ~n11691 ) | ( x11 & n11690 ) | ( ~n11691 & n11690 ) ;
  assign n11694 = ( n11691 & ~n11692 ) | ( n11691 & n11693 ) | ( ~n11692 & n11693 ) ;
  assign n11695 = ( n11450 & n11451 ) | ( n11450 & n11666 ) | ( n11451 & n11666 ) ;
  assign n11699 = x117 &  n942 ;
  assign n11696 = ( x119 & ~n896 ) | ( x119 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n11697 = x118 &  n891 ;
  assign n11698 = n11696 | n11697 ;
  assign n11700 = ( x117 & ~n11699 ) | ( x117 & n11698 ) | ( ~n11699 & n11698 ) ;
  assign n11701 = ~n899 & n7648 ;
  assign n11702 = n11700 | n11701 ;
  assign n11703 = ( n11461 & ~n11663 ) | ( n11461 & n11662 ) | ( ~n11663 & n11662 ) ;
  assign n11704 = ( x17 & n11702 ) | ( x17 & n11703 ) | ( n11702 & n11703 ) ;
  assign n11705 = ( x17 & ~n11702 ) | ( x17 & n11703 ) | ( ~n11702 & n11703 ) ;
  assign n11706 = ( n11702 & ~n11704 ) | ( n11702 & n11705 ) | ( ~n11704 & n11705 ) ;
  assign n11707 = ( n11462 & n11472 ) | ( n11462 & n11659 ) | ( n11472 & n11659 ) ;
  assign n11711 = x114 &  n1227 ;
  assign n11708 = ( x116 & ~n1154 ) | ( x116 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n11709 = x115 &  n1149 ;
  assign n11710 = n11708 | n11709 ;
  assign n11712 = ( x114 & ~n11711 ) | ( x114 & n11710 ) | ( ~n11711 & n11710 ) ;
  assign n11713 = n1157 | n6885 ;
  assign n11714 = ~n11712 & n11713 ;
  assign n11715 = x20 &  n11714 ;
  assign n11716 = x20 | n11714 ;
  assign n11717 = ~n11715 & n11716 ;
  assign n11721 = x111 &  n1551 ;
  assign n11718 = ( x113 & ~n1451 ) | ( x113 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n11719 = x112 &  n1446 ;
  assign n11720 = n11718 | n11719 ;
  assign n11722 = ( x111 & ~n11721 ) | ( x111 & n11720 ) | ( ~n11721 & n11720 ) ;
  assign n11723 = n1454 | n6169 ;
  assign n11724 = ~n11722 & n11723 ;
  assign n11725 = x23 &  n11724 ;
  assign n11726 = x23 | n11724 ;
  assign n11727 = ~n11725 & n11726 ;
  assign n11731 = x108 &  n1894 ;
  assign n11728 = ( x110 & ~n1816 ) | ( x110 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n11729 = x109 &  n1811 ;
  assign n11730 = n11728 | n11729 ;
  assign n11732 = ( x108 & ~n11731 ) | ( x108 & n11730 ) | ( ~n11731 & n11730 ) ;
  assign n11733 = ~n1819 & n5283 ;
  assign n11734 = ( n1819 & ~n11732 ) | ( n1819 & n11733 ) | ( ~n11732 & n11733 ) ;
  assign n11736 = x26 &  n11734 ;
  assign n11735 = ~x26 & n11734 ;
  assign n11737 = ( x26 & ~n11736 ) | ( x26 & n11735 ) | ( ~n11736 & n11735 ) ;
  assign n11748 = ( n11635 & ~n11646 ) | ( n11635 & n11636 ) | ( ~n11646 & n11636 ) ;
  assign n11759 = ( n11621 & n11622 ) | ( n11621 & n11632 ) | ( n11622 & n11632 ) ;
  assign n11773 = x96 &  n3756 ;
  assign n11770 = ( x98 & ~n3602 ) | ( x98 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n11771 = x97 &  n3597 ;
  assign n11772 = n11770 | n11771 ;
  assign n11774 = ( x96 & ~n11773 ) | ( x96 & n11772 ) | ( ~n11773 & n11772 ) ;
  assign n11775 = ( n3170 & ~n3605 ) | ( n3170 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n11776 = n11774 | n11775 ;
  assign n11777 = ( x38 & ~n11776 ) | ( x38 & 1'b0 ) | ( ~n11776 & 1'b0 ) ;
  assign n11778 = ~x38 & n11776 ;
  assign n11779 = n11777 | n11778 ;
  assign n11780 = ( n11607 & n11608 ) | ( n11607 & n11618 ) | ( n11608 & n11618 ) ;
  assign n11781 = ( n11589 & n11590 ) | ( n11589 & n11600 ) | ( n11590 & n11600 ) ;
  assign n11782 = ( n11575 & n11576 ) | ( n11575 & n11586 ) | ( n11576 & n11586 ) ;
  assign n11783 = ( n11534 & n11567 ) | ( n11534 & n11568 ) | ( n11567 & n11568 ) ;
  assign n11784 = ( n11220 & n11551 ) | ( n11220 & n11561 ) | ( n11551 & n11561 ) ;
  assign n11809 = x59 | n11784 ;
  assign n11810 = ~x59 & n11784 ;
  assign n11811 = ( n11809 & ~n11784 ) | ( n11809 & n11810 ) | ( ~n11784 & n11810 ) ;
  assign n11785 = x70 &  n10104 ;
  assign n11786 = ( x71 & ~n9760 ) | ( x71 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n11787 = n11785 | n11786 ;
  assign n11788 = ( x2 & ~n11548 ) | ( x2 & x5 ) | ( ~n11548 & x5 ) ;
  assign n11792 = x72 &  n9457 ;
  assign n11789 = ( x74 & ~n9150 ) | ( x74 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n11790 = x73 &  n9145 ;
  assign n11791 = n11789 | n11790 ;
  assign n11793 = ( x72 & ~n11792 ) | ( x72 & n11791 ) | ( ~n11792 & n11791 ) ;
  assign n11794 = ( n482 & ~n11793 ) | ( n482 & n9153 ) | ( ~n11793 & n9153 ) ;
  assign n11795 = ~n9153 & n11794 ;
  assign n11796 = ( x62 & n11793 ) | ( x62 & n11795 ) | ( n11793 & n11795 ) ;
  assign n11797 = ( x62 & ~n11795 ) | ( x62 & n11793 ) | ( ~n11795 & n11793 ) ;
  assign n11798 = ( n11795 & ~n11796 ) | ( n11795 & n11797 ) | ( ~n11796 & n11797 ) ;
  assign n11799 = ( n11787 & n11788 ) | ( n11787 & n11798 ) | ( n11788 & n11798 ) ;
  assign n11800 = ( n11788 & ~n11787 ) | ( n11788 & n11798 ) | ( ~n11787 & n11798 ) ;
  assign n11801 = ( n11787 & ~n11799 ) | ( n11787 & n11800 ) | ( ~n11799 & n11800 ) ;
  assign n11805 = x75 &  n8558 ;
  assign n11802 = ( x77 & ~n8314 ) | ( x77 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n11803 = x76 &  n8309 ;
  assign n11804 = n11802 | n11803 ;
  assign n11806 = ( x75 & ~n11805 ) | ( x75 & n11804 ) | ( ~n11805 & n11804 ) ;
  assign n11807 = ( n677 & ~n8317 ) | ( n677 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n11808 = n11806 | n11807 ;
  assign n11813 = ( n11801 & n11808 ) | ( n11801 & n11811 ) | ( n11808 & n11811 ) ;
  assign n11812 = ( n11801 & ~n11811 ) | ( n11801 & n11808 ) | ( ~n11811 & n11808 ) ;
  assign n11814 = ( n11811 & ~n11813 ) | ( n11811 & n11812 ) | ( ~n11813 & n11812 ) ;
  assign n11818 = x78 &  n7731 ;
  assign n11815 = ( x80 & ~n7538 ) | ( x80 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n11816 = x79 &  n7533 ;
  assign n11817 = n11815 | n11816 ;
  assign n11819 = ( x78 & ~n11818 ) | ( x78 & n11817 ) | ( ~n11818 & n11817 ) ;
  assign n11820 = ( n842 & ~n7541 ) | ( n842 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n11821 = n11819 | n11820 ;
  assign n11822 = ( x56 & ~n11821 ) | ( x56 & 1'b0 ) | ( ~n11821 & 1'b0 ) ;
  assign n11823 = ~x56 & n11821 ;
  assign n11824 = n11822 | n11823 ;
  assign n11825 = ( n11566 & ~n11814 ) | ( n11566 & n11824 ) | ( ~n11814 & n11824 ) ;
  assign n11826 = ( n11566 & ~n11824 ) | ( n11566 & n11814 ) | ( ~n11824 & n11814 ) ;
  assign n11827 = ( n11825 & ~n11566 ) | ( n11825 & n11826 ) | ( ~n11566 & n11826 ) ;
  assign n11831 = x81 &  n6982 ;
  assign n11828 = ( x83 & ~n6727 ) | ( x83 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n11829 = x82 &  n6722 ;
  assign n11830 = n11828 | n11829 ;
  assign n11832 = ( x81 & ~n11831 ) | ( x81 & n11830 ) | ( ~n11831 & n11830 ) ;
  assign n11833 = ( n1100 & ~n6730 ) | ( n1100 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n11834 = n11832 | n11833 ;
  assign n11835 = ( x53 & ~n11834 ) | ( x53 & 1'b0 ) | ( ~n11834 & 1'b0 ) ;
  assign n11836 = ~x53 & n11834 ;
  assign n11837 = n11835 | n11836 ;
  assign n11838 = ( n11783 & ~n11827 ) | ( n11783 & n11837 ) | ( ~n11827 & n11837 ) ;
  assign n11839 = ( n11783 & ~n11837 ) | ( n11783 & n11827 ) | ( ~n11837 & n11827 ) ;
  assign n11840 = ( n11838 & ~n11783 ) | ( n11838 & n11839 ) | ( ~n11783 & n11839 ) ;
  assign n11844 = x84 &  n6288 ;
  assign n11841 = ( x86 & ~n6032 ) | ( x86 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n11842 = x85 &  n6027 ;
  assign n11843 = n11841 | n11842 ;
  assign n11845 = ( x84 & ~n11844 ) | ( x84 & n11843 ) | ( ~n11844 & n11843 ) ;
  assign n11846 = ( n1496 & ~n6035 ) | ( n1496 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n11847 = n11845 | n11846 ;
  assign n11848 = ( x50 & ~n11847 ) | ( x50 & 1'b0 ) | ( ~n11847 & 1'b0 ) ;
  assign n11849 = ~x50 & n11847 ;
  assign n11850 = n11848 | n11849 ;
  assign n11851 = ( n11573 & ~n11840 ) | ( n11573 & n11850 ) | ( ~n11840 & n11850 ) ;
  assign n11852 = ( n11573 & ~n11850 ) | ( n11573 & n11840 ) | ( ~n11850 & n11840 ) ;
  assign n11853 = ( n11851 & ~n11573 ) | ( n11851 & n11852 ) | ( ~n11573 & n11852 ) ;
  assign n11857 = x87 &  n5586 ;
  assign n11854 = ( x89 & ~n5389 ) | ( x89 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n11855 = x88 &  n5384 ;
  assign n11856 = n11854 | n11855 ;
  assign n11858 = ( x87 & ~n11857 ) | ( x87 & n11856 ) | ( ~n11857 & n11856 ) ;
  assign n11859 = ( n1741 & ~n5392 ) | ( n1741 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n11860 = n11858 | n11859 ;
  assign n11861 = ( x47 & ~n11860 ) | ( x47 & 1'b0 ) | ( ~n11860 & 1'b0 ) ;
  assign n11862 = ~x47 & n11860 ;
  assign n11863 = n11861 | n11862 ;
  assign n11864 = ( n11782 & ~n11853 ) | ( n11782 & n11863 ) | ( ~n11853 & n11863 ) ;
  assign n11865 = ( n11782 & ~n11863 ) | ( n11782 & n11853 ) | ( ~n11863 & n11853 ) ;
  assign n11866 = ( n11864 & ~n11782 ) | ( n11864 & n11865 ) | ( ~n11782 & n11865 ) ;
  assign n11870 = x90 &  n4934 ;
  assign n11867 = ( x92 & ~n4725 ) | ( x92 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n11868 = x91 &  n4720 ;
  assign n11869 = n11867 | n11868 ;
  assign n11871 = ( x90 & ~n11870 ) | ( x90 & n11869 ) | ( ~n11870 & n11869 ) ;
  assign n11872 = ( n2248 & ~n4728 ) | ( n2248 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n11873 = n11871 | n11872 ;
  assign n11874 = ( x44 & ~n11873 ) | ( x44 & 1'b0 ) | ( ~n11873 & 1'b0 ) ;
  assign n11875 = ~x44 & n11873 ;
  assign n11876 = n11874 | n11875 ;
  assign n11877 = ( n11781 & ~n11866 ) | ( n11781 & n11876 ) | ( ~n11866 & n11876 ) ;
  assign n11878 = ( n11781 & ~n11876 ) | ( n11781 & n11866 ) | ( ~n11876 & n11866 ) ;
  assign n11879 = ( n11877 & ~n11781 ) | ( n11877 & n11878 ) | ( ~n11781 & n11878 ) ;
  assign n11883 = x93 &  n4344 ;
  assign n11880 = ( x95 & ~n4143 ) | ( x95 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n11881 = x94 &  n4138 ;
  assign n11882 = n11880 | n11881 ;
  assign n11884 = ( x93 & ~n11883 ) | ( x93 & n11882 ) | ( ~n11883 & n11882 ) ;
  assign n11885 = ( n2547 & ~n4146 ) | ( n2547 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n11886 = n11884 | n11885 ;
  assign n11887 = ( x41 & ~n11886 ) | ( x41 & 1'b0 ) | ( ~n11886 & 1'b0 ) ;
  assign n11888 = ~x41 & n11886 ;
  assign n11889 = n11887 | n11888 ;
  assign n11890 = ( n11605 & ~n11879 ) | ( n11605 & n11889 ) | ( ~n11879 & n11889 ) ;
  assign n11891 = ( n11605 & ~n11889 ) | ( n11605 & n11879 ) | ( ~n11889 & n11879 ) ;
  assign n11892 = ( n11890 & ~n11605 ) | ( n11890 & n11891 ) | ( ~n11605 & n11891 ) ;
  assign n11894 = ( n11779 & n11780 ) | ( n11779 & n11892 ) | ( n11780 & n11892 ) ;
  assign n11893 = ( n11780 & ~n11779 ) | ( n11780 & n11892 ) | ( ~n11779 & n11892 ) ;
  assign n11895 = ( n11779 & ~n11894 ) | ( n11779 & n11893 ) | ( ~n11894 & n11893 ) ;
  assign n11763 = x99 &  n3214 ;
  assign n11760 = ( x101 & ~n3087 ) | ( x101 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n11761 = x100 &  n3082 ;
  assign n11762 = n11760 | n11761 ;
  assign n11764 = ( x99 & ~n11763 ) | ( x99 & n11762 ) | ( ~n11763 & n11762 ) ;
  assign n11765 = n3090 | n3694 ;
  assign n11766 = ~n11764 & n11765 ;
  assign n11767 = x35 &  n11766 ;
  assign n11768 = x35 | n11766 ;
  assign n11769 = ~n11767 & n11768 ;
  assign n11896 = ( n11759 & ~n11895 ) | ( n11759 & n11769 ) | ( ~n11895 & n11769 ) ;
  assign n11897 = ( n11759 & ~n11769 ) | ( n11759 & n11895 ) | ( ~n11769 & n11895 ) ;
  assign n11898 = ( n11896 & ~n11759 ) | ( n11896 & n11897 ) | ( ~n11759 & n11897 ) ;
  assign n11752 = x102 &  n2718 ;
  assign n11749 = ( x104 & ~n2642 ) | ( x104 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n11750 = x103 &  n2637 ;
  assign n11751 = n11749 | n11750 ;
  assign n11753 = ( x102 & ~n11752 ) | ( x102 & n11751 ) | ( ~n11752 & n11751 ) ;
  assign n11754 = n2645 | n4249 ;
  assign n11755 = ~n11753 & n11754 ;
  assign n11756 = x32 | n11755 ;
  assign n11757 = ( x32 & ~n11755 ) | ( x32 & 1'b0 ) | ( ~n11755 & 1'b0 ) ;
  assign n11758 = ( n11756 & ~x32 ) | ( n11756 & n11757 ) | ( ~x32 & n11757 ) ;
  assign n11899 = ( n11748 & ~n11898 ) | ( n11748 & n11758 ) | ( ~n11898 & n11758 ) ;
  assign n11900 = ( n11748 & ~n11758 ) | ( n11748 & n11898 ) | ( ~n11758 & n11898 ) ;
  assign n11901 = ( n11899 & ~n11748 ) | ( n11899 & n11900 ) | ( ~n11748 & n11900 ) ;
  assign n11741 = x105 &  n2312 ;
  assign n11738 = ( x107 & ~n2195 ) | ( x107 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n11739 = x106 &  n2190 ;
  assign n11740 = n11738 | n11739 ;
  assign n11742 = ( x105 & ~n11741 ) | ( x105 & n11740 ) | ( ~n11741 & n11740 ) ;
  assign n11743 = ~n2198 & n4848 ;
  assign n11744 = n11742 | n11743 ;
  assign n11745 = ( x29 & ~n11744 ) | ( x29 & 1'b0 ) | ( ~n11744 & 1'b0 ) ;
  assign n11746 = ~x29 & n11744 ;
  assign n11747 = n11745 | n11746 ;
  assign n11902 = ( n11651 & ~n11901 ) | ( n11651 & n11747 ) | ( ~n11901 & n11747 ) ;
  assign n11903 = ( n11651 & ~n11747 ) | ( n11651 & n11901 ) | ( ~n11747 & n11901 ) ;
  assign n11904 = ( n11902 & ~n11651 ) | ( n11902 & n11903 ) | ( ~n11651 & n11903 ) ;
  assign n11905 = ( n11655 & n11737 ) | ( n11655 & n11904 ) | ( n11737 & n11904 ) ;
  assign n11906 = ( n11655 & ~n11737 ) | ( n11655 & n11904 ) | ( ~n11737 & n11904 ) ;
  assign n11907 = ( n11737 & ~n11905 ) | ( n11737 & n11906 ) | ( ~n11905 & n11906 ) ;
  assign n11909 = ( n11658 & n11727 ) | ( n11658 & n11907 ) | ( n11727 & n11907 ) ;
  assign n11908 = ( n11727 & ~n11658 ) | ( n11727 & n11907 ) | ( ~n11658 & n11907 ) ;
  assign n11910 = ( n11658 & ~n11909 ) | ( n11658 & n11908 ) | ( ~n11909 & n11908 ) ;
  assign n11911 = ( n11707 & n11717 ) | ( n11707 & n11910 ) | ( n11717 & n11910 ) ;
  assign n11912 = ( n11717 & ~n11707 ) | ( n11717 & n11910 ) | ( ~n11707 & n11910 ) ;
  assign n11913 = ( n11707 & ~n11911 ) | ( n11707 & n11912 ) | ( ~n11911 & n11912 ) ;
  assign n11914 = ( n11706 & ~n11913 ) | ( n11706 & 1'b0 ) | ( ~n11913 & 1'b0 ) ;
  assign n11915 = ~n11706 & n11913 ;
  assign n11916 = n11914 | n11915 ;
  assign n11920 = x120 &  n713 ;
  assign n11917 = ( x122 & ~n641 ) | ( x122 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n11918 = x121 &  n636 ;
  assign n11919 = n11917 | n11918 ;
  assign n11921 = ( x120 & ~n11920 ) | ( x120 & n11919 ) | ( ~n11920 & n11919 ) ;
  assign n11922 = ( n644 & n9987 ) | ( n644 & n11921 ) | ( n9987 & n11921 ) ;
  assign n11923 = ( n9987 & ~n11922 ) | ( n9987 & 1'b0 ) | ( ~n11922 & 1'b0 ) ;
  assign n11924 = ( x14 & n11921 ) | ( x14 & n11923 ) | ( n11921 & n11923 ) ;
  assign n11925 = ( x14 & ~n11923 ) | ( x14 & n11921 ) | ( ~n11923 & n11921 ) ;
  assign n11926 = ( n11923 & ~n11924 ) | ( n11923 & n11925 ) | ( ~n11924 & n11925 ) ;
  assign n11928 = ( n11695 & n11916 ) | ( n11695 & n11926 ) | ( n11916 & n11926 ) ;
  assign n11927 = ( n11916 & ~n11695 ) | ( n11916 & n11926 ) | ( ~n11695 & n11926 ) ;
  assign n11929 = ( n11695 & ~n11928 ) | ( n11695 & n11927 ) | ( ~n11928 & n11927 ) ;
  assign n11930 = n11694 &  n11929 ;
  assign n11931 = n11694 | n11929 ;
  assign n11932 = ~n11930 & n11931 ;
  assign n11933 = ( x126 & ~n353 ) | ( x126 & 1'b0 ) | ( ~n353 & 1'b0 ) ;
  assign n11934 = x127 &  n308 ;
  assign n11935 = n11933 | n11934 ;
  assign n11936 = n316 | n9960 ;
  assign n11937 = ( n11935 & ~n316 ) | ( n11935 & n11936 ) | ( ~n316 & n11936 ) ;
  assign n11938 = x8 | n11937 ;
  assign n11939 = ( x8 & ~n11937 ) | ( x8 & 1'b0 ) | ( ~n11937 & 1'b0 ) ;
  assign n11940 = ( n11938 & ~x8 ) | ( n11938 & n11939 ) | ( ~x8 & n11939 ) ;
  assign n11941 = ( n11683 & ~n11932 ) | ( n11683 & n11940 ) | ( ~n11932 & n11940 ) ;
  assign n11942 = ( n11683 & ~n11940 ) | ( n11683 & n11932 ) | ( ~n11940 & n11932 ) ;
  assign n11943 = ( n11941 & ~n11683 ) | ( n11941 & n11942 ) | ( ~n11683 & n11942 ) ;
  assign n11944 = ( n11405 & ~n11408 ) | ( n11405 & n11679 ) | ( ~n11408 & n11679 ) ;
  assign n11945 = ( n11677 & n11943 ) | ( n11677 & n11944 ) | ( n11943 & n11944 ) ;
  assign n11946 = ( n11943 & ~n11677 ) | ( n11943 & n11944 ) | ( ~n11677 & n11944 ) ;
  assign n11947 = ( n11677 & ~n11945 ) | ( n11677 & n11946 ) | ( ~n11945 & n11946 ) ;
  assign n11948 = ( n11683 & n11932 ) | ( n11683 & n11940 ) | ( n11932 & n11940 ) ;
  assign n11954 = ( x127 & ~n353 ) | ( x127 & 1'b0 ) | ( ~n353 & 1'b0 ) ;
  assign n11955 = n316 | n10258 ;
  assign n11956 = ~n11954 & n11955 ;
  assign n11950 = ( x11 & ~n11690 ) | ( x11 & 1'b0 ) | ( ~n11690 & 1'b0 ) ;
  assign n11951 = ~x11 & n11690 ;
  assign n11952 = n11950 | n11951 ;
  assign n11953 = ( n11691 & n11929 ) | ( n11691 & n11952 ) | ( n11929 & n11952 ) ;
  assign n11957 = ( x8 & ~n11956 ) | ( x8 & n11953 ) | ( ~n11956 & n11953 ) ;
  assign n11958 = ( n11953 & ~x8 ) | ( n11953 & n11956 ) | ( ~x8 & n11956 ) ;
  assign n11959 = ( n11957 & ~n11953 ) | ( n11957 & n11958 ) | ( ~n11953 & n11958 ) ;
  assign n11960 = ( n11695 & ~n11926 ) | ( n11695 & n11916 ) | ( ~n11926 & n11916 ) ;
  assign n11964 = x121 &  n713 ;
  assign n11961 = ( x123 & ~n641 ) | ( x123 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n11962 = x122 &  n636 ;
  assign n11963 = n11961 | n11962 ;
  assign n11965 = ( x121 & ~n11964 ) | ( x121 & n11963 ) | ( ~n11964 & n11963 ) ;
  assign n11966 = ~n644 & n8472 ;
  assign n11967 = n11965 | n11966 ;
  assign n11968 = ( x14 & ~n11967 ) | ( x14 & 1'b0 ) | ( ~n11967 & 1'b0 ) ;
  assign n11969 = ~x14 & n11967 ;
  assign n11970 = n11968 | n11969 ;
  assign n11971 = ( n11707 & ~n11717 ) | ( n11707 & n11910 ) | ( ~n11717 & n11910 ) ;
  assign n11975 = x118 &  n942 ;
  assign n11972 = ( x120 & ~n896 ) | ( x120 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n11973 = x119 &  n891 ;
  assign n11974 = n11972 | n11973 ;
  assign n11976 = ( x118 & ~n11975 ) | ( x118 & n11974 ) | ( ~n11975 & n11974 ) ;
  assign n11977 = ~n899 & n9364 ;
  assign n11978 = n11976 | n11977 ;
  assign n11979 = ( x17 & ~n11978 ) | ( x17 & 1'b0 ) | ( ~n11978 & 1'b0 ) ;
  assign n11980 = ~x17 & n11978 ;
  assign n11981 = n11979 | n11980 ;
  assign n11982 = ( n11658 & ~n11907 ) | ( n11658 & n11727 ) | ( ~n11907 & n11727 ) ;
  assign n11983 = ( n11737 & ~n11655 ) | ( n11737 & n11904 ) | ( ~n11655 & n11904 ) ;
  assign n11987 = x112 &  n1551 ;
  assign n11984 = ( x114 & ~n1451 ) | ( x114 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n11985 = x113 &  n1446 ;
  assign n11986 = n11984 | n11985 ;
  assign n11988 = ( x112 & ~n11987 ) | ( x112 & n11986 ) | ( ~n11987 & n11986 ) ;
  assign n11989 = n1454 | n6185 ;
  assign n11990 = ~n11988 & n11989 ;
  assign n11991 = x23 &  n11990 ;
  assign n11992 = x23 | n11990 ;
  assign n11993 = ~n11991 & n11992 ;
  assign n11994 = ( n11747 & ~n11651 ) | ( n11747 & n11901 ) | ( ~n11651 & n11901 ) ;
  assign n11998 = x109 &  n1894 ;
  assign n11995 = ( x111 & ~n1816 ) | ( x111 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n11996 = x110 &  n1811 ;
  assign n11997 = n11995 | n11996 ;
  assign n11999 = ( x109 & ~n11998 ) | ( x109 & n11997 ) | ( ~n11998 & n11997 ) ;
  assign n12000 = n1819 | n5711 ;
  assign n12001 = ~n11999 & n12000 ;
  assign n12002 = x26 &  n12001 ;
  assign n12003 = x26 | n12001 ;
  assign n12004 = ~n12002 & n12003 ;
  assign n12005 = ( n11758 & ~n11748 ) | ( n11758 & n11898 ) | ( ~n11748 & n11898 ) ;
  assign n12016 = ( n11781 & n11866 ) | ( n11781 & n11876 ) | ( n11866 & n11876 ) ;
  assign n12017 = ( n11782 & n11853 ) | ( n11782 & n11863 ) | ( n11853 & n11863 ) ;
  assign n12018 = ( n11573 & n11840 ) | ( n11573 & n11850 ) | ( n11840 & n11850 ) ;
  assign n12022 = x88 &  n5586 ;
  assign n12019 = ( x90 & ~n5389 ) | ( x90 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n12020 = x89 &  n5384 ;
  assign n12021 = n12019 | n12020 ;
  assign n12023 = ( x88 & ~n12022 ) | ( x88 & n12021 ) | ( ~n12022 & n12021 ) ;
  assign n12024 = ( n1976 & ~n5392 ) | ( n1976 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n12025 = n12023 | n12024 ;
  assign n12026 = ( x47 & ~n12025 ) | ( x47 & 1'b0 ) | ( ~n12025 & 1'b0 ) ;
  assign n12027 = ~x47 & n12025 ;
  assign n12028 = n12026 | n12027 ;
  assign n12029 = ( n11783 & n11827 ) | ( n11783 & n11837 ) | ( n11827 & n11837 ) ;
  assign n12033 = x85 &  n6288 ;
  assign n12030 = ( x87 & ~n6032 ) | ( x87 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n12031 = x86 &  n6027 ;
  assign n12032 = n12030 | n12031 ;
  assign n12034 = ( x85 & ~n12033 ) | ( x85 & n12032 ) | ( ~n12033 & n12032 ) ;
  assign n12035 = ( n1512 & ~n6035 ) | ( n1512 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n12036 = n12034 | n12035 ;
  assign n12037 = ( x50 & ~n12036 ) | ( x50 & 1'b0 ) | ( ~n12036 & 1'b0 ) ;
  assign n12038 = ~x50 & n12036 ;
  assign n12039 = n12037 | n12038 ;
  assign n12040 = ( n11566 & n11814 ) | ( n11566 & n11824 ) | ( n11814 & n11824 ) ;
  assign n12044 = x73 &  n9457 ;
  assign n12041 = ( x75 & ~n9150 ) | ( x75 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n12042 = x74 &  n9145 ;
  assign n12043 = n12041 | n12042 ;
  assign n12045 = ( x73 & ~n12044 ) | ( x73 & n12043 ) | ( ~n12044 & n12043 ) ;
  assign n12046 = ( n540 & ~n9153 ) | ( n540 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n12047 = n12045 | n12046 ;
  assign n12048 = ( x62 & ~n12047 ) | ( x62 & 1'b0 ) | ( ~n12047 & 1'b0 ) ;
  assign n12049 = ~x62 & n12047 ;
  assign n12050 = n12048 | n12049 ;
  assign n12051 = ( n11787 & ~n11798 ) | ( n11787 & n11788 ) | ( ~n11798 & n11788 ) ;
  assign n12052 = x71 &  n10104 ;
  assign n12053 = ( x72 & ~n9760 ) | ( x72 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n12054 = n12052 | n12053 ;
  assign n12056 = ( n11787 & n12051 ) | ( n11787 & n12054 ) | ( n12051 & n12054 ) ;
  assign n12055 = ( n11787 & ~n12051 ) | ( n11787 & n12054 ) | ( ~n12051 & n12054 ) ;
  assign n12057 = ( n12051 & ~n12056 ) | ( n12051 & n12055 ) | ( ~n12056 & n12055 ) ;
  assign n12061 = x76 &  n8558 ;
  assign n12058 = ( x78 & ~n8314 ) | ( x78 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n12059 = x77 &  n8309 ;
  assign n12060 = n12058 | n12059 ;
  assign n12062 = ( x76 & ~n12061 ) | ( x76 & n12060 ) | ( ~n12061 & n12060 ) ;
  assign n12063 = ( n693 & ~n8317 ) | ( n693 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n12064 = n12062 | n12063 ;
  assign n12065 = ( x59 & ~n12064 ) | ( x59 & 1'b0 ) | ( ~n12064 & 1'b0 ) ;
  assign n12066 = ~x59 & n12064 ;
  assign n12067 = n12065 | n12066 ;
  assign n12068 = ( n12050 & ~n12057 ) | ( n12050 & n12067 ) | ( ~n12057 & n12067 ) ;
  assign n12069 = ( n12050 & ~n12067 ) | ( n12050 & n12057 ) | ( ~n12067 & n12057 ) ;
  assign n12070 = ( n12068 & ~n12050 ) | ( n12068 & n12069 ) | ( ~n12050 & n12069 ) ;
  assign n12078 = x79 &  n7731 ;
  assign n12075 = ( x81 & ~n7538 ) | ( x81 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n12076 = x80 &  n7533 ;
  assign n12077 = n12075 | n12076 ;
  assign n12079 = ( x79 & ~n12078 ) | ( x79 & n12077 ) | ( ~n12078 & n12077 ) ;
  assign n12080 = ( n994 & ~n7541 ) | ( n994 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n12081 = n12079 | n12080 ;
  assign n12082 = ( x56 & ~n12081 ) | ( x56 & 1'b0 ) | ( ~n12081 & 1'b0 ) ;
  assign n12083 = ~x56 & n12081 ;
  assign n12084 = n12082 | n12083 ;
  assign n12071 = ( x59 & ~n11808 ) | ( x59 & 1'b0 ) | ( ~n11808 & 1'b0 ) ;
  assign n12072 = ~x59 & n11808 ;
  assign n12073 = n12071 | n12072 ;
  assign n12074 = ( n11784 & n11801 ) | ( n11784 & n12073 ) | ( n11801 & n12073 ) ;
  assign n12085 = ( n12070 & ~n12084 ) | ( n12070 & n12074 ) | ( ~n12084 & n12074 ) ;
  assign n12086 = ( n12070 & ~n12074 ) | ( n12070 & n12084 ) | ( ~n12074 & n12084 ) ;
  assign n12087 = ( n12085 & ~n12070 ) | ( n12085 & n12086 ) | ( ~n12070 & n12086 ) ;
  assign n12091 = x82 &  n6982 ;
  assign n12088 = ( x84 & ~n6727 ) | ( x84 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n12089 = x83 &  n6722 ;
  assign n12090 = n12088 | n12089 ;
  assign n12092 = ( x82 & ~n12091 ) | ( x82 & n12090 ) | ( ~n12091 & n12090 ) ;
  assign n12093 = ( n1199 & ~n6730 ) | ( n1199 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n12094 = n12092 | n12093 ;
  assign n12095 = ( x53 & ~n12094 ) | ( x53 & 1'b0 ) | ( ~n12094 & 1'b0 ) ;
  assign n12096 = ~x53 & n12094 ;
  assign n12097 = n12095 | n12096 ;
  assign n12098 = ( n12040 & ~n12087 ) | ( n12040 & n12097 ) | ( ~n12087 & n12097 ) ;
  assign n12099 = ( n12040 & ~n12097 ) | ( n12040 & n12087 ) | ( ~n12097 & n12087 ) ;
  assign n12100 = ( n12098 & ~n12040 ) | ( n12098 & n12099 ) | ( ~n12040 & n12099 ) ;
  assign n12102 = ( n12029 & n12039 ) | ( n12029 & n12100 ) | ( n12039 & n12100 ) ;
  assign n12101 = ( n12039 & ~n12029 ) | ( n12039 & n12100 ) | ( ~n12029 & n12100 ) ;
  assign n12103 = ( n12029 & ~n12102 ) | ( n12029 & n12101 ) | ( ~n12102 & n12101 ) ;
  assign n12105 = ( n12018 & n12028 ) | ( n12018 & n12103 ) | ( n12028 & n12103 ) ;
  assign n12104 = ( n12028 & ~n12018 ) | ( n12028 & n12103 ) | ( ~n12018 & n12103 ) ;
  assign n12106 = ( n12018 & ~n12105 ) | ( n12018 & n12104 ) | ( ~n12105 & n12104 ) ;
  assign n12110 = x91 &  n4934 ;
  assign n12107 = ( x93 & ~n4725 ) | ( x93 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n12108 = x92 &  n4720 ;
  assign n12109 = n12107 | n12108 ;
  assign n12111 = ( x91 & ~n12110 ) | ( x91 & n12109 ) | ( ~n12110 & n12109 ) ;
  assign n12112 = n2264 | n4728 ;
  assign n12113 = ~n12111 & n12112 ;
  assign n12114 = x44 &  n12113 ;
  assign n12115 = x44 | n12113 ;
  assign n12116 = ~n12114 & n12115 ;
  assign n12118 = ( n12017 & n12106 ) | ( n12017 & n12116 ) | ( n12106 & n12116 ) ;
  assign n12117 = ( n12106 & ~n12017 ) | ( n12106 & n12116 ) | ( ~n12017 & n12116 ) ;
  assign n12119 = ( n12017 & ~n12118 ) | ( n12017 & n12117 ) | ( ~n12118 & n12117 ) ;
  assign n12123 = x94 &  n4344 ;
  assign n12120 = ( x96 & ~n4143 ) | ( x96 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n12121 = x95 &  n4138 ;
  assign n12122 = n12120 | n12121 ;
  assign n12124 = ( x94 & ~n12123 ) | ( x94 & n12122 ) | ( ~n12123 & n12122 ) ;
  assign n12125 = ( n2836 & ~n4146 ) | ( n2836 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n12126 = n12124 | n12125 ;
  assign n12127 = ( x41 & ~n12126 ) | ( x41 & 1'b0 ) | ( ~n12126 & 1'b0 ) ;
  assign n12128 = ~x41 & n12126 ;
  assign n12129 = n12127 | n12128 ;
  assign n12130 = ( n12016 & n12119 ) | ( n12016 & n12129 ) | ( n12119 & n12129 ) ;
  assign n12131 = ( n12119 & ~n12016 ) | ( n12119 & n12129 ) | ( ~n12016 & n12129 ) ;
  assign n12132 = ( n12016 & ~n12130 ) | ( n12016 & n12131 ) | ( ~n12130 & n12131 ) ;
  assign n12136 = x97 &  n3756 ;
  assign n12133 = ( x99 & ~n3602 ) | ( x99 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n12134 = x98 &  n3597 ;
  assign n12135 = n12133 | n12134 ;
  assign n12137 = ( x97 & ~n12136 ) | ( x97 & n12135 ) | ( ~n12136 & n12135 ) ;
  assign n12138 = ( n3338 & ~n3605 ) | ( n3338 & 1'b0 ) | ( ~n3605 & 1'b0 ) ;
  assign n12139 = n12137 | n12138 ;
  assign n12140 = ( x38 & ~n12139 ) | ( x38 & 1'b0 ) | ( ~n12139 & 1'b0 ) ;
  assign n12141 = ~x38 & n12139 ;
  assign n12142 = n12140 | n12141 ;
  assign n12143 = ( n11605 & n11879 ) | ( n11605 & n11889 ) | ( n11879 & n11889 ) ;
  assign n12144 = ( n12132 & ~n12142 ) | ( n12132 & n12143 ) | ( ~n12142 & n12143 ) ;
  assign n12145 = ( n12132 & ~n12143 ) | ( n12132 & n12142 ) | ( ~n12143 & n12142 ) ;
  assign n12146 = ( n12144 & ~n12132 ) | ( n12144 & n12145 ) | ( ~n12132 & n12145 ) ;
  assign n12150 = x100 &  n3214 ;
  assign n12147 = ( x102 & ~n3087 ) | ( x102 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n12148 = x101 &  n3082 ;
  assign n12149 = n12147 | n12148 ;
  assign n12151 = ( x100 & ~n12150 ) | ( x100 & n12149 ) | ( ~n12150 & n12149 ) ;
  assign n12152 = n3090 | n3872 ;
  assign n12153 = ~n12151 & n12152 ;
  assign n12154 = x35 &  n12153 ;
  assign n12155 = x35 | n12153 ;
  assign n12156 = ~n12154 & n12155 ;
  assign n12158 = ( n11894 & n12146 ) | ( n11894 & n12156 ) | ( n12146 & n12156 ) ;
  assign n12157 = ( n11894 & ~n12146 ) | ( n11894 & n12156 ) | ( ~n12146 & n12156 ) ;
  assign n12159 = ( n12146 & ~n12158 ) | ( n12146 & n12157 ) | ( ~n12158 & n12157 ) ;
  assign n12009 = x103 &  n2718 ;
  assign n12006 = ( x105 & ~n2642 ) | ( x105 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n12007 = x104 &  n2637 ;
  assign n12008 = n12006 | n12007 ;
  assign n12010 = ( x103 & ~n12009 ) | ( x103 & n12008 ) | ( ~n12009 & n12008 ) ;
  assign n12011 = ~n2645 & n4442 ;
  assign n12012 = n12010 | n12011 ;
  assign n12013 = ( x32 & ~n12012 ) | ( x32 & 1'b0 ) | ( ~n12012 & 1'b0 ) ;
  assign n12014 = ~x32 & n12012 ;
  assign n12015 = n12013 | n12014 ;
  assign n12160 = ( n11897 & ~n12159 ) | ( n11897 & n12015 ) | ( ~n12159 & n12015 ) ;
  assign n12161 = ( n12015 & ~n11897 ) | ( n12015 & n12159 ) | ( ~n11897 & n12159 ) ;
  assign n12162 = ( n12160 & ~n12015 ) | ( n12160 & n12161 ) | ( ~n12015 & n12161 ) ;
  assign n12166 = x106 &  n2312 ;
  assign n12163 = ( x108 & ~n2195 ) | ( x108 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n12164 = x107 &  n2190 ;
  assign n12165 = n12163 | n12164 ;
  assign n12167 = ( x106 & ~n12166 ) | ( x106 & n12165 ) | ( ~n12166 & n12165 ) ;
  assign n12168 = ( n2198 & ~n5055 ) | ( n2198 & n12167 ) | ( ~n5055 & n12167 ) ;
  assign n12169 = n5055 | n12168 ;
  assign n12171 = ( x29 & n12167 ) | ( x29 & n12169 ) | ( n12167 & n12169 ) ;
  assign n12170 = ( x29 & ~n12169 ) | ( x29 & n12167 ) | ( ~n12169 & n12167 ) ;
  assign n12172 = ( n12169 & ~n12171 ) | ( n12169 & n12170 ) | ( ~n12171 & n12170 ) ;
  assign n12173 = ( n12005 & n12162 ) | ( n12005 & n12172 ) | ( n12162 & n12172 ) ;
  assign n12174 = ( n12162 & ~n12005 ) | ( n12162 & n12172 ) | ( ~n12005 & n12172 ) ;
  assign n12175 = ( n12005 & ~n12173 ) | ( n12005 & n12174 ) | ( ~n12173 & n12174 ) ;
  assign n12176 = ( n11994 & n12004 ) | ( n11994 & n12175 ) | ( n12004 & n12175 ) ;
  assign n12177 = ( n12004 & ~n11994 ) | ( n12004 & n12175 ) | ( ~n11994 & n12175 ) ;
  assign n12178 = ( n11994 & ~n12176 ) | ( n11994 & n12177 ) | ( ~n12176 & n12177 ) ;
  assign n12179 = ( n11983 & ~n11993 ) | ( n11983 & n12178 ) | ( ~n11993 & n12178 ) ;
  assign n12180 = ( n11983 & ~n12178 ) | ( n11983 & n11993 ) | ( ~n12178 & n11993 ) ;
  assign n12181 = ( n12179 & ~n11983 ) | ( n12179 & n12180 ) | ( ~n11983 & n12180 ) ;
  assign n12185 = x115 &  n1227 ;
  assign n12182 = ( x117 & ~n1154 ) | ( x117 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n12183 = x116 &  n1149 ;
  assign n12184 = n12182 | n12183 ;
  assign n12186 = ( x115 & ~n12185 ) | ( x115 & n12184 ) | ( ~n12185 & n12184 ) ;
  assign n12187 = ( n1157 & ~n7136 ) | ( n1157 & n12186 ) | ( ~n7136 & n12186 ) ;
  assign n12188 = n7136 | n12187 ;
  assign n12190 = ( x20 & n12186 ) | ( x20 & n12188 ) | ( n12186 & n12188 ) ;
  assign n12189 = ( x20 & ~n12188 ) | ( x20 & n12186 ) | ( ~n12188 & n12186 ) ;
  assign n12191 = ( n12188 & ~n12190 ) | ( n12188 & n12189 ) | ( ~n12190 & n12189 ) ;
  assign n12192 = ( n11982 & n12181 ) | ( n11982 & n12191 ) | ( n12181 & n12191 ) ;
  assign n12193 = ( n12181 & ~n11982 ) | ( n12181 & n12191 ) | ( ~n11982 & n12191 ) ;
  assign n12194 = ( n11982 & ~n12192 ) | ( n11982 & n12193 ) | ( ~n12192 & n12193 ) ;
  assign n12196 = ( n11971 & n11981 ) | ( n11971 & n12194 ) | ( n11981 & n12194 ) ;
  assign n12195 = ( n11981 & ~n11971 ) | ( n11981 & n12194 ) | ( ~n11971 & n12194 ) ;
  assign n12197 = ( n11971 & ~n12196 ) | ( n11971 & n12195 ) | ( ~n12196 & n12195 ) ;
  assign n12198 = x17 &  n11702 ;
  assign n12199 = ( n11704 & ~n12198 ) | ( n11704 & n11914 ) | ( ~n12198 & n11914 ) ;
  assign n12200 = ( n11970 & n12197 ) | ( n11970 & n12199 ) | ( n12197 & n12199 ) ;
  assign n12201 = ( n12197 & ~n11970 ) | ( n12197 & n12199 ) | ( ~n11970 & n12199 ) ;
  assign n12202 = ( n11970 & ~n12200 ) | ( n11970 & n12201 ) | ( ~n12200 & n12201 ) ;
  assign n12206 = x124 &  n503 ;
  assign n12203 = ( x126 & ~n450 ) | ( x126 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n12204 = x125 &  n445 ;
  assign n12205 = n12203 | n12204 ;
  assign n12207 = ( x124 & ~n12206 ) | ( x124 & n12205 ) | ( ~n12206 & n12205 ) ;
  assign n12208 = ( n453 & ~n9349 ) | ( n453 & n12207 ) | ( ~n9349 & n12207 ) ;
  assign n12209 = n9349 | n12208 ;
  assign n12211 = ( x11 & n12207 ) | ( x11 & n12209 ) | ( n12207 & n12209 ) ;
  assign n12210 = ( x11 & ~n12209 ) | ( x11 & n12207 ) | ( ~n12209 & n12207 ) ;
  assign n12212 = ( n12209 & ~n12211 ) | ( n12209 & n12210 ) | ( ~n12211 & n12210 ) ;
  assign n12213 = ( n11960 & ~n12202 ) | ( n11960 & n12212 ) | ( ~n12202 & n12212 ) ;
  assign n12214 = ( n11960 & ~n12212 ) | ( n11960 & n12202 ) | ( ~n12212 & n12202 ) ;
  assign n12215 = ( n12213 & ~n11960 ) | ( n12213 & n12214 ) | ( ~n11960 & n12214 ) ;
  assign n12216 = n11959 | n12215 ;
  assign n12217 = n11959 &  n12215 ;
  assign n12218 = ( n12216 & ~n12217 ) | ( n12216 & 1'b0 ) | ( ~n12217 & 1'b0 ) ;
  assign n11949 = ( n11677 & ~n11943 ) | ( n11677 & n11944 ) | ( ~n11943 & n11944 ) ;
  assign n12219 = ( n11948 & ~n12218 ) | ( n11948 & n11949 ) | ( ~n12218 & n11949 ) ;
  assign n12220 = ( n11948 & ~n11949 ) | ( n11948 & n12218 ) | ( ~n11949 & n12218 ) ;
  assign n12221 = ( n12219 & ~n11948 ) | ( n12219 & n12220 ) | ( ~n11948 & n12220 ) ;
  assign n12222 = ~x8 & n11956 ;
  assign n12223 = ( n12216 & ~n11958 ) | ( n12216 & n12222 ) | ( ~n11958 & n12222 ) ;
  assign n12227 = x125 &  n503 ;
  assign n12224 = ( x127 & ~n450 ) | ( x127 & 1'b0 ) | ( ~n450 & 1'b0 ) ;
  assign n12225 = x126 &  n445 ;
  assign n12226 = n12224 | n12225 ;
  assign n12228 = ( x125 & ~n12227 ) | ( x125 & n12226 ) | ( ~n12227 & n12226 ) ;
  assign n12229 = n453 | n9941 ;
  assign n12230 = ~n12228 & n12229 ;
  assign n12231 = x11 &  n12230 ;
  assign n12232 = x11 | n12230 ;
  assign n12233 = ~n12231 & n12232 ;
  assign n12234 = ( n11960 & n12202 ) | ( n11960 & n12212 ) | ( n12202 & n12212 ) ;
  assign n12235 = ( n11970 & ~n12197 ) | ( n11970 & n12199 ) | ( ~n12197 & n12199 ) ;
  assign n12239 = x119 &  n942 ;
  assign n12236 = ( x121 & ~n896 ) | ( x121 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n12237 = x120 &  n891 ;
  assign n12238 = n12236 | n12237 ;
  assign n12240 = ( x119 & ~n12239 ) | ( x119 & n12238 ) | ( ~n12239 & n12238 ) ;
  assign n12241 = ~n899 & n8176 ;
  assign n12242 = n12240 | n12241 ;
  assign n12457 = x17 | n12242 ;
  assign n12458 = ~x17 & n12242 ;
  assign n12459 = ( n12457 & ~n12242 ) | ( n12457 & n12458 ) | ( ~n12242 & n12458 ) ;
  assign n12243 = ( n11971 & ~n12194 ) | ( n11971 & n11981 ) | ( ~n12194 & n11981 ) ;
  assign n12247 = x116 &  n1227 ;
  assign n12244 = ( x118 & ~n1154 ) | ( x118 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n12245 = x117 &  n1149 ;
  assign n12246 = n12244 | n12245 ;
  assign n12248 = ( x116 & ~n12247 ) | ( x116 & n12246 ) | ( ~n12247 & n12246 ) ;
  assign n12249 = n1157 | n7152 ;
  assign n12250 = ~n12248 & n12249 ;
  assign n12251 = x20 &  n12250 ;
  assign n12252 = x20 | n12250 ;
  assign n12253 = ~n12251 & n12252 ;
  assign n12257 = x113 &  n1551 ;
  assign n12254 = ( x115 & ~n1451 ) | ( x115 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n12255 = x114 &  n1446 ;
  assign n12256 = n12254 | n12255 ;
  assign n12258 = ( x113 & ~n12257 ) | ( x113 & n12256 ) | ( ~n12257 & n12256 ) ;
  assign n12259 = ~n1454 & n6420 ;
  assign n12260 = n12258 | n12259 ;
  assign n12261 = ( x23 & ~n12260 ) | ( x23 & 1'b0 ) | ( ~n12260 & 1'b0 ) ;
  assign n12262 = ~x23 & n12260 ;
  assign n12263 = n12261 | n12262 ;
  assign n12264 = ( n11994 & ~n12004 ) | ( n11994 & n12175 ) | ( ~n12004 & n12175 ) ;
  assign n12268 = x110 &  n1894 ;
  assign n12265 = ( x112 & ~n1816 ) | ( x112 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n12266 = x111 &  n1811 ;
  assign n12267 = n12265 | n12266 ;
  assign n12269 = ( x110 & ~n12268 ) | ( x110 & n12267 ) | ( ~n12268 & n12267 ) ;
  assign n12270 = ~n1819 & n5727 ;
  assign n12271 = n12269 | n12270 ;
  assign n12272 = ( x26 & ~n12271 ) | ( x26 & 1'b0 ) | ( ~n12271 & 1'b0 ) ;
  assign n12273 = ~x26 & n12271 ;
  assign n12274 = n12272 | n12273 ;
  assign n12278 = x107 &  n2312 ;
  assign n12275 = ( x109 & ~n2195 ) | ( x109 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n12276 = x108 &  n2190 ;
  assign n12277 = n12275 | n12276 ;
  assign n12279 = ( x107 & ~n12278 ) | ( x107 & n12277 ) | ( ~n12278 & n12277 ) ;
  assign n12280 = ~n2198 & n5267 ;
  assign n12281 = n12279 | n12280 ;
  assign n12282 = ( x29 & ~n12281 ) | ( x29 & 1'b0 ) | ( ~n12281 & 1'b0 ) ;
  assign n12283 = ~x29 & n12281 ;
  assign n12284 = n12282 | n12283 ;
  assign n12289 = x104 &  n2718 ;
  assign n12286 = ( x106 & ~n2642 ) | ( x106 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n12287 = x105 &  n2637 ;
  assign n12288 = n12286 | n12287 ;
  assign n12290 = ( x104 & ~n12289 ) | ( x104 & n12288 ) | ( ~n12289 & n12288 ) ;
  assign n12291 = ~n2645 & n4458 ;
  assign n12292 = n12290 | n12291 ;
  assign n12293 = ( x32 & ~n12292 ) | ( x32 & 1'b0 ) | ( ~n12292 & 1'b0 ) ;
  assign n12294 = ~x32 & n12292 ;
  assign n12295 = n12293 | n12294 ;
  assign n12296 = ( n11897 & n12015 ) | ( n11897 & n12159 ) | ( n12015 & n12159 ) ;
  assign n12300 = x101 &  n3214 ;
  assign n12297 = ( x103 & ~n3087 ) | ( x103 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n12298 = x102 &  n3082 ;
  assign n12299 = n12297 | n12298 ;
  assign n12301 = ( x101 & ~n12300 ) | ( x101 & n12299 ) | ( ~n12300 & n12299 ) ;
  assign n12302 = n3090 | n4056 ;
  assign n12303 = ~n12301 & n12302 ;
  assign n12304 = x35 &  n12303 ;
  assign n12305 = x35 | n12303 ;
  assign n12306 = ~n12304 & n12305 ;
  assign n12320 = x86 &  n6288 ;
  assign n12317 = ( x88 & ~n6032 ) | ( x88 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n12318 = x87 &  n6027 ;
  assign n12319 = n12317 | n12318 ;
  assign n12321 = ( x86 & ~n12320 ) | ( x86 & n12319 ) | ( ~n12320 & n12319 ) ;
  assign n12322 = ( n1624 & ~n6035 ) | ( n1624 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n12323 = n12321 | n12322 ;
  assign n12324 = ( x50 & ~n12323 ) | ( x50 & 1'b0 ) | ( ~n12323 & 1'b0 ) ;
  assign n12325 = ~x50 & n12323 ;
  assign n12326 = n12324 | n12325 ;
  assign n12330 = x83 &  n6982 ;
  assign n12327 = ( x85 & ~n6727 ) | ( x85 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n12328 = x84 &  n6722 ;
  assign n12329 = n12327 | n12328 ;
  assign n12331 = ( x83 & ~n12330 ) | ( x83 & n12329 ) | ( ~n12330 & n12329 ) ;
  assign n12332 = ( n1295 & ~n6730 ) | ( n1295 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n12333 = n12331 | n12332 ;
  assign n12334 = ( x53 & ~n12333 ) | ( x53 & 1'b0 ) | ( ~n12333 & 1'b0 ) ;
  assign n12335 = ~x53 & n12333 ;
  assign n12336 = n12334 | n12335 ;
  assign n12340 = x74 &  n9457 ;
  assign n12337 = ( x76 & ~n9150 ) | ( x76 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n12338 = x75 &  n9145 ;
  assign n12339 = n12337 | n12338 ;
  assign n12341 = ( x74 & ~n12340 ) | ( x74 & n12339 ) | ( ~n12340 & n12339 ) ;
  assign n12342 = ( n603 & ~n9153 ) | ( n603 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n12343 = n12341 | n12342 ;
  assign n12344 = ( x62 & ~n12343 ) | ( x62 & 1'b0 ) | ( ~n12343 & 1'b0 ) ;
  assign n12345 = ~x62 & n12343 ;
  assign n12346 = n12344 | n12345 ;
  assign n12347 = ( n12051 & ~n11787 ) | ( n12051 & n12054 ) | ( ~n11787 & n12054 ) ;
  assign n12348 = x72 &  n10104 ;
  assign n12349 = ( x73 & ~n9760 ) | ( x73 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n12350 = n12348 | n12349 ;
  assign n12351 = ( x8 & n12054 ) | ( x8 & n12350 ) | ( n12054 & n12350 ) ;
  assign n12352 = ( x8 & ~n12054 ) | ( x8 & n12350 ) | ( ~n12054 & n12350 ) ;
  assign n12353 = ( n12054 & ~n12351 ) | ( n12054 & n12352 ) | ( ~n12351 & n12352 ) ;
  assign n12354 = ( n12346 & n12347 ) | ( n12346 & n12353 ) | ( n12347 & n12353 ) ;
  assign n12355 = ( n12347 & ~n12346 ) | ( n12347 & n12353 ) | ( ~n12346 & n12353 ) ;
  assign n12356 = ( n12346 & ~n12354 ) | ( n12346 & n12355 ) | ( ~n12354 & n12355 ) ;
  assign n12357 = ( n12050 & n12057 ) | ( n12050 & n12067 ) | ( n12057 & n12067 ) ;
  assign n12361 = x77 &  n8558 ;
  assign n12358 = ( x79 & ~n8314 ) | ( x79 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n12359 = x78 &  n8309 ;
  assign n12360 = n12358 | n12359 ;
  assign n12362 = ( x77 & ~n12361 ) | ( x77 & n12360 ) | ( ~n12361 & n12360 ) ;
  assign n12363 = ( n766 & ~n8317 ) | ( n766 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n12364 = n12362 | n12363 ;
  assign n12365 = ( x59 & ~n12364 ) | ( x59 & 1'b0 ) | ( ~n12364 & 1'b0 ) ;
  assign n12366 = ~x59 & n12364 ;
  assign n12367 = n12365 | n12366 ;
  assign n12368 = ( n12356 & ~n12357 ) | ( n12356 & n12367 ) | ( ~n12357 & n12367 ) ;
  assign n12369 = ( n12356 & ~n12367 ) | ( n12356 & n12357 ) | ( ~n12367 & n12357 ) ;
  assign n12370 = ( n12368 & ~n12356 ) | ( n12368 & n12369 ) | ( ~n12356 & n12369 ) ;
  assign n12381 = ( n12070 & n12074 ) | ( n12070 & n12084 ) | ( n12074 & n12084 ) ;
  assign n12374 = x80 &  n7731 ;
  assign n12371 = ( x82 & ~n7538 ) | ( x82 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n12372 = x81 &  n7533 ;
  assign n12373 = n12371 | n12372 ;
  assign n12375 = ( x80 & ~n12374 ) | ( x80 & n12373 ) | ( ~n12374 & n12373 ) ;
  assign n12376 = ( n1084 & ~n7541 ) | ( n1084 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n12377 = n12375 | n12376 ;
  assign n12378 = ( x56 & ~n12377 ) | ( x56 & 1'b0 ) | ( ~n12377 & 1'b0 ) ;
  assign n12379 = ~x56 & n12377 ;
  assign n12380 = n12378 | n12379 ;
  assign n12382 = ( n12370 & ~n12381 ) | ( n12370 & n12380 ) | ( ~n12381 & n12380 ) ;
  assign n12383 = ( n12370 & ~n12380 ) | ( n12370 & n12381 ) | ( ~n12380 & n12381 ) ;
  assign n12384 = ( n12382 & ~n12370 ) | ( n12382 & n12383 ) | ( ~n12370 & n12383 ) ;
  assign n12385 = ( n12040 & n12087 ) | ( n12040 & n12097 ) | ( n12087 & n12097 ) ;
  assign n12386 = ( n12336 & n12384 ) | ( n12336 & n12385 ) | ( n12384 & n12385 ) ;
  assign n12387 = ( n12384 & ~n12336 ) | ( n12384 & n12385 ) | ( ~n12336 & n12385 ) ;
  assign n12388 = ( n12336 & ~n12386 ) | ( n12336 & n12387 ) | ( ~n12386 & n12387 ) ;
  assign n12390 = ( n12102 & n12326 ) | ( n12102 & n12388 ) | ( n12326 & n12388 ) ;
  assign n12389 = ( n12102 & ~n12326 ) | ( n12102 & n12388 ) | ( ~n12326 & n12388 ) ;
  assign n12391 = ( n12326 & ~n12390 ) | ( n12326 & n12389 ) | ( ~n12390 & n12389 ) ;
  assign n12310 = x89 &  n5586 ;
  assign n12307 = ( x91 & ~n5389 ) | ( x91 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n12308 = x90 &  n5384 ;
  assign n12309 = n12307 | n12308 ;
  assign n12311 = ( x89 & ~n12310 ) | ( x89 & n12309 ) | ( ~n12310 & n12309 ) ;
  assign n12312 = ( n2108 & ~n5392 ) | ( n2108 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n12313 = n12311 | n12312 ;
  assign n12314 = ( x47 & ~n12313 ) | ( x47 & 1'b0 ) | ( ~n12313 & 1'b0 ) ;
  assign n12315 = ~x47 & n12313 ;
  assign n12316 = n12314 | n12315 ;
  assign n12392 = ( n12105 & ~n12391 ) | ( n12105 & n12316 ) | ( ~n12391 & n12316 ) ;
  assign n12393 = ( n12316 & ~n12105 ) | ( n12316 & n12391 ) | ( ~n12105 & n12391 ) ;
  assign n12394 = ( n12392 & ~n12316 ) | ( n12392 & n12393 ) | ( ~n12316 & n12393 ) ;
  assign n12399 = x92 &  n4934 ;
  assign n12396 = ( x94 & ~n4725 ) | ( x94 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n12397 = x93 &  n4720 ;
  assign n12398 = n12396 | n12397 ;
  assign n12400 = ( x92 & ~n12399 ) | ( x92 & n12398 ) | ( ~n12399 & n12398 ) ;
  assign n12401 = ( n2401 & ~n4728 ) | ( n2401 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n12402 = n12400 | n12401 ;
  assign n12403 = ( x44 & ~n12402 ) | ( x44 & 1'b0 ) | ( ~n12402 & 1'b0 ) ;
  assign n12404 = ~x44 & n12402 ;
  assign n12405 = n12403 | n12404 ;
  assign n12395 = ( n12017 & ~n12116 ) | ( n12017 & n12106 ) | ( ~n12116 & n12106 ) ;
  assign n12406 = ( n12394 & ~n12405 ) | ( n12394 & n12395 ) | ( ~n12405 & n12395 ) ;
  assign n12407 = ( n12394 & ~n12395 ) | ( n12394 & n12405 ) | ( ~n12395 & n12405 ) ;
  assign n12408 = ( n12406 & ~n12394 ) | ( n12406 & n12407 ) | ( ~n12394 & n12407 ) ;
  assign n12409 = ( n12016 & ~n12119 ) | ( n12016 & n12129 ) | ( ~n12119 & n12129 ) ;
  assign n12413 = x95 &  n4344 ;
  assign n12410 = ( x97 & ~n4143 ) | ( x97 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n12411 = x96 &  n4138 ;
  assign n12412 = n12410 | n12411 ;
  assign n12414 = ( x95 & ~n12413 ) | ( x95 & n12412 ) | ( ~n12413 & n12412 ) ;
  assign n12415 = ( n2999 & ~n4146 ) | ( n2999 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n12416 = n12414 | n12415 ;
  assign n12417 = ( x41 & ~n12416 ) | ( x41 & 1'b0 ) | ( ~n12416 & 1'b0 ) ;
  assign n12418 = ~x41 & n12416 ;
  assign n12419 = n12417 | n12418 ;
  assign n12420 = ( n12408 & ~n12409 ) | ( n12408 & n12419 ) | ( ~n12409 & n12419 ) ;
  assign n12421 = ( n12408 & ~n12419 ) | ( n12408 & n12409 ) | ( ~n12419 & n12409 ) ;
  assign n12422 = ( n12420 & ~n12408 ) | ( n12420 & n12421 ) | ( ~n12408 & n12421 ) ;
  assign n12423 = ( n12142 & ~n12132 ) | ( n12142 & n12143 ) | ( ~n12132 & n12143 ) ;
  assign n12427 = x98 &  n3756 ;
  assign n12424 = ( x100 & ~n3602 ) | ( x100 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n12425 = x99 &  n3597 ;
  assign n12426 = n12424 | n12425 ;
  assign n12428 = ( x98 & ~n12427 ) | ( x98 & n12426 ) | ( ~n12427 & n12426 ) ;
  assign n12429 = n3354 | n3605 ;
  assign n12430 = ~n12428 & n12429 ;
  assign n12431 = x38 &  n12430 ;
  assign n12432 = x38 | n12430 ;
  assign n12433 = ~n12431 & n12432 ;
  assign n12435 = ( n12422 & n12423 ) | ( n12422 & n12433 ) | ( n12423 & n12433 ) ;
  assign n12434 = ( n12423 & ~n12422 ) | ( n12423 & n12433 ) | ( ~n12422 & n12433 ) ;
  assign n12436 = ( n12422 & ~n12435 ) | ( n12422 & n12434 ) | ( ~n12435 & n12434 ) ;
  assign n12437 = ( n12146 & ~n11894 ) | ( n12146 & n12156 ) | ( ~n11894 & n12156 ) ;
  assign n12438 = ( n12306 & n12436 ) | ( n12306 & n12437 ) | ( n12436 & n12437 ) ;
  assign n12439 = ( n12436 & ~n12306 ) | ( n12436 & n12437 ) | ( ~n12306 & n12437 ) ;
  assign n12440 = ( n12306 & ~n12438 ) | ( n12306 & n12439 ) | ( ~n12438 & n12439 ) ;
  assign n12442 = ( n12295 & n12296 ) | ( n12295 & n12440 ) | ( n12296 & n12440 ) ;
  assign n12441 = ( n12296 & ~n12295 ) | ( n12296 & n12440 ) | ( ~n12295 & n12440 ) ;
  assign n12443 = ( n12295 & ~n12442 ) | ( n12295 & n12441 ) | ( ~n12442 & n12441 ) ;
  assign n12285 = ( n12005 & ~n12162 ) | ( n12005 & n12172 ) | ( ~n12162 & n12172 ) ;
  assign n12444 = ( n12284 & ~n12443 ) | ( n12284 & n12285 ) | ( ~n12443 & n12285 ) ;
  assign n12445 = ( n12284 & ~n12285 ) | ( n12284 & n12443 ) | ( ~n12285 & n12443 ) ;
  assign n12446 = ( n12444 & ~n12284 ) | ( n12444 & n12445 ) | ( ~n12284 & n12445 ) ;
  assign n12447 = ( n12264 & ~n12274 ) | ( n12264 & n12446 ) | ( ~n12274 & n12446 ) ;
  assign n12448 = ( n12264 & ~n12446 ) | ( n12264 & n12274 ) | ( ~n12446 & n12274 ) ;
  assign n12449 = ( n12447 & ~n12264 ) | ( n12447 & n12448 ) | ( ~n12264 & n12448 ) ;
  assign n12450 = ( n11983 & n11993 ) | ( n11983 & n12178 ) | ( n11993 & n12178 ) ;
  assign n12452 = ( n12263 & n12449 ) | ( n12263 & n12450 ) | ( n12449 & n12450 ) ;
  assign n12451 = ( n12449 & ~n12263 ) | ( n12449 & n12450 ) | ( ~n12263 & n12450 ) ;
  assign n12453 = ( n12263 & ~n12452 ) | ( n12263 & n12451 ) | ( ~n12452 & n12451 ) ;
  assign n12454 = ( n12253 & ~n12192 ) | ( n12253 & n12453 ) | ( ~n12192 & n12453 ) ;
  assign n12455 = ( n12192 & ~n12453 ) | ( n12192 & n12253 ) | ( ~n12453 & n12253 ) ;
  assign n12456 = ( n12454 & ~n12253 ) | ( n12454 & n12455 ) | ( ~n12253 & n12455 ) ;
  assign n12461 = ( n12243 & n12456 ) | ( n12243 & n12459 ) | ( n12456 & n12459 ) ;
  assign n12460 = ( n12243 & ~n12459 ) | ( n12243 & n12456 ) | ( ~n12459 & n12456 ) ;
  assign n12462 = ( n12459 & ~n12461 ) | ( n12459 & n12460 ) | ( ~n12461 & n12460 ) ;
  assign n12466 = x122 &  n713 ;
  assign n12463 = ( x124 & ~n641 ) | ( x124 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n12464 = x123 &  n636 ;
  assign n12465 = n12463 | n12464 ;
  assign n12467 = ( x122 & ~n12466 ) | ( x122 & n12465 ) | ( ~n12466 & n12465 ) ;
  assign n12468 = ~n644 & n8755 ;
  assign n12469 = n12467 | n12468 ;
  assign n12470 = ( x14 & ~n12469 ) | ( x14 & 1'b0 ) | ( ~n12469 & 1'b0 ) ;
  assign n12471 = ~x14 & n12469 ;
  assign n12472 = n12470 | n12471 ;
  assign n12473 = ( n12235 & n12462 ) | ( n12235 & n12472 ) | ( n12462 & n12472 ) ;
  assign n12474 = ( n12462 & ~n12235 ) | ( n12462 & n12472 ) | ( ~n12235 & n12472 ) ;
  assign n12475 = ( n12235 & ~n12473 ) | ( n12235 & n12474 ) | ( ~n12473 & n12474 ) ;
  assign n12476 = ( n12233 & ~n12234 ) | ( n12233 & n12475 ) | ( ~n12234 & n12475 ) ;
  assign n12477 = ( n12233 & ~n12475 ) | ( n12233 & n12234 ) | ( ~n12475 & n12234 ) ;
  assign n12478 = ( n12476 & ~n12233 ) | ( n12476 & n12477 ) | ( ~n12233 & n12477 ) ;
  assign n12479 = ( n12220 & n12223 ) | ( n12220 & n12478 ) | ( n12223 & n12478 ) ;
  assign n12480 = ( n12220 & ~n12223 ) | ( n12220 & n12478 ) | ( ~n12223 & n12478 ) ;
  assign n12481 = ( n12223 & ~n12479 ) | ( n12223 & n12480 ) | ( ~n12479 & n12480 ) ;
  assign n12482 = ( n12233 & n12234 ) | ( n12233 & n12475 ) | ( n12234 & n12475 ) ;
  assign n12483 = ( n12223 & ~n12220 ) | ( n12223 & n12478 ) | ( ~n12220 & n12478 ) ;
  assign n12484 = ( n12235 & ~n12462 ) | ( n12235 & n12472 ) | ( ~n12462 & n12472 ) ;
  assign n12485 = ( x17 & ~n12242 ) | ( x17 & 1'b0 ) | ( ~n12242 & 1'b0 ) ;
  assign n12486 = n12458 | n12485 ;
  assign n12487 = ( n12243 & ~n12456 ) | ( n12243 & n12486 ) | ( ~n12456 & n12486 ) ;
  assign n12491 = x123 &  n713 ;
  assign n12488 = ( x125 & ~n641 ) | ( x125 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n12489 = x124 &  n636 ;
  assign n12490 = n12488 | n12489 ;
  assign n12492 = ( x123 & ~n12491 ) | ( x123 & n12490 ) | ( ~n12491 & n12490 ) ;
  assign n12493 = ~n644 & n9324 ;
  assign n12494 = n12492 | n12493 ;
  assign n12496 = x14 &  n12494 ;
  assign n12495 = ~x14 & n12494 ;
  assign n12497 = ( x14 & ~n12496 ) | ( x14 & n12495 ) | ( ~n12496 & n12495 ) ;
  assign n12498 = ( n12192 & n12253 ) | ( n12192 & n12453 ) | ( n12253 & n12453 ) ;
  assign n12502 = x117 &  n1227 ;
  assign n12499 = ( x119 & ~n1154 ) | ( x119 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n12500 = x118 &  n1149 ;
  assign n12501 = n12499 | n12500 ;
  assign n12503 = ( x117 & ~n12502 ) | ( x117 & n12501 ) | ( ~n12502 & n12501 ) ;
  assign n12504 = ~n1157 & n7648 ;
  assign n12505 = n12503 | n12504 ;
  assign n12506 = ( x20 & ~n12505 ) | ( x20 & 1'b0 ) | ( ~n12505 & 1'b0 ) ;
  assign n12507 = ~x20 & n12505 ;
  assign n12508 = n12506 | n12507 ;
  assign n12512 = x114 &  n1551 ;
  assign n12509 = ( x116 & ~n1451 ) | ( x116 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n12510 = x115 &  n1446 ;
  assign n12511 = n12509 | n12510 ;
  assign n12513 = ( x114 & ~n12512 ) | ( x114 & n12511 ) | ( ~n12512 & n12511 ) ;
  assign n12514 = n1454 | n6885 ;
  assign n12515 = ~n12513 & n12514 ;
  assign n12516 = ( n12264 & n12274 ) | ( n12264 & n12446 ) | ( n12274 & n12446 ) ;
  assign n12518 = ( x23 & n12515 ) | ( x23 & n12516 ) | ( n12515 & n12516 ) ;
  assign n12517 = ( x23 & ~n12515 ) | ( x23 & n12516 ) | ( ~n12515 & n12516 ) ;
  assign n12519 = ( n12515 & ~n12518 ) | ( n12515 & n12517 ) | ( ~n12518 & n12517 ) ;
  assign n12520 = ( n12285 & ~n12284 ) | ( n12285 & n12443 ) | ( ~n12284 & n12443 ) ;
  assign n12524 = x111 &  n1894 ;
  assign n12521 = ( x113 & ~n1816 ) | ( x113 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n12522 = x112 &  n1811 ;
  assign n12523 = n12521 | n12522 ;
  assign n12525 = ( x111 & ~n12524 ) | ( x111 & n12523 ) | ( ~n12524 & n12523 ) ;
  assign n12526 = n1819 | n6169 ;
  assign n12527 = ~n12525 & n12526 ;
  assign n12528 = x26 | n12527 ;
  assign n12529 = ( x26 & ~n12527 ) | ( x26 & 1'b0 ) | ( ~n12527 & 1'b0 ) ;
  assign n12530 = ( n12528 & ~x26 ) | ( n12528 & n12529 ) | ( ~x26 & n12529 ) ;
  assign n12531 = ( n12295 & ~n12440 ) | ( n12295 & n12296 ) | ( ~n12440 & n12296 ) ;
  assign n12688 = x108 &  n2312 ;
  assign n12685 = ( x110 & ~n2195 ) | ( x110 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n12686 = x109 &  n2190 ;
  assign n12687 = n12685 | n12686 ;
  assign n12689 = ( x108 & ~n12688 ) | ( x108 & n12687 ) | ( ~n12688 & n12687 ) ;
  assign n12690 = ( n2198 & ~n5283 ) | ( n2198 & n12689 ) | ( ~n5283 & n12689 ) ;
  assign n12691 = n5283 | n12690 ;
  assign n12693 = ( x29 & n12689 ) | ( x29 & n12691 ) | ( n12689 & n12691 ) ;
  assign n12692 = ( x29 & ~n12691 ) | ( x29 & n12689 ) | ( ~n12691 & n12689 ) ;
  assign n12694 = ( n12691 & ~n12693 ) | ( n12691 & n12692 ) | ( ~n12693 & n12692 ) ;
  assign n12542 = ( n12422 & ~n12433 ) | ( n12422 & n12423 ) | ( ~n12433 & n12423 ) ;
  assign n12546 = x102 &  n3214 ;
  assign n12543 = ( x104 & ~n3087 ) | ( x104 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n12544 = x103 &  n3082 ;
  assign n12545 = n12543 | n12544 ;
  assign n12547 = ( x102 & ~n12546 ) | ( x102 & n12545 ) | ( ~n12546 & n12545 ) ;
  assign n12548 = n3090 | n4249 ;
  assign n12549 = ~n12547 & n12548 ;
  assign n12550 = x35 &  n12549 ;
  assign n12551 = x35 | n12549 ;
  assign n12552 = ~n12550 & n12551 ;
  assign n12553 = ( n12408 & n12409 ) | ( n12408 & n12419 ) | ( n12409 & n12419 ) ;
  assign n12567 = x96 &  n4344 ;
  assign n12564 = ( x98 & ~n4143 ) | ( x98 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n12565 = x97 &  n4138 ;
  assign n12566 = n12564 | n12565 ;
  assign n12568 = ( x96 & ~n12567 ) | ( x96 & n12566 ) | ( ~n12567 & n12566 ) ;
  assign n12569 = ( n3170 & ~n4146 ) | ( n3170 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n12570 = n12568 | n12569 ;
  assign n12571 = ( x41 & ~n12570 ) | ( x41 & 1'b0 ) | ( ~n12570 & 1'b0 ) ;
  assign n12572 = ~x41 & n12570 ;
  assign n12573 = n12571 | n12572 ;
  assign n12574 = ( n12394 & n12395 ) | ( n12394 & n12405 ) | ( n12395 & n12405 ) ;
  assign n12575 = ( n12105 & n12316 ) | ( n12105 & n12391 ) | ( n12316 & n12391 ) ;
  assign n12576 = ( n12370 & n12380 ) | ( n12370 & n12381 ) | ( n12380 & n12381 ) ;
  assign n12577 = ( n12356 & n12357 ) | ( n12356 & n12367 ) | ( n12357 & n12367 ) ;
  assign n12578 = ( n12054 & ~x8 ) | ( n12054 & n12350 ) | ( ~x8 & n12350 ) ;
  assign n12582 = x75 &  n9457 ;
  assign n12579 = ( x77 & ~n9150 ) | ( x77 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n12580 = x76 &  n9145 ;
  assign n12581 = n12579 | n12580 ;
  assign n12583 = ( x75 & ~n12582 ) | ( x75 & n12581 ) | ( ~n12582 & n12581 ) ;
  assign n12584 = ( n677 & ~n9153 ) | ( n677 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n12585 = n12583 | n12584 ;
  assign n12586 = ( x62 & ~n12585 ) | ( x62 & 1'b0 ) | ( ~n12585 & 1'b0 ) ;
  assign n12587 = ~x62 & n12585 ;
  assign n12588 = n12586 | n12587 ;
  assign n12589 = x73 &  n10104 ;
  assign n12590 = ( x74 & ~n9760 ) | ( x74 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n12591 = n12589 | n12590 ;
  assign n12592 = ( n12578 & ~n12588 ) | ( n12578 & n12591 ) | ( ~n12588 & n12591 ) ;
  assign n12593 = ( n12588 & ~n12578 ) | ( n12588 & n12591 ) | ( ~n12578 & n12591 ) ;
  assign n12594 = ( n12592 & ~n12591 ) | ( n12592 & n12593 ) | ( ~n12591 & n12593 ) ;
  assign n12598 = x78 &  n8558 ;
  assign n12595 = ( x80 & ~n8314 ) | ( x80 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n12596 = x79 &  n8309 ;
  assign n12597 = n12595 | n12596 ;
  assign n12599 = ( x78 & ~n12598 ) | ( x78 & n12597 ) | ( ~n12598 & n12597 ) ;
  assign n12600 = ( n842 & ~n8317 ) | ( n842 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n12601 = n12599 | n12600 ;
  assign n12602 = ( x59 & ~n12601 ) | ( x59 & 1'b0 ) | ( ~n12601 & 1'b0 ) ;
  assign n12603 = ~x59 & n12601 ;
  assign n12604 = n12602 | n12603 ;
  assign n12606 = ( n12355 & n12594 ) | ( n12355 & n12604 ) | ( n12594 & n12604 ) ;
  assign n12605 = ( n12594 & ~n12355 ) | ( n12594 & n12604 ) | ( ~n12355 & n12604 ) ;
  assign n12607 = ( n12355 & ~n12606 ) | ( n12355 & n12605 ) | ( ~n12606 & n12605 ) ;
  assign n12611 = x81 &  n7731 ;
  assign n12608 = ( x83 & ~n7538 ) | ( x83 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n12609 = x82 &  n7533 ;
  assign n12610 = n12608 | n12609 ;
  assign n12612 = ( x81 & ~n12611 ) | ( x81 & n12610 ) | ( ~n12611 & n12610 ) ;
  assign n12613 = ( n1100 & ~n7541 ) | ( n1100 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n12614 = n12612 | n12613 ;
  assign n12615 = ( x56 & ~n12614 ) | ( x56 & 1'b0 ) | ( ~n12614 & 1'b0 ) ;
  assign n12616 = ~x56 & n12614 ;
  assign n12617 = n12615 | n12616 ;
  assign n12618 = ( n12577 & ~n12607 ) | ( n12577 & n12617 ) | ( ~n12607 & n12617 ) ;
  assign n12619 = ( n12577 & ~n12617 ) | ( n12577 & n12607 ) | ( ~n12617 & n12607 ) ;
  assign n12620 = ( n12618 & ~n12577 ) | ( n12618 & n12619 ) | ( ~n12577 & n12619 ) ;
  assign n12624 = x84 &  n6982 ;
  assign n12621 = ( x86 & ~n6727 ) | ( x86 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n12622 = x85 &  n6722 ;
  assign n12623 = n12621 | n12622 ;
  assign n12625 = ( x84 & ~n12624 ) | ( x84 & n12623 ) | ( ~n12624 & n12623 ) ;
  assign n12626 = ( n1496 & ~n6730 ) | ( n1496 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n12627 = n12625 | n12626 ;
  assign n12628 = ( x53 & ~n12627 ) | ( x53 & 1'b0 ) | ( ~n12627 & 1'b0 ) ;
  assign n12629 = ~x53 & n12627 ;
  assign n12630 = n12628 | n12629 ;
  assign n12631 = ( n12576 & ~n12620 ) | ( n12576 & n12630 ) | ( ~n12620 & n12630 ) ;
  assign n12632 = ( n12576 & ~n12630 ) | ( n12576 & n12620 ) | ( ~n12630 & n12620 ) ;
  assign n12633 = ( n12631 & ~n12576 ) | ( n12631 & n12632 ) | ( ~n12576 & n12632 ) ;
  assign n12637 = x87 &  n6288 ;
  assign n12634 = ( x89 & ~n6032 ) | ( x89 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n12635 = x88 &  n6027 ;
  assign n12636 = n12634 | n12635 ;
  assign n12638 = ( x87 & ~n12637 ) | ( x87 & n12636 ) | ( ~n12637 & n12636 ) ;
  assign n12639 = ( n1741 & ~n6035 ) | ( n1741 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n12640 = n12638 | n12639 ;
  assign n12641 = ( x50 & ~n12640 ) | ( x50 & 1'b0 ) | ( ~n12640 & 1'b0 ) ;
  assign n12642 = ~x50 & n12640 ;
  assign n12643 = n12641 | n12642 ;
  assign n12644 = ( n12386 & ~n12633 ) | ( n12386 & n12643 ) | ( ~n12633 & n12643 ) ;
  assign n12645 = ( n12386 & ~n12643 ) | ( n12386 & n12633 ) | ( ~n12643 & n12633 ) ;
  assign n12646 = ( n12644 & ~n12386 ) | ( n12644 & n12645 ) | ( ~n12386 & n12645 ) ;
  assign n12650 = x90 &  n5586 ;
  assign n12647 = ( x92 & ~n5389 ) | ( x92 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n12648 = x91 &  n5384 ;
  assign n12649 = n12647 | n12648 ;
  assign n12651 = ( x90 & ~n12650 ) | ( x90 & n12649 ) | ( ~n12650 & n12649 ) ;
  assign n12652 = ( n2248 & ~n5392 ) | ( n2248 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n12653 = n12651 | n12652 ;
  assign n12654 = ( x47 & ~n12653 ) | ( x47 & 1'b0 ) | ( ~n12653 & 1'b0 ) ;
  assign n12655 = ~x47 & n12653 ;
  assign n12656 = n12654 | n12655 ;
  assign n12657 = ( n12390 & ~n12646 ) | ( n12390 & n12656 ) | ( ~n12646 & n12656 ) ;
  assign n12658 = ( n12390 & ~n12656 ) | ( n12390 & n12646 ) | ( ~n12656 & n12646 ) ;
  assign n12659 = ( n12657 & ~n12390 ) | ( n12657 & n12658 ) | ( ~n12390 & n12658 ) ;
  assign n12663 = x93 &  n4934 ;
  assign n12660 = ( x95 & ~n4725 ) | ( x95 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n12661 = x94 &  n4720 ;
  assign n12662 = n12660 | n12661 ;
  assign n12664 = ( x93 & ~n12663 ) | ( x93 & n12662 ) | ( ~n12663 & n12662 ) ;
  assign n12665 = ( n2547 & ~n4728 ) | ( n2547 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n12666 = n12664 | n12665 ;
  assign n12667 = ( x44 & ~n12666 ) | ( x44 & 1'b0 ) | ( ~n12666 & 1'b0 ) ;
  assign n12668 = ~x44 & n12666 ;
  assign n12669 = n12667 | n12668 ;
  assign n12670 = ( n12575 & ~n12659 ) | ( n12575 & n12669 ) | ( ~n12659 & n12669 ) ;
  assign n12671 = ( n12575 & ~n12669 ) | ( n12575 & n12659 ) | ( ~n12669 & n12659 ) ;
  assign n12672 = ( n12670 & ~n12575 ) | ( n12670 & n12671 ) | ( ~n12575 & n12671 ) ;
  assign n12674 = ( n12573 & n12574 ) | ( n12573 & n12672 ) | ( n12574 & n12672 ) ;
  assign n12673 = ( n12574 & ~n12573 ) | ( n12574 & n12672 ) | ( ~n12573 & n12672 ) ;
  assign n12675 = ( n12573 & ~n12674 ) | ( n12573 & n12673 ) | ( ~n12674 & n12673 ) ;
  assign n12557 = x99 &  n3756 ;
  assign n12554 = ( x101 & ~n3602 ) | ( x101 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n12555 = x100 &  n3597 ;
  assign n12556 = n12554 | n12555 ;
  assign n12558 = ( x99 & ~n12557 ) | ( x99 & n12556 ) | ( ~n12557 & n12556 ) ;
  assign n12559 = n3605 | n3694 ;
  assign n12560 = ~n12558 & n12559 ;
  assign n12561 = x38 &  n12560 ;
  assign n12562 = x38 | n12560 ;
  assign n12563 = ~n12561 & n12562 ;
  assign n12676 = ( n12553 & ~n12675 ) | ( n12553 & n12563 ) | ( ~n12675 & n12563 ) ;
  assign n12677 = ( n12553 & ~n12563 ) | ( n12553 & n12675 ) | ( ~n12563 & n12675 ) ;
  assign n12678 = ( n12676 & ~n12553 ) | ( n12676 & n12677 ) | ( ~n12553 & n12677 ) ;
  assign n12679 = ( n12542 & n12552 ) | ( n12542 & n12678 ) | ( n12552 & n12678 ) ;
  assign n12680 = ( n12552 & ~n12542 ) | ( n12552 & n12678 ) | ( ~n12542 & n12678 ) ;
  assign n12681 = ( n12542 & ~n12679 ) | ( n12542 & n12680 ) | ( ~n12679 & n12680 ) ;
  assign n12535 = x105 &  n2718 ;
  assign n12532 = ( x107 & ~n2642 ) | ( x107 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n12533 = x106 &  n2637 ;
  assign n12534 = n12532 | n12533 ;
  assign n12536 = ( x105 & ~n12535 ) | ( x105 & n12534 ) | ( ~n12535 & n12534 ) ;
  assign n12537 = ~n2645 & n4848 ;
  assign n12538 = n12536 | n12537 ;
  assign n12539 = ( x32 & ~n12538 ) | ( x32 & 1'b0 ) | ( ~n12538 & 1'b0 ) ;
  assign n12540 = ~x32 & n12538 ;
  assign n12541 = n12539 | n12540 ;
  assign n12682 = ( n12438 & ~n12681 ) | ( n12438 & n12541 ) | ( ~n12681 & n12541 ) ;
  assign n12683 = ( n12438 & ~n12541 ) | ( n12438 & n12681 ) | ( ~n12541 & n12681 ) ;
  assign n12684 = ( n12682 & ~n12438 ) | ( n12682 & n12683 ) | ( ~n12438 & n12683 ) ;
  assign n12695 = ( n12531 & ~n12694 ) | ( n12531 & n12684 ) | ( ~n12694 & n12684 ) ;
  assign n12696 = ( n12531 & ~n12684 ) | ( n12531 & n12694 ) | ( ~n12684 & n12694 ) ;
  assign n12697 = ( n12695 & ~n12531 ) | ( n12695 & n12696 ) | ( ~n12531 & n12696 ) ;
  assign n12699 = ( n12520 & n12530 ) | ( n12520 & n12697 ) | ( n12530 & n12697 ) ;
  assign n12698 = ( n12530 & ~n12520 ) | ( n12530 & n12697 ) | ( ~n12520 & n12697 ) ;
  assign n12700 = ( n12520 & ~n12699 ) | ( n12520 & n12698 ) | ( ~n12699 & n12698 ) ;
  assign n12701 = ~n12519 & n12700 ;
  assign n12702 = ( n12519 & ~n12700 ) | ( n12519 & 1'b0 ) | ( ~n12700 & 1'b0 ) ;
  assign n12703 = n12701 | n12702 ;
  assign n12704 = ( n12263 & ~n12450 ) | ( n12263 & n12449 ) | ( ~n12450 & n12449 ) ;
  assign n12705 = ( n12508 & n12703 ) | ( n12508 & n12704 ) | ( n12703 & n12704 ) ;
  assign n12706 = ( n12703 & ~n12508 ) | ( n12703 & n12704 ) | ( ~n12508 & n12704 ) ;
  assign n12707 = ( n12508 & ~n12705 ) | ( n12508 & n12706 ) | ( ~n12705 & n12706 ) ;
  assign n12711 = x120 &  n942 ;
  assign n12708 = ( x122 & ~n896 ) | ( x122 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n12709 = x121 &  n891 ;
  assign n12710 = n12708 | n12709 ;
  assign n12712 = ( x120 & ~n12711 ) | ( x120 & n12710 ) | ( ~n12711 & n12710 ) ;
  assign n12713 = ( n899 & n9987 ) | ( n899 & n12712 ) | ( n9987 & n12712 ) ;
  assign n12714 = ( n9987 & ~n12713 ) | ( n9987 & 1'b0 ) | ( ~n12713 & 1'b0 ) ;
  assign n12715 = ( x17 & n12712 ) | ( x17 & n12714 ) | ( n12712 & n12714 ) ;
  assign n12716 = ( x17 & ~n12714 ) | ( x17 & n12712 ) | ( ~n12714 & n12712 ) ;
  assign n12717 = ( n12714 & ~n12715 ) | ( n12714 & n12716 ) | ( ~n12715 & n12716 ) ;
  assign n12719 = ( n12498 & n12707 ) | ( n12498 & n12717 ) | ( n12707 & n12717 ) ;
  assign n12718 = ( n12707 & ~n12498 ) | ( n12707 & n12717 ) | ( ~n12498 & n12717 ) ;
  assign n12720 = ( n12498 & ~n12719 ) | ( n12498 & n12718 ) | ( ~n12719 & n12718 ) ;
  assign n12721 = ( n12487 & ~n12497 ) | ( n12487 & n12720 ) | ( ~n12497 & n12720 ) ;
  assign n12722 = ( n12487 & ~n12720 ) | ( n12487 & n12497 ) | ( ~n12720 & n12497 ) ;
  assign n12723 = ( n12721 & ~n12487 ) | ( n12721 & n12722 ) | ( ~n12487 & n12722 ) ;
  assign n12724 = ( x126 & ~n503 ) | ( x126 & 1'b0 ) | ( ~n503 & 1'b0 ) ;
  assign n12725 = x127 &  n445 ;
  assign n12726 = n12724 | n12725 ;
  assign n12727 = n453 | n9960 ;
  assign n12728 = ( n12726 & ~n453 ) | ( n12726 & n12727 ) | ( ~n453 & n12727 ) ;
  assign n12729 = x11 | n12728 ;
  assign n12730 = ( x11 & ~n12728 ) | ( x11 & 1'b0 ) | ( ~n12728 & 1'b0 ) ;
  assign n12731 = ( n12729 & ~x11 ) | ( n12729 & n12730 ) | ( ~x11 & n12730 ) ;
  assign n12732 = ( n12484 & ~n12723 ) | ( n12484 & n12731 ) | ( ~n12723 & n12731 ) ;
  assign n12733 = ( n12484 & ~n12731 ) | ( n12484 & n12723 ) | ( ~n12731 & n12723 ) ;
  assign n12734 = ( n12732 & ~n12484 ) | ( n12732 & n12733 ) | ( ~n12484 & n12733 ) ;
  assign n12735 = ( n12482 & ~n12483 ) | ( n12482 & n12734 ) | ( ~n12483 & n12734 ) ;
  assign n12736 = ( n12482 & ~n12734 ) | ( n12482 & n12483 ) | ( ~n12734 & n12483 ) ;
  assign n12737 = ( n12735 & ~n12482 ) | ( n12735 & n12736 ) | ( ~n12482 & n12736 ) ;
  assign n12738 = ( n12484 & n12723 ) | ( n12484 & n12731 ) | ( n12723 & n12731 ) ;
  assign n12739 = ( x127 & ~n503 ) | ( x127 & 1'b0 ) | ( ~n503 & 1'b0 ) ;
  assign n12740 = n453 | n10258 ;
  assign n12741 = ~n12739 & n12740 ;
  assign n12742 = ~x11 & n12741 ;
  assign n12743 = ( x11 & ~n12741 ) | ( x11 & 1'b0 ) | ( ~n12741 & 1'b0 ) ;
  assign n12744 = n12742 | n12743 ;
  assign n12745 = ( n12487 & n12497 ) | ( n12487 & n12720 ) | ( n12497 & n12720 ) ;
  assign n12746 = ( n12498 & ~n12717 ) | ( n12498 & n12707 ) | ( ~n12717 & n12707 ) ;
  assign n12750 = x121 &  n942 ;
  assign n12747 = ( x123 & ~n896 ) | ( x123 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n12748 = x122 &  n891 ;
  assign n12749 = n12747 | n12748 ;
  assign n12751 = ( x121 & ~n12750 ) | ( x121 & n12749 ) | ( ~n12750 & n12749 ) ;
  assign n12752 = ~n899 & n8472 ;
  assign n12753 = n12751 | n12752 ;
  assign n12754 = ( n12508 & ~n12703 ) | ( n12508 & n12704 ) | ( ~n12703 & n12704 ) ;
  assign n12755 = ( x17 & n12753 ) | ( x17 & n12754 ) | ( n12753 & n12754 ) ;
  assign n12756 = ( x17 & ~n12753 ) | ( x17 & n12754 ) | ( ~n12753 & n12754 ) ;
  assign n12757 = ( n12753 & ~n12755 ) | ( n12753 & n12756 ) | ( ~n12755 & n12756 ) ;
  assign n12758 = ( x23 & ~n12515 ) | ( x23 & 1'b0 ) | ( ~n12515 & 1'b0 ) ;
  assign n12759 = ( n12517 & ~n12758 ) | ( n12517 & n12701 ) | ( ~n12758 & n12701 ) ;
  assign n12763 = x118 &  n1227 ;
  assign n12760 = ( x120 & ~n1154 ) | ( x120 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n12761 = x119 &  n1149 ;
  assign n12762 = n12760 | n12761 ;
  assign n12764 = ( x118 & ~n12763 ) | ( x118 & n12762 ) | ( ~n12763 & n12762 ) ;
  assign n12765 = ~n1157 & n9364 ;
  assign n12766 = n12764 | n12765 ;
  assign n12767 = ( x20 & ~n12766 ) | ( x20 & 1'b0 ) | ( ~n12766 & 1'b0 ) ;
  assign n12768 = ~x20 & n12766 ;
  assign n12769 = n12767 | n12768 ;
  assign n12770 = ( n12520 & ~n12697 ) | ( n12520 & n12530 ) | ( ~n12697 & n12530 ) ;
  assign n12771 = ( n12684 & ~n12531 ) | ( n12684 & n12694 ) | ( ~n12531 & n12694 ) ;
  assign n12775 = x109 &  n2312 ;
  assign n12772 = ( x111 & ~n2195 ) | ( x111 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n12773 = x110 &  n2190 ;
  assign n12774 = n12772 | n12773 ;
  assign n12776 = ( x109 & ~n12775 ) | ( x109 & n12774 ) | ( ~n12775 & n12774 ) ;
  assign n12777 = n2198 | n5711 ;
  assign n12778 = ~n12776 & n12777 ;
  assign n12779 = ( n12541 & ~n12438 ) | ( n12541 & n12681 ) | ( ~n12438 & n12681 ) ;
  assign n12781 = ( x29 & n12778 ) | ( x29 & n12779 ) | ( n12778 & n12779 ) ;
  assign n12780 = ( x29 & ~n12778 ) | ( x29 & n12779 ) | ( ~n12778 & n12779 ) ;
  assign n12782 = ( n12778 & ~n12781 ) | ( n12778 & n12780 ) | ( ~n12781 & n12780 ) ;
  assign n12786 = x106 &  n2718 ;
  assign n12783 = ( x108 & ~n2642 ) | ( x108 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n12784 = x107 &  n2637 ;
  assign n12785 = n12783 | n12784 ;
  assign n12787 = ( x106 & ~n12786 ) | ( x106 & n12785 ) | ( ~n12786 & n12785 ) ;
  assign n12788 = ( n2645 & ~n5055 ) | ( n2645 & n12787 ) | ( ~n5055 & n12787 ) ;
  assign n12789 = n5055 | n12788 ;
  assign n12791 = ( x32 & n12787 ) | ( x32 & n12789 ) | ( n12787 & n12789 ) ;
  assign n12790 = ( x32 & ~n12789 ) | ( x32 & n12787 ) | ( ~n12789 & n12787 ) ;
  assign n12792 = ( n12789 & ~n12791 ) | ( n12789 & n12790 ) | ( ~n12791 & n12790 ) ;
  assign n12796 = x103 &  n3214 ;
  assign n12793 = ( x105 & ~n3087 ) | ( x105 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n12794 = x104 &  n3082 ;
  assign n12795 = n12793 | n12794 ;
  assign n12797 = ( x103 & ~n12796 ) | ( x103 & n12795 ) | ( ~n12796 & n12795 ) ;
  assign n12798 = ~n3090 & n4442 ;
  assign n12799 = n12797 | n12798 ;
  assign n12800 = ( x35 & ~n12799 ) | ( x35 & 1'b0 ) | ( ~n12799 & 1'b0 ) ;
  assign n12801 = ~x35 & n12799 ;
  assign n12802 = n12800 | n12801 ;
  assign n12920 = x100 &  n3756 ;
  assign n12917 = ( x102 & ~n3602 ) | ( x102 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n12918 = x101 &  n3597 ;
  assign n12919 = n12917 | n12918 ;
  assign n12921 = ( x100 & ~n12920 ) | ( x100 & n12919 ) | ( ~n12920 & n12919 ) ;
  assign n12922 = n3605 | n3872 ;
  assign n12923 = ~n12921 & n12922 ;
  assign n12924 = x38 &  n12923 ;
  assign n12925 = x38 | n12923 ;
  assign n12926 = ~n12924 & n12925 ;
  assign n12803 = ( n12390 & n12646 ) | ( n12390 & n12656 ) | ( n12646 & n12656 ) ;
  assign n12804 = ( n12576 & n12620 ) | ( n12576 & n12630 ) | ( n12620 & n12630 ) ;
  assign n12808 = x88 &  n6288 ;
  assign n12805 = ( x90 & ~n6032 ) | ( x90 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n12806 = x89 &  n6027 ;
  assign n12807 = n12805 | n12806 ;
  assign n12809 = ( x88 & ~n12808 ) | ( x88 & n12807 ) | ( ~n12808 & n12807 ) ;
  assign n12810 = ( n1976 & ~n6035 ) | ( n1976 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n12811 = n12809 | n12810 ;
  assign n12812 = ( x50 & ~n12811 ) | ( x50 & 1'b0 ) | ( ~n12811 & 1'b0 ) ;
  assign n12813 = ~x50 & n12811 ;
  assign n12814 = n12812 | n12813 ;
  assign n12815 = ( n12577 & n12607 ) | ( n12577 & n12617 ) | ( n12607 & n12617 ) ;
  assign n12819 = x85 &  n6982 ;
  assign n12816 = ( x87 & ~n6727 ) | ( x87 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n12817 = x86 &  n6722 ;
  assign n12818 = n12816 | n12817 ;
  assign n12820 = ( x85 & ~n12819 ) | ( x85 & n12818 ) | ( ~n12819 & n12818 ) ;
  assign n12821 = ( n1512 & ~n6730 ) | ( n1512 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n12822 = n12820 | n12821 ;
  assign n12823 = ( x53 & ~n12822 ) | ( x53 & 1'b0 ) | ( ~n12822 & 1'b0 ) ;
  assign n12824 = ~x53 & n12822 ;
  assign n12825 = n12823 | n12824 ;
  assign n12826 = ( n12355 & ~n12604 ) | ( n12355 & n12594 ) | ( ~n12604 & n12594 ) ;
  assign n12830 = x76 &  n9457 ;
  assign n12827 = ( x78 & ~n9150 ) | ( x78 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n12828 = x77 &  n9145 ;
  assign n12829 = n12827 | n12828 ;
  assign n12831 = ( x76 & ~n12830 ) | ( x76 & n12829 ) | ( ~n12830 & n12829 ) ;
  assign n12832 = ( n693 & ~n9153 ) | ( n693 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n12833 = n12831 | n12832 ;
  assign n12834 = ( x62 & ~n12833 ) | ( x62 & 1'b0 ) | ( ~n12833 & 1'b0 ) ;
  assign n12835 = ~x62 & n12833 ;
  assign n12836 = n12834 | n12835 ;
  assign n12837 = ( n12578 & ~n12591 ) | ( n12578 & n12588 ) | ( ~n12591 & n12588 ) ;
  assign n12838 = x74 &  n10104 ;
  assign n12839 = ( x75 & ~n9760 ) | ( x75 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n12840 = n12838 | n12839 ;
  assign n12841 = ( n12837 & ~n12591 ) | ( n12837 & n12840 ) | ( ~n12591 & n12840 ) ;
  assign n12842 = ( n12591 & ~n12840 ) | ( n12591 & n12837 ) | ( ~n12840 & n12837 ) ;
  assign n12843 = ( n12841 & ~n12837 ) | ( n12841 & n12842 ) | ( ~n12837 & n12842 ) ;
  assign n12847 = x79 &  n8558 ;
  assign n12844 = ( x81 & ~n8314 ) | ( x81 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n12845 = x80 &  n8309 ;
  assign n12846 = n12844 | n12845 ;
  assign n12848 = ( x79 & ~n12847 ) | ( x79 & n12846 ) | ( ~n12847 & n12846 ) ;
  assign n12849 = ( n994 & ~n8317 ) | ( n994 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n12850 = n12848 | n12849 ;
  assign n12851 = ( x59 & ~n12850 ) | ( x59 & 1'b0 ) | ( ~n12850 & 1'b0 ) ;
  assign n12852 = ~x59 & n12850 ;
  assign n12853 = n12851 | n12852 ;
  assign n12854 = ( n12836 & n12843 ) | ( n12836 & n12853 ) | ( n12843 & n12853 ) ;
  assign n12855 = ( n12843 & ~n12836 ) | ( n12843 & n12853 ) | ( ~n12836 & n12853 ) ;
  assign n12856 = ( n12836 & ~n12854 ) | ( n12836 & n12855 ) | ( ~n12854 & n12855 ) ;
  assign n12860 = x82 &  n7731 ;
  assign n12857 = ( x84 & ~n7538 ) | ( x84 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n12858 = x83 &  n7533 ;
  assign n12859 = n12857 | n12858 ;
  assign n12861 = ( x82 & ~n12860 ) | ( x82 & n12859 ) | ( ~n12860 & n12859 ) ;
  assign n12862 = ( n1199 & ~n7541 ) | ( n1199 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n12863 = n12861 | n12862 ;
  assign n12864 = ( x56 & ~n12863 ) | ( x56 & 1'b0 ) | ( ~n12863 & 1'b0 ) ;
  assign n12865 = ~x56 & n12863 ;
  assign n12866 = n12864 | n12865 ;
  assign n12868 = ( n12826 & n12856 ) | ( n12826 & n12866 ) | ( n12856 & n12866 ) ;
  assign n12867 = ( n12856 & ~n12826 ) | ( n12856 & n12866 ) | ( ~n12826 & n12866 ) ;
  assign n12869 = ( n12826 & ~n12868 ) | ( n12826 & n12867 ) | ( ~n12868 & n12867 ) ;
  assign n12871 = ( n12815 & n12825 ) | ( n12815 & n12869 ) | ( n12825 & n12869 ) ;
  assign n12870 = ( n12825 & ~n12815 ) | ( n12825 & n12869 ) | ( ~n12815 & n12869 ) ;
  assign n12872 = ( n12815 & ~n12871 ) | ( n12815 & n12870 ) | ( ~n12871 & n12870 ) ;
  assign n12874 = ( n12804 & n12814 ) | ( n12804 & n12872 ) | ( n12814 & n12872 ) ;
  assign n12873 = ( n12814 & ~n12804 ) | ( n12814 & n12872 ) | ( ~n12804 & n12872 ) ;
  assign n12875 = ( n12804 & ~n12874 ) | ( n12804 & n12873 ) | ( ~n12874 & n12873 ) ;
  assign n12876 = ( n12386 & n12633 ) | ( n12386 & n12643 ) | ( n12633 & n12643 ) ;
  assign n12880 = x91 &  n5586 ;
  assign n12877 = ( x93 & ~n5389 ) | ( x93 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n12878 = x92 &  n5384 ;
  assign n12879 = n12877 | n12878 ;
  assign n12881 = ( x91 & ~n12880 ) | ( x91 & n12879 ) | ( ~n12880 & n12879 ) ;
  assign n12882 = n2264 | n5392 ;
  assign n12883 = ~n12881 & n12882 ;
  assign n12884 = x47 &  n12883 ;
  assign n12885 = x47 | n12883 ;
  assign n12886 = ~n12884 & n12885 ;
  assign n12887 = ( n12875 & n12876 ) | ( n12875 & n12886 ) | ( n12876 & n12886 ) ;
  assign n12888 = ( n12876 & ~n12875 ) | ( n12876 & n12886 ) | ( ~n12875 & n12886 ) ;
  assign n12889 = ( n12875 & ~n12887 ) | ( n12875 & n12888 ) | ( ~n12887 & n12888 ) ;
  assign n12893 = x94 &  n4934 ;
  assign n12890 = ( x96 & ~n4725 ) | ( x96 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n12891 = x95 &  n4720 ;
  assign n12892 = n12890 | n12891 ;
  assign n12894 = ( x94 & ~n12893 ) | ( x94 & n12892 ) | ( ~n12893 & n12892 ) ;
  assign n12895 = ( n2836 & ~n4728 ) | ( n2836 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n12896 = n12894 | n12895 ;
  assign n12897 = ( x44 & ~n12896 ) | ( x44 & 1'b0 ) | ( ~n12896 & 1'b0 ) ;
  assign n12898 = ~x44 & n12896 ;
  assign n12899 = n12897 | n12898 ;
  assign n12900 = ( n12803 & n12889 ) | ( n12803 & n12899 ) | ( n12889 & n12899 ) ;
  assign n12901 = ( n12889 & ~n12803 ) | ( n12889 & n12899 ) | ( ~n12803 & n12899 ) ;
  assign n12902 = ( n12803 & ~n12900 ) | ( n12803 & n12901 ) | ( ~n12900 & n12901 ) ;
  assign n12906 = x97 &  n4344 ;
  assign n12903 = ( x99 & ~n4143 ) | ( x99 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n12904 = x98 &  n4138 ;
  assign n12905 = n12903 | n12904 ;
  assign n12907 = ( x97 & ~n12906 ) | ( x97 & n12905 ) | ( ~n12906 & n12905 ) ;
  assign n12908 = ( n3338 & ~n4146 ) | ( n3338 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n12909 = n12907 | n12908 ;
  assign n12910 = ( x41 & ~n12909 ) | ( x41 & 1'b0 ) | ( ~n12909 & 1'b0 ) ;
  assign n12911 = ~x41 & n12909 ;
  assign n12912 = n12910 | n12911 ;
  assign n12913 = ( n12575 & n12659 ) | ( n12575 & n12669 ) | ( n12659 & n12669 ) ;
  assign n12914 = ( n12902 & ~n12912 ) | ( n12902 & n12913 ) | ( ~n12912 & n12913 ) ;
  assign n12915 = ( n12902 & ~n12913 ) | ( n12902 & n12912 ) | ( ~n12913 & n12912 ) ;
  assign n12916 = ( n12914 & ~n12902 ) | ( n12914 & n12915 ) | ( ~n12902 & n12915 ) ;
  assign n12927 = ( n12674 & ~n12926 ) | ( n12674 & n12916 ) | ( ~n12926 & n12916 ) ;
  assign n12928 = ( n12674 & ~n12916 ) | ( n12674 & n12926 ) | ( ~n12916 & n12926 ) ;
  assign n12929 = ( n12927 & ~n12674 ) | ( n12927 & n12928 ) | ( ~n12674 & n12928 ) ;
  assign n12931 = ( n12677 & n12802 ) | ( n12677 & n12929 ) | ( n12802 & n12929 ) ;
  assign n12930 = ( n12802 & ~n12677 ) | ( n12802 & n12929 ) | ( ~n12677 & n12929 ) ;
  assign n12932 = ( n12677 & ~n12931 ) | ( n12677 & n12930 ) | ( ~n12931 & n12930 ) ;
  assign n12934 = ( n12680 & n12792 ) | ( n12680 & n12932 ) | ( n12792 & n12932 ) ;
  assign n12933 = ( n12680 & ~n12792 ) | ( n12680 & n12932 ) | ( ~n12792 & n12932 ) ;
  assign n12935 = ( n12792 & ~n12934 ) | ( n12792 & n12933 ) | ( ~n12934 & n12933 ) ;
  assign n12936 = ~n12782 & n12935 ;
  assign n12937 = ( n12782 & ~n12935 ) | ( n12782 & 1'b0 ) | ( ~n12935 & 1'b0 ) ;
  assign n12938 = n12936 | n12937 ;
  assign n12942 = x112 &  n1894 ;
  assign n12939 = ( x114 & ~n1816 ) | ( x114 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n12940 = x113 &  n1811 ;
  assign n12941 = n12939 | n12940 ;
  assign n12943 = ( x112 & ~n12942 ) | ( x112 & n12941 ) | ( ~n12942 & n12941 ) ;
  assign n12944 = ( n1819 & ~n6185 ) | ( n1819 & n12943 ) | ( ~n6185 & n12943 ) ;
  assign n12945 = n6185 | n12944 ;
  assign n12947 = ( x26 & n12943 ) | ( x26 & n12945 ) | ( n12943 & n12945 ) ;
  assign n12946 = ( x26 & ~n12945 ) | ( x26 & n12943 ) | ( ~n12945 & n12943 ) ;
  assign n12948 = ( n12945 & ~n12947 ) | ( n12945 & n12946 ) | ( ~n12947 & n12946 ) ;
  assign n12949 = ( n12771 & ~n12938 ) | ( n12771 & n12948 ) | ( ~n12938 & n12948 ) ;
  assign n12950 = ( n12771 & ~n12948 ) | ( n12771 & n12938 ) | ( ~n12948 & n12938 ) ;
  assign n12951 = ( n12949 & ~n12771 ) | ( n12949 & n12950 ) | ( ~n12771 & n12950 ) ;
  assign n12955 = x115 &  n1551 ;
  assign n12952 = ( x117 & ~n1451 ) | ( x117 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n12953 = x116 &  n1446 ;
  assign n12954 = n12952 | n12953 ;
  assign n12956 = ( x115 & ~n12955 ) | ( x115 & n12954 ) | ( ~n12955 & n12954 ) ;
  assign n12957 = ( n1454 & ~n7136 ) | ( n1454 & n12956 ) | ( ~n7136 & n12956 ) ;
  assign n12958 = n7136 | n12957 ;
  assign n12960 = ( x23 & n12956 ) | ( x23 & n12958 ) | ( n12956 & n12958 ) ;
  assign n12959 = ( x23 & ~n12958 ) | ( x23 & n12956 ) | ( ~n12958 & n12956 ) ;
  assign n12961 = ( n12958 & ~n12960 ) | ( n12958 & n12959 ) | ( ~n12960 & n12959 ) ;
  assign n12962 = ( n12770 & ~n12951 ) | ( n12770 & n12961 ) | ( ~n12951 & n12961 ) ;
  assign n12963 = ( n12770 & ~n12961 ) | ( n12770 & n12951 ) | ( ~n12961 & n12951 ) ;
  assign n12964 = ( n12962 & ~n12770 ) | ( n12962 & n12963 ) | ( ~n12770 & n12963 ) ;
  assign n12966 = ( n12759 & n12769 ) | ( n12759 & n12964 ) | ( n12769 & n12964 ) ;
  assign n12965 = ( n12769 & ~n12759 ) | ( n12769 & n12964 ) | ( ~n12759 & n12964 ) ;
  assign n12967 = ( n12759 & ~n12966 ) | ( n12759 & n12965 ) | ( ~n12966 & n12965 ) ;
  assign n12968 = ( n12757 & ~n12967 ) | ( n12757 & 1'b0 ) | ( ~n12967 & 1'b0 ) ;
  assign n12969 = ~n12757 & n12967 ;
  assign n12970 = n12968 | n12969 ;
  assign n12974 = x124 &  n713 ;
  assign n12971 = ( x126 & ~n641 ) | ( x126 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n12972 = x125 &  n636 ;
  assign n12973 = n12971 | n12972 ;
  assign n12975 = ( x124 & ~n12974 ) | ( x124 & n12973 ) | ( ~n12974 & n12973 ) ;
  assign n12976 = ( n644 & ~n9349 ) | ( n644 & n12975 ) | ( ~n9349 & n12975 ) ;
  assign n12977 = n9349 | n12976 ;
  assign n12979 = ( x14 & n12975 ) | ( x14 & n12977 ) | ( n12975 & n12977 ) ;
  assign n12978 = ( x14 & ~n12977 ) | ( x14 & n12975 ) | ( ~n12977 & n12975 ) ;
  assign n12980 = ( n12977 & ~n12979 ) | ( n12977 & n12978 ) | ( ~n12979 & n12978 ) ;
  assign n12981 = ( n12746 & ~n12970 ) | ( n12746 & n12980 ) | ( ~n12970 & n12980 ) ;
  assign n12982 = ( n12746 & ~n12980 ) | ( n12746 & n12970 ) | ( ~n12980 & n12970 ) ;
  assign n12983 = ( n12981 & ~n12746 ) | ( n12981 & n12982 ) | ( ~n12746 & n12982 ) ;
  assign n12984 = ( n12744 & n12745 ) | ( n12744 & n12983 ) | ( n12745 & n12983 ) ;
  assign n12985 = ( n12745 & ~n12744 ) | ( n12745 & n12983 ) | ( ~n12744 & n12983 ) ;
  assign n12986 = ( n12744 & ~n12984 ) | ( n12744 & n12985 ) | ( ~n12984 & n12985 ) ;
  assign n12987 = ( n12736 & n12738 ) | ( n12736 & n12986 ) | ( n12738 & n12986 ) ;
  assign n12988 = ( n12736 & ~n12738 ) | ( n12736 & n12986 ) | ( ~n12738 & n12986 ) ;
  assign n12989 = ( n12738 & ~n12987 ) | ( n12738 & n12988 ) | ( ~n12987 & n12988 ) ;
  assign n12990 = ( n12744 & ~n12745 ) | ( n12744 & n12983 ) | ( ~n12745 & n12983 ) ;
  assign n12991 = ( n12738 & ~n12736 ) | ( n12738 & n12986 ) | ( ~n12736 & n12986 ) ;
  assign n12995 = x125 &  n713 ;
  assign n12992 = ( x127 & ~n641 ) | ( x127 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n12993 = x126 &  n636 ;
  assign n12994 = n12992 | n12993 ;
  assign n12996 = ( x125 & ~n12995 ) | ( x125 & n12994 ) | ( ~n12995 & n12994 ) ;
  assign n12997 = n644 | n9941 ;
  assign n12998 = ~n12996 & n12997 ;
  assign n12999 = x14 &  n12998 ;
  assign n13000 = x14 | n12998 ;
  assign n13001 = ~n12999 & n13000 ;
  assign n13002 = ( n12746 & n12970 ) | ( n12746 & n12980 ) | ( n12970 & n12980 ) ;
  assign n13003 = x17 &  n12753 ;
  assign n13004 = ( n12755 & ~n13003 ) | ( n12755 & n12968 ) | ( ~n13003 & n12968 ) ;
  assign n13008 = x119 &  n1227 ;
  assign n13005 = ( x121 & ~n1154 ) | ( x121 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n13006 = x120 &  n1149 ;
  assign n13007 = n13005 | n13006 ;
  assign n13009 = ( x119 & ~n13008 ) | ( x119 & n13007 ) | ( ~n13008 & n13007 ) ;
  assign n13010 = ~n1157 & n8176 ;
  assign n13011 = n13009 | n13010 ;
  assign n13212 = x20 | n13011 ;
  assign n13213 = ~x20 & n13011 ;
  assign n13214 = ( n13212 & ~n13011 ) | ( n13212 & n13213 ) | ( ~n13011 & n13213 ) ;
  assign n13012 = ( n12759 & ~n12964 ) | ( n12759 & n12769 ) | ( ~n12964 & n12769 ) ;
  assign n13013 = ( n12770 & n12951 ) | ( n12770 & n12961 ) | ( n12951 & n12961 ) ;
  assign n13021 = ( n12771 & n12938 ) | ( n12771 & n12948 ) | ( n12938 & n12948 ) ;
  assign n13022 = ( x29 & ~n12778 ) | ( x29 & 1'b0 ) | ( ~n12778 & 1'b0 ) ;
  assign n13023 = ( n12780 & ~n13022 ) | ( n12780 & n12936 ) | ( ~n13022 & n12936 ) ;
  assign n13166 = ( n12680 & ~n12932 ) | ( n12680 & n12792 ) | ( ~n12932 & n12792 ) ;
  assign n13170 = x107 &  n2718 ;
  assign n13167 = ( x109 & ~n2642 ) | ( x109 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n13168 = x108 &  n2637 ;
  assign n13169 = n13167 | n13168 ;
  assign n13171 = ( x107 & ~n13170 ) | ( x107 & n13169 ) | ( ~n13170 & n13169 ) ;
  assign n13172 = ~n2645 & n5267 ;
  assign n13173 = n13171 | n13172 ;
  assign n13156 = x104 &  n3214 ;
  assign n13153 = ( x106 & ~n3087 ) | ( x106 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n13154 = x105 &  n3082 ;
  assign n13155 = n13153 | n13154 ;
  assign n13157 = ( x104 & ~n13156 ) | ( x104 & n13155 ) | ( ~n13156 & n13155 ) ;
  assign n13158 = ~n3090 & n4458 ;
  assign n13159 = n13157 | n13158 ;
  assign n13160 = ( x35 & ~n13159 ) | ( x35 & 1'b0 ) | ( ~n13159 & 1'b0 ) ;
  assign n13161 = ~x35 & n13159 ;
  assign n13162 = n13160 | n13161 ;
  assign n13037 = x86 &  n6982 ;
  assign n13034 = ( x88 & ~n6727 ) | ( x88 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n13035 = x87 &  n6722 ;
  assign n13036 = n13034 | n13035 ;
  assign n13038 = ( x86 & ~n13037 ) | ( x86 & n13036 ) | ( ~n13037 & n13036 ) ;
  assign n13039 = ( n1624 & ~n6730 ) | ( n1624 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n13040 = n13038 | n13039 ;
  assign n13041 = ( x53 & ~n13040 ) | ( x53 & 1'b0 ) | ( ~n13040 & 1'b0 ) ;
  assign n13042 = ~x53 & n13040 ;
  assign n13043 = n13041 | n13042 ;
  assign n13047 = x83 &  n7731 ;
  assign n13044 = ( x85 & ~n7538 ) | ( x85 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n13045 = x84 &  n7533 ;
  assign n13046 = n13044 | n13045 ;
  assign n13048 = ( x83 & ~n13047 ) | ( x83 & n13046 ) | ( ~n13047 & n13046 ) ;
  assign n13049 = ( n1295 & ~n7541 ) | ( n1295 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n13050 = n13048 | n13049 ;
  assign n13051 = ( x56 & ~n13050 ) | ( x56 & 1'b0 ) | ( ~n13050 & 1'b0 ) ;
  assign n13052 = ~x56 & n13050 ;
  assign n13053 = n13051 | n13052 ;
  assign n13057 = x80 &  n8558 ;
  assign n13054 = ( x82 & ~n8314 ) | ( x82 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n13055 = x81 &  n8309 ;
  assign n13056 = n13054 | n13055 ;
  assign n13058 = ( x80 & ~n13057 ) | ( x80 & n13056 ) | ( ~n13057 & n13056 ) ;
  assign n13059 = ( n1084 & ~n8317 ) | ( n1084 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n13060 = n13058 | n13059 ;
  assign n13061 = ( x59 & ~n13060 ) | ( x59 & 1'b0 ) | ( ~n13060 & 1'b0 ) ;
  assign n13062 = ~x59 & n13060 ;
  assign n13063 = n13061 | n13062 ;
  assign n13067 = x77 &  n9457 ;
  assign n13064 = ( x79 & ~n9150 ) | ( x79 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n13065 = x78 &  n9145 ;
  assign n13066 = n13064 | n13065 ;
  assign n13068 = ( x77 & ~n13067 ) | ( x77 & n13066 ) | ( ~n13067 & n13066 ) ;
  assign n13069 = ( n766 & ~n9153 ) | ( n766 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n13070 = n13068 | n13069 ;
  assign n13071 = ( x62 & ~n13070 ) | ( x62 & 1'b0 ) | ( ~n13070 & 1'b0 ) ;
  assign n13072 = ~x62 & n13070 ;
  assign n13073 = n13071 | n13072 ;
  assign n13074 = x75 &  n10104 ;
  assign n13075 = ( x76 & ~n9760 ) | ( x76 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n13076 = n13074 | n13075 ;
  assign n13077 = ( x11 & n12591 ) | ( x11 & n13076 ) | ( n12591 & n13076 ) ;
  assign n13078 = ( x11 & ~n12591 ) | ( x11 & n13076 ) | ( ~n12591 & n13076 ) ;
  assign n13079 = ( n12591 & ~n13077 ) | ( n12591 & n13078 ) | ( ~n13077 & n13078 ) ;
  assign n13080 = ( n13073 & ~n12841 ) | ( n13073 & n13079 ) | ( ~n12841 & n13079 ) ;
  assign n13081 = ( n12841 & ~n13079 ) | ( n12841 & n13073 ) | ( ~n13079 & n13073 ) ;
  assign n13082 = ( n13080 & ~n13073 ) | ( n13080 & n13081 ) | ( ~n13073 & n13081 ) ;
  assign n13083 = ( n12836 & ~n12843 ) | ( n12836 & n12853 ) | ( ~n12843 & n12853 ) ;
  assign n13084 = ( n13063 & n13082 ) | ( n13063 & n13083 ) | ( n13082 & n13083 ) ;
  assign n13085 = ( n13082 & ~n13063 ) | ( n13082 & n13083 ) | ( ~n13063 & n13083 ) ;
  assign n13086 = ( n13063 & ~n13084 ) | ( n13063 & n13085 ) | ( ~n13084 & n13085 ) ;
  assign n13087 = ( n12826 & ~n12866 ) | ( n12826 & n12856 ) | ( ~n12866 & n12856 ) ;
  assign n13089 = ( n13053 & n13086 ) | ( n13053 & n13087 ) | ( n13086 & n13087 ) ;
  assign n13088 = ( n13086 & ~n13053 ) | ( n13086 & n13087 ) | ( ~n13053 & n13087 ) ;
  assign n13090 = ( n13053 & ~n13089 ) | ( n13053 & n13088 ) | ( ~n13089 & n13088 ) ;
  assign n13092 = ( n12871 & n13043 ) | ( n12871 & n13090 ) | ( n13043 & n13090 ) ;
  assign n13091 = ( n12871 & ~n13043 ) | ( n12871 & n13090 ) | ( ~n13043 & n13090 ) ;
  assign n13093 = ( n13043 & ~n13092 ) | ( n13043 & n13091 ) | ( ~n13092 & n13091 ) ;
  assign n13027 = x89 &  n6288 ;
  assign n13024 = ( x91 & ~n6032 ) | ( x91 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n13025 = x90 &  n6027 ;
  assign n13026 = n13024 | n13025 ;
  assign n13028 = ( x89 & ~n13027 ) | ( x89 & n13026 ) | ( ~n13027 & n13026 ) ;
  assign n13029 = ( n2108 & ~n6035 ) | ( n2108 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n13030 = n13028 | n13029 ;
  assign n13031 = ( x50 & ~n13030 ) | ( x50 & 1'b0 ) | ( ~n13030 & 1'b0 ) ;
  assign n13032 = ~x50 & n13030 ;
  assign n13033 = n13031 | n13032 ;
  assign n13094 = ( n12874 & ~n13093 ) | ( n12874 & n13033 ) | ( ~n13093 & n13033 ) ;
  assign n13095 = ( n13033 & ~n12874 ) | ( n13033 & n13093 ) | ( ~n12874 & n13093 ) ;
  assign n13096 = ( n13094 & ~n13033 ) | ( n13094 & n13095 ) | ( ~n13033 & n13095 ) ;
  assign n13101 = x92 &  n5586 ;
  assign n13098 = ( x94 & ~n5389 ) | ( x94 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n13099 = x93 &  n5384 ;
  assign n13100 = n13098 | n13099 ;
  assign n13102 = ( x92 & ~n13101 ) | ( x92 & n13100 ) | ( ~n13101 & n13100 ) ;
  assign n13103 = ( n2401 & ~n5392 ) | ( n2401 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n13104 = n13102 | n13103 ;
  assign n13105 = ( x47 & ~n13104 ) | ( x47 & 1'b0 ) | ( ~n13104 & 1'b0 ) ;
  assign n13106 = ~x47 & n13104 ;
  assign n13107 = n13105 | n13106 ;
  assign n13097 = ( n12875 & ~n12886 ) | ( n12875 & n12876 ) | ( ~n12886 & n12876 ) ;
  assign n13108 = ( n13096 & ~n13107 ) | ( n13096 & n13097 ) | ( ~n13107 & n13097 ) ;
  assign n13109 = ( n13096 & ~n13097 ) | ( n13096 & n13107 ) | ( ~n13097 & n13107 ) ;
  assign n13110 = ( n13108 & ~n13096 ) | ( n13108 & n13109 ) | ( ~n13096 & n13109 ) ;
  assign n13111 = ( n12803 & ~n12889 ) | ( n12803 & n12899 ) | ( ~n12889 & n12899 ) ;
  assign n13115 = x95 &  n4934 ;
  assign n13112 = ( x97 & ~n4725 ) | ( x97 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n13113 = x96 &  n4720 ;
  assign n13114 = n13112 | n13113 ;
  assign n13116 = ( x95 & ~n13115 ) | ( x95 & n13114 ) | ( ~n13115 & n13114 ) ;
  assign n13117 = ( n2999 & ~n4728 ) | ( n2999 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n13118 = n13116 | n13117 ;
  assign n13119 = ( x44 & ~n13118 ) | ( x44 & 1'b0 ) | ( ~n13118 & 1'b0 ) ;
  assign n13120 = ~x44 & n13118 ;
  assign n13121 = n13119 | n13120 ;
  assign n13122 = ( n13110 & ~n13111 ) | ( n13110 & n13121 ) | ( ~n13111 & n13121 ) ;
  assign n13123 = ( n13110 & ~n13121 ) | ( n13110 & n13111 ) | ( ~n13121 & n13111 ) ;
  assign n13124 = ( n13122 & ~n13110 ) | ( n13122 & n13123 ) | ( ~n13110 & n13123 ) ;
  assign n13125 = ( n12912 & ~n12902 ) | ( n12912 & n12913 ) | ( ~n12902 & n12913 ) ;
  assign n13129 = x98 &  n4344 ;
  assign n13126 = ( x100 & ~n4143 ) | ( x100 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n13127 = x99 &  n4138 ;
  assign n13128 = n13126 | n13127 ;
  assign n13130 = ( x98 & ~n13129 ) | ( x98 & n13128 ) | ( ~n13129 & n13128 ) ;
  assign n13131 = n3354 | n4146 ;
  assign n13132 = ~n13130 & n13131 ;
  assign n13133 = x41 &  n13132 ;
  assign n13134 = x41 | n13132 ;
  assign n13135 = ~n13133 & n13134 ;
  assign n13137 = ( n13124 & n13125 ) | ( n13124 & n13135 ) | ( n13125 & n13135 ) ;
  assign n13136 = ( n13125 & ~n13124 ) | ( n13125 & n13135 ) | ( ~n13124 & n13135 ) ;
  assign n13138 = ( n13124 & ~n13137 ) | ( n13124 & n13136 ) | ( ~n13137 & n13136 ) ;
  assign n13143 = x101 &  n3756 ;
  assign n13140 = ( x103 & ~n3602 ) | ( x103 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n13141 = x102 &  n3597 ;
  assign n13142 = n13140 | n13141 ;
  assign n13144 = ( x101 & ~n13143 ) | ( x101 & n13142 ) | ( ~n13143 & n13142 ) ;
  assign n13145 = n3605 | n4056 ;
  assign n13146 = ~n13144 & n13145 ;
  assign n13147 = x38 &  n13146 ;
  assign n13148 = x38 | n13146 ;
  assign n13149 = ~n13147 & n13148 ;
  assign n13139 = ( n12916 & ~n12674 ) | ( n12916 & n12926 ) | ( ~n12674 & n12926 ) ;
  assign n13150 = ( n13138 & ~n13149 ) | ( n13138 & n13139 ) | ( ~n13149 & n13139 ) ;
  assign n13151 = ( n13138 & ~n13139 ) | ( n13138 & n13149 ) | ( ~n13139 & n13149 ) ;
  assign n13152 = ( n13150 & ~n13138 ) | ( n13150 & n13151 ) | ( ~n13138 & n13151 ) ;
  assign n13163 = ( n12931 & ~n13162 ) | ( n12931 & n13152 ) | ( ~n13162 & n13152 ) ;
  assign n13164 = ( n13152 & ~n12931 ) | ( n13152 & n13162 ) | ( ~n12931 & n13162 ) ;
  assign n13165 = ( n13163 & ~n13152 ) | ( n13163 & n13164 ) | ( ~n13152 & n13164 ) ;
  assign n13174 = x32 | n13165 ;
  assign n13175 = ~x32 & n13165 ;
  assign n13176 = ( n13174 & ~n13165 ) | ( n13174 & n13175 ) | ( ~n13165 & n13175 ) ;
  assign n13177 = ( n13166 & ~n13173 ) | ( n13166 & n13176 ) | ( ~n13173 & n13176 ) ;
  assign n13178 = ( n13173 & ~n13166 ) | ( n13173 & n13176 ) | ( ~n13166 & n13176 ) ;
  assign n13179 = ( n13177 & ~n13176 ) | ( n13177 & n13178 ) | ( ~n13176 & n13178 ) ;
  assign n13183 = x110 &  n2312 ;
  assign n13180 = ( x112 & ~n2195 ) | ( x112 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n13181 = x111 &  n2190 ;
  assign n13182 = n13180 | n13181 ;
  assign n13184 = ( x110 & ~n13183 ) | ( x110 & n13182 ) | ( ~n13183 & n13182 ) ;
  assign n13185 = ~n2198 & n5727 ;
  assign n13186 = n13184 | n13185 ;
  assign n13187 = ( x29 & ~n13186 ) | ( x29 & 1'b0 ) | ( ~n13186 & 1'b0 ) ;
  assign n13188 = ~x29 & n13186 ;
  assign n13189 = n13187 | n13188 ;
  assign n13190 = ( n13023 & ~n13179 ) | ( n13023 & n13189 ) | ( ~n13179 & n13189 ) ;
  assign n13191 = ( n13023 & ~n13189 ) | ( n13023 & n13179 ) | ( ~n13189 & n13179 ) ;
  assign n13192 = ( n13190 & ~n13023 ) | ( n13190 & n13191 ) | ( ~n13023 & n13191 ) ;
  assign n13017 = x113 &  n1894 ;
  assign n13014 = ( x115 & ~n1816 ) | ( x115 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n13015 = x114 &  n1811 ;
  assign n13016 = n13014 | n13015 ;
  assign n13018 = ( x113 & ~n13017 ) | ( x113 & n13016 ) | ( ~n13017 & n13016 ) ;
  assign n13019 = ~n1819 & n6420 ;
  assign n13020 = n13018 | n13019 ;
  assign n13193 = x26 | n13020 ;
  assign n13194 = ~x26 & n13020 ;
  assign n13195 = ( n13193 & ~n13020 ) | ( n13193 & n13194 ) | ( ~n13020 & n13194 ) ;
  assign n13196 = ( n13021 & ~n13192 ) | ( n13021 & n13195 ) | ( ~n13192 & n13195 ) ;
  assign n13197 = ( n13192 & ~n13021 ) | ( n13192 & n13195 ) | ( ~n13021 & n13195 ) ;
  assign n13198 = ( n13196 & ~n13195 ) | ( n13196 & n13197 ) | ( ~n13195 & n13197 ) ;
  assign n13202 = x116 &  n1551 ;
  assign n13199 = ( x118 & ~n1451 ) | ( x118 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n13200 = x117 &  n1446 ;
  assign n13201 = n13199 | n13200 ;
  assign n13203 = ( x116 & ~n13202 ) | ( x116 & n13201 ) | ( ~n13202 & n13201 ) ;
  assign n13204 = n1454 | n7152 ;
  assign n13205 = ~n13203 & n13204 ;
  assign n13206 = x23 &  n13205 ;
  assign n13207 = x23 | n13205 ;
  assign n13208 = ~n13206 & n13207 ;
  assign n13209 = ( n13013 & ~n13198 ) | ( n13013 & n13208 ) | ( ~n13198 & n13208 ) ;
  assign n13210 = ( n13013 & ~n13208 ) | ( n13013 & n13198 ) | ( ~n13208 & n13198 ) ;
  assign n13211 = ( n13209 & ~n13013 ) | ( n13209 & n13210 ) | ( ~n13013 & n13210 ) ;
  assign n13216 = ( n13012 & n13211 ) | ( n13012 & n13214 ) | ( n13211 & n13214 ) ;
  assign n13215 = ( n13012 & ~n13214 ) | ( n13012 & n13211 ) | ( ~n13214 & n13211 ) ;
  assign n13217 = ( n13214 & ~n13216 ) | ( n13214 & n13215 ) | ( ~n13216 & n13215 ) ;
  assign n13221 = x122 &  n942 ;
  assign n13218 = ( x124 & ~n896 ) | ( x124 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n13219 = x123 &  n891 ;
  assign n13220 = n13218 | n13219 ;
  assign n13222 = ( x122 & ~n13221 ) | ( x122 & n13220 ) | ( ~n13221 & n13220 ) ;
  assign n13223 = ~n899 & n8755 ;
  assign n13224 = n13222 | n13223 ;
  assign n13225 = ( x17 & ~n13224 ) | ( x17 & 1'b0 ) | ( ~n13224 & 1'b0 ) ;
  assign n13226 = ~x17 & n13224 ;
  assign n13227 = n13225 | n13226 ;
  assign n13228 = ( n13004 & n13217 ) | ( n13004 & n13227 ) | ( n13217 & n13227 ) ;
  assign n13229 = ( n13217 & ~n13004 ) | ( n13217 & n13227 ) | ( ~n13004 & n13227 ) ;
  assign n13230 = ( n13004 & ~n13228 ) | ( n13004 & n13229 ) | ( ~n13228 & n13229 ) ;
  assign n13231 = ( n13001 & ~n13002 ) | ( n13001 & n13230 ) | ( ~n13002 & n13230 ) ;
  assign n13232 = ( n13001 & ~n13230 ) | ( n13001 & n13002 ) | ( ~n13230 & n13002 ) ;
  assign n13233 = ( n13231 & ~n13001 ) | ( n13231 & n13232 ) | ( ~n13001 & n13232 ) ;
  assign n13234 = ( n12990 & n12991 ) | ( n12990 & n13233 ) | ( n12991 & n13233 ) ;
  assign n13235 = ( n12991 & ~n12990 ) | ( n12991 & n13233 ) | ( ~n12990 & n13233 ) ;
  assign n13236 = ( n12990 & ~n13234 ) | ( n12990 & n13235 ) | ( ~n13234 & n13235 ) ;
  assign n13237 = ( n13001 & n13002 ) | ( n13001 & n13230 ) | ( n13002 & n13230 ) ;
  assign n13238 = ( n12990 & ~n12991 ) | ( n12990 & n13233 ) | ( ~n12991 & n13233 ) ;
  assign n13239 = ( n13004 & ~n13217 ) | ( n13004 & n13227 ) | ( ~n13217 & n13227 ) ;
  assign n13240 = ( x20 & ~n13011 ) | ( x20 & 1'b0 ) | ( ~n13011 & 1'b0 ) ;
  assign n13241 = n13213 | n13240 ;
  assign n13242 = ( n13012 & ~n13211 ) | ( n13012 & n13241 ) | ( ~n13211 & n13241 ) ;
  assign n13246 = x123 &  n942 ;
  assign n13243 = ( x125 & ~n896 ) | ( x125 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n13244 = x124 &  n891 ;
  assign n13245 = n13243 | n13244 ;
  assign n13247 = ( x123 & ~n13246 ) | ( x123 & n13245 ) | ( ~n13246 & n13245 ) ;
  assign n13248 = ~n899 & n9324 ;
  assign n13249 = n13247 | n13248 ;
  assign n13250 = ( x17 & ~n13249 ) | ( x17 & 1'b0 ) | ( ~n13249 & 1'b0 ) ;
  assign n13251 = ~x17 & n13249 ;
  assign n13252 = n13250 | n13251 ;
  assign n13253 = ( n13013 & n13198 ) | ( n13013 & n13208 ) | ( n13198 & n13208 ) ;
  assign n13254 = x26 &  n13020 ;
  assign n13255 = ( n13193 & ~n13254 ) | ( n13193 & 1'b0 ) | ( ~n13254 & 1'b0 ) ;
  assign n13256 = ( n13192 & ~n13021 ) | ( n13192 & n13255 ) | ( ~n13021 & n13255 ) ;
  assign n13260 = x117 &  n1551 ;
  assign n13257 = ( x119 & ~n1451 ) | ( x119 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n13258 = x118 &  n1446 ;
  assign n13259 = n13257 | n13258 ;
  assign n13261 = ( x117 & ~n13260 ) | ( x117 & n13259 ) | ( ~n13260 & n13259 ) ;
  assign n13262 = ~n1454 & n7648 ;
  assign n13263 = n13261 | n13262 ;
  assign n13265 = x23 &  n13263 ;
  assign n13264 = ~x23 & n13263 ;
  assign n13266 = ( x23 & ~n13265 ) | ( x23 & n13264 ) | ( ~n13265 & n13264 ) ;
  assign n13267 = ( n13023 & n13179 ) | ( n13023 & n13189 ) | ( n13179 & n13189 ) ;
  assign n13268 = ( x32 & ~n13173 ) | ( x32 & 1'b0 ) | ( ~n13173 & 1'b0 ) ;
  assign n13269 = ~x32 & n13173 ;
  assign n13270 = n13268 | n13269 ;
  assign n13271 = ( n13165 & ~n13270 ) | ( n13165 & n13166 ) | ( ~n13270 & n13166 ) ;
  assign n13275 = x111 &  n2312 ;
  assign n13272 = ( x113 & ~n2195 ) | ( x113 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n13273 = x112 &  n2190 ;
  assign n13274 = n13272 | n13273 ;
  assign n13276 = ( x111 & ~n13275 ) | ( x111 & n13274 ) | ( ~n13275 & n13274 ) ;
  assign n13277 = n2198 | n6169 ;
  assign n13278 = ~n13276 & n13277 ;
  assign n13279 = x29 | n13278 ;
  assign n13280 = ( x29 & ~n13278 ) | ( x29 & 1'b0 ) | ( ~n13278 & 1'b0 ) ;
  assign n13281 = ( n13279 & ~x29 ) | ( n13279 & n13280 ) | ( ~x29 & n13280 ) ;
  assign n13282 = ( n12931 & ~n13152 ) | ( n12931 & n13162 ) | ( ~n13152 & n13162 ) ;
  assign n13426 = x108 &  n2718 ;
  assign n13423 = ( x110 & ~n2642 ) | ( x110 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n13424 = x109 &  n2637 ;
  assign n13425 = n13423 | n13424 ;
  assign n13427 = ( x108 & ~n13426 ) | ( x108 & n13425 ) | ( ~n13426 & n13425 ) ;
  assign n13428 = ~n2645 & n5283 ;
  assign n13429 = ( n2645 & ~n13427 ) | ( n2645 & n13428 ) | ( ~n13427 & n13428 ) ;
  assign n13431 = x32 &  n13429 ;
  assign n13430 = ~x32 & n13429 ;
  assign n13432 = ( x32 & ~n13431 ) | ( x32 & n13430 ) | ( ~n13431 & n13430 ) ;
  assign n13283 = ( n13138 & n13139 ) | ( n13138 & n13149 ) | ( n13139 & n13149 ) ;
  assign n13287 = x105 &  n3214 ;
  assign n13284 = ( x107 & ~n3087 ) | ( x107 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n13285 = x106 &  n3082 ;
  assign n13286 = n13284 | n13285 ;
  assign n13288 = ( x105 & ~n13287 ) | ( x105 & n13286 ) | ( ~n13287 & n13286 ) ;
  assign n13289 = ~n3090 & n4848 ;
  assign n13290 = n13288 | n13289 ;
  assign n13291 = ( x35 & ~n13290 ) | ( x35 & 1'b0 ) | ( ~n13290 & 1'b0 ) ;
  assign n13292 = ~x35 & n13290 ;
  assign n13293 = n13291 | n13292 ;
  assign n13294 = ( n13124 & ~n13135 ) | ( n13124 & n13125 ) | ( ~n13135 & n13125 ) ;
  assign n13298 = x102 &  n3756 ;
  assign n13295 = ( x104 & ~n3602 ) | ( x104 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n13296 = x103 &  n3597 ;
  assign n13297 = n13295 | n13296 ;
  assign n13299 = ( x102 & ~n13298 ) | ( x102 & n13297 ) | ( ~n13298 & n13297 ) ;
  assign n13300 = n3605 | n4249 ;
  assign n13301 = ~n13299 & n13300 ;
  assign n13302 = x38 &  n13301 ;
  assign n13303 = x38 | n13301 ;
  assign n13304 = ~n13302 & n13303 ;
  assign n13305 = ( n13110 & n13111 ) | ( n13110 & n13121 ) | ( n13111 & n13121 ) ;
  assign n13319 = x96 &  n4934 ;
  assign n13316 = ( x98 & ~n4725 ) | ( x98 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n13317 = x97 &  n4720 ;
  assign n13318 = n13316 | n13317 ;
  assign n13320 = ( x96 & ~n13319 ) | ( x96 & n13318 ) | ( ~n13319 & n13318 ) ;
  assign n13321 = ( n3170 & ~n4728 ) | ( n3170 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n13322 = n13320 | n13321 ;
  assign n13323 = ( x44 & ~n13322 ) | ( x44 & 1'b0 ) | ( ~n13322 & 1'b0 ) ;
  assign n13324 = ~x44 & n13322 ;
  assign n13325 = n13323 | n13324 ;
  assign n13326 = ( n13096 & n13097 ) | ( n13096 & n13107 ) | ( n13097 & n13107 ) ;
  assign n13327 = ( n12874 & n13033 ) | ( n12874 & n13093 ) | ( n13033 & n13093 ) ;
  assign n13331 = x93 &  n5586 ;
  assign n13328 = ( x95 & ~n5389 ) | ( x95 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n13329 = x94 &  n5384 ;
  assign n13330 = n13328 | n13329 ;
  assign n13332 = ( x93 & ~n13331 ) | ( x93 & n13330 ) | ( ~n13331 & n13330 ) ;
  assign n13333 = ( n2547 & ~n5392 ) | ( n2547 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n13334 = n13332 | n13333 ;
  assign n13335 = ( x47 & ~n13334 ) | ( x47 & 1'b0 ) | ( ~n13334 & 1'b0 ) ;
  assign n13336 = ~x47 & n13334 ;
  assign n13337 = n13335 | n13336 ;
  assign n13338 = ( n13063 & ~n13082 ) | ( n13063 & n13083 ) | ( ~n13082 & n13083 ) ;
  assign n13339 = ( n12591 & ~x11 ) | ( n12591 & n13076 ) | ( ~x11 & n13076 ) ;
  assign n13340 = x76 &  n10104 ;
  assign n13341 = ( x77 & ~n9760 ) | ( x77 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n13342 = n13340 | n13341 ;
  assign n13346 = x78 &  n9457 ;
  assign n13343 = ( x80 & ~n9150 ) | ( x80 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n13344 = x79 &  n9145 ;
  assign n13345 = n13343 | n13344 ;
  assign n13347 = ( x78 & ~n13346 ) | ( x78 & n13345 ) | ( ~n13346 & n13345 ) ;
  assign n13348 = ( n842 & ~n9153 ) | ( n842 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n13349 = n13347 | n13348 ;
  assign n13350 = ( x62 & ~n13349 ) | ( x62 & 1'b0 ) | ( ~n13349 & 1'b0 ) ;
  assign n13351 = ~x62 & n13349 ;
  assign n13352 = n13350 | n13351 ;
  assign n13353 = ( n13339 & ~n13342 ) | ( n13339 & n13352 ) | ( ~n13342 & n13352 ) ;
  assign n13354 = ( n13339 & ~n13352 ) | ( n13339 & n13342 ) | ( ~n13352 & n13342 ) ;
  assign n13355 = ( n13353 & ~n13339 ) | ( n13353 & n13354 ) | ( ~n13339 & n13354 ) ;
  assign n13359 = x81 &  n8558 ;
  assign n13356 = ( x83 & ~n8314 ) | ( x83 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n13357 = x82 &  n8309 ;
  assign n13358 = n13356 | n13357 ;
  assign n13360 = ( x81 & ~n13359 ) | ( x81 & n13358 ) | ( ~n13359 & n13358 ) ;
  assign n13361 = ( n1100 & ~n8317 ) | ( n1100 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n13362 = n13360 | n13361 ;
  assign n13363 = ( x59 & ~n13362 ) | ( x59 & 1'b0 ) | ( ~n13362 & 1'b0 ) ;
  assign n13364 = ~x59 & n13362 ;
  assign n13365 = n13363 | n13364 ;
  assign n13366 = ( n13081 & n13355 ) | ( n13081 & n13365 ) | ( n13355 & n13365 ) ;
  assign n13367 = ( n13355 & ~n13081 ) | ( n13355 & n13365 ) | ( ~n13081 & n13365 ) ;
  assign n13368 = ( n13081 & ~n13366 ) | ( n13081 & n13367 ) | ( ~n13366 & n13367 ) ;
  assign n13372 = x84 &  n7731 ;
  assign n13369 = ( x86 & ~n7538 ) | ( x86 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n13370 = x85 &  n7533 ;
  assign n13371 = n13369 | n13370 ;
  assign n13373 = ( x84 & ~n13372 ) | ( x84 & n13371 ) | ( ~n13372 & n13371 ) ;
  assign n13374 = ( n1496 & ~n7541 ) | ( n1496 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n13375 = n13373 | n13374 ;
  assign n13376 = ( x56 & ~n13375 ) | ( x56 & 1'b0 ) | ( ~n13375 & 1'b0 ) ;
  assign n13377 = ~x56 & n13375 ;
  assign n13378 = n13376 | n13377 ;
  assign n13379 = ( n13338 & n13368 ) | ( n13338 & n13378 ) | ( n13368 & n13378 ) ;
  assign n13380 = ( n13368 & ~n13338 ) | ( n13368 & n13378 ) | ( ~n13338 & n13378 ) ;
  assign n13381 = ( n13338 & ~n13379 ) | ( n13338 & n13380 ) | ( ~n13379 & n13380 ) ;
  assign n13385 = x87 &  n6982 ;
  assign n13382 = ( x89 & ~n6727 ) | ( x89 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n13383 = x88 &  n6722 ;
  assign n13384 = n13382 | n13383 ;
  assign n13386 = ( x87 & ~n13385 ) | ( x87 & n13384 ) | ( ~n13385 & n13384 ) ;
  assign n13387 = ( n1741 & ~n6730 ) | ( n1741 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n13388 = n13386 | n13387 ;
  assign n13389 = ( x53 & ~n13388 ) | ( x53 & 1'b0 ) | ( ~n13388 & 1'b0 ) ;
  assign n13390 = ~x53 & n13388 ;
  assign n13391 = n13389 | n13390 ;
  assign n13393 = ( n13088 & n13381 ) | ( n13088 & n13391 ) | ( n13381 & n13391 ) ;
  assign n13392 = ( n13381 & ~n13088 ) | ( n13381 & n13391 ) | ( ~n13088 & n13391 ) ;
  assign n13394 = ( n13088 & ~n13393 ) | ( n13088 & n13392 ) | ( ~n13393 & n13392 ) ;
  assign n13398 = x90 &  n6288 ;
  assign n13395 = ( x92 & ~n6032 ) | ( x92 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n13396 = x91 &  n6027 ;
  assign n13397 = n13395 | n13396 ;
  assign n13399 = ( x90 & ~n13398 ) | ( x90 & n13397 ) | ( ~n13398 & n13397 ) ;
  assign n13400 = ( n2248 & ~n6035 ) | ( n2248 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n13401 = n13399 | n13400 ;
  assign n13402 = ( x50 & ~n13401 ) | ( x50 & 1'b0 ) | ( ~n13401 & 1'b0 ) ;
  assign n13403 = ~x50 & n13401 ;
  assign n13404 = n13402 | n13403 ;
  assign n13405 = ( n13092 & ~n13394 ) | ( n13092 & n13404 ) | ( ~n13394 & n13404 ) ;
  assign n13406 = ( n13092 & ~n13404 ) | ( n13092 & n13394 ) | ( ~n13404 & n13394 ) ;
  assign n13407 = ( n13405 & ~n13092 ) | ( n13405 & n13406 ) | ( ~n13092 & n13406 ) ;
  assign n13409 = ( n13327 & n13337 ) | ( n13327 & n13407 ) | ( n13337 & n13407 ) ;
  assign n13408 = ( n13337 & ~n13327 ) | ( n13337 & n13407 ) | ( ~n13327 & n13407 ) ;
  assign n13410 = ( n13327 & ~n13409 ) | ( n13327 & n13408 ) | ( ~n13409 & n13408 ) ;
  assign n13412 = ( n13325 & n13326 ) | ( n13325 & n13410 ) | ( n13326 & n13410 ) ;
  assign n13411 = ( n13326 & ~n13325 ) | ( n13326 & n13410 ) | ( ~n13325 & n13410 ) ;
  assign n13413 = ( n13325 & ~n13412 ) | ( n13325 & n13411 ) | ( ~n13412 & n13411 ) ;
  assign n13309 = x99 &  n4344 ;
  assign n13306 = ( x101 & ~n4143 ) | ( x101 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n13307 = x100 &  n4138 ;
  assign n13308 = n13306 | n13307 ;
  assign n13310 = ( x99 & ~n13309 ) | ( x99 & n13308 ) | ( ~n13309 & n13308 ) ;
  assign n13311 = n3694 | n4146 ;
  assign n13312 = ~n13310 & n13311 ;
  assign n13313 = x41 &  n13312 ;
  assign n13314 = x41 | n13312 ;
  assign n13315 = ~n13313 & n13314 ;
  assign n13414 = ( n13305 & ~n13413 ) | ( n13305 & n13315 ) | ( ~n13413 & n13315 ) ;
  assign n13415 = ( n13305 & ~n13315 ) | ( n13305 & n13413 ) | ( ~n13315 & n13413 ) ;
  assign n13416 = ( n13414 & ~n13305 ) | ( n13414 & n13415 ) | ( ~n13305 & n13415 ) ;
  assign n13417 = ( n13294 & n13304 ) | ( n13294 & n13416 ) | ( n13304 & n13416 ) ;
  assign n13418 = ( n13304 & ~n13294 ) | ( n13304 & n13416 ) | ( ~n13294 & n13416 ) ;
  assign n13419 = ( n13294 & ~n13417 ) | ( n13294 & n13418 ) | ( ~n13417 & n13418 ) ;
  assign n13420 = ( n13283 & n13293 ) | ( n13283 & n13419 ) | ( n13293 & n13419 ) ;
  assign n13421 = ( n13293 & ~n13283 ) | ( n13293 & n13419 ) | ( ~n13283 & n13419 ) ;
  assign n13422 = ( n13283 & ~n13420 ) | ( n13283 & n13421 ) | ( ~n13420 & n13421 ) ;
  assign n13433 = ( n13282 & ~n13432 ) | ( n13282 & n13422 ) | ( ~n13432 & n13422 ) ;
  assign n13434 = ( n13282 & ~n13422 ) | ( n13282 & n13432 ) | ( ~n13422 & n13432 ) ;
  assign n13435 = ( n13433 & ~n13282 ) | ( n13433 & n13434 ) | ( ~n13282 & n13434 ) ;
  assign n13437 = ( n13271 & n13281 ) | ( n13271 & n13435 ) | ( n13281 & n13435 ) ;
  assign n13436 = ( n13281 & ~n13271 ) | ( n13281 & n13435 ) | ( ~n13271 & n13435 ) ;
  assign n13438 = ( n13271 & ~n13437 ) | ( n13271 & n13436 ) | ( ~n13437 & n13436 ) ;
  assign n13442 = x114 &  n1894 ;
  assign n13439 = ( x116 & ~n1816 ) | ( x116 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n13440 = x115 &  n1811 ;
  assign n13441 = n13439 | n13440 ;
  assign n13443 = ( x114 & ~n13442 ) | ( x114 & n13441 ) | ( ~n13442 & n13441 ) ;
  assign n13444 = ( n1819 & ~n6885 ) | ( n1819 & n13443 ) | ( ~n6885 & n13443 ) ;
  assign n13445 = n6885 | n13444 ;
  assign n13447 = ( x26 & n13443 ) | ( x26 & n13445 ) | ( n13443 & n13445 ) ;
  assign n13446 = ( x26 & ~n13445 ) | ( x26 & n13443 ) | ( ~n13445 & n13443 ) ;
  assign n13448 = ( n13445 & ~n13447 ) | ( n13445 & n13446 ) | ( ~n13447 & n13446 ) ;
  assign n13450 = ( n13267 & n13438 ) | ( n13267 & n13448 ) | ( n13438 & n13448 ) ;
  assign n13449 = ( n13438 & ~n13267 ) | ( n13438 & n13448 ) | ( ~n13267 & n13448 ) ;
  assign n13451 = ( n13267 & ~n13450 ) | ( n13267 & n13449 ) | ( ~n13450 & n13449 ) ;
  assign n13453 = ( n13256 & n13266 ) | ( n13256 & n13451 ) | ( n13266 & n13451 ) ;
  assign n13452 = ( n13266 & ~n13256 ) | ( n13266 & n13451 ) | ( ~n13256 & n13451 ) ;
  assign n13454 = ( n13256 & ~n13453 ) | ( n13256 & n13452 ) | ( ~n13453 & n13452 ) ;
  assign n13458 = x120 &  n1227 ;
  assign n13455 = ( x122 & ~n1154 ) | ( x122 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n13456 = x121 &  n1149 ;
  assign n13457 = n13455 | n13456 ;
  assign n13459 = ( x120 & ~n13458 ) | ( x120 & n13457 ) | ( ~n13458 & n13457 ) ;
  assign n13460 = ( n1157 & n9987 ) | ( n1157 & n13459 ) | ( n9987 & n13459 ) ;
  assign n13461 = ( n9987 & ~n13460 ) | ( n9987 & 1'b0 ) | ( ~n13460 & 1'b0 ) ;
  assign n13462 = ( x20 & n13459 ) | ( x20 & n13461 ) | ( n13459 & n13461 ) ;
  assign n13463 = ( x20 & ~n13461 ) | ( x20 & n13459 ) | ( ~n13461 & n13459 ) ;
  assign n13464 = ( n13461 & ~n13462 ) | ( n13461 & n13463 ) | ( ~n13462 & n13463 ) ;
  assign n13466 = ( n13253 & n13454 ) | ( n13253 & n13464 ) | ( n13454 & n13464 ) ;
  assign n13465 = ( n13454 & ~n13253 ) | ( n13454 & n13464 ) | ( ~n13253 & n13464 ) ;
  assign n13467 = ( n13253 & ~n13466 ) | ( n13253 & n13465 ) | ( ~n13466 & n13465 ) ;
  assign n13468 = ( n13242 & ~n13252 ) | ( n13242 & n13467 ) | ( ~n13252 & n13467 ) ;
  assign n13469 = ( n13242 & ~n13467 ) | ( n13242 & n13252 ) | ( ~n13467 & n13252 ) ;
  assign n13470 = ( n13468 & ~n13242 ) | ( n13468 & n13469 ) | ( ~n13242 & n13469 ) ;
  assign n13471 = ( x126 & ~n713 ) | ( x126 & 1'b0 ) | ( ~n713 & 1'b0 ) ;
  assign n13472 = x127 &  n636 ;
  assign n13473 = n13471 | n13472 ;
  assign n13474 = n644 | n9960 ;
  assign n13475 = ( n13473 & ~n644 ) | ( n13473 & n13474 ) | ( ~n644 & n13474 ) ;
  assign n13476 = x14 | n13475 ;
  assign n13477 = ( x14 & ~n13475 ) | ( x14 & 1'b0 ) | ( ~n13475 & 1'b0 ) ;
  assign n13478 = ( n13476 & ~x14 ) | ( n13476 & n13477 ) | ( ~x14 & n13477 ) ;
  assign n13479 = ( n13239 & ~n13470 ) | ( n13239 & n13478 ) | ( ~n13470 & n13478 ) ;
  assign n13480 = ( n13239 & ~n13478 ) | ( n13239 & n13470 ) | ( ~n13478 & n13470 ) ;
  assign n13481 = ( n13479 & ~n13239 ) | ( n13479 & n13480 ) | ( ~n13239 & n13480 ) ;
  assign n13482 = ( n13237 & ~n13238 ) | ( n13237 & n13481 ) | ( ~n13238 & n13481 ) ;
  assign n13483 = ( n13237 & ~n13481 ) | ( n13237 & n13238 ) | ( ~n13481 & n13238 ) ;
  assign n13484 = ( n13482 & ~n13237 ) | ( n13482 & n13483 ) | ( ~n13237 & n13483 ) ;
  assign n13486 = ( x127 & ~n713 ) | ( x127 & 1'b0 ) | ( ~n713 & 1'b0 ) ;
  assign n13487 = n644 | n10258 ;
  assign n13488 = ~n13486 & n13487 ;
  assign n13489 = ~x14 & n13488 ;
  assign n13490 = ( x14 & ~n13488 ) | ( x14 & 1'b0 ) | ( ~n13488 & 1'b0 ) ;
  assign n13491 = n13489 | n13490 ;
  assign n13493 = ( n13253 & ~n13464 ) | ( n13253 & n13454 ) | ( ~n13464 & n13454 ) ;
  assign n13497 = x121 &  n1227 ;
  assign n13494 = ( x123 & ~n1154 ) | ( x123 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n13495 = x122 &  n1149 ;
  assign n13496 = n13494 | n13495 ;
  assign n13498 = ( x121 & ~n13497 ) | ( x121 & n13496 ) | ( ~n13497 & n13496 ) ;
  assign n13499 = ~n1157 & n8472 ;
  assign n13500 = n13498 | n13499 ;
  assign n13501 = ( x20 & ~n13500 ) | ( x20 & 1'b0 ) | ( ~n13500 & 1'b0 ) ;
  assign n13502 = ~x20 & n13500 ;
  assign n13503 = n13501 | n13502 ;
  assign n13511 = ( n13267 & ~n13448 ) | ( n13267 & n13438 ) | ( ~n13448 & n13438 ) ;
  assign n13507 = x118 &  n1551 ;
  assign n13504 = ( x120 & ~n1451 ) | ( x120 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n13505 = x119 &  n1446 ;
  assign n13506 = n13504 | n13505 ;
  assign n13508 = ( x118 & ~n13507 ) | ( x118 & n13506 ) | ( ~n13507 & n13506 ) ;
  assign n13509 = ~n1454 & n9364 ;
  assign n13510 = n13508 | n13509 ;
  assign n13512 = ( x23 & n13510 ) | ( x23 & n13511 ) | ( n13510 & n13511 ) ;
  assign n13513 = ( x23 & ~n13511 ) | ( x23 & n13510 ) | ( ~n13511 & n13510 ) ;
  assign n13514 = ( n13511 & ~n13512 ) | ( n13511 & n13513 ) | ( ~n13512 & n13513 ) ;
  assign n13515 = ( n13271 & ~n13435 ) | ( n13271 & n13281 ) | ( ~n13435 & n13281 ) ;
  assign n13519 = x115 &  n1894 ;
  assign n13516 = ( x117 & ~n1816 ) | ( x117 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n13517 = x116 &  n1811 ;
  assign n13518 = n13516 | n13517 ;
  assign n13520 = ( x115 & ~n13519 ) | ( x115 & n13518 ) | ( ~n13519 & n13518 ) ;
  assign n13521 = n1819 | n7136 ;
  assign n13522 = ~n13520 & n13521 ;
  assign n13523 = x26 &  n13522 ;
  assign n13524 = x26 | n13522 ;
  assign n13525 = ~n13523 & n13524 ;
  assign n13526 = ( n13422 & ~n13282 ) | ( n13422 & n13432 ) | ( ~n13282 & n13432 ) ;
  assign n13540 = x106 &  n3214 ;
  assign n13537 = ( x108 & ~n3087 ) | ( x108 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n13538 = x107 &  n3082 ;
  assign n13539 = n13537 | n13538 ;
  assign n13541 = ( x106 & ~n13540 ) | ( x106 & n13539 ) | ( ~n13540 & n13539 ) ;
  assign n13542 = n3090 | n5055 ;
  assign n13543 = ~n13541 & n13542 ;
  assign n13544 = x35 &  n13543 ;
  assign n13545 = x35 | n13543 ;
  assign n13546 = ~n13544 & n13545 ;
  assign n13550 = x103 &  n3756 ;
  assign n13547 = ( x105 & ~n3602 ) | ( x105 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n13548 = x104 &  n3597 ;
  assign n13549 = n13547 | n13548 ;
  assign n13551 = ( x103 & ~n13550 ) | ( x103 & n13549 ) | ( ~n13550 & n13549 ) ;
  assign n13552 = ~n3605 & n4442 ;
  assign n13553 = n13551 | n13552 ;
  assign n13554 = ( x38 & ~n13553 ) | ( x38 & 1'b0 ) | ( ~n13553 & 1'b0 ) ;
  assign n13555 = ~x38 & n13553 ;
  assign n13556 = n13554 | n13555 ;
  assign n13658 = x100 &  n4344 ;
  assign n13655 = ( x102 & ~n4143 ) | ( x102 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n13656 = x101 &  n4138 ;
  assign n13657 = n13655 | n13656 ;
  assign n13659 = ( x100 & ~n13658 ) | ( x100 & n13657 ) | ( ~n13658 & n13657 ) ;
  assign n13660 = n3872 | n4146 ;
  assign n13661 = ~n13659 & n13660 ;
  assign n13662 = x41 &  n13661 ;
  assign n13663 = x41 | n13661 ;
  assign n13664 = ~n13662 & n13663 ;
  assign n13645 = x97 &  n4934 ;
  assign n13642 = ( x99 & ~n4725 ) | ( x99 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n13643 = x98 &  n4720 ;
  assign n13644 = n13642 | n13643 ;
  assign n13646 = ( x97 & ~n13645 ) | ( x97 & n13644 ) | ( ~n13645 & n13644 ) ;
  assign n13647 = ( n3338 & ~n4728 ) | ( n3338 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n13648 = n13646 | n13647 ;
  assign n13649 = ( x44 & ~n13648 ) | ( x44 & 1'b0 ) | ( ~n13648 & 1'b0 ) ;
  assign n13650 = ~x44 & n13648 ;
  assign n13651 = n13649 | n13650 ;
  assign n13557 = ( n13092 & n13394 ) | ( n13092 & n13404 ) | ( n13394 & n13404 ) ;
  assign n13558 = ( n13338 & ~n13368 ) | ( n13338 & n13378 ) | ( ~n13368 & n13378 ) ;
  assign n13562 = x88 &  n6982 ;
  assign n13559 = ( x90 & ~n6727 ) | ( x90 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n13560 = x89 &  n6722 ;
  assign n13561 = n13559 | n13560 ;
  assign n13563 = ( x88 & ~n13562 ) | ( x88 & n13561 ) | ( ~n13562 & n13561 ) ;
  assign n13564 = ( n1976 & ~n6730 ) | ( n1976 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n13565 = n13563 | n13564 ;
  assign n13566 = ( x53 & ~n13565 ) | ( x53 & 1'b0 ) | ( ~n13565 & 1'b0 ) ;
  assign n13567 = ~x53 & n13565 ;
  assign n13568 = n13566 | n13567 ;
  assign n13569 = ( n13081 & ~n13355 ) | ( n13081 & n13365 ) | ( ~n13355 & n13365 ) ;
  assign n13570 = x77 &  n10104 ;
  assign n13571 = ( x78 & ~n9760 ) | ( x78 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n13572 = n13570 | n13571 ;
  assign n13576 = x79 &  n9457 ;
  assign n13573 = ( x81 & ~n9150 ) | ( x81 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n13574 = x80 &  n9145 ;
  assign n13575 = n13573 | n13574 ;
  assign n13577 = ( x79 & ~n13576 ) | ( x79 & n13575 ) | ( ~n13576 & n13575 ) ;
  assign n13578 = ( n994 & ~n13577 ) | ( n994 & n9153 ) | ( ~n13577 & n9153 ) ;
  assign n13579 = ~n9153 & n13578 ;
  assign n13580 = ( x62 & n13577 ) | ( x62 & n13579 ) | ( n13577 & n13579 ) ;
  assign n13581 = ( x62 & ~n13579 ) | ( x62 & n13577 ) | ( ~n13579 & n13577 ) ;
  assign n13582 = ( n13579 & ~n13580 ) | ( n13579 & n13581 ) | ( ~n13580 & n13581 ) ;
  assign n13583 = ( n13572 & ~n13342 ) | ( n13572 & n13582 ) | ( ~n13342 & n13582 ) ;
  assign n13584 = ( n13342 & ~n13582 ) | ( n13342 & n13572 ) | ( ~n13582 & n13572 ) ;
  assign n13585 = ( n13583 & ~n13572 ) | ( n13583 & n13584 ) | ( ~n13572 & n13584 ) ;
  assign n13589 = x82 &  n8558 ;
  assign n13586 = ( x84 & ~n8314 ) | ( x84 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n13587 = x83 &  n8309 ;
  assign n13588 = n13586 | n13587 ;
  assign n13590 = ( x82 & ~n13589 ) | ( x82 & n13588 ) | ( ~n13589 & n13588 ) ;
  assign n13591 = ( n1199 & ~n8317 ) | ( n1199 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n13592 = n13590 | n13591 ;
  assign n13593 = ( x59 & ~n13592 ) | ( x59 & 1'b0 ) | ( ~n13592 & 1'b0 ) ;
  assign n13594 = ~x59 & n13592 ;
  assign n13595 = n13593 | n13594 ;
  assign n13596 = ( n13585 & ~n13353 ) | ( n13585 & n13595 ) | ( ~n13353 & n13595 ) ;
  assign n13597 = ( n13353 & ~n13595 ) | ( n13353 & n13585 ) | ( ~n13595 & n13585 ) ;
  assign n13598 = ( n13596 & ~n13585 ) | ( n13596 & n13597 ) | ( ~n13585 & n13597 ) ;
  assign n13602 = x85 &  n7731 ;
  assign n13599 = ( x87 & ~n7538 ) | ( x87 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n13600 = x86 &  n7533 ;
  assign n13601 = n13599 | n13600 ;
  assign n13603 = ( x85 & ~n13602 ) | ( x85 & n13601 ) | ( ~n13602 & n13601 ) ;
  assign n13604 = ( n1512 & ~n7541 ) | ( n1512 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n13605 = n13603 | n13604 ;
  assign n13606 = ( x56 & ~n13605 ) | ( x56 & 1'b0 ) | ( ~n13605 & 1'b0 ) ;
  assign n13607 = ~x56 & n13605 ;
  assign n13608 = n13606 | n13607 ;
  assign n13609 = ( n13569 & n13598 ) | ( n13569 & n13608 ) | ( n13598 & n13608 ) ;
  assign n13610 = ( n13598 & ~n13569 ) | ( n13598 & n13608 ) | ( ~n13569 & n13608 ) ;
  assign n13611 = ( n13569 & ~n13609 ) | ( n13569 & n13610 ) | ( ~n13609 & n13610 ) ;
  assign n13612 = ( n13558 & ~n13568 ) | ( n13558 & n13611 ) | ( ~n13568 & n13611 ) ;
  assign n13613 = ( n13558 & ~n13611 ) | ( n13558 & n13568 ) | ( ~n13611 & n13568 ) ;
  assign n13614 = ( n13612 & ~n13558 ) | ( n13612 & n13613 ) | ( ~n13558 & n13613 ) ;
  assign n13619 = x91 &  n6288 ;
  assign n13616 = ( x93 & ~n6032 ) | ( x93 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n13617 = x92 &  n6027 ;
  assign n13618 = n13616 | n13617 ;
  assign n13620 = ( x91 & ~n13619 ) | ( x91 & n13618 ) | ( ~n13619 & n13618 ) ;
  assign n13621 = n2264 | n6035 ;
  assign n13622 = ~n13620 & n13621 ;
  assign n13623 = x50 &  n13622 ;
  assign n13624 = x50 | n13622 ;
  assign n13625 = ~n13623 & n13624 ;
  assign n13615 = ( n13088 & ~n13391 ) | ( n13088 & n13381 ) | ( ~n13391 & n13381 ) ;
  assign n13626 = ( n13614 & ~n13625 ) | ( n13614 & n13615 ) | ( ~n13625 & n13615 ) ;
  assign n13627 = ( n13614 & ~n13615 ) | ( n13614 & n13625 ) | ( ~n13615 & n13625 ) ;
  assign n13628 = ( n13626 & ~n13614 ) | ( n13626 & n13627 ) | ( ~n13614 & n13627 ) ;
  assign n13632 = x94 &  n5586 ;
  assign n13629 = ( x96 & ~n5389 ) | ( x96 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n13630 = x95 &  n5384 ;
  assign n13631 = n13629 | n13630 ;
  assign n13633 = ( x94 & ~n13632 ) | ( x94 & n13631 ) | ( ~n13632 & n13631 ) ;
  assign n13634 = ( n2836 & ~n5392 ) | ( n2836 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n13635 = n13633 | n13634 ;
  assign n13636 = ( x47 & ~n13635 ) | ( x47 & 1'b0 ) | ( ~n13635 & 1'b0 ) ;
  assign n13637 = ~x47 & n13635 ;
  assign n13638 = n13636 | n13637 ;
  assign n13639 = ( n13557 & n13628 ) | ( n13557 & n13638 ) | ( n13628 & n13638 ) ;
  assign n13640 = ( n13628 & ~n13557 ) | ( n13628 & n13638 ) | ( ~n13557 & n13638 ) ;
  assign n13641 = ( n13557 & ~n13639 ) | ( n13557 & n13640 ) | ( ~n13639 & n13640 ) ;
  assign n13652 = ( n13409 & ~n13651 ) | ( n13409 & n13641 ) | ( ~n13651 & n13641 ) ;
  assign n13653 = ( n13641 & ~n13409 ) | ( n13641 & n13651 ) | ( ~n13409 & n13651 ) ;
  assign n13654 = ( n13652 & ~n13641 ) | ( n13652 & n13653 ) | ( ~n13641 & n13653 ) ;
  assign n13665 = ( n13412 & ~n13664 ) | ( n13412 & n13654 ) | ( ~n13664 & n13654 ) ;
  assign n13666 = ( n13412 & ~n13654 ) | ( n13412 & n13664 ) | ( ~n13654 & n13664 ) ;
  assign n13667 = ( n13665 & ~n13412 ) | ( n13665 & n13666 ) | ( ~n13412 & n13666 ) ;
  assign n13669 = ( n13415 & n13556 ) | ( n13415 & n13667 ) | ( n13556 & n13667 ) ;
  assign n13668 = ( n13556 & ~n13415 ) | ( n13556 & n13667 ) | ( ~n13415 & n13667 ) ;
  assign n13670 = ( n13415 & ~n13669 ) | ( n13415 & n13668 ) | ( ~n13669 & n13668 ) ;
  assign n13671 = ( n13418 & ~n13546 ) | ( n13418 & n13670 ) | ( ~n13546 & n13670 ) ;
  assign n13672 = ( n13418 & ~n13670 ) | ( n13418 & n13546 ) | ( ~n13670 & n13546 ) ;
  assign n13673 = ( n13671 & ~n13418 ) | ( n13671 & n13672 ) | ( ~n13418 & n13672 ) ;
  assign n13530 = x109 &  n2718 ;
  assign n13527 = ( x111 & ~n2642 ) | ( x111 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n13528 = x110 &  n2637 ;
  assign n13529 = n13527 | n13528 ;
  assign n13531 = ( x109 & ~n13530 ) | ( x109 & n13529 ) | ( ~n13530 & n13529 ) ;
  assign n13532 = ( n2645 & ~n5711 ) | ( n2645 & n13531 ) | ( ~n5711 & n13531 ) ;
  assign n13533 = n5711 | n13532 ;
  assign n13535 = ( x32 & n13531 ) | ( x32 & n13533 ) | ( n13531 & n13533 ) ;
  assign n13534 = ( x32 & ~n13533 ) | ( x32 & n13531 ) | ( ~n13533 & n13531 ) ;
  assign n13536 = ( n13533 & ~n13535 ) | ( n13533 & n13534 ) | ( ~n13535 & n13534 ) ;
  assign n13674 = ( n13421 & ~n13673 ) | ( n13421 & n13536 ) | ( ~n13673 & n13536 ) ;
  assign n13675 = ( n13536 & ~n13421 ) | ( n13536 & n13673 ) | ( ~n13421 & n13673 ) ;
  assign n13676 = ( n13674 & ~n13536 ) | ( n13674 & n13675 ) | ( ~n13536 & n13675 ) ;
  assign n13680 = x112 &  n2312 ;
  assign n13677 = ( x114 & ~n2195 ) | ( x114 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n13678 = x113 &  n2190 ;
  assign n13679 = n13677 | n13678 ;
  assign n13681 = ( x112 & ~n13680 ) | ( x112 & n13679 ) | ( ~n13680 & n13679 ) ;
  assign n13682 = ( n2198 & ~n6185 ) | ( n2198 & n13681 ) | ( ~n6185 & n13681 ) ;
  assign n13683 = n6185 | n13682 ;
  assign n13685 = ( x29 & n13681 ) | ( x29 & n13683 ) | ( n13681 & n13683 ) ;
  assign n13684 = ( x29 & ~n13683 ) | ( x29 & n13681 ) | ( ~n13683 & n13681 ) ;
  assign n13686 = ( n13683 & ~n13685 ) | ( n13683 & n13684 ) | ( ~n13685 & n13684 ) ;
  assign n13687 = ( n13526 & ~n13676 ) | ( n13526 & n13686 ) | ( ~n13676 & n13686 ) ;
  assign n13688 = ( n13526 & ~n13686 ) | ( n13526 & n13676 ) | ( ~n13686 & n13676 ) ;
  assign n13689 = ( n13687 & ~n13526 ) | ( n13687 & n13688 ) | ( ~n13526 & n13688 ) ;
  assign n13690 = ( n13515 & ~n13525 ) | ( n13515 & n13689 ) | ( ~n13525 & n13689 ) ;
  assign n13691 = ( n13515 & ~n13689 ) | ( n13515 & n13525 ) | ( ~n13689 & n13525 ) ;
  assign n13692 = ( n13690 & ~n13515 ) | ( n13690 & n13691 ) | ( ~n13515 & n13691 ) ;
  assign n13693 = ( n13514 & ~n13692 ) | ( n13514 & 1'b0 ) | ( ~n13692 & 1'b0 ) ;
  assign n13694 = ~n13514 & n13692 ;
  assign n13695 = n13693 | n13694 ;
  assign n13696 = ( n13256 & ~n13451 ) | ( n13256 & n13266 ) | ( ~n13451 & n13266 ) ;
  assign n13697 = ( n13503 & n13695 ) | ( n13503 & n13696 ) | ( n13695 & n13696 ) ;
  assign n13698 = ( n13695 & ~n13503 ) | ( n13695 & n13696 ) | ( ~n13503 & n13696 ) ;
  assign n13699 = ( n13503 & ~n13697 ) | ( n13503 & n13698 ) | ( ~n13697 & n13698 ) ;
  assign n13703 = x124 &  n942 ;
  assign n13700 = ( x126 & ~n896 ) | ( x126 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n13701 = x125 &  n891 ;
  assign n13702 = n13700 | n13701 ;
  assign n13704 = ( x124 & ~n13703 ) | ( x124 & n13702 ) | ( ~n13703 & n13702 ) ;
  assign n13705 = ( n899 & ~n9349 ) | ( n899 & n13704 ) | ( ~n9349 & n13704 ) ;
  assign n13706 = n9349 | n13705 ;
  assign n13708 = ( x17 & n13704 ) | ( x17 & n13706 ) | ( n13704 & n13706 ) ;
  assign n13707 = ( x17 & ~n13706 ) | ( x17 & n13704 ) | ( ~n13706 & n13704 ) ;
  assign n13709 = ( n13706 & ~n13708 ) | ( n13706 & n13707 ) | ( ~n13708 & n13707 ) ;
  assign n13710 = ( n13493 & ~n13699 ) | ( n13493 & n13709 ) | ( ~n13699 & n13709 ) ;
  assign n13711 = ( n13493 & ~n13709 ) | ( n13493 & n13699 ) | ( ~n13709 & n13699 ) ;
  assign n13712 = ( n13710 & ~n13493 ) | ( n13710 & n13711 ) | ( ~n13493 & n13711 ) ;
  assign n13492 = ( n13242 & n13252 ) | ( n13242 & n13467 ) | ( n13252 & n13467 ) ;
  assign n13713 = ( n13491 & ~n13712 ) | ( n13491 & n13492 ) | ( ~n13712 & n13492 ) ;
  assign n13714 = ( n13491 & ~n13492 ) | ( n13491 & n13712 ) | ( ~n13492 & n13712 ) ;
  assign n13715 = ( n13713 & ~n13491 ) | ( n13713 & n13714 ) | ( ~n13491 & n13714 ) ;
  assign n13485 = ( n13239 & n13470 ) | ( n13239 & n13478 ) | ( n13470 & n13478 ) ;
  assign n13716 = ( n13483 & ~n13715 ) | ( n13483 & n13485 ) | ( ~n13715 & n13485 ) ;
  assign n13717 = ( n13485 & ~n13483 ) | ( n13485 & n13715 ) | ( ~n13483 & n13715 ) ;
  assign n13718 = ( n13716 & ~n13485 ) | ( n13716 & n13717 ) | ( ~n13485 & n13717 ) ;
  assign n13719 = ( n13493 & n13699 ) | ( n13493 & n13709 ) | ( n13699 & n13709 ) ;
  assign n13728 = ( x23 & ~n13510 ) | ( x23 & 1'b0 ) | ( ~n13510 & 1'b0 ) ;
  assign n13729 = ~x23 & n13510 ;
  assign n13730 = n13728 | n13729 ;
  assign n13731 = ( n13511 & ~n13692 ) | ( n13511 & n13730 ) | ( ~n13692 & n13730 ) ;
  assign n13743 = x113 &  n2312 ;
  assign n13740 = ( x115 & ~n2195 ) | ( x115 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n13741 = x114 &  n2190 ;
  assign n13742 = n13740 | n13741 ;
  assign n13744 = ( x113 & ~n13743 ) | ( x113 & n13742 ) | ( ~n13743 & n13742 ) ;
  assign n13745 = ~n2198 & n6420 ;
  assign n13746 = n13744 | n13745 ;
  assign n13747 = ( x29 & ~n13746 ) | ( x29 & 1'b0 ) | ( ~n13746 & 1'b0 ) ;
  assign n13748 = ~x29 & n13746 ;
  assign n13749 = n13747 | n13748 ;
  assign n13753 = x107 &  n3214 ;
  assign n13750 = ( x109 & ~n3087 ) | ( x109 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n13751 = x108 &  n3082 ;
  assign n13752 = n13750 | n13751 ;
  assign n13754 = ( x107 & ~n13753 ) | ( x107 & n13752 ) | ( ~n13753 & n13752 ) ;
  assign n13755 = ~n3090 & n5267 ;
  assign n13756 = n13754 | n13755 ;
  assign n13757 = ( x35 & ~n13756 ) | ( x35 & 1'b0 ) | ( ~n13756 & 1'b0 ) ;
  assign n13758 = ~x35 & n13756 ;
  assign n13759 = n13757 | n13758 ;
  assign n13879 = x104 &  n3756 ;
  assign n13876 = ( x106 & ~n3602 ) | ( x106 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n13877 = x105 &  n3597 ;
  assign n13878 = n13876 | n13877 ;
  assign n13880 = ( x104 & ~n13879 ) | ( x104 & n13878 ) | ( ~n13879 & n13878 ) ;
  assign n13881 = ~n3605 & n4458 ;
  assign n13882 = n13880 | n13881 ;
  assign n13883 = ( x38 & ~n13882 ) | ( x38 & 1'b0 ) | ( ~n13882 & 1'b0 ) ;
  assign n13884 = ~x38 & n13882 ;
  assign n13885 = n13883 | n13884 ;
  assign n13763 = x92 &  n6288 ;
  assign n13760 = ( x94 & ~n6032 ) | ( x94 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n13761 = x93 &  n6027 ;
  assign n13762 = n13760 | n13761 ;
  assign n13764 = ( x92 & ~n13763 ) | ( x92 & n13762 ) | ( ~n13763 & n13762 ) ;
  assign n13765 = ( n2401 & ~n6035 ) | ( n2401 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n13766 = n13764 | n13765 ;
  assign n13767 = ( x50 & ~n13766 ) | ( x50 & 1'b0 ) | ( ~n13766 & 1'b0 ) ;
  assign n13768 = ~x50 & n13766 ;
  assign n13769 = n13767 | n13768 ;
  assign n13773 = x89 &  n6982 ;
  assign n13770 = ( x91 & ~n6727 ) | ( x91 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n13771 = x90 &  n6722 ;
  assign n13772 = n13770 | n13771 ;
  assign n13774 = ( x89 & ~n13773 ) | ( x89 & n13772 ) | ( ~n13773 & n13772 ) ;
  assign n13775 = ( n2108 & ~n6730 ) | ( n2108 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n13776 = n13774 | n13775 ;
  assign n13777 = ( x53 & ~n13776 ) | ( x53 & 1'b0 ) | ( ~n13776 & 1'b0 ) ;
  assign n13778 = ~x53 & n13776 ;
  assign n13779 = n13777 | n13778 ;
  assign n13783 = x83 &  n8558 ;
  assign n13780 = ( x85 & ~n8314 ) | ( x85 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n13781 = x84 &  n8309 ;
  assign n13782 = n13780 | n13781 ;
  assign n13784 = ( x83 & ~n13783 ) | ( x83 & n13782 ) | ( ~n13783 & n13782 ) ;
  assign n13785 = ( n1295 & ~n8317 ) | ( n1295 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n13786 = n13784 | n13785 ;
  assign n13787 = ( x59 & ~n13786 ) | ( x59 & 1'b0 ) | ( ~n13786 & 1'b0 ) ;
  assign n13788 = ~x59 & n13786 ;
  assign n13789 = n13787 | n13788 ;
  assign n13793 = x80 &  n9457 ;
  assign n13790 = ( x82 & ~n9150 ) | ( x82 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n13791 = x81 &  n9145 ;
  assign n13792 = n13790 | n13791 ;
  assign n13794 = ( x80 & ~n13793 ) | ( x80 & n13792 ) | ( ~n13793 & n13792 ) ;
  assign n13795 = ( n1084 & ~n9153 ) | ( n1084 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n13796 = n13794 | n13795 ;
  assign n13797 = ( x62 & ~n13796 ) | ( x62 & 1'b0 ) | ( ~n13796 & 1'b0 ) ;
  assign n13798 = ~x62 & n13796 ;
  assign n13799 = n13797 | n13798 ;
  assign n13800 = x78 &  n10104 ;
  assign n13801 = ( x79 & ~n9760 ) | ( x79 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n13802 = n13800 | n13801 ;
  assign n13803 = ( x14 & n13342 ) | ( x14 & n13802 ) | ( n13342 & n13802 ) ;
  assign n13804 = ( x14 & ~n13342 ) | ( x14 & n13802 ) | ( ~n13342 & n13802 ) ;
  assign n13805 = ( n13342 & ~n13803 ) | ( n13342 & n13804 ) | ( ~n13803 & n13804 ) ;
  assign n13806 = ( n13583 & n13799 ) | ( n13583 & n13805 ) | ( n13799 & n13805 ) ;
  assign n13807 = ( n13583 & ~n13799 ) | ( n13583 & n13805 ) | ( ~n13799 & n13805 ) ;
  assign n13808 = ( n13799 & ~n13806 ) | ( n13799 & n13807 ) | ( ~n13806 & n13807 ) ;
  assign n13809 = ( n13353 & ~n13585 ) | ( n13353 & n13595 ) | ( ~n13585 & n13595 ) ;
  assign n13810 = ( n13789 & ~n13808 ) | ( n13789 & n13809 ) | ( ~n13808 & n13809 ) ;
  assign n13811 = ( n13789 & ~n13809 ) | ( n13789 & n13808 ) | ( ~n13809 & n13808 ) ;
  assign n13812 = ( n13810 & ~n13789 ) | ( n13810 & n13811 ) | ( ~n13789 & n13811 ) ;
  assign n13813 = ( n13569 & ~n13598 ) | ( n13569 & n13608 ) | ( ~n13598 & n13608 ) ;
  assign n13817 = x86 &  n7731 ;
  assign n13814 = ( x88 & ~n7538 ) | ( x88 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n13815 = x87 &  n7533 ;
  assign n13816 = n13814 | n13815 ;
  assign n13818 = ( x86 & ~n13817 ) | ( x86 & n13816 ) | ( ~n13817 & n13816 ) ;
  assign n13819 = ( n1624 & ~n7541 ) | ( n1624 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n13820 = n13818 | n13819 ;
  assign n13821 = ( x56 & ~n13820 ) | ( x56 & 1'b0 ) | ( ~n13820 & 1'b0 ) ;
  assign n13822 = ~x56 & n13820 ;
  assign n13823 = n13821 | n13822 ;
  assign n13824 = ( n13812 & ~n13813 ) | ( n13812 & n13823 ) | ( ~n13813 & n13823 ) ;
  assign n13825 = ( n13812 & ~n13823 ) | ( n13812 & n13813 ) | ( ~n13823 & n13813 ) ;
  assign n13826 = ( n13824 & ~n13812 ) | ( n13824 & n13825 ) | ( ~n13812 & n13825 ) ;
  assign n13827 = ( n13613 & n13779 ) | ( n13613 & n13826 ) | ( n13779 & n13826 ) ;
  assign n13828 = ( n13613 & ~n13779 ) | ( n13613 & n13826 ) | ( ~n13779 & n13826 ) ;
  assign n13829 = ( n13779 & ~n13827 ) | ( n13779 & n13828 ) | ( ~n13827 & n13828 ) ;
  assign n13830 = ( n13614 & n13615 ) | ( n13614 & n13625 ) | ( n13615 & n13625 ) ;
  assign n13832 = ( n13769 & n13829 ) | ( n13769 & n13830 ) | ( n13829 & n13830 ) ;
  assign n13831 = ( n13829 & ~n13769 ) | ( n13829 & n13830 ) | ( ~n13769 & n13830 ) ;
  assign n13833 = ( n13769 & ~n13832 ) | ( n13769 & n13831 ) | ( ~n13832 & n13831 ) ;
  assign n13838 = x95 &  n5586 ;
  assign n13835 = ( x97 & ~n5389 ) | ( x97 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n13836 = x96 &  n5384 ;
  assign n13837 = n13835 | n13836 ;
  assign n13839 = ( x95 & ~n13838 ) | ( x95 & n13837 ) | ( ~n13838 & n13837 ) ;
  assign n13840 = ( n2999 & ~n5392 ) | ( n2999 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n13841 = n13839 | n13840 ;
  assign n13842 = ( x47 & ~n13841 ) | ( x47 & 1'b0 ) | ( ~n13841 & 1'b0 ) ;
  assign n13843 = ~x47 & n13841 ;
  assign n13844 = n13842 | n13843 ;
  assign n13834 = ( n13557 & ~n13628 ) | ( n13557 & n13638 ) | ( ~n13628 & n13638 ) ;
  assign n13845 = ( n13833 & ~n13844 ) | ( n13833 & n13834 ) | ( ~n13844 & n13834 ) ;
  assign n13846 = ( n13833 & ~n13834 ) | ( n13833 & n13844 ) | ( ~n13834 & n13844 ) ;
  assign n13847 = ( n13845 & ~n13833 ) | ( n13845 & n13846 ) | ( ~n13833 & n13846 ) ;
  assign n13848 = ( n13409 & ~n13641 ) | ( n13409 & n13651 ) | ( ~n13641 & n13651 ) ;
  assign n13852 = x98 &  n4934 ;
  assign n13849 = ( x100 & ~n4725 ) | ( x100 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n13850 = x99 &  n4720 ;
  assign n13851 = n13849 | n13850 ;
  assign n13853 = ( x98 & ~n13852 ) | ( x98 & n13851 ) | ( ~n13852 & n13851 ) ;
  assign n13854 = n3354 | n4728 ;
  assign n13855 = ~n13853 & n13854 ;
  assign n13856 = x44 &  n13855 ;
  assign n13857 = x44 | n13855 ;
  assign n13858 = ~n13856 & n13857 ;
  assign n13860 = ( n13847 & n13848 ) | ( n13847 & n13858 ) | ( n13848 & n13858 ) ;
  assign n13859 = ( n13848 & ~n13847 ) | ( n13848 & n13858 ) | ( ~n13847 & n13858 ) ;
  assign n13861 = ( n13847 & ~n13860 ) | ( n13847 & n13859 ) | ( ~n13860 & n13859 ) ;
  assign n13866 = x101 &  n4344 ;
  assign n13863 = ( x103 & ~n4143 ) | ( x103 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n13864 = x102 &  n4138 ;
  assign n13865 = n13863 | n13864 ;
  assign n13867 = ( x101 & ~n13866 ) | ( x101 & n13865 ) | ( ~n13866 & n13865 ) ;
  assign n13868 = n4056 | n4146 ;
  assign n13869 = ~n13867 & n13868 ;
  assign n13870 = x41 &  n13869 ;
  assign n13871 = x41 | n13869 ;
  assign n13872 = ~n13870 & n13871 ;
  assign n13862 = ( n13654 & ~n13412 ) | ( n13654 & n13664 ) | ( ~n13412 & n13664 ) ;
  assign n13873 = ( n13861 & ~n13872 ) | ( n13861 & n13862 ) | ( ~n13872 & n13862 ) ;
  assign n13874 = ( n13861 & ~n13862 ) | ( n13861 & n13872 ) | ( ~n13862 & n13872 ) ;
  assign n13875 = ( n13873 & ~n13861 ) | ( n13873 & n13874 ) | ( ~n13861 & n13874 ) ;
  assign n13886 = ( n13669 & ~n13885 ) | ( n13669 & n13875 ) | ( ~n13885 & n13875 ) ;
  assign n13887 = ( n13875 & ~n13669 ) | ( n13875 & n13885 ) | ( ~n13669 & n13885 ) ;
  assign n13888 = ( n13886 & ~n13875 ) | ( n13886 & n13887 ) | ( ~n13875 & n13887 ) ;
  assign n13890 = ( n13672 & n13759 ) | ( n13672 & n13888 ) | ( n13759 & n13888 ) ;
  assign n13889 = ( n13672 & ~n13759 ) | ( n13672 & n13888 ) | ( ~n13759 & n13888 ) ;
  assign n13891 = ( n13759 & ~n13890 ) | ( n13759 & n13889 ) | ( ~n13890 & n13889 ) ;
  assign n13900 = x32 | n13891 ;
  assign n13901 = ~x32 & n13891 ;
  assign n13902 = ( n13900 & ~n13891 ) | ( n13900 & n13901 ) | ( ~n13891 & n13901 ) ;
  assign n13892 = ( n13421 & ~n13536 ) | ( n13421 & n13673 ) | ( ~n13536 & n13673 ) ;
  assign n13896 = x110 &  n2718 ;
  assign n13893 = ( x112 & ~n2642 ) | ( x112 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n13894 = x111 &  n2637 ;
  assign n13895 = n13893 | n13894 ;
  assign n13897 = ( x110 & ~n13896 ) | ( x110 & n13895 ) | ( ~n13896 & n13895 ) ;
  assign n13898 = ~n2645 & n5727 ;
  assign n13899 = n13897 | n13898 ;
  assign n13904 = ( n13892 & n13899 ) | ( n13892 & n13902 ) | ( n13899 & n13902 ) ;
  assign n13903 = ( n13892 & ~n13902 ) | ( n13892 & n13899 ) | ( ~n13902 & n13899 ) ;
  assign n13905 = ( n13902 & ~n13904 ) | ( n13902 & n13903 ) | ( ~n13904 & n13903 ) ;
  assign n13906 = ( n13526 & n13676 ) | ( n13526 & n13686 ) | ( n13676 & n13686 ) ;
  assign n13908 = ( n13749 & n13905 ) | ( n13749 & n13906 ) | ( n13905 & n13906 ) ;
  assign n13907 = ( n13905 & ~n13749 ) | ( n13905 & n13906 ) | ( ~n13749 & n13906 ) ;
  assign n13909 = ( n13749 & ~n13908 ) | ( n13749 & n13907 ) | ( ~n13908 & n13907 ) ;
  assign n13739 = ( n13515 & n13525 ) | ( n13515 & n13689 ) | ( n13525 & n13689 ) ;
  assign n13735 = x116 &  n1894 ;
  assign n13732 = ( x118 & ~n1816 ) | ( x118 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n13733 = x117 &  n1811 ;
  assign n13734 = n13732 | n13733 ;
  assign n13736 = ( x116 & ~n13735 ) | ( x116 & n13734 ) | ( ~n13735 & n13734 ) ;
  assign n13737 = n1819 | n7152 ;
  assign n13738 = ~n13736 & n13737 ;
  assign n13910 = ~x26 & n13738 ;
  assign n13911 = x26 | n13738 ;
  assign n13912 = ( n13910 & ~n13738 ) | ( n13910 & n13911 ) | ( ~n13738 & n13911 ) ;
  assign n13913 = ( n13909 & ~n13739 ) | ( n13909 & n13912 ) | ( ~n13739 & n13912 ) ;
  assign n13914 = ( n13739 & ~n13909 ) | ( n13739 & n13912 ) | ( ~n13909 & n13912 ) ;
  assign n13915 = ( n13913 & ~n13912 ) | ( n13913 & n13914 ) | ( ~n13912 & n13914 ) ;
  assign n13919 = x119 &  n1551 ;
  assign n13916 = ( x121 & ~n1451 ) | ( x121 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n13917 = x120 &  n1446 ;
  assign n13918 = n13916 | n13917 ;
  assign n13920 = ( x119 & ~n13919 ) | ( x119 & n13918 ) | ( ~n13919 & n13918 ) ;
  assign n13921 = ~n1454 & n8176 ;
  assign n13922 = n13920 | n13921 ;
  assign n13923 = ( x23 & ~n13922 ) | ( x23 & 1'b0 ) | ( ~n13922 & 1'b0 ) ;
  assign n13924 = ~x23 & n13922 ;
  assign n13925 = n13923 | n13924 ;
  assign n13926 = ( n13731 & n13915 ) | ( n13731 & n13925 ) | ( n13915 & n13925 ) ;
  assign n13927 = ( n13915 & ~n13731 ) | ( n13915 & n13925 ) | ( ~n13731 & n13925 ) ;
  assign n13928 = ( n13731 & ~n13926 ) | ( n13731 & n13927 ) | ( ~n13926 & n13927 ) ;
  assign n13727 = ( n13503 & ~n13695 ) | ( n13503 & n13696 ) | ( ~n13695 & n13696 ) ;
  assign n13723 = x122 &  n1227 ;
  assign n13720 = ( x124 & ~n1154 ) | ( x124 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n13721 = x123 &  n1149 ;
  assign n13722 = n13720 | n13721 ;
  assign n13724 = ( x122 & ~n13723 ) | ( x122 & n13722 ) | ( ~n13723 & n13722 ) ;
  assign n13725 = ~n1157 & n8755 ;
  assign n13726 = n13724 | n13725 ;
  assign n13929 = x20 | n13726 ;
  assign n13930 = ~x20 & n13726 ;
  assign n13931 = ( n13929 & ~n13726 ) | ( n13929 & n13930 ) | ( ~n13726 & n13930 ) ;
  assign n13932 = ( n13928 & ~n13727 ) | ( n13928 & n13931 ) | ( ~n13727 & n13931 ) ;
  assign n13933 = ( n13727 & ~n13928 ) | ( n13727 & n13931 ) | ( ~n13928 & n13931 ) ;
  assign n13934 = ( n13932 & ~n13931 ) | ( n13932 & n13933 ) | ( ~n13931 & n13933 ) ;
  assign n13938 = x125 &  n942 ;
  assign n13935 = ( x127 & ~n896 ) | ( x127 & 1'b0 ) | ( ~n896 & 1'b0 ) ;
  assign n13936 = x126 &  n891 ;
  assign n13937 = n13935 | n13936 ;
  assign n13939 = ( x125 & ~n13938 ) | ( x125 & n13937 ) | ( ~n13938 & n13937 ) ;
  assign n13940 = n899 | n9941 ;
  assign n13941 = ~n13939 & n13940 ;
  assign n13942 = x17 &  n13941 ;
  assign n13943 = x17 | n13941 ;
  assign n13944 = ~n13942 & n13943 ;
  assign n13945 = ( n13719 & ~n13934 ) | ( n13719 & n13944 ) | ( ~n13934 & n13944 ) ;
  assign n13946 = ( n13719 & ~n13944 ) | ( n13719 & n13934 ) | ( ~n13944 & n13934 ) ;
  assign n13947 = ( n13945 & ~n13719 ) | ( n13945 & n13946 ) | ( ~n13719 & n13946 ) ;
  assign n13949 = ( n13714 & n13717 ) | ( n13714 & n13947 ) | ( n13717 & n13947 ) ;
  assign n13948 = ( n13717 & ~n13714 ) | ( n13717 & n13947 ) | ( ~n13714 & n13947 ) ;
  assign n13950 = ( n13714 & ~n13949 ) | ( n13714 & n13948 ) | ( ~n13949 & n13948 ) ;
  assign n13951 = ( n13719 & n13934 ) | ( n13719 & n13944 ) | ( n13934 & n13944 ) ;
  assign n13952 = x20 &  n13726 ;
  assign n13953 = ( n13929 & ~n13952 ) | ( n13929 & 1'b0 ) | ( ~n13952 & 1'b0 ) ;
  assign n13954 = ( n13727 & ~n13928 ) | ( n13727 & n13953 ) | ( ~n13928 & n13953 ) ;
  assign n13962 = ( n13731 & ~n13915 ) | ( n13731 & n13925 ) | ( ~n13915 & n13925 ) ;
  assign n13958 = x123 &  n1227 ;
  assign n13955 = ( x125 & ~n1154 ) | ( x125 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n13956 = x124 &  n1149 ;
  assign n13957 = n13955 | n13956 ;
  assign n13959 = ( x123 & ~n13958 ) | ( x123 & n13957 ) | ( ~n13958 & n13957 ) ;
  assign n13960 = ~n1157 & n9324 ;
  assign n13961 = n13959 | n13960 ;
  assign n13963 = ( x20 & n13961 ) | ( x20 & n13962 ) | ( n13961 & n13962 ) ;
  assign n13964 = ( x20 & ~n13962 ) | ( x20 & n13961 ) | ( ~n13962 & n13961 ) ;
  assign n13965 = ( n13962 & ~n13963 ) | ( n13962 & n13964 ) | ( ~n13963 & n13964 ) ;
  assign n13966 = x26 &  n13738 ;
  assign n13967 = ( n13911 & ~n13966 ) | ( n13911 & 1'b0 ) | ( ~n13966 & 1'b0 ) ;
  assign n13968 = ( n13739 & n13909 ) | ( n13739 & n13967 ) | ( n13909 & n13967 ) ;
  assign n13972 = x117 &  n1894 ;
  assign n13969 = ( x119 & ~n1816 ) | ( x119 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n13970 = x118 &  n1811 ;
  assign n13971 = n13969 | n13970 ;
  assign n13973 = ( x117 & ~n13972 ) | ( x117 & n13971 ) | ( ~n13972 & n13971 ) ;
  assign n13974 = ~n1819 & n7648 ;
  assign n13975 = n13973 | n13974 ;
  assign n13976 = ( n13749 & ~n13906 ) | ( n13749 & n13905 ) | ( ~n13906 & n13905 ) ;
  assign n13977 = ( x26 & n13975 ) | ( x26 & n13976 ) | ( n13975 & n13976 ) ;
  assign n13978 = ( x26 & ~n13975 ) | ( x26 & n13976 ) | ( ~n13975 & n13976 ) ;
  assign n13979 = ( n13975 & ~n13977 ) | ( n13975 & n13978 ) | ( ~n13977 & n13978 ) ;
  assign n13983 = x114 &  n2312 ;
  assign n13980 = ( x116 & ~n2195 ) | ( x116 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n13981 = x115 &  n2190 ;
  assign n13982 = n13980 | n13981 ;
  assign n13984 = ( x114 & ~n13983 ) | ( x114 & n13982 ) | ( ~n13983 & n13982 ) ;
  assign n13985 = n2198 | n6885 ;
  assign n13986 = ~n13984 & n13985 ;
  assign n13987 = x29 &  n13986 ;
  assign n13988 = x29 | n13986 ;
  assign n13989 = ~n13987 & n13988 ;
  assign n14144 = ( x32 & ~n13899 ) | ( x32 & 1'b0 ) | ( ~n13899 & 1'b0 ) ;
  assign n14145 = ~x32 & n13899 ;
  assign n14146 = n14144 | n14145 ;
  assign n14147 = ( n13891 & n13892 ) | ( n13891 & n14146 ) | ( n13892 & n14146 ) ;
  assign n14138 = x32 | n13889 ;
  assign n14139 = ~x32 & n13889 ;
  assign n14140 = ( n14138 & ~n13889 ) | ( n14138 & n14139 ) | ( ~n13889 & n14139 ) ;
  assign n13993 = x111 &  n2718 ;
  assign n13990 = ( x113 & ~n2642 ) | ( x113 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n13991 = x112 &  n2637 ;
  assign n13992 = n13990 | n13991 ;
  assign n13994 = ( x111 & ~n13993 ) | ( x111 & n13992 ) | ( ~n13993 & n13992 ) ;
  assign n13995 = n2645 | n6169 ;
  assign n13996 = ~n13994 & n13995 ;
  assign n13997 = ( n13669 & ~n13875 ) | ( n13669 & n13885 ) | ( ~n13875 & n13885 ) ;
  assign n14128 = x108 &  n3214 ;
  assign n14125 = ( x110 & ~n3087 ) | ( x110 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n14126 = x109 &  n3082 ;
  assign n14127 = n14125 | n14126 ;
  assign n14129 = ( x108 & ~n14128 ) | ( x108 & n14127 ) | ( ~n14128 & n14127 ) ;
  assign n14130 = n3090 | n5283 ;
  assign n14131 = ~n14129 & n14130 ;
  assign n14132 = x35 &  n14131 ;
  assign n14133 = x35 | n14131 ;
  assign n14134 = ~n14132 & n14133 ;
  assign n13998 = ( n13861 & n13862 ) | ( n13861 & n13872 ) | ( n13862 & n13872 ) ;
  assign n14002 = x105 &  n3756 ;
  assign n13999 = ( x107 & ~n3602 ) | ( x107 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n14000 = x106 &  n3597 ;
  assign n14001 = n13999 | n14000 ;
  assign n14003 = ( x105 & ~n14002 ) | ( x105 & n14001 ) | ( ~n14002 & n14001 ) ;
  assign n14004 = ~n3605 & n4848 ;
  assign n14005 = n14003 | n14004 ;
  assign n14006 = ( x38 & ~n14005 ) | ( x38 & 1'b0 ) | ( ~n14005 & 1'b0 ) ;
  assign n14007 = ~x38 & n14005 ;
  assign n14008 = n14006 | n14007 ;
  assign n14009 = ( n13847 & ~n13858 ) | ( n13847 & n13848 ) | ( ~n13858 & n13848 ) ;
  assign n14013 = x102 &  n4344 ;
  assign n14010 = ( x104 & ~n4143 ) | ( x104 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n14011 = x103 &  n4138 ;
  assign n14012 = n14010 | n14011 ;
  assign n14014 = ( x102 & ~n14013 ) | ( x102 & n14012 ) | ( ~n14013 & n14012 ) ;
  assign n14015 = n4146 | n4249 ;
  assign n14016 = ~n14014 & n14015 ;
  assign n14017 = x41 &  n14016 ;
  assign n14018 = x41 | n14016 ;
  assign n14019 = ~n14017 & n14018 ;
  assign n14020 = ( n13833 & n13834 ) | ( n13833 & n13844 ) | ( n13834 & n13844 ) ;
  assign n14032 = ( n13342 & ~x14 ) | ( n13342 & n13802 ) | ( ~x14 & n13802 ) ;
  assign n14033 = x79 &  n10104 ;
  assign n14034 = ( x80 & ~n9760 ) | ( x80 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n14035 = n14033 | n14034 ;
  assign n14039 = x81 &  n9457 ;
  assign n14036 = ( x83 & ~n9150 ) | ( x83 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n14037 = x82 &  n9145 ;
  assign n14038 = n14036 | n14037 ;
  assign n14040 = ( x81 & ~n14039 ) | ( x81 & n14038 ) | ( ~n14039 & n14038 ) ;
  assign n14041 = ( n1100 & ~n14040 ) | ( n1100 & n9153 ) | ( ~n14040 & n9153 ) ;
  assign n14042 = ~n9153 & n14041 ;
  assign n14043 = ( x62 & n14040 ) | ( x62 & n14042 ) | ( n14040 & n14042 ) ;
  assign n14044 = ( x62 & ~n14042 ) | ( x62 & n14040 ) | ( ~n14042 & n14040 ) ;
  assign n14045 = ( n14042 & ~n14043 ) | ( n14042 & n14044 ) | ( ~n14043 & n14044 ) ;
  assign n14046 = ( n14032 & ~n14035 ) | ( n14032 & n14045 ) | ( ~n14035 & n14045 ) ;
  assign n14047 = ( n14032 & ~n14045 ) | ( n14032 & n14035 ) | ( ~n14045 & n14035 ) ;
  assign n14048 = ( n14046 & ~n14032 ) | ( n14046 & n14047 ) | ( ~n14032 & n14047 ) ;
  assign n14052 = x84 &  n8558 ;
  assign n14049 = ( x86 & ~n8314 ) | ( x86 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n14050 = x85 &  n8309 ;
  assign n14051 = n14049 | n14050 ;
  assign n14053 = ( x84 & ~n14052 ) | ( x84 & n14051 ) | ( ~n14052 & n14051 ) ;
  assign n14054 = ( n1496 & ~n8317 ) | ( n1496 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n14055 = n14053 | n14054 ;
  assign n14031 = ( n13583 & ~n13805 ) | ( n13583 & n13799 ) | ( ~n13805 & n13799 ) ;
  assign n14056 = x59 | n14031 ;
  assign n14057 = ~x59 & n14031 ;
  assign n14058 = ( n14056 & ~n14031 ) | ( n14056 & n14057 ) | ( ~n14031 & n14057 ) ;
  assign n14059 = ( n14048 & ~n14055 ) | ( n14048 & n14058 ) | ( ~n14055 & n14058 ) ;
  assign n14060 = ( n14055 & ~n14048 ) | ( n14055 & n14058 ) | ( ~n14048 & n14058 ) ;
  assign n14061 = ( n14059 & ~n14058 ) | ( n14059 & n14060 ) | ( ~n14058 & n14060 ) ;
  assign n14065 = x87 &  n7731 ;
  assign n14062 = ( x89 & ~n7538 ) | ( x89 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n14063 = x88 &  n7533 ;
  assign n14064 = n14062 | n14063 ;
  assign n14066 = ( x87 & ~n14065 ) | ( x87 & n14064 ) | ( ~n14065 & n14064 ) ;
  assign n14067 = ( n1741 & ~n7541 ) | ( n1741 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n14068 = n14066 | n14067 ;
  assign n14069 = ( x56 & ~n14068 ) | ( x56 & 1'b0 ) | ( ~n14068 & 1'b0 ) ;
  assign n14070 = ~x56 & n14068 ;
  assign n14071 = n14069 | n14070 ;
  assign n14072 = ( n13810 & n14061 ) | ( n13810 & n14071 ) | ( n14061 & n14071 ) ;
  assign n14073 = ( n14061 & ~n13810 ) | ( n14061 & n14071 ) | ( ~n13810 & n14071 ) ;
  assign n14074 = ( n13810 & ~n14072 ) | ( n13810 & n14073 ) | ( ~n14072 & n14073 ) ;
  assign n14079 = x90 &  n6982 ;
  assign n14076 = ( x92 & ~n6727 ) | ( x92 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n14077 = x91 &  n6722 ;
  assign n14078 = n14076 | n14077 ;
  assign n14080 = ( x90 & ~n14079 ) | ( x90 & n14078 ) | ( ~n14079 & n14078 ) ;
  assign n14081 = ( n2248 & ~n6730 ) | ( n2248 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n14082 = n14080 | n14081 ;
  assign n14083 = ( x53 & ~n14082 ) | ( x53 & 1'b0 ) | ( ~n14082 & 1'b0 ) ;
  assign n14084 = ~x53 & n14082 ;
  assign n14085 = n14083 | n14084 ;
  assign n14075 = ( n13813 & ~n13812 ) | ( n13813 & n13823 ) | ( ~n13812 & n13823 ) ;
  assign n14086 = ( n14074 & ~n14085 ) | ( n14074 & n14075 ) | ( ~n14085 & n14075 ) ;
  assign n14087 = ( n14074 & ~n14075 ) | ( n14074 & n14085 ) | ( ~n14075 & n14085 ) ;
  assign n14088 = ( n14086 & ~n14074 ) | ( n14086 & n14087 ) | ( ~n14074 & n14087 ) ;
  assign n14092 = x93 &  n6288 ;
  assign n14089 = ( x95 & ~n6032 ) | ( x95 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n14090 = x94 &  n6027 ;
  assign n14091 = n14089 | n14090 ;
  assign n14093 = ( x93 & ~n14092 ) | ( x93 & n14091 ) | ( ~n14092 & n14091 ) ;
  assign n14094 = ( n2547 & ~n6035 ) | ( n2547 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n14095 = n14093 | n14094 ;
  assign n14096 = ( x50 & ~n14095 ) | ( x50 & 1'b0 ) | ( ~n14095 & 1'b0 ) ;
  assign n14097 = ~x50 & n14095 ;
  assign n14098 = n14096 | n14097 ;
  assign n14099 = ( n13613 & ~n13826 ) | ( n13613 & n13779 ) | ( ~n13826 & n13779 ) ;
  assign n14100 = ( n14088 & ~n14098 ) | ( n14088 & n14099 ) | ( ~n14098 & n14099 ) ;
  assign n14101 = ( n14088 & ~n14099 ) | ( n14088 & n14098 ) | ( ~n14099 & n14098 ) ;
  assign n14102 = ( n14100 & ~n14088 ) | ( n14100 & n14101 ) | ( ~n14088 & n14101 ) ;
  assign n14106 = x96 &  n5586 ;
  assign n14103 = ( x98 & ~n5389 ) | ( x98 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n14104 = x97 &  n5384 ;
  assign n14105 = n14103 | n14104 ;
  assign n14107 = ( x96 & ~n14106 ) | ( x96 & n14105 ) | ( ~n14106 & n14105 ) ;
  assign n14108 = ( n3170 & ~n5392 ) | ( n3170 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n14109 = n14107 | n14108 ;
  assign n14110 = ( x47 & ~n14109 ) | ( x47 & 1'b0 ) | ( ~n14109 & 1'b0 ) ;
  assign n14111 = ~x47 & n14109 ;
  assign n14112 = n14110 | n14111 ;
  assign n14114 = ( n13831 & n14102 ) | ( n13831 & n14112 ) | ( n14102 & n14112 ) ;
  assign n14113 = ( n14102 & ~n13831 ) | ( n14102 & n14112 ) | ( ~n13831 & n14112 ) ;
  assign n14115 = ( n13831 & ~n14114 ) | ( n13831 & n14113 ) | ( ~n14114 & n14113 ) ;
  assign n14024 = x99 &  n4934 ;
  assign n14021 = ( x101 & ~n4725 ) | ( x101 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n14022 = x100 &  n4720 ;
  assign n14023 = n14021 | n14022 ;
  assign n14025 = ( x99 & ~n14024 ) | ( x99 & n14023 ) | ( ~n14024 & n14023 ) ;
  assign n14026 = n3694 | n4728 ;
  assign n14027 = ~n14025 & n14026 ;
  assign n14028 = x44 &  n14027 ;
  assign n14029 = x44 | n14027 ;
  assign n14030 = ~n14028 & n14029 ;
  assign n14116 = ( n14020 & ~n14115 ) | ( n14020 & n14030 ) | ( ~n14115 & n14030 ) ;
  assign n14117 = ( n14020 & ~n14030 ) | ( n14020 & n14115 ) | ( ~n14030 & n14115 ) ;
  assign n14118 = ( n14116 & ~n14020 ) | ( n14116 & n14117 ) | ( ~n14020 & n14117 ) ;
  assign n14119 = ( n14009 & n14019 ) | ( n14009 & n14118 ) | ( n14019 & n14118 ) ;
  assign n14120 = ( n14019 & ~n14009 ) | ( n14019 & n14118 ) | ( ~n14009 & n14118 ) ;
  assign n14121 = ( n14009 & ~n14119 ) | ( n14009 & n14120 ) | ( ~n14119 & n14120 ) ;
  assign n14122 = ( n13998 & n14008 ) | ( n13998 & n14121 ) | ( n14008 & n14121 ) ;
  assign n14123 = ( n14008 & ~n13998 ) | ( n14008 & n14121 ) | ( ~n13998 & n14121 ) ;
  assign n14124 = ( n13998 & ~n14122 ) | ( n13998 & n14123 ) | ( ~n14122 & n14123 ) ;
  assign n14135 = ( n13997 & ~n14134 ) | ( n13997 & n14124 ) | ( ~n14134 & n14124 ) ;
  assign n14136 = ( n13997 & ~n14124 ) | ( n13997 & n14134 ) | ( ~n14124 & n14134 ) ;
  assign n14137 = ( n14135 & ~n13997 ) | ( n14135 & n14136 ) | ( ~n13997 & n14136 ) ;
  assign n14142 = ( n13996 & n14137 ) | ( n13996 & n14140 ) | ( n14137 & n14140 ) ;
  assign n14141 = ( n13996 & ~n14140 ) | ( n13996 & n14137 ) | ( ~n14140 & n14137 ) ;
  assign n14143 = ( n14140 & ~n14142 ) | ( n14140 & n14141 ) | ( ~n14142 & n14141 ) ;
  assign n14148 = ( n13989 & ~n14147 ) | ( n13989 & n14143 ) | ( ~n14147 & n14143 ) ;
  assign n14149 = ( n13989 & ~n14143 ) | ( n13989 & n14147 ) | ( ~n14143 & n14147 ) ;
  assign n14150 = ( n14148 & ~n13989 ) | ( n14148 & n14149 ) | ( ~n13989 & n14149 ) ;
  assign n14151 = ( n13979 & ~n14150 ) | ( n13979 & 1'b0 ) | ( ~n14150 & 1'b0 ) ;
  assign n14152 = ~n13979 & n14150 ;
  assign n14153 = n14151 | n14152 ;
  assign n14157 = x120 &  n1551 ;
  assign n14154 = ( x122 & ~n1451 ) | ( x122 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n14155 = x121 &  n1446 ;
  assign n14156 = n14154 | n14155 ;
  assign n14158 = ( x120 & ~n14157 ) | ( x120 & n14156 ) | ( ~n14157 & n14156 ) ;
  assign n14159 = ( n1454 & n9987 ) | ( n1454 & n14158 ) | ( n9987 & n14158 ) ;
  assign n14160 = ( n9987 & ~n14159 ) | ( n9987 & 1'b0 ) | ( ~n14159 & 1'b0 ) ;
  assign n14161 = ( x23 & n14158 ) | ( x23 & n14160 ) | ( n14158 & n14160 ) ;
  assign n14162 = ( x23 & ~n14160 ) | ( x23 & n14158 ) | ( ~n14160 & n14158 ) ;
  assign n14163 = ( n14160 & ~n14161 ) | ( n14160 & n14162 ) | ( ~n14161 & n14162 ) ;
  assign n14165 = ( n13968 & n14153 ) | ( n13968 & n14163 ) | ( n14153 & n14163 ) ;
  assign n14164 = ( n14153 & ~n13968 ) | ( n14153 & n14163 ) | ( ~n13968 & n14163 ) ;
  assign n14166 = ( n13968 & ~n14165 ) | ( n13968 & n14164 ) | ( ~n14165 & n14164 ) ;
  assign n14167 = n13965 &  n14166 ;
  assign n14168 = n13965 | n14166 ;
  assign n14169 = ~n14167 & n14168 ;
  assign n14170 = ( x126 & ~n942 ) | ( x126 & 1'b0 ) | ( ~n942 & 1'b0 ) ;
  assign n14171 = x127 &  n891 ;
  assign n14172 = n14170 | n14171 ;
  assign n14173 = n899 | n9960 ;
  assign n14174 = ( n14172 & ~n899 ) | ( n14172 & n14173 ) | ( ~n899 & n14173 ) ;
  assign n14175 = x17 | n14174 ;
  assign n14176 = ( x17 & ~n14174 ) | ( x17 & 1'b0 ) | ( ~n14174 & 1'b0 ) ;
  assign n14177 = ( n14175 & ~x17 ) | ( n14175 & n14176 ) | ( ~x17 & n14176 ) ;
  assign n14178 = ( n13954 & ~n14169 ) | ( n13954 & n14177 ) | ( ~n14169 & n14177 ) ;
  assign n14179 = ( n13954 & ~n14177 ) | ( n13954 & n14169 ) | ( ~n14177 & n14169 ) ;
  assign n14180 = ( n14178 & ~n13954 ) | ( n14178 & n14179 ) | ( ~n13954 & n14179 ) ;
  assign n14181 = ( n13714 & ~n13717 ) | ( n13714 & n13947 ) | ( ~n13717 & n13947 ) ;
  assign n14182 = ( n13951 & n14180 ) | ( n13951 & n14181 ) | ( n14180 & n14181 ) ;
  assign n14183 = ( n14180 & ~n13951 ) | ( n14180 & n14181 ) | ( ~n13951 & n14181 ) ;
  assign n14184 = ( n13951 & ~n14182 ) | ( n13951 & n14183 ) | ( ~n14182 & n14183 ) ;
  assign n14185 = ( n13954 & n14169 ) | ( n13954 & n14177 ) | ( n14169 & n14177 ) ;
  assign n14191 = ( x127 & ~n942 ) | ( x127 & 1'b0 ) | ( ~n942 & 1'b0 ) ;
  assign n14192 = n899 | n10258 ;
  assign n14193 = ~n14191 & n14192 ;
  assign n14187 = ( x20 & ~n13961 ) | ( x20 & 1'b0 ) | ( ~n13961 & 1'b0 ) ;
  assign n14188 = ~x20 & n13961 ;
  assign n14189 = n14187 | n14188 ;
  assign n14190 = ( n13962 & n14166 ) | ( n13962 & n14189 ) | ( n14166 & n14189 ) ;
  assign n14194 = ( x17 & ~n14193 ) | ( x17 & n14190 ) | ( ~n14193 & n14190 ) ;
  assign n14195 = ( n14190 & ~x17 ) | ( n14190 & n14193 ) | ( ~x17 & n14193 ) ;
  assign n14196 = ( n14194 & ~n14190 ) | ( n14194 & n14195 ) | ( ~n14190 & n14195 ) ;
  assign n14197 = ( n13968 & ~n14163 ) | ( n13968 & n14153 ) | ( ~n14163 & n14153 ) ;
  assign n14201 = x124 &  n1227 ;
  assign n14198 = ( x126 & ~n1154 ) | ( x126 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n14199 = x125 &  n1149 ;
  assign n14200 = n14198 | n14199 ;
  assign n14202 = ( x124 & ~n14201 ) | ( x124 & n14200 ) | ( ~n14201 & n14200 ) ;
  assign n14203 = n1157 | n9349 ;
  assign n14204 = ~n14202 & n14203 ;
  assign n14205 = x20 &  n14204 ;
  assign n14206 = x20 | n14204 ;
  assign n14207 = ~n14205 & n14206 ;
  assign n14211 = x121 &  n1551 ;
  assign n14208 = ( x123 & ~n1451 ) | ( x123 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n14209 = x122 &  n1446 ;
  assign n14210 = n14208 | n14209 ;
  assign n14212 = ( x121 & ~n14211 ) | ( x121 & n14210 ) | ( ~n14211 & n14210 ) ;
  assign n14213 = ~n1454 & n8472 ;
  assign n14214 = n14212 | n14213 ;
  assign n14215 = ( x23 & ~n14214 ) | ( x23 & 1'b0 ) | ( ~n14214 & 1'b0 ) ;
  assign n14216 = ~x23 & n14214 ;
  assign n14217 = n14215 | n14216 ;
  assign n14221 = x118 &  n1894 ;
  assign n14218 = ( x120 & ~n1816 ) | ( x120 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n14219 = x119 &  n1811 ;
  assign n14220 = n14218 | n14219 ;
  assign n14222 = ( x118 & ~n14221 ) | ( x118 & n14220 ) | ( ~n14221 & n14220 ) ;
  assign n14223 = ~n1819 & n9364 ;
  assign n14224 = n14222 | n14223 ;
  assign n14225 = ( n14143 & ~n13989 ) | ( n14143 & n14147 ) | ( ~n13989 & n14147 ) ;
  assign n14226 = ( x26 & n14224 ) | ( x26 & n14225 ) | ( n14224 & n14225 ) ;
  assign n14227 = ( x26 & ~n14224 ) | ( x26 & n14225 ) | ( ~n14224 & n14225 ) ;
  assign n14228 = ( n14224 & ~n14226 ) | ( n14224 & n14227 ) | ( ~n14226 & n14227 ) ;
  assign n14232 = x115 &  n2312 ;
  assign n14229 = ( x117 & ~n2195 ) | ( x117 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n14230 = x116 &  n2190 ;
  assign n14231 = n14229 | n14230 ;
  assign n14233 = ( x115 & ~n14232 ) | ( x115 & n14231 ) | ( ~n14232 & n14231 ) ;
  assign n14234 = n2198 | n7136 ;
  assign n14235 = ~n14233 & n14234 ;
  assign n14236 = x29 &  n14235 ;
  assign n14237 = x29 | n14235 ;
  assign n14238 = ~n14236 & n14237 ;
  assign n14242 = x112 &  n2718 ;
  assign n14239 = ( x114 & ~n2642 ) | ( x114 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n14240 = x113 &  n2637 ;
  assign n14241 = n14239 | n14240 ;
  assign n14243 = ( x112 & ~n14242 ) | ( x112 & n14241 ) | ( ~n14242 & n14241 ) ;
  assign n14244 = n2645 | n6185 ;
  assign n14245 = ~n14243 & n14244 ;
  assign n14246 = ( n14124 & ~n13997 ) | ( n14124 & n14134 ) | ( ~n13997 & n14134 ) ;
  assign n14247 = ( n14245 & ~x32 ) | ( n14245 & n14246 ) | ( ~x32 & n14246 ) ;
  assign n14248 = ( x32 & ~n14246 ) | ( x32 & n14245 ) | ( ~n14246 & n14245 ) ;
  assign n14249 = ( n14247 & ~n14245 ) | ( n14247 & n14248 ) | ( ~n14245 & n14248 ) ;
  assign n14253 = x106 &  n3756 ;
  assign n14250 = ( x108 & ~n3602 ) | ( x108 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n14251 = x107 &  n3597 ;
  assign n14252 = n14250 | n14251 ;
  assign n14254 = ( x106 & ~n14253 ) | ( x106 & n14252 ) | ( ~n14253 & n14252 ) ;
  assign n14255 = n3605 | n5055 ;
  assign n14256 = ~n14254 & n14255 ;
  assign n14257 = x38 &  n14256 ;
  assign n14258 = x38 | n14256 ;
  assign n14259 = ~n14257 & n14258 ;
  assign n14263 = x103 &  n4344 ;
  assign n14260 = ( x105 & ~n4143 ) | ( x105 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n14261 = x104 &  n4138 ;
  assign n14262 = n14260 | n14261 ;
  assign n14264 = ( x103 & ~n14263 ) | ( x103 & n14262 ) | ( ~n14263 & n14262 ) ;
  assign n14265 = ~n4146 & n4442 ;
  assign n14266 = n14264 | n14265 ;
  assign n14267 = ( x41 & ~n14266 ) | ( x41 & 1'b0 ) | ( ~n14266 & 1'b0 ) ;
  assign n14268 = ~x41 & n14266 ;
  assign n14269 = n14267 | n14268 ;
  assign n14270 = ( n13831 & ~n14112 ) | ( n13831 & n14102 ) | ( ~n14112 & n14102 ) ;
  assign n14271 = ( n14098 & ~n14088 ) | ( n14098 & n14099 ) | ( ~n14088 & n14099 ) ;
  assign n14272 = ( n14075 & ~n14074 ) | ( n14075 & n14085 ) | ( ~n14074 & n14085 ) ;
  assign n14273 = ( x59 & ~n14055 ) | ( x59 & 1'b0 ) | ( ~n14055 & 1'b0 ) ;
  assign n14274 = ~x59 & n14055 ;
  assign n14275 = n14273 | n14274 ;
  assign n14276 = ( n14031 & ~n14048 ) | ( n14031 & n14275 ) | ( ~n14048 & n14275 ) ;
  assign n14280 = x88 &  n7731 ;
  assign n14277 = ( x90 & ~n7538 ) | ( x90 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n14278 = x89 &  n7533 ;
  assign n14279 = n14277 | n14278 ;
  assign n14281 = ( x88 & ~n14280 ) | ( x88 & n14279 ) | ( ~n14280 & n14279 ) ;
  assign n14282 = ( n1976 & ~n7541 ) | ( n1976 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n14283 = n14281 | n14282 ;
  assign n14284 = ( x56 & ~n14283 ) | ( x56 & 1'b0 ) | ( ~n14283 & 1'b0 ) ;
  assign n14285 = ~x56 & n14283 ;
  assign n14286 = n14284 | n14285 ;
  assign n14290 = x82 &  n9457 ;
  assign n14287 = ( x84 & ~n9150 ) | ( x84 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n14288 = x83 &  n9145 ;
  assign n14289 = n14287 | n14288 ;
  assign n14291 = ( x82 & ~n14290 ) | ( x82 & n14289 ) | ( ~n14290 & n14289 ) ;
  assign n14292 = ( n1199 & ~n9153 ) | ( n1199 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n14293 = n14291 | n14292 ;
  assign n14294 = ( x62 & ~n14293 ) | ( x62 & 1'b0 ) | ( ~n14293 & 1'b0 ) ;
  assign n14295 = ~x62 & n14293 ;
  assign n14296 = n14294 | n14295 ;
  assign n14297 = x80 &  n10104 ;
  assign n14298 = ( x81 & ~n9760 ) | ( x81 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n14299 = n14297 | n14298 ;
  assign n14300 = ( n14035 & n14296 ) | ( n14035 & n14299 ) | ( n14296 & n14299 ) ;
  assign n14301 = ( n14035 & ~n14296 ) | ( n14035 & n14299 ) | ( ~n14296 & n14299 ) ;
  assign n14302 = ( n14296 & ~n14300 ) | ( n14296 & n14301 ) | ( ~n14300 & n14301 ) ;
  assign n14306 = x85 &  n8558 ;
  assign n14303 = ( x87 & ~n8314 ) | ( x87 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n14304 = x86 &  n8309 ;
  assign n14305 = n14303 | n14304 ;
  assign n14307 = ( x85 & ~n14306 ) | ( x85 & n14305 ) | ( ~n14306 & n14305 ) ;
  assign n14308 = ( n1512 & ~n8317 ) | ( n1512 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n14309 = n14307 | n14308 ;
  assign n14310 = ( x59 & ~n14309 ) | ( x59 & 1'b0 ) | ( ~n14309 & 1'b0 ) ;
  assign n14311 = ~x59 & n14309 ;
  assign n14312 = n14310 | n14311 ;
  assign n14313 = ( n14046 & n14302 ) | ( n14046 & n14312 ) | ( n14302 & n14312 ) ;
  assign n14314 = ( n14302 & ~n14046 ) | ( n14302 & n14312 ) | ( ~n14046 & n14312 ) ;
  assign n14315 = ( n14046 & ~n14313 ) | ( n14046 & n14314 ) | ( ~n14313 & n14314 ) ;
  assign n14316 = ( n14276 & ~n14286 ) | ( n14276 & n14315 ) | ( ~n14286 & n14315 ) ;
  assign n14317 = ( n14276 & ~n14315 ) | ( n14276 & n14286 ) | ( ~n14315 & n14286 ) ;
  assign n14318 = ( n14316 & ~n14276 ) | ( n14316 & n14317 ) | ( ~n14276 & n14317 ) ;
  assign n14319 = ( n13810 & ~n14061 ) | ( n13810 & n14071 ) | ( ~n14061 & n14071 ) ;
  assign n14323 = x91 &  n6982 ;
  assign n14320 = ( x93 & ~n6727 ) | ( x93 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n14321 = x92 &  n6722 ;
  assign n14322 = n14320 | n14321 ;
  assign n14324 = ( x91 & ~n14323 ) | ( x91 & n14322 ) | ( ~n14323 & n14322 ) ;
  assign n14325 = n2264 | n6730 ;
  assign n14326 = ~n14324 & n14325 ;
  assign n14327 = x53 &  n14326 ;
  assign n14328 = x53 | n14326 ;
  assign n14329 = ~n14327 & n14328 ;
  assign n14331 = ( n14318 & n14319 ) | ( n14318 & n14329 ) | ( n14319 & n14329 ) ;
  assign n14330 = ( n14319 & ~n14318 ) | ( n14319 & n14329 ) | ( ~n14318 & n14329 ) ;
  assign n14332 = ( n14318 & ~n14331 ) | ( n14318 & n14330 ) | ( ~n14331 & n14330 ) ;
  assign n14336 = x94 &  n6288 ;
  assign n14333 = ( x96 & ~n6032 ) | ( x96 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n14334 = x95 &  n6027 ;
  assign n14335 = n14333 | n14334 ;
  assign n14337 = ( x94 & ~n14336 ) | ( x94 & n14335 ) | ( ~n14336 & n14335 ) ;
  assign n14338 = ( n2836 & ~n6035 ) | ( n2836 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n14339 = n14337 | n14338 ;
  assign n14340 = ( x50 & ~n14339 ) | ( x50 & 1'b0 ) | ( ~n14339 & 1'b0 ) ;
  assign n14341 = ~x50 & n14339 ;
  assign n14342 = n14340 | n14341 ;
  assign n14343 = ( n14272 & ~n14332 ) | ( n14272 & n14342 ) | ( ~n14332 & n14342 ) ;
  assign n14344 = ( n14272 & ~n14342 ) | ( n14272 & n14332 ) | ( ~n14342 & n14332 ) ;
  assign n14345 = ( n14343 & ~n14272 ) | ( n14343 & n14344 ) | ( ~n14272 & n14344 ) ;
  assign n14349 = x97 &  n5586 ;
  assign n14346 = ( x99 & ~n5389 ) | ( x99 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n14347 = x98 &  n5384 ;
  assign n14348 = n14346 | n14347 ;
  assign n14350 = ( x97 & ~n14349 ) | ( x97 & n14348 ) | ( ~n14349 & n14348 ) ;
  assign n14351 = ( n3338 & ~n5392 ) | ( n3338 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n14352 = n14350 | n14351 ;
  assign n14353 = ( x47 & ~n14352 ) | ( x47 & 1'b0 ) | ( ~n14352 & 1'b0 ) ;
  assign n14354 = ~x47 & n14352 ;
  assign n14355 = n14353 | n14354 ;
  assign n14356 = ( n14271 & ~n14345 ) | ( n14271 & n14355 ) | ( ~n14345 & n14355 ) ;
  assign n14357 = ( n14271 & ~n14355 ) | ( n14271 & n14345 ) | ( ~n14355 & n14345 ) ;
  assign n14358 = ( n14356 & ~n14271 ) | ( n14356 & n14357 ) | ( ~n14271 & n14357 ) ;
  assign n14362 = x100 &  n4934 ;
  assign n14359 = ( x102 & ~n4725 ) | ( x102 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n14360 = x101 &  n4720 ;
  assign n14361 = n14359 | n14360 ;
  assign n14363 = ( x100 & ~n14362 ) | ( x100 & n14361 ) | ( ~n14362 & n14361 ) ;
  assign n14364 = n3872 | n4728 ;
  assign n14365 = ~n14363 & n14364 ;
  assign n14366 = x44 &  n14365 ;
  assign n14367 = x44 | n14365 ;
  assign n14368 = ~n14366 & n14367 ;
  assign n14369 = ( n14270 & n14358 ) | ( n14270 & n14368 ) | ( n14358 & n14368 ) ;
  assign n14370 = ( n14358 & ~n14270 ) | ( n14358 & n14368 ) | ( ~n14270 & n14368 ) ;
  assign n14371 = ( n14270 & ~n14369 ) | ( n14270 & n14370 ) | ( ~n14369 & n14370 ) ;
  assign n14372 = ( n14117 & ~n14269 ) | ( n14117 & n14371 ) | ( ~n14269 & n14371 ) ;
  assign n14373 = ( n14117 & ~n14371 ) | ( n14117 & n14269 ) | ( ~n14371 & n14269 ) ;
  assign n14374 = ( n14372 & ~n14117 ) | ( n14372 & n14373 ) | ( ~n14117 & n14373 ) ;
  assign n14375 = ( n14120 & ~n14259 ) | ( n14120 & n14374 ) | ( ~n14259 & n14374 ) ;
  assign n14376 = ( n14120 & ~n14374 ) | ( n14120 & n14259 ) | ( ~n14374 & n14259 ) ;
  assign n14377 = ( n14375 & ~n14120 ) | ( n14375 & n14376 ) | ( ~n14120 & n14376 ) ;
  assign n14381 = x109 &  n3214 ;
  assign n14378 = ( x111 & ~n3087 ) | ( x111 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n14379 = x110 &  n3082 ;
  assign n14380 = n14378 | n14379 ;
  assign n14382 = ( x109 & ~n14381 ) | ( x109 & n14380 ) | ( ~n14381 & n14380 ) ;
  assign n14383 = n3090 | n5711 ;
  assign n14384 = ~n14382 & n14383 ;
  assign n14385 = x35 &  n14384 ;
  assign n14386 = x35 | n14384 ;
  assign n14387 = ~n14385 & n14386 ;
  assign n14388 = ( n14123 & n14377 ) | ( n14123 & n14387 ) | ( n14377 & n14387 ) ;
  assign n14389 = ( n14123 & ~n14377 ) | ( n14123 & n14387 ) | ( ~n14377 & n14387 ) ;
  assign n14390 = ( n14377 & ~n14388 ) | ( n14377 & n14389 ) | ( ~n14388 & n14389 ) ;
  assign n14391 = ( n14249 & ~n14390 ) | ( n14249 & 1'b0 ) | ( ~n14390 & 1'b0 ) ;
  assign n14392 = ~n14249 & n14390 ;
  assign n14393 = n14391 | n14392 ;
  assign n14394 = ~x32 & n13996 ;
  assign n14395 = ( x32 & ~n13996 ) | ( x32 & 1'b0 ) | ( ~n13996 & 1'b0 ) ;
  assign n14396 = n14394 | n14395 ;
  assign n14397 = ( n13889 & ~n14137 ) | ( n13889 & n14396 ) | ( ~n14137 & n14396 ) ;
  assign n14398 = ( n14238 & ~n14393 ) | ( n14238 & n14397 ) | ( ~n14393 & n14397 ) ;
  assign n14399 = ( n14238 & ~n14397 ) | ( n14238 & n14393 ) | ( ~n14397 & n14393 ) ;
  assign n14400 = ( n14398 & ~n14238 ) | ( n14398 & n14399 ) | ( ~n14238 & n14399 ) ;
  assign n14401 = ( n14228 & ~n14400 ) | ( n14228 & 1'b0 ) | ( ~n14400 & 1'b0 ) ;
  assign n14402 = ~n14228 & n14400 ;
  assign n14403 = n14401 | n14402 ;
  assign n14404 = x26 &  n13975 ;
  assign n14405 = ( n13977 & ~n14404 ) | ( n13977 & n14151 ) | ( ~n14404 & n14151 ) ;
  assign n14406 = ( n14217 & n14403 ) | ( n14217 & n14405 ) | ( n14403 & n14405 ) ;
  assign n14407 = ( n14403 & ~n14217 ) | ( n14403 & n14405 ) | ( ~n14217 & n14405 ) ;
  assign n14408 = ( n14217 & ~n14406 ) | ( n14217 & n14407 ) | ( ~n14406 & n14407 ) ;
  assign n14409 = ( n14197 & ~n14207 ) | ( n14197 & n14408 ) | ( ~n14207 & n14408 ) ;
  assign n14410 = ( n14197 & ~n14408 ) | ( n14197 & n14207 ) | ( ~n14408 & n14207 ) ;
  assign n14411 = ( n14409 & ~n14197 ) | ( n14409 & n14410 ) | ( ~n14197 & n14410 ) ;
  assign n14412 = n14196 | n14411 ;
  assign n14413 = n14196 &  n14411 ;
  assign n14414 = ( n14412 & ~n14413 ) | ( n14412 & 1'b0 ) | ( ~n14413 & 1'b0 ) ;
  assign n14186 = ( n13951 & ~n14180 ) | ( n13951 & n14181 ) | ( ~n14180 & n14181 ) ;
  assign n14415 = ( n14185 & ~n14414 ) | ( n14185 & n14186 ) | ( ~n14414 & n14186 ) ;
  assign n14416 = ( n14185 & ~n14186 ) | ( n14185 & n14414 ) | ( ~n14186 & n14414 ) ;
  assign n14417 = ( n14415 & ~n14185 ) | ( n14415 & n14416 ) | ( ~n14185 & n14416 ) ;
  assign n14418 = ~x17 & n14193 ;
  assign n14419 = ( n14412 & ~n14195 ) | ( n14412 & n14418 ) | ( ~n14195 & n14418 ) ;
  assign n14423 = x125 &  n1227 ;
  assign n14420 = ( x127 & ~n1154 ) | ( x127 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n14421 = x126 &  n1149 ;
  assign n14422 = n14420 | n14421 ;
  assign n14424 = ( x125 & ~n14423 ) | ( x125 & n14422 ) | ( ~n14423 & n14422 ) ;
  assign n14425 = n1157 | n9941 ;
  assign n14426 = ~n14424 & n14425 ;
  assign n14427 = x20 &  n14426 ;
  assign n14428 = x20 | n14426 ;
  assign n14429 = ~n14427 & n14428 ;
  assign n14430 = ( n14197 & n14207 ) | ( n14197 & n14408 ) | ( n14207 & n14408 ) ;
  assign n14431 = ( n14217 & ~n14403 ) | ( n14217 & n14405 ) | ( ~n14403 & n14405 ) ;
  assign n14435 = x122 &  n1551 ;
  assign n14432 = ( x124 & ~n1451 ) | ( x124 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n14433 = x123 &  n1446 ;
  assign n14434 = n14432 | n14433 ;
  assign n14436 = ( x122 & ~n14435 ) | ( x122 & n14434 ) | ( ~n14435 & n14434 ) ;
  assign n14437 = ~n1454 & n8755 ;
  assign n14438 = n14436 | n14437 ;
  assign n14440 = x23 &  n14438 ;
  assign n14439 = ~x23 & n14438 ;
  assign n14441 = ( x23 & ~n14440 ) | ( x23 & n14439 ) | ( ~n14440 & n14439 ) ;
  assign n14445 = x119 &  n1894 ;
  assign n14442 = ( x121 & ~n1816 ) | ( x121 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n14443 = x120 &  n1811 ;
  assign n14444 = n14442 | n14443 ;
  assign n14446 = ( x119 & ~n14445 ) | ( x119 & n14444 ) | ( ~n14445 & n14444 ) ;
  assign n14447 = ~n1819 & n8176 ;
  assign n14448 = n14446 | n14447 ;
  assign n14449 = ( x26 & ~n14448 ) | ( x26 & 1'b0 ) | ( ~n14448 & 1'b0 ) ;
  assign n14450 = ~x26 & n14448 ;
  assign n14451 = n14449 | n14450 ;
  assign n14452 = ( n14238 & n14393 ) | ( n14238 & n14397 ) | ( n14393 & n14397 ) ;
  assign n14456 = x116 &  n2312 ;
  assign n14453 = ( x118 & ~n2195 ) | ( x118 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n14454 = x117 &  n2190 ;
  assign n14455 = n14453 | n14454 ;
  assign n14457 = ( x116 & ~n14456 ) | ( x116 & n14455 ) | ( ~n14456 & n14455 ) ;
  assign n14458 = n2198 | n7152 ;
  assign n14459 = ~n14457 & n14458 ;
  assign n14460 = x29 &  n14459 ;
  assign n14461 = x29 | n14459 ;
  assign n14462 = ~n14460 & n14461 ;
  assign n14466 = x113 &  n2718 ;
  assign n14463 = ( x115 & ~n2642 ) | ( x115 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n14464 = x114 &  n2637 ;
  assign n14465 = n14463 | n14464 ;
  assign n14467 = ( x113 & ~n14466 ) | ( x113 & n14465 ) | ( ~n14466 & n14465 ) ;
  assign n14468 = ~n2645 & n6420 ;
  assign n14469 = n14467 | n14468 ;
  assign n14470 = ( x32 & ~n14469 ) | ( x32 & 1'b0 ) | ( ~n14469 & 1'b0 ) ;
  assign n14471 = ~x32 & n14469 ;
  assign n14472 = n14470 | n14471 ;
  assign n14617 = ( x32 & ~n14245 ) | ( x32 & 1'b0 ) | ( ~n14245 & 1'b0 ) ;
  assign n14618 = ( n14247 & ~n14391 ) | ( n14247 & n14617 ) | ( ~n14391 & n14617 ) ;
  assign n14476 = x110 &  n3214 ;
  assign n14473 = ( x112 & ~n3087 ) | ( x112 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n14474 = x111 &  n3082 ;
  assign n14475 = n14473 | n14474 ;
  assign n14477 = ( x110 & ~n14476 ) | ( x110 & n14475 ) | ( ~n14476 & n14475 ) ;
  assign n14478 = ~n3090 & n5727 ;
  assign n14479 = n14477 | n14478 ;
  assign n14480 = ( x35 & ~n14479 ) | ( x35 & 1'b0 ) | ( ~n14479 & 1'b0 ) ;
  assign n14481 = ~x35 & n14479 ;
  assign n14482 = n14480 | n14481 ;
  assign n14486 = x107 &  n3756 ;
  assign n14483 = ( x109 & ~n3602 ) | ( x109 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n14484 = x108 &  n3597 ;
  assign n14485 = n14483 | n14484 ;
  assign n14487 = ( x107 & ~n14486 ) | ( x107 & n14485 ) | ( ~n14486 & n14485 ) ;
  assign n14488 = ~n3605 & n5267 ;
  assign n14489 = n14487 | n14488 ;
  assign n14490 = ( x38 & ~n14489 ) | ( x38 & 1'b0 ) | ( ~n14489 & 1'b0 ) ;
  assign n14491 = ~x38 & n14489 ;
  assign n14492 = n14490 | n14491 ;
  assign n14496 = x95 &  n6288 ;
  assign n14493 = ( x97 & ~n6032 ) | ( x97 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n14494 = x96 &  n6027 ;
  assign n14495 = n14493 | n14494 ;
  assign n14497 = ( x95 & ~n14496 ) | ( x95 & n14495 ) | ( ~n14496 & n14495 ) ;
  assign n14498 = ( n2999 & ~n6035 ) | ( n2999 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n14499 = n14497 | n14498 ;
  assign n14500 = ( x50 & ~n14499 ) | ( x50 & 1'b0 ) | ( ~n14499 & 1'b0 ) ;
  assign n14501 = ~x50 & n14499 ;
  assign n14502 = n14500 | n14501 ;
  assign n14506 = x92 &  n6982 ;
  assign n14503 = ( x94 & ~n6727 ) | ( x94 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n14504 = x93 &  n6722 ;
  assign n14505 = n14503 | n14504 ;
  assign n14507 = ( x92 & ~n14506 ) | ( x92 & n14505 ) | ( ~n14506 & n14505 ) ;
  assign n14508 = ( n2401 & ~n6730 ) | ( n2401 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n14509 = n14507 | n14508 ;
  assign n14510 = ( x53 & ~n14509 ) | ( x53 & 1'b0 ) | ( ~n14509 & 1'b0 ) ;
  assign n14511 = ~x53 & n14509 ;
  assign n14512 = n14510 | n14511 ;
  assign n14550 = x89 &  n7731 ;
  assign n14547 = ( x91 & ~n7538 ) | ( x91 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n14548 = x90 &  n7533 ;
  assign n14549 = n14547 | n14548 ;
  assign n14551 = ( x89 & ~n14550 ) | ( x89 & n14549 ) | ( ~n14550 & n14549 ) ;
  assign n14552 = ( n2108 & ~n7541 ) | ( n2108 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n14553 = n14551 | n14552 ;
  assign n14554 = ( x56 & ~n14553 ) | ( x56 & 1'b0 ) | ( ~n14553 & 1'b0 ) ;
  assign n14555 = ~x56 & n14553 ;
  assign n14556 = n14554 | n14555 ;
  assign n14516 = x83 &  n9457 ;
  assign n14513 = ( x85 & ~n9150 ) | ( x85 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n14514 = x84 &  n9145 ;
  assign n14515 = n14513 | n14514 ;
  assign n14517 = ( x83 & ~n14516 ) | ( x83 & n14515 ) | ( ~n14516 & n14515 ) ;
  assign n14518 = ( n1295 & ~n9153 ) | ( n1295 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n14519 = n14517 | n14518 ;
  assign n14521 = x62 &  n14519 ;
  assign n14520 = ~x62 & n14519 ;
  assign n14522 = ( x62 & ~n14521 ) | ( x62 & n14520 ) | ( ~n14521 & n14520 ) ;
  assign n14523 = ( n14035 & ~n14299 ) | ( n14035 & n14296 ) | ( ~n14299 & n14296 ) ;
  assign n14524 = x81 &  n10104 ;
  assign n14525 = ( x82 & ~n9760 ) | ( x82 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n14526 = n14524 | n14525 ;
  assign n14527 = ( x17 & n14299 ) | ( x17 & n14526 ) | ( n14299 & n14526 ) ;
  assign n14528 = ( x17 & ~n14299 ) | ( x17 & n14526 ) | ( ~n14299 & n14526 ) ;
  assign n14529 = ( n14299 & ~n14527 ) | ( n14299 & n14528 ) | ( ~n14527 & n14528 ) ;
  assign n14530 = ( n14522 & ~n14523 ) | ( n14522 & n14529 ) | ( ~n14523 & n14529 ) ;
  assign n14531 = ( n14522 & ~n14529 ) | ( n14522 & n14523 ) | ( ~n14529 & n14523 ) ;
  assign n14532 = ( n14530 & ~n14522 ) | ( n14530 & n14531 ) | ( ~n14522 & n14531 ) ;
  assign n14537 = x86 &  n8558 ;
  assign n14534 = ( x88 & ~n8314 ) | ( x88 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n14535 = x87 &  n8309 ;
  assign n14536 = n14534 | n14535 ;
  assign n14538 = ( x86 & ~n14537 ) | ( x86 & n14536 ) | ( ~n14537 & n14536 ) ;
  assign n14539 = ( n1624 & ~n8317 ) | ( n1624 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n14540 = n14538 | n14539 ;
  assign n14541 = ( x59 & ~n14540 ) | ( x59 & 1'b0 ) | ( ~n14540 & 1'b0 ) ;
  assign n14542 = ~x59 & n14540 ;
  assign n14543 = n14541 | n14542 ;
  assign n14533 = ( n14046 & ~n14302 ) | ( n14046 & n14312 ) | ( ~n14302 & n14312 ) ;
  assign n14544 = ( n14532 & ~n14543 ) | ( n14532 & n14533 ) | ( ~n14543 & n14533 ) ;
  assign n14545 = ( n14532 & ~n14533 ) | ( n14532 & n14543 ) | ( ~n14533 & n14543 ) ;
  assign n14546 = ( n14544 & ~n14532 ) | ( n14544 & n14545 ) | ( ~n14532 & n14545 ) ;
  assign n14557 = ( n14317 & ~n14556 ) | ( n14317 & n14546 ) | ( ~n14556 & n14546 ) ;
  assign n14558 = ( n14546 & ~n14317 ) | ( n14546 & n14556 ) | ( ~n14317 & n14556 ) ;
  assign n14559 = ( n14557 & ~n14546 ) | ( n14557 & n14558 ) | ( ~n14546 & n14558 ) ;
  assign n14560 = ( n14318 & ~n14319 ) | ( n14318 & n14329 ) | ( ~n14319 & n14329 ) ;
  assign n14562 = ( n14512 & n14559 ) | ( n14512 & n14560 ) | ( n14559 & n14560 ) ;
  assign n14561 = ( n14559 & ~n14512 ) | ( n14559 & n14560 ) | ( ~n14512 & n14560 ) ;
  assign n14563 = ( n14512 & ~n14562 ) | ( n14512 & n14561 ) | ( ~n14562 & n14561 ) ;
  assign n14564 = ( n14272 & n14332 ) | ( n14272 & n14342 ) | ( n14332 & n14342 ) ;
  assign n14565 = ( n14502 & n14563 ) | ( n14502 & n14564 ) | ( n14563 & n14564 ) ;
  assign n14566 = ( n14563 & ~n14502 ) | ( n14563 & n14564 ) | ( ~n14502 & n14564 ) ;
  assign n14567 = ( n14502 & ~n14565 ) | ( n14502 & n14566 ) | ( ~n14565 & n14566 ) ;
  assign n14568 = ( n14271 & n14345 ) | ( n14271 & n14355 ) | ( n14345 & n14355 ) ;
  assign n14572 = x98 &  n5586 ;
  assign n14569 = ( x100 & ~n5389 ) | ( x100 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n14570 = x99 &  n5384 ;
  assign n14571 = n14569 | n14570 ;
  assign n14573 = ( x98 & ~n14572 ) | ( x98 & n14571 ) | ( ~n14572 & n14571 ) ;
  assign n14574 = n3354 | n5392 ;
  assign n14575 = ~n14573 & n14574 ;
  assign n14576 = x47 &  n14575 ;
  assign n14577 = x47 | n14575 ;
  assign n14578 = ~n14576 & n14577 ;
  assign n14580 = ( n14567 & n14568 ) | ( n14567 & n14578 ) | ( n14568 & n14578 ) ;
  assign n14579 = ( n14568 & ~n14567 ) | ( n14568 & n14578 ) | ( ~n14567 & n14578 ) ;
  assign n14581 = ( n14567 & ~n14580 ) | ( n14567 & n14579 ) | ( ~n14580 & n14579 ) ;
  assign n14586 = x101 &  n4934 ;
  assign n14583 = ( x103 & ~n4725 ) | ( x103 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n14584 = x102 &  n4720 ;
  assign n14585 = n14583 | n14584 ;
  assign n14587 = ( x101 & ~n14586 ) | ( x101 & n14585 ) | ( ~n14586 & n14585 ) ;
  assign n14588 = n4056 | n4728 ;
  assign n14589 = ~n14587 & n14588 ;
  assign n14590 = x44 &  n14589 ;
  assign n14591 = x44 | n14589 ;
  assign n14592 = ~n14590 & n14591 ;
  assign n14582 = ( n14270 & ~n14358 ) | ( n14270 & n14368 ) | ( ~n14358 & n14368 ) ;
  assign n14593 = ( n14581 & ~n14592 ) | ( n14581 & n14582 ) | ( ~n14592 & n14582 ) ;
  assign n14594 = ( n14581 & ~n14582 ) | ( n14581 & n14592 ) | ( ~n14582 & n14592 ) ;
  assign n14595 = ( n14593 & ~n14581 ) | ( n14593 & n14594 ) | ( ~n14581 & n14594 ) ;
  assign n14600 = x104 &  n4344 ;
  assign n14597 = ( x106 & ~n4143 ) | ( x106 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n14598 = x105 &  n4138 ;
  assign n14599 = n14597 | n14598 ;
  assign n14601 = ( x104 & ~n14600 ) | ( x104 & n14599 ) | ( ~n14600 & n14599 ) ;
  assign n14602 = ~n4146 & n4458 ;
  assign n14603 = n14601 | n14602 ;
  assign n14604 = ( x41 & ~n14603 ) | ( x41 & 1'b0 ) | ( ~n14603 & 1'b0 ) ;
  assign n14605 = ~x41 & n14603 ;
  assign n14606 = n14604 | n14605 ;
  assign n14596 = ( n14117 & n14269 ) | ( n14117 & n14371 ) | ( n14269 & n14371 ) ;
  assign n14607 = ( n14595 & ~n14606 ) | ( n14595 & n14596 ) | ( ~n14606 & n14596 ) ;
  assign n14608 = ( n14595 & ~n14596 ) | ( n14595 & n14606 ) | ( ~n14596 & n14606 ) ;
  assign n14609 = ( n14607 & ~n14595 ) | ( n14607 & n14608 ) | ( ~n14595 & n14608 ) ;
  assign n14611 = ( n14376 & n14492 ) | ( n14376 & n14609 ) | ( n14492 & n14609 ) ;
  assign n14610 = ( n14376 & ~n14492 ) | ( n14376 & n14609 ) | ( ~n14492 & n14609 ) ;
  assign n14612 = ( n14492 & ~n14611 ) | ( n14492 & n14610 ) | ( ~n14611 & n14610 ) ;
  assign n14613 = ( n14123 & ~n14387 ) | ( n14123 & n14377 ) | ( ~n14387 & n14377 ) ;
  assign n14614 = ( n14482 & n14612 ) | ( n14482 & n14613 ) | ( n14612 & n14613 ) ;
  assign n14615 = ( n14612 & ~n14482 ) | ( n14612 & n14613 ) | ( ~n14482 & n14613 ) ;
  assign n14616 = ( n14482 & ~n14614 ) | ( n14482 & n14615 ) | ( ~n14614 & n14615 ) ;
  assign n14619 = ( n14472 & ~n14618 ) | ( n14472 & n14616 ) | ( ~n14618 & n14616 ) ;
  assign n14620 = ( n14472 & ~n14616 ) | ( n14472 & n14618 ) | ( ~n14616 & n14618 ) ;
  assign n14621 = ( n14619 & ~n14472 ) | ( n14619 & n14620 ) | ( ~n14472 & n14620 ) ;
  assign n14622 = ( n14452 & ~n14462 ) | ( n14452 & n14621 ) | ( ~n14462 & n14621 ) ;
  assign n14623 = ( n14452 & ~n14621 ) | ( n14452 & n14462 ) | ( ~n14621 & n14462 ) ;
  assign n14624 = ( n14622 & ~n14452 ) | ( n14622 & n14623 ) | ( ~n14452 & n14623 ) ;
  assign n14625 = x26 &  n14224 ;
  assign n14626 = ( n14226 & ~n14625 ) | ( n14226 & n14401 ) | ( ~n14625 & n14401 ) ;
  assign n14627 = ( n14451 & n14624 ) | ( n14451 & n14626 ) | ( n14624 & n14626 ) ;
  assign n14628 = ( n14624 & ~n14451 ) | ( n14624 & n14626 ) | ( ~n14451 & n14626 ) ;
  assign n14629 = ( n14451 & ~n14627 ) | ( n14451 & n14628 ) | ( ~n14627 & n14628 ) ;
  assign n14631 = ( n14431 & n14441 ) | ( n14431 & n14629 ) | ( n14441 & n14629 ) ;
  assign n14630 = ( n14441 & ~n14431 ) | ( n14441 & n14629 ) | ( ~n14431 & n14629 ) ;
  assign n14632 = ( n14431 & ~n14631 ) | ( n14431 & n14630 ) | ( ~n14631 & n14630 ) ;
  assign n14633 = ( n14429 & ~n14430 ) | ( n14429 & n14632 ) | ( ~n14430 & n14632 ) ;
  assign n14634 = ( n14429 & ~n14632 ) | ( n14429 & n14430 ) | ( ~n14632 & n14430 ) ;
  assign n14635 = ( n14633 & ~n14429 ) | ( n14633 & n14634 ) | ( ~n14429 & n14634 ) ;
  assign n14636 = ( n14416 & n14419 ) | ( n14416 & n14635 ) | ( n14419 & n14635 ) ;
  assign n14637 = ( n14416 & ~n14419 ) | ( n14416 & n14635 ) | ( ~n14419 & n14635 ) ;
  assign n14638 = ( n14419 & ~n14636 ) | ( n14419 & n14637 ) | ( ~n14636 & n14637 ) ;
  assign n14639 = ( n14429 & n14430 ) | ( n14429 & n14632 ) | ( n14430 & n14632 ) ;
  assign n14640 = ( n14419 & ~n14416 ) | ( n14419 & n14635 ) | ( ~n14416 & n14635 ) ;
  assign n14641 = ( n14431 & ~n14629 ) | ( n14431 & n14441 ) | ( ~n14629 & n14441 ) ;
  assign n14645 = x123 &  n1551 ;
  assign n14642 = ( x125 & ~n1451 ) | ( x125 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n14643 = x124 &  n1446 ;
  assign n14644 = n14642 | n14643 ;
  assign n14646 = ( x123 & ~n14645 ) | ( x123 & n14644 ) | ( ~n14645 & n14644 ) ;
  assign n14647 = ~n1454 & n9324 ;
  assign n14648 = n14646 | n14647 ;
  assign n14649 = ( x23 & ~n14648 ) | ( x23 & 1'b0 ) | ( ~n14648 & 1'b0 ) ;
  assign n14650 = ~x23 & n14648 ;
  assign n14651 = n14649 | n14650 ;
  assign n14659 = ( n14452 & n14462 ) | ( n14452 & n14621 ) | ( n14462 & n14621 ) ;
  assign n14655 = x120 &  n1894 ;
  assign n14652 = ( x122 & ~n1816 ) | ( x122 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n14653 = x121 &  n1811 ;
  assign n14654 = n14652 | n14653 ;
  assign n14656 = ( x120 & ~n14655 ) | ( x120 & n14654 ) | ( ~n14655 & n14654 ) ;
  assign n14657 = ~n1819 & n9987 ;
  assign n14658 = n14656 | n14657 ;
  assign n14660 = ( x26 & ~n14659 ) | ( x26 & n14658 ) | ( ~n14659 & n14658 ) ;
  assign n14661 = ( n14658 & ~x26 ) | ( n14658 & n14659 ) | ( ~x26 & n14659 ) ;
  assign n14662 = ( n14660 & ~n14658 ) | ( n14660 & n14661 ) | ( ~n14658 & n14661 ) ;
  assign n14666 = x117 &  n2312 ;
  assign n14663 = ( x119 & ~n2195 ) | ( x119 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n14664 = x118 &  n2190 ;
  assign n14665 = n14663 | n14664 ;
  assign n14667 = ( x117 & ~n14666 ) | ( x117 & n14665 ) | ( ~n14666 & n14665 ) ;
  assign n14668 = ~n2198 & n7648 ;
  assign n14669 = n14667 | n14668 ;
  assign n14670 = ( x29 & ~n14669 ) | ( x29 & 1'b0 ) | ( ~n14669 & 1'b0 ) ;
  assign n14671 = ~x29 & n14669 ;
  assign n14672 = n14670 | n14671 ;
  assign n14819 = ~x32 & n14614 ;
  assign n14820 = x32 | n14614 ;
  assign n14821 = ( n14819 & ~n14614 ) | ( n14819 & n14820 ) | ( ~n14614 & n14820 ) ;
  assign n14676 = x114 &  n2718 ;
  assign n14673 = ( x116 & ~n2642 ) | ( x116 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n14674 = x115 &  n2637 ;
  assign n14675 = n14673 | n14674 ;
  assign n14677 = ( x114 & ~n14676 ) | ( x114 & n14675 ) | ( ~n14676 & n14675 ) ;
  assign n14678 = n2645 | n6885 ;
  assign n14679 = ~n14677 & n14678 ;
  assign n14680 = ( n14596 & ~n14595 ) | ( n14596 & n14606 ) | ( ~n14595 & n14606 ) ;
  assign n14796 = x108 &  n3756 ;
  assign n14793 = ( x110 & ~n3602 ) | ( x110 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n14794 = x109 &  n3597 ;
  assign n14795 = n14793 | n14794 ;
  assign n14797 = ( x108 & ~n14796 ) | ( x108 & n14795 ) | ( ~n14796 & n14795 ) ;
  assign n14798 = n3605 | n5283 ;
  assign n14799 = ~n14797 & n14798 ;
  assign n14800 = x38 &  n14799 ;
  assign n14801 = x38 | n14799 ;
  assign n14802 = ~n14800 & n14801 ;
  assign n14681 = ( n14581 & n14582 ) | ( n14581 & n14592 ) | ( n14582 & n14592 ) ;
  assign n14685 = x105 &  n4344 ;
  assign n14682 = ( x107 & ~n4143 ) | ( x107 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n14683 = x106 &  n4138 ;
  assign n14684 = n14682 | n14683 ;
  assign n14686 = ( x105 & ~n14685 ) | ( x105 & n14684 ) | ( ~n14685 & n14684 ) ;
  assign n14687 = ~n4146 & n4848 ;
  assign n14688 = n14686 | n14687 ;
  assign n14689 = ( x41 & ~n14688 ) | ( x41 & 1'b0 ) | ( ~n14688 & 1'b0 ) ;
  assign n14690 = ~x41 & n14688 ;
  assign n14691 = n14689 | n14690 ;
  assign n14692 = ( n14567 & ~n14578 ) | ( n14567 & n14568 ) | ( ~n14578 & n14568 ) ;
  assign n14696 = x102 &  n4934 ;
  assign n14693 = ( x104 & ~n4725 ) | ( x104 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n14694 = x103 &  n4720 ;
  assign n14695 = n14693 | n14694 ;
  assign n14697 = ( x102 & ~n14696 ) | ( x102 & n14695 ) | ( ~n14696 & n14695 ) ;
  assign n14698 = n4249 | n4728 ;
  assign n14699 = ~n14697 & n14698 ;
  assign n14700 = x44 &  n14699 ;
  assign n14701 = x44 | n14699 ;
  assign n14702 = ~n14700 & n14701 ;
  assign n14723 = x87 &  n8558 ;
  assign n14720 = ( x89 & ~n8314 ) | ( x89 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n14721 = x88 &  n8309 ;
  assign n14722 = n14720 | n14721 ;
  assign n14724 = ( x87 & ~n14723 ) | ( x87 & n14722 ) | ( ~n14723 & n14722 ) ;
  assign n14725 = ( n1741 & ~n8317 ) | ( n1741 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n14726 = n14724 | n14725 ;
  assign n14727 = ( x59 & ~n14726 ) | ( x59 & 1'b0 ) | ( ~n14726 & 1'b0 ) ;
  assign n14728 = ~x59 & n14726 ;
  assign n14729 = n14727 | n14728 ;
  assign n14703 = ( n14299 & ~x17 ) | ( n14299 & n14526 ) | ( ~x17 & n14526 ) ;
  assign n14707 = x84 &  n9457 ;
  assign n14704 = ( x86 & ~n9150 ) | ( x86 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n14705 = x85 &  n9145 ;
  assign n14706 = n14704 | n14705 ;
  assign n14708 = ( x84 & ~n14707 ) | ( x84 & n14706 ) | ( ~n14707 & n14706 ) ;
  assign n14709 = ( n1496 & ~n9153 ) | ( n1496 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n14710 = n14708 | n14709 ;
  assign n14711 = ( x62 & ~n14710 ) | ( x62 & 1'b0 ) | ( ~n14710 & 1'b0 ) ;
  assign n14712 = ~x62 & n14710 ;
  assign n14713 = n14711 | n14712 ;
  assign n14714 = x82 &  n10104 ;
  assign n14715 = ( x83 & ~n9760 ) | ( x83 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n14716 = n14714 | n14715 ;
  assign n14718 = ( n14703 & n14713 ) | ( n14703 & n14716 ) | ( n14713 & n14716 ) ;
  assign n14717 = ( n14713 & ~n14703 ) | ( n14713 & n14716 ) | ( ~n14703 & n14716 ) ;
  assign n14719 = ( n14703 & ~n14718 ) | ( n14703 & n14717 ) | ( ~n14718 & n14717 ) ;
  assign n14730 = ( n14531 & ~n14729 ) | ( n14531 & n14719 ) | ( ~n14729 & n14719 ) ;
  assign n14731 = ( n14719 & ~n14531 ) | ( n14719 & n14729 ) | ( ~n14531 & n14729 ) ;
  assign n14732 = ( n14730 & ~n14719 ) | ( n14730 & n14731 ) | ( ~n14719 & n14731 ) ;
  assign n14737 = x90 &  n7731 ;
  assign n14734 = ( x92 & ~n7538 ) | ( x92 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n14735 = x91 &  n7533 ;
  assign n14736 = n14734 | n14735 ;
  assign n14738 = ( x90 & ~n14737 ) | ( x90 & n14736 ) | ( ~n14737 & n14736 ) ;
  assign n14739 = ( n2248 & ~n7541 ) | ( n2248 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n14740 = n14738 | n14739 ;
  assign n14741 = ( x56 & ~n14740 ) | ( x56 & 1'b0 ) | ( ~n14740 & 1'b0 ) ;
  assign n14742 = ~x56 & n14740 ;
  assign n14743 = n14741 | n14742 ;
  assign n14733 = ( n14533 & ~n14532 ) | ( n14533 & n14543 ) | ( ~n14532 & n14543 ) ;
  assign n14744 = ( n14732 & ~n14743 ) | ( n14732 & n14733 ) | ( ~n14743 & n14733 ) ;
  assign n14745 = ( n14732 & ~n14733 ) | ( n14732 & n14743 ) | ( ~n14733 & n14743 ) ;
  assign n14746 = ( n14744 & ~n14732 ) | ( n14744 & n14745 ) | ( ~n14732 & n14745 ) ;
  assign n14750 = x93 &  n6982 ;
  assign n14747 = ( x95 & ~n6727 ) | ( x95 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n14748 = x94 &  n6722 ;
  assign n14749 = n14747 | n14748 ;
  assign n14751 = ( x93 & ~n14750 ) | ( x93 & n14749 ) | ( ~n14750 & n14749 ) ;
  assign n14752 = ( n2547 & ~n6730 ) | ( n2547 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n14753 = n14751 | n14752 ;
  assign n14754 = ( x53 & ~n14753 ) | ( x53 & 1'b0 ) | ( ~n14753 & 1'b0 ) ;
  assign n14755 = ~x53 & n14753 ;
  assign n14756 = n14754 | n14755 ;
  assign n14757 = ( n14317 & ~n14546 ) | ( n14317 & n14556 ) | ( ~n14546 & n14556 ) ;
  assign n14758 = ( n14746 & ~n14756 ) | ( n14746 & n14757 ) | ( ~n14756 & n14757 ) ;
  assign n14759 = ( n14746 & ~n14757 ) | ( n14746 & n14756 ) | ( ~n14757 & n14756 ) ;
  assign n14760 = ( n14758 & ~n14746 ) | ( n14758 & n14759 ) | ( ~n14746 & n14759 ) ;
  assign n14764 = x96 &  n6288 ;
  assign n14761 = ( x98 & ~n6032 ) | ( x98 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n14762 = x97 &  n6027 ;
  assign n14763 = n14761 | n14762 ;
  assign n14765 = ( x96 & ~n14764 ) | ( x96 & n14763 ) | ( ~n14764 & n14763 ) ;
  assign n14766 = ( n3170 & ~n6035 ) | ( n3170 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n14767 = n14765 | n14766 ;
  assign n14768 = ( x50 & ~n14767 ) | ( x50 & 1'b0 ) | ( ~n14767 & 1'b0 ) ;
  assign n14769 = ~x50 & n14767 ;
  assign n14770 = n14768 | n14769 ;
  assign n14772 = ( n14561 & n14760 ) | ( n14561 & n14770 ) | ( n14760 & n14770 ) ;
  assign n14771 = ( n14760 & ~n14561 ) | ( n14760 & n14770 ) | ( ~n14561 & n14770 ) ;
  assign n14773 = ( n14561 & ~n14772 ) | ( n14561 & n14771 ) | ( ~n14772 & n14771 ) ;
  assign n14777 = x99 &  n5586 ;
  assign n14774 = ( x101 & ~n5389 ) | ( x101 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n14775 = x100 &  n5384 ;
  assign n14776 = n14774 | n14775 ;
  assign n14778 = ( x99 & ~n14777 ) | ( x99 & n14776 ) | ( ~n14777 & n14776 ) ;
  assign n14779 = n3694 | n5392 ;
  assign n14780 = ~n14778 & n14779 ;
  assign n14781 = x47 &  n14780 ;
  assign n14782 = x47 | n14780 ;
  assign n14783 = ~n14781 & n14782 ;
  assign n14785 = ( n14565 & n14773 ) | ( n14565 & n14783 ) | ( n14773 & n14783 ) ;
  assign n14784 = ( n14773 & ~n14565 ) | ( n14773 & n14783 ) | ( ~n14565 & n14783 ) ;
  assign n14786 = ( n14565 & ~n14785 ) | ( n14565 & n14784 ) | ( ~n14785 & n14784 ) ;
  assign n14787 = ( n14692 & n14702 ) | ( n14692 & n14786 ) | ( n14702 & n14786 ) ;
  assign n14788 = ( n14702 & ~n14692 ) | ( n14702 & n14786 ) | ( ~n14692 & n14786 ) ;
  assign n14789 = ( n14692 & ~n14787 ) | ( n14692 & n14788 ) | ( ~n14787 & n14788 ) ;
  assign n14790 = ( n14681 & n14691 ) | ( n14681 & n14789 ) | ( n14691 & n14789 ) ;
  assign n14791 = ( n14691 & ~n14681 ) | ( n14691 & n14789 ) | ( ~n14681 & n14789 ) ;
  assign n14792 = ( n14681 & ~n14790 ) | ( n14681 & n14791 ) | ( ~n14790 & n14791 ) ;
  assign n14803 = ( n14680 & ~n14802 ) | ( n14680 & n14792 ) | ( ~n14802 & n14792 ) ;
  assign n14804 = ( n14680 & ~n14792 ) | ( n14680 & n14802 ) | ( ~n14792 & n14802 ) ;
  assign n14805 = ( n14803 & ~n14680 ) | ( n14803 & n14804 ) | ( ~n14680 & n14804 ) ;
  assign n14809 = x111 &  n3214 ;
  assign n14806 = ( x113 & ~n3087 ) | ( x113 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n14807 = x112 &  n3082 ;
  assign n14808 = n14806 | n14807 ;
  assign n14810 = ( x111 & ~n14809 ) | ( x111 & n14808 ) | ( ~n14809 & n14808 ) ;
  assign n14811 = n3090 | n6169 ;
  assign n14812 = ~n14810 & n14811 ;
  assign n14813 = x35 &  n14812 ;
  assign n14814 = x35 | n14812 ;
  assign n14815 = ~n14813 & n14814 ;
  assign n14816 = ( n14610 & n14805 ) | ( n14610 & n14815 ) | ( n14805 & n14815 ) ;
  assign n14817 = ( n14805 & ~n14610 ) | ( n14805 & n14815 ) | ( ~n14610 & n14815 ) ;
  assign n14818 = ( n14610 & ~n14816 ) | ( n14610 & n14817 ) | ( ~n14816 & n14817 ) ;
  assign n14822 = ( n14679 & n14818 ) | ( n14679 & n14821 ) | ( n14818 & n14821 ) ;
  assign n14823 = ( n14679 & ~n14821 ) | ( n14679 & n14818 ) | ( ~n14821 & n14818 ) ;
  assign n14824 = ( n14821 & ~n14822 ) | ( n14821 & n14823 ) | ( ~n14822 & n14823 ) ;
  assign n14825 = ( n14619 & n14672 ) | ( n14619 & n14824 ) | ( n14672 & n14824 ) ;
  assign n14826 = ( n14619 & ~n14672 ) | ( n14619 & n14824 ) | ( ~n14672 & n14824 ) ;
  assign n14827 = ( n14672 & ~n14825 ) | ( n14672 & n14826 ) | ( ~n14825 & n14826 ) ;
  assign n14828 = n14662 | n14827 ;
  assign n14829 = n14662 &  n14827 ;
  assign n14830 = ( n14828 & ~n14829 ) | ( n14828 & 1'b0 ) | ( ~n14829 & 1'b0 ) ;
  assign n14831 = ( n14451 & ~n14624 ) | ( n14451 & n14626 ) | ( ~n14624 & n14626 ) ;
  assign n14832 = ( n14651 & ~n14830 ) | ( n14651 & n14831 ) | ( ~n14830 & n14831 ) ;
  assign n14833 = ( n14651 & ~n14831 ) | ( n14651 & n14830 ) | ( ~n14831 & n14830 ) ;
  assign n14834 = ( n14832 & ~n14651 ) | ( n14832 & n14833 ) | ( ~n14651 & n14833 ) ;
  assign n14835 = ( x126 & ~n1227 ) | ( x126 & 1'b0 ) | ( ~n1227 & 1'b0 ) ;
  assign n14836 = x127 &  n1149 ;
  assign n14837 = n14835 | n14836 ;
  assign n14838 = n1157 | n9960 ;
  assign n14839 = ( n14837 & ~n1157 ) | ( n14837 & n14838 ) | ( ~n1157 & n14838 ) ;
  assign n14840 = x20 | n14839 ;
  assign n14841 = ( x20 & ~n14839 ) | ( x20 & 1'b0 ) | ( ~n14839 & 1'b0 ) ;
  assign n14842 = ( n14840 & ~x20 ) | ( n14840 & n14841 ) | ( ~x20 & n14841 ) ;
  assign n14843 = ( n14641 & ~n14834 ) | ( n14641 & n14842 ) | ( ~n14834 & n14842 ) ;
  assign n14844 = ( n14641 & ~n14842 ) | ( n14641 & n14834 ) | ( ~n14842 & n14834 ) ;
  assign n14845 = ( n14843 & ~n14641 ) | ( n14843 & n14844 ) | ( ~n14641 & n14844 ) ;
  assign n14846 = ( n14639 & ~n14640 ) | ( n14639 & n14845 ) | ( ~n14640 & n14845 ) ;
  assign n14847 = ( n14639 & ~n14845 ) | ( n14639 & n14640 ) | ( ~n14845 & n14640 ) ;
  assign n14848 = ( n14846 & ~n14639 ) | ( n14846 & n14847 ) | ( ~n14639 & n14847 ) ;
  assign n14850 = ( x127 & ~n1227 ) | ( x127 & 1'b0 ) | ( ~n1227 & 1'b0 ) ;
  assign n14851 = n1157 | n10258 ;
  assign n14852 = ~n14850 & n14851 ;
  assign n14853 = ~x20 & n14852 ;
  assign n14854 = ( x20 & ~n14852 ) | ( x20 & 1'b0 ) | ( ~n14852 & 1'b0 ) ;
  assign n14855 = n14853 | n14854 ;
  assign n14856 = ( n14651 & n14830 ) | ( n14651 & n14831 ) | ( n14830 & n14831 ) ;
  assign n14857 = x26 &  n14658 ;
  assign n14858 = ( n14828 & ~n14660 ) | ( n14828 & n14857 ) | ( ~n14660 & n14857 ) ;
  assign n14862 = x124 &  n1551 ;
  assign n14859 = ( x126 & ~n1451 ) | ( x126 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n14860 = x125 &  n1446 ;
  assign n14861 = n14859 | n14860 ;
  assign n14863 = ( x124 & ~n14862 ) | ( x124 & n14861 ) | ( ~n14862 & n14861 ) ;
  assign n14864 = n1454 | n9349 ;
  assign n14865 = ~n14863 & n14864 ;
  assign n14866 = x23 &  n14865 ;
  assign n14867 = x23 | n14865 ;
  assign n14868 = ~n14866 & n14867 ;
  assign n14869 = ( n14619 & ~n14824 ) | ( n14619 & n14672 ) | ( ~n14824 & n14672 ) ;
  assign n14873 = x121 &  n1894 ;
  assign n14870 = ( x123 & ~n1816 ) | ( x123 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n14871 = x122 &  n1811 ;
  assign n14872 = n14870 | n14871 ;
  assign n14874 = ( x121 & ~n14873 ) | ( x121 & n14872 ) | ( ~n14873 & n14872 ) ;
  assign n14875 = ~n1819 & n8472 ;
  assign n14876 = n14874 | n14875 ;
  assign n14877 = ( x26 & ~n14876 ) | ( x26 & 1'b0 ) | ( ~n14876 & 1'b0 ) ;
  assign n14878 = ~x26 & n14876 ;
  assign n14879 = n14877 | n14878 ;
  assign n14880 = ~x32 & n14679 ;
  assign n14881 = ( x32 & ~n14679 ) | ( x32 & 1'b0 ) | ( ~n14679 & 1'b0 ) ;
  assign n14882 = n14880 | n14881 ;
  assign n14883 = ( n14614 & ~n14882 ) | ( n14614 & n14818 ) | ( ~n14882 & n14818 ) ;
  assign n14887 = x118 &  n2312 ;
  assign n14884 = ( x120 & ~n2195 ) | ( x120 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n14885 = x119 &  n2190 ;
  assign n14886 = n14884 | n14885 ;
  assign n14888 = ( x118 & ~n14887 ) | ( x118 & n14886 ) | ( ~n14887 & n14886 ) ;
  assign n14889 = ~n2198 & n9364 ;
  assign n14890 = n14888 | n14889 ;
  assign n14891 = ( x29 & ~n14890 ) | ( x29 & 1'b0 ) | ( ~n14890 & 1'b0 ) ;
  assign n14892 = ~x29 & n14890 ;
  assign n14893 = n14891 | n14892 ;
  assign n14897 = x115 &  n2718 ;
  assign n14894 = ( x117 & ~n2642 ) | ( x117 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n14895 = x116 &  n2637 ;
  assign n14896 = n14894 | n14895 ;
  assign n14898 = ( x115 & ~n14897 ) | ( x115 & n14896 ) | ( ~n14897 & n14896 ) ;
  assign n14899 = n2645 | n7136 ;
  assign n14900 = ~n14898 & n14899 ;
  assign n14901 = x32 &  n14900 ;
  assign n14902 = x32 | n14900 ;
  assign n14903 = ~n14901 & n14902 ;
  assign n14908 = x106 &  n4344 ;
  assign n14905 = ( x108 & ~n4143 ) | ( x108 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n14906 = x107 &  n4138 ;
  assign n14907 = n14905 | n14906 ;
  assign n14909 = ( x106 & ~n14908 ) | ( x106 & n14907 ) | ( ~n14908 & n14907 ) ;
  assign n14910 = n4146 | n5055 ;
  assign n14911 = ~n14909 & n14910 ;
  assign n14912 = x41 &  n14911 ;
  assign n14913 = x41 | n14911 ;
  assign n14914 = ~n14912 & n14913 ;
  assign n14915 = ( n14565 & ~n14783 ) | ( n14565 & n14773 ) | ( ~n14783 & n14773 ) ;
  assign n14919 = x103 &  n4934 ;
  assign n14916 = ( x105 & ~n4725 ) | ( x105 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n14917 = x104 &  n4720 ;
  assign n14918 = n14916 | n14917 ;
  assign n14920 = ( x103 & ~n14919 ) | ( x103 & n14918 ) | ( ~n14919 & n14918 ) ;
  assign n14921 = ( n4442 & ~n4728 ) | ( n4442 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n14922 = n14920 | n14921 ;
  assign n14923 = ( x44 & ~n14922 ) | ( x44 & 1'b0 ) | ( ~n14922 & 1'b0 ) ;
  assign n14924 = ~x44 & n14922 ;
  assign n14925 = n14923 | n14924 ;
  assign n14926 = ( n14561 & ~n14770 ) | ( n14561 & n14760 ) | ( ~n14770 & n14760 ) ;
  assign n14930 = x100 &  n5586 ;
  assign n14927 = ( x102 & ~n5389 ) | ( x102 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n14928 = x101 &  n5384 ;
  assign n14929 = n14927 | n14928 ;
  assign n14931 = ( x100 & ~n14930 ) | ( x100 & n14929 ) | ( ~n14930 & n14929 ) ;
  assign n14932 = n3872 | n5392 ;
  assign n14933 = ~n14931 & n14932 ;
  assign n14934 = x47 &  n14933 ;
  assign n14935 = x47 | n14933 ;
  assign n14936 = ~n14934 & n14935 ;
  assign n14937 = ( n14756 & ~n14746 ) | ( n14756 & n14757 ) | ( ~n14746 & n14757 ) ;
  assign n14941 = x97 &  n6288 ;
  assign n14938 = ( x99 & ~n6032 ) | ( x99 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n14939 = x98 &  n6027 ;
  assign n14940 = n14938 | n14939 ;
  assign n14942 = ( x97 & ~n14941 ) | ( x97 & n14940 ) | ( ~n14941 & n14940 ) ;
  assign n14943 = ( n3338 & ~n6035 ) | ( n3338 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n14944 = n14942 | n14943 ;
  assign n14945 = ( x50 & ~n14944 ) | ( x50 & 1'b0 ) | ( ~n14944 & 1'b0 ) ;
  assign n14946 = ~x50 & n14944 ;
  assign n14947 = n14945 | n14946 ;
  assign n14948 = ( n14733 & ~n14732 ) | ( n14733 & n14743 ) | ( ~n14732 & n14743 ) ;
  assign n14949 = ( n14703 & ~n14716 ) | ( n14703 & n14713 ) | ( ~n14716 & n14713 ) ;
  assign n14953 = x88 &  n8558 ;
  assign n14950 = ( x90 & ~n8314 ) | ( x90 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n14951 = x89 &  n8309 ;
  assign n14952 = n14950 | n14951 ;
  assign n14954 = ( x88 & ~n14953 ) | ( x88 & n14952 ) | ( ~n14953 & n14952 ) ;
  assign n14955 = ( n1976 & ~n8317 ) | ( n1976 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n14956 = n14954 | n14955 ;
  assign n14957 = ( x59 & ~n14956 ) | ( x59 & 1'b0 ) | ( ~n14956 & 1'b0 ) ;
  assign n14958 = ~x59 & n14956 ;
  assign n14959 = n14957 | n14958 ;
  assign n14960 = x83 &  n10104 ;
  assign n14961 = ( x84 & ~n9760 ) | ( x84 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n14962 = n14960 | n14961 ;
  assign n14966 = x85 &  n9457 ;
  assign n14963 = ( x87 & ~n9150 ) | ( x87 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n14964 = x86 &  n9145 ;
  assign n14965 = n14963 | n14964 ;
  assign n14967 = ( x85 & ~n14966 ) | ( x85 & n14965 ) | ( ~n14966 & n14965 ) ;
  assign n14968 = ( n1512 & ~n14967 ) | ( n1512 & n9153 ) | ( ~n14967 & n9153 ) ;
  assign n14969 = ~n9153 & n14968 ;
  assign n14970 = ( x62 & n14967 ) | ( x62 & n14969 ) | ( n14967 & n14969 ) ;
  assign n14971 = ( x62 & ~n14969 ) | ( x62 & n14967 ) | ( ~n14969 & n14967 ) ;
  assign n14972 = ( n14969 & ~n14970 ) | ( n14969 & n14971 ) | ( ~n14970 & n14971 ) ;
  assign n14973 = ( n14962 & ~n14716 ) | ( n14962 & n14972 ) | ( ~n14716 & n14972 ) ;
  assign n14974 = ( n14716 & ~n14972 ) | ( n14716 & n14962 ) | ( ~n14972 & n14962 ) ;
  assign n14975 = ( n14973 & ~n14962 ) | ( n14973 & n14974 ) | ( ~n14962 & n14974 ) ;
  assign n14976 = ( n14949 & ~n14959 ) | ( n14949 & n14975 ) | ( ~n14959 & n14975 ) ;
  assign n14977 = ( n14949 & ~n14975 ) | ( n14949 & n14959 ) | ( ~n14975 & n14959 ) ;
  assign n14978 = ( n14976 & ~n14949 ) | ( n14976 & n14977 ) | ( ~n14949 & n14977 ) ;
  assign n14979 = ( n14531 & ~n14719 ) | ( n14531 & n14729 ) | ( ~n14719 & n14729 ) ;
  assign n14983 = x91 &  n7731 ;
  assign n14980 = ( x93 & ~n7538 ) | ( x93 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n14981 = x92 &  n7533 ;
  assign n14982 = n14980 | n14981 ;
  assign n14984 = ( x91 & ~n14983 ) | ( x91 & n14982 ) | ( ~n14983 & n14982 ) ;
  assign n14985 = n2264 | n7541 ;
  assign n14986 = ~n14984 & n14985 ;
  assign n14987 = x56 &  n14986 ;
  assign n14988 = x56 | n14986 ;
  assign n14989 = ~n14987 & n14988 ;
  assign n14991 = ( n14978 & n14979 ) | ( n14978 & n14989 ) | ( n14979 & n14989 ) ;
  assign n14990 = ( n14979 & ~n14978 ) | ( n14979 & n14989 ) | ( ~n14978 & n14989 ) ;
  assign n14992 = ( n14978 & ~n14991 ) | ( n14978 & n14990 ) | ( ~n14991 & n14990 ) ;
  assign n14996 = x94 &  n6982 ;
  assign n14993 = ( x96 & ~n6727 ) | ( x96 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n14994 = x95 &  n6722 ;
  assign n14995 = n14993 | n14994 ;
  assign n14997 = ( x94 & ~n14996 ) | ( x94 & n14995 ) | ( ~n14996 & n14995 ) ;
  assign n14998 = ( n2836 & ~n6730 ) | ( n2836 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n14999 = n14997 | n14998 ;
  assign n15000 = ( x53 & ~n14999 ) | ( x53 & 1'b0 ) | ( ~n14999 & 1'b0 ) ;
  assign n15001 = ~x53 & n14999 ;
  assign n15002 = n15000 | n15001 ;
  assign n15003 = ( n14948 & ~n14992 ) | ( n14948 & n15002 ) | ( ~n14992 & n15002 ) ;
  assign n15004 = ( n14948 & ~n15002 ) | ( n14948 & n14992 ) | ( ~n15002 & n14992 ) ;
  assign n15005 = ( n15003 & ~n14948 ) | ( n15003 & n15004 ) | ( ~n14948 & n15004 ) ;
  assign n15006 = ( n14937 & ~n14947 ) | ( n14937 & n15005 ) | ( ~n14947 & n15005 ) ;
  assign n15007 = ( n14937 & ~n15005 ) | ( n14937 & n14947 ) | ( ~n15005 & n14947 ) ;
  assign n15008 = ( n15006 & ~n14937 ) | ( n15006 & n15007 ) | ( ~n14937 & n15007 ) ;
  assign n15009 = ( n14926 & ~n14936 ) | ( n14926 & n15008 ) | ( ~n14936 & n15008 ) ;
  assign n15010 = ( n14926 & ~n15008 ) | ( n14926 & n14936 ) | ( ~n15008 & n14936 ) ;
  assign n15011 = ( n15009 & ~n14926 ) | ( n15009 & n15010 ) | ( ~n14926 & n15010 ) ;
  assign n15013 = ( n14915 & n14925 ) | ( n14915 & n15011 ) | ( n14925 & n15011 ) ;
  assign n15012 = ( n14925 & ~n14915 ) | ( n14925 & n15011 ) | ( ~n14915 & n15011 ) ;
  assign n15014 = ( n14915 & ~n15013 ) | ( n14915 & n15012 ) | ( ~n15013 & n15012 ) ;
  assign n15015 = ( n14788 & ~n14914 ) | ( n14788 & n15014 ) | ( ~n14914 & n15014 ) ;
  assign n15016 = ( n14788 & ~n15014 ) | ( n14788 & n14914 ) | ( ~n15014 & n14914 ) ;
  assign n15017 = ( n15015 & ~n14788 ) | ( n15015 & n15016 ) | ( ~n14788 & n15016 ) ;
  assign n15021 = x109 &  n3756 ;
  assign n15018 = ( x111 & ~n3602 ) | ( x111 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n15019 = x110 &  n3597 ;
  assign n15020 = n15018 | n15019 ;
  assign n15022 = ( x109 & ~n15021 ) | ( x109 & n15020 ) | ( ~n15021 & n15020 ) ;
  assign n15023 = n3605 | n5711 ;
  assign n15024 = ~n15022 & n15023 ;
  assign n15025 = x38 &  n15024 ;
  assign n15026 = x38 | n15024 ;
  assign n15027 = ~n15025 & n15026 ;
  assign n15028 = ( n14791 & n15017 ) | ( n14791 & n15027 ) | ( n15017 & n15027 ) ;
  assign n15029 = ( n14791 & ~n15017 ) | ( n14791 & n15027 ) | ( ~n15017 & n15027 ) ;
  assign n15030 = ( n15017 & ~n15028 ) | ( n15017 & n15029 ) | ( ~n15028 & n15029 ) ;
  assign n14904 = ( n14792 & ~n14680 ) | ( n14792 & n14802 ) | ( ~n14680 & n14802 ) ;
  assign n15034 = x112 &  n3214 ;
  assign n15031 = ( x114 & ~n3087 ) | ( x114 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n15032 = x113 &  n3082 ;
  assign n15033 = n15031 | n15032 ;
  assign n15035 = ( x112 & ~n15034 ) | ( x112 & n15033 ) | ( ~n15034 & n15033 ) ;
  assign n15036 = n3090 | n6185 ;
  assign n15037 = ~n15035 & n15036 ;
  assign n15038 = x35 &  n15037 ;
  assign n15039 = x35 | n15037 ;
  assign n15040 = ~n15038 & n15039 ;
  assign n15042 = ( n14904 & n15030 ) | ( n14904 & n15040 ) | ( n15030 & n15040 ) ;
  assign n15041 = ( n14904 & ~n15030 ) | ( n14904 & n15040 ) | ( ~n15030 & n15040 ) ;
  assign n15043 = ( n15030 & ~n15042 ) | ( n15030 & n15041 ) | ( ~n15042 & n15041 ) ;
  assign n15044 = ( n14610 & ~n14805 ) | ( n14610 & n14815 ) | ( ~n14805 & n14815 ) ;
  assign n15045 = ( n14903 & ~n15043 ) | ( n14903 & n15044 ) | ( ~n15043 & n15044 ) ;
  assign n15046 = ( n14903 & ~n15044 ) | ( n14903 & n15043 ) | ( ~n15044 & n15043 ) ;
  assign n15047 = ( n15045 & ~n14903 ) | ( n15045 & n15046 ) | ( ~n14903 & n15046 ) ;
  assign n15049 = ( n14883 & n14893 ) | ( n14883 & n15047 ) | ( n14893 & n15047 ) ;
  assign n15048 = ( n14893 & ~n14883 ) | ( n14893 & n15047 ) | ( ~n14883 & n15047 ) ;
  assign n15050 = ( n14883 & ~n15049 ) | ( n14883 & n15048 ) | ( ~n15049 & n15048 ) ;
  assign n15052 = ( n14869 & n14879 ) | ( n14869 & n15050 ) | ( n14879 & n15050 ) ;
  assign n15051 = ( n14879 & ~n14869 ) | ( n14879 & n15050 ) | ( ~n14869 & n15050 ) ;
  assign n15053 = ( n14869 & ~n15052 ) | ( n14869 & n15051 ) | ( ~n15052 & n15051 ) ;
  assign n15054 = ( n14858 & ~n14868 ) | ( n14858 & n15053 ) | ( ~n14868 & n15053 ) ;
  assign n15055 = ( n14858 & ~n15053 ) | ( n14858 & n14868 ) | ( ~n15053 & n14868 ) ;
  assign n15056 = ( n15054 & ~n14858 ) | ( n15054 & n15055 ) | ( ~n14858 & n15055 ) ;
  assign n15057 = ( n14855 & n14856 ) | ( n14855 & n15056 ) | ( n14856 & n15056 ) ;
  assign n15058 = ( n14856 & ~n14855 ) | ( n14856 & n15056 ) | ( ~n14855 & n15056 ) ;
  assign n15059 = ( n14855 & ~n15057 ) | ( n14855 & n15058 ) | ( ~n15057 & n15058 ) ;
  assign n14849 = ( n14641 & n14834 ) | ( n14641 & n14842 ) | ( n14834 & n14842 ) ;
  assign n15060 = ( n14847 & ~n15059 ) | ( n14847 & n14849 ) | ( ~n15059 & n14849 ) ;
  assign n15061 = ( n14849 & ~n14847 ) | ( n14849 & n15059 ) | ( ~n14847 & n15059 ) ;
  assign n15062 = ( n15060 & ~n14849 ) | ( n15060 & n15061 ) | ( ~n14849 & n15061 ) ;
  assign n15063 = ( n14855 & ~n14856 ) | ( n14855 & n15056 ) | ( ~n14856 & n15056 ) ;
  assign n15064 = ( n14858 & n14868 ) | ( n14858 & n15053 ) | ( n14868 & n15053 ) ;
  assign n15068 = x122 &  n1894 ;
  assign n15065 = ( x124 & ~n1816 ) | ( x124 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n15066 = x123 &  n1811 ;
  assign n15067 = n15065 | n15066 ;
  assign n15069 = ( x122 & ~n15068 ) | ( x122 & n15067 ) | ( ~n15068 & n15067 ) ;
  assign n15070 = ~n1819 & n8755 ;
  assign n15071 = n15069 | n15070 ;
  assign n15242 = x26 | n15071 ;
  assign n15243 = ~x26 & n15071 ;
  assign n15244 = ( n15242 & ~n15071 ) | ( n15242 & n15243 ) | ( ~n15071 & n15243 ) ;
  assign n15072 = ( n14869 & ~n15050 ) | ( n14869 & n14879 ) | ( ~n15050 & n14879 ) ;
  assign n15073 = ( n14883 & ~n15047 ) | ( n14883 & n14893 ) | ( ~n15047 & n14893 ) ;
  assign n15077 = x116 &  n2718 ;
  assign n15074 = ( x118 & ~n2642 ) | ( x118 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n15075 = x117 &  n2637 ;
  assign n15076 = n15074 | n15075 ;
  assign n15078 = ( x116 & ~n15077 ) | ( x116 & n15076 ) | ( ~n15077 & n15076 ) ;
  assign n15079 = n2645 | n7152 ;
  assign n15080 = ~n15078 & n15079 ;
  assign n15223 = ~x32 & n15080 ;
  assign n15224 = x32 | n15080 ;
  assign n15225 = ( n15223 & ~n15080 ) | ( n15223 & n15224 ) | ( ~n15080 & n15224 ) ;
  assign n15081 = ( n14903 & n15043 ) | ( n14903 & n15044 ) | ( n15043 & n15044 ) ;
  assign n15085 = x110 &  n3756 ;
  assign n15082 = ( x112 & ~n3602 ) | ( x112 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n15083 = x111 &  n3597 ;
  assign n15084 = n15082 | n15083 ;
  assign n15086 = ( x110 & ~n15085 ) | ( x110 & n15084 ) | ( ~n15085 & n15084 ) ;
  assign n15087 = ~n3605 & n5727 ;
  assign n15088 = n15086 | n15087 ;
  assign n15089 = ( x38 & ~n15088 ) | ( x38 & 1'b0 ) | ( ~n15088 & 1'b0 ) ;
  assign n15090 = ~x38 & n15088 ;
  assign n15091 = n15089 | n15090 ;
  assign n15095 = x107 &  n4344 ;
  assign n15092 = ( x109 & ~n4143 ) | ( x109 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n15093 = x108 &  n4138 ;
  assign n15094 = n15092 | n15093 ;
  assign n15096 = ( x107 & ~n15095 ) | ( x107 & n15094 ) | ( ~n15095 & n15094 ) ;
  assign n15097 = ~n4146 & n5267 ;
  assign n15098 = n15096 | n15097 ;
  assign n15099 = ( x41 & ~n15098 ) | ( x41 & 1'b0 ) | ( ~n15098 & 1'b0 ) ;
  assign n15100 = ~x41 & n15098 ;
  assign n15101 = n15099 | n15100 ;
  assign n15115 = x101 &  n5586 ;
  assign n15112 = ( x103 & ~n5389 ) | ( x103 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n15113 = x102 &  n5384 ;
  assign n15114 = n15112 | n15113 ;
  assign n15116 = ( x101 & ~n15115 ) | ( x101 & n15114 ) | ( ~n15115 & n15114 ) ;
  assign n15117 = n4056 | n5392 ;
  assign n15118 = ~n15116 & n15117 ;
  assign n15119 = x47 &  n15118 ;
  assign n15120 = x47 | n15118 ;
  assign n15121 = ~n15119 & n15120 ;
  assign n15125 = x95 &  n6982 ;
  assign n15122 = ( x97 & ~n6727 ) | ( x97 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n15123 = x96 &  n6722 ;
  assign n15124 = n15122 | n15123 ;
  assign n15126 = ( x95 & ~n15125 ) | ( x95 & n15124 ) | ( ~n15125 & n15124 ) ;
  assign n15127 = ( n2999 & ~n6730 ) | ( n2999 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n15128 = n15126 | n15127 ;
  assign n15129 = ( x53 & ~n15128 ) | ( x53 & 1'b0 ) | ( ~n15128 & 1'b0 ) ;
  assign n15130 = ~x53 & n15128 ;
  assign n15131 = n15129 | n15130 ;
  assign n15135 = x92 &  n7731 ;
  assign n15132 = ( x94 & ~n7538 ) | ( x94 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n15133 = x93 &  n7533 ;
  assign n15134 = n15132 | n15133 ;
  assign n15136 = ( x92 & ~n15135 ) | ( x92 & n15134 ) | ( ~n15135 & n15134 ) ;
  assign n15137 = ( n2401 & ~n7541 ) | ( n2401 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n15138 = n15136 | n15137 ;
  assign n15139 = ( x56 & ~n15138 ) | ( x56 & 1'b0 ) | ( ~n15138 & 1'b0 ) ;
  assign n15140 = ~x56 & n15138 ;
  assign n15141 = n15139 | n15140 ;
  assign n15145 = x89 &  n8558 ;
  assign n15142 = ( x91 & ~n8314 ) | ( x91 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n15143 = x90 &  n8309 ;
  assign n15144 = n15142 | n15143 ;
  assign n15146 = ( x89 & ~n15145 ) | ( x89 & n15144 ) | ( ~n15145 & n15144 ) ;
  assign n15147 = ( n2108 & ~n8317 ) | ( n2108 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n15148 = n15146 | n15147 ;
  assign n15149 = ( x59 & ~n15148 ) | ( x59 & 1'b0 ) | ( ~n15148 & 1'b0 ) ;
  assign n15150 = ~x59 & n15148 ;
  assign n15151 = n15149 | n15150 ;
  assign n15155 = x86 &  n9457 ;
  assign n15152 = ( x88 & ~n9150 ) | ( x88 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n15153 = x87 &  n9145 ;
  assign n15154 = n15152 | n15153 ;
  assign n15156 = ( x86 & ~n15155 ) | ( x86 & n15154 ) | ( ~n15155 & n15154 ) ;
  assign n15157 = ( n1624 & ~n9153 ) | ( n1624 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n15158 = n15156 | n15157 ;
  assign n15159 = ( x62 & ~n15158 ) | ( x62 & 1'b0 ) | ( ~n15158 & 1'b0 ) ;
  assign n15160 = ~x62 & n15158 ;
  assign n15161 = n15159 | n15160 ;
  assign n15162 = x84 &  n10104 ;
  assign n15163 = ( x85 & ~n9760 ) | ( x85 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n15164 = n15162 | n15163 ;
  assign n15165 = ( x20 & n14962 ) | ( x20 & n15164 ) | ( n14962 & n15164 ) ;
  assign n15166 = ( x20 & ~n14962 ) | ( x20 & n15164 ) | ( ~n14962 & n15164 ) ;
  assign n15167 = ( n14962 & ~n15165 ) | ( n14962 & n15166 ) | ( ~n15165 & n15166 ) ;
  assign n15168 = ( n14716 & ~n14962 ) | ( n14716 & n14972 ) | ( ~n14962 & n14972 ) ;
  assign n15169 = ( n15161 & ~n15167 ) | ( n15161 & n15168 ) | ( ~n15167 & n15168 ) ;
  assign n15170 = ( n15161 & ~n15168 ) | ( n15161 & n15167 ) | ( ~n15168 & n15167 ) ;
  assign n15171 = ( n15169 & ~n15161 ) | ( n15169 & n15170 ) | ( ~n15161 & n15170 ) ;
  assign n15172 = ( n14977 & n15151 ) | ( n14977 & n15171 ) | ( n15151 & n15171 ) ;
  assign n15173 = ( n14977 & ~n15151 ) | ( n14977 & n15171 ) | ( ~n15151 & n15171 ) ;
  assign n15174 = ( n15151 & ~n15172 ) | ( n15151 & n15173 ) | ( ~n15172 & n15173 ) ;
  assign n15175 = ( n14978 & ~n14979 ) | ( n14978 & n14989 ) | ( ~n14979 & n14989 ) ;
  assign n15177 = ( n15141 & n15174 ) | ( n15141 & n15175 ) | ( n15174 & n15175 ) ;
  assign n15176 = ( n15174 & ~n15141 ) | ( n15174 & n15175 ) | ( ~n15141 & n15175 ) ;
  assign n15178 = ( n15141 & ~n15177 ) | ( n15141 & n15176 ) | ( ~n15177 & n15176 ) ;
  assign n15179 = ( n14948 & n14992 ) | ( n14948 & n15002 ) | ( n14992 & n15002 ) ;
  assign n15180 = ( n15131 & n15178 ) | ( n15131 & n15179 ) | ( n15178 & n15179 ) ;
  assign n15181 = ( n15178 & ~n15131 ) | ( n15178 & n15179 ) | ( ~n15131 & n15179 ) ;
  assign n15182 = ( n15131 & ~n15180 ) | ( n15131 & n15181 ) | ( ~n15180 & n15181 ) ;
  assign n15183 = ( n14937 & n14947 ) | ( n14937 & n15005 ) | ( n14947 & n15005 ) ;
  assign n15187 = x98 &  n6288 ;
  assign n15184 = ( x100 & ~n6032 ) | ( x100 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n15185 = x99 &  n6027 ;
  assign n15186 = n15184 | n15185 ;
  assign n15188 = ( x98 & ~n15187 ) | ( x98 & n15186 ) | ( ~n15187 & n15186 ) ;
  assign n15189 = n3354 | n6035 ;
  assign n15190 = ~n15188 & n15189 ;
  assign n15191 = x50 &  n15190 ;
  assign n15192 = x50 | n15190 ;
  assign n15193 = ~n15191 & n15192 ;
  assign n15195 = ( n15182 & n15183 ) | ( n15182 & n15193 ) | ( n15183 & n15193 ) ;
  assign n15194 = ( n15183 & ~n15182 ) | ( n15183 & n15193 ) | ( ~n15182 & n15193 ) ;
  assign n15196 = ( n15182 & ~n15195 ) | ( n15182 & n15194 ) | ( ~n15195 & n15194 ) ;
  assign n15197 = ( n15010 & n15121 ) | ( n15010 & n15196 ) | ( n15121 & n15196 ) ;
  assign n15198 = ( n15010 & ~n15121 ) | ( n15010 & n15196 ) | ( ~n15121 & n15196 ) ;
  assign n15199 = ( n15121 & ~n15197 ) | ( n15121 & n15198 ) | ( ~n15197 & n15198 ) ;
  assign n15105 = x104 &  n4934 ;
  assign n15102 = ( x106 & ~n4725 ) | ( x106 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n15103 = x105 &  n4720 ;
  assign n15104 = n15102 | n15103 ;
  assign n15106 = ( x104 & ~n15105 ) | ( x104 & n15104 ) | ( ~n15105 & n15104 ) ;
  assign n15107 = ( n4458 & ~n4728 ) | ( n4458 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n15108 = n15106 | n15107 ;
  assign n15109 = ( x44 & ~n15108 ) | ( x44 & 1'b0 ) | ( ~n15108 & 1'b0 ) ;
  assign n15110 = ~x44 & n15108 ;
  assign n15111 = n15109 | n15110 ;
  assign n15200 = ( n15013 & ~n15199 ) | ( n15013 & n15111 ) | ( ~n15199 & n15111 ) ;
  assign n15201 = ( n15111 & ~n15013 ) | ( n15111 & n15199 ) | ( ~n15013 & n15199 ) ;
  assign n15202 = ( n15200 & ~n15111 ) | ( n15200 & n15201 ) | ( ~n15111 & n15201 ) ;
  assign n15204 = ( n15016 & n15101 ) | ( n15016 & n15202 ) | ( n15101 & n15202 ) ;
  assign n15203 = ( n15016 & ~n15101 ) | ( n15016 & n15202 ) | ( ~n15101 & n15202 ) ;
  assign n15205 = ( n15101 & ~n15204 ) | ( n15101 & n15203 ) | ( ~n15204 & n15203 ) ;
  assign n15206 = ( n14791 & ~n15027 ) | ( n14791 & n15017 ) | ( ~n15027 & n15017 ) ;
  assign n15207 = ( n15091 & n15205 ) | ( n15091 & n15206 ) | ( n15205 & n15206 ) ;
  assign n15208 = ( n15205 & ~n15091 ) | ( n15205 & n15206 ) | ( ~n15091 & n15206 ) ;
  assign n15209 = ( n15091 & ~n15207 ) | ( n15091 & n15208 ) | ( ~n15207 & n15208 ) ;
  assign n15213 = x113 &  n3214 ;
  assign n15210 = ( x115 & ~n3087 ) | ( x115 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n15211 = x114 &  n3082 ;
  assign n15212 = n15210 | n15211 ;
  assign n15214 = ( x113 & ~n15213 ) | ( x113 & n15212 ) | ( ~n15213 & n15212 ) ;
  assign n15215 = ~n3090 & n6420 ;
  assign n15216 = n15214 | n15215 ;
  assign n15217 = ( x35 & ~n15216 ) | ( x35 & 1'b0 ) | ( ~n15216 & 1'b0 ) ;
  assign n15218 = ~x35 & n15216 ;
  assign n15219 = n15217 | n15218 ;
  assign n15221 = ( n15042 & n15209 ) | ( n15042 & n15219 ) | ( n15209 & n15219 ) ;
  assign n15220 = ( n15042 & ~n15209 ) | ( n15042 & n15219 ) | ( ~n15209 & n15219 ) ;
  assign n15222 = ( n15209 & ~n15221 ) | ( n15209 & n15220 ) | ( ~n15221 & n15220 ) ;
  assign n15227 = ( n15081 & n15222 ) | ( n15081 & n15225 ) | ( n15222 & n15225 ) ;
  assign n15226 = ( n15081 & ~n15225 ) | ( n15081 & n15222 ) | ( ~n15225 & n15222 ) ;
  assign n15228 = ( n15225 & ~n15227 ) | ( n15225 & n15226 ) | ( ~n15227 & n15226 ) ;
  assign n15232 = x119 &  n2312 ;
  assign n15229 = ( x121 & ~n2195 ) | ( x121 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n15230 = x120 &  n2190 ;
  assign n15231 = n15229 | n15230 ;
  assign n15233 = ( x119 & ~n15232 ) | ( x119 & n15231 ) | ( ~n15232 & n15231 ) ;
  assign n15234 = ~n2198 & n8176 ;
  assign n15235 = n15233 | n15234 ;
  assign n15236 = ( x29 & ~n15235 ) | ( x29 & 1'b0 ) | ( ~n15235 & 1'b0 ) ;
  assign n15237 = ~x29 & n15235 ;
  assign n15238 = n15236 | n15237 ;
  assign n15239 = ( n15073 & n15228 ) | ( n15073 & n15238 ) | ( n15228 & n15238 ) ;
  assign n15240 = ( n15228 & ~n15073 ) | ( n15228 & n15238 ) | ( ~n15073 & n15238 ) ;
  assign n15241 = ( n15073 & ~n15239 ) | ( n15073 & n15240 ) | ( ~n15239 & n15240 ) ;
  assign n15246 = ( n15072 & n15241 ) | ( n15072 & n15244 ) | ( n15241 & n15244 ) ;
  assign n15245 = ( n15072 & ~n15244 ) | ( n15072 & n15241 ) | ( ~n15244 & n15241 ) ;
  assign n15247 = ( n15244 & ~n15246 ) | ( n15244 & n15245 ) | ( ~n15246 & n15245 ) ;
  assign n15251 = x125 &  n1551 ;
  assign n15248 = ( x127 & ~n1451 ) | ( x127 & 1'b0 ) | ( ~n1451 & 1'b0 ) ;
  assign n15249 = x126 &  n1446 ;
  assign n15250 = n15248 | n15249 ;
  assign n15252 = ( x125 & ~n15251 ) | ( x125 & n15250 ) | ( ~n15251 & n15250 ) ;
  assign n15253 = n1454 | n9941 ;
  assign n15254 = ~n15252 & n15253 ;
  assign n15255 = x23 &  n15254 ;
  assign n15256 = x23 | n15254 ;
  assign n15257 = ~n15255 & n15256 ;
  assign n15258 = ( n15064 & ~n15247 ) | ( n15064 & n15257 ) | ( ~n15247 & n15257 ) ;
  assign n15259 = ( n15064 & ~n15257 ) | ( n15064 & n15247 ) | ( ~n15257 & n15247 ) ;
  assign n15260 = ( n15258 & ~n15064 ) | ( n15258 & n15259 ) | ( ~n15064 & n15259 ) ;
  assign n15262 = ( n15061 & n15063 ) | ( n15061 & n15260 ) | ( n15063 & n15260 ) ;
  assign n15261 = ( n15061 & ~n15063 ) | ( n15061 & n15260 ) | ( ~n15063 & n15260 ) ;
  assign n15263 = ( n15063 & ~n15262 ) | ( n15063 & n15261 ) | ( ~n15262 & n15261 ) ;
  assign n15264 = ( n15064 & n15247 ) | ( n15064 & n15257 ) | ( n15247 & n15257 ) ;
  assign n15265 = ( x26 & ~n15071 ) | ( x26 & 1'b0 ) | ( ~n15071 & 1'b0 ) ;
  assign n15266 = n15243 | n15265 ;
  assign n15267 = ( n15072 & ~n15241 ) | ( n15072 & n15266 ) | ( ~n15241 & n15266 ) ;
  assign n15271 = x123 &  n1894 ;
  assign n15268 = ( x125 & ~n1816 ) | ( x125 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n15269 = x124 &  n1811 ;
  assign n15270 = n15268 | n15269 ;
  assign n15272 = ( x123 & ~n15271 ) | ( x123 & n15270 ) | ( ~n15271 & n15270 ) ;
  assign n15273 = ~n1819 & n9324 ;
  assign n15274 = n15272 | n15273 ;
  assign n15275 = ( n15073 & ~n15228 ) | ( n15073 & n15238 ) | ( ~n15228 & n15238 ) ;
  assign n15276 = ( x26 & n15274 ) | ( x26 & n15275 ) | ( n15274 & n15275 ) ;
  assign n15277 = ( x26 & ~n15274 ) | ( x26 & n15275 ) | ( ~n15274 & n15275 ) ;
  assign n15278 = ( n15274 & ~n15276 ) | ( n15274 & n15277 ) | ( ~n15276 & n15277 ) ;
  assign n15296 = x120 &  n2312 ;
  assign n15293 = ( x122 & ~n2195 ) | ( x122 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n15294 = x121 &  n2190 ;
  assign n15295 = n15293 | n15294 ;
  assign n15297 = ( x120 & ~n15296 ) | ( x120 & n15295 ) | ( ~n15296 & n15295 ) ;
  assign n15298 = ( n2198 & n9987 ) | ( n2198 & n15297 ) | ( n9987 & n15297 ) ;
  assign n15299 = ( n9987 & ~n15298 ) | ( n9987 & 1'b0 ) | ( ~n15298 & 1'b0 ) ;
  assign n15300 = ( x29 & n15297 ) | ( x29 & n15299 ) | ( n15297 & n15299 ) ;
  assign n15301 = ( x29 & ~n15299 ) | ( x29 & n15297 ) | ( ~n15299 & n15297 ) ;
  assign n15302 = ( n15299 & ~n15300 ) | ( n15299 & n15301 ) | ( ~n15300 & n15301 ) ;
  assign n15403 = x108 &  n4344 ;
  assign n15400 = ( x110 & ~n4143 ) | ( x110 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n15401 = x109 &  n4138 ;
  assign n15402 = n15400 | n15401 ;
  assign n15404 = ( x108 & ~n15403 ) | ( x108 & n15402 ) | ( ~n15403 & n15402 ) ;
  assign n15405 = n4146 | n5283 ;
  assign n15406 = ~n15404 & n15405 ;
  assign n15407 = x41 &  n15406 ;
  assign n15408 = x41 | n15406 ;
  assign n15409 = ~n15407 & n15408 ;
  assign n15306 = x105 &  n4934 ;
  assign n15303 = ( x107 & ~n4725 ) | ( x107 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n15304 = x106 &  n4720 ;
  assign n15305 = n15303 | n15304 ;
  assign n15307 = ( x105 & ~n15306 ) | ( x105 & n15305 ) | ( ~n15306 & n15305 ) ;
  assign n15308 = ~n4728 & n4848 ;
  assign n15309 = n15307 | n15308 ;
  assign n15310 = ( x44 & ~n15309 ) | ( x44 & 1'b0 ) | ( ~n15309 & 1'b0 ) ;
  assign n15311 = ~x44 & n15309 ;
  assign n15312 = n15310 | n15311 ;
  assign n15313 = ( n15182 & ~n15193 ) | ( n15182 & n15183 ) | ( ~n15193 & n15183 ) ;
  assign n15317 = x102 &  n5586 ;
  assign n15314 = ( x104 & ~n5389 ) | ( x104 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n15315 = x103 &  n5384 ;
  assign n15316 = n15314 | n15315 ;
  assign n15318 = ( x102 & ~n15317 ) | ( x102 & n15316 ) | ( ~n15317 & n15316 ) ;
  assign n15319 = n4249 | n5392 ;
  assign n15320 = ~n15318 & n15319 ;
  assign n15321 = x47 &  n15320 ;
  assign n15322 = x47 | n15320 ;
  assign n15323 = ~n15321 & n15322 ;
  assign n15327 = x90 &  n8558 ;
  assign n15324 = ( x92 & ~n8314 ) | ( x92 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n15325 = x91 &  n8309 ;
  assign n15326 = n15324 | n15325 ;
  assign n15328 = ( x90 & ~n15327 ) | ( x90 & n15326 ) | ( ~n15327 & n15326 ) ;
  assign n15329 = ( n2248 & ~n8317 ) | ( n2248 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n15330 = n15328 | n15329 ;
  assign n15331 = ( x59 & ~n15330 ) | ( x59 & 1'b0 ) | ( ~n15330 & 1'b0 ) ;
  assign n15332 = ~x59 & n15330 ;
  assign n15333 = n15331 | n15332 ;
  assign n15334 = ( n14962 & ~x20 ) | ( n14962 & n15164 ) | ( ~x20 & n15164 ) ;
  assign n15338 = x87 &  n9457 ;
  assign n15335 = ( x89 & ~n9150 ) | ( x89 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n15336 = x88 &  n9145 ;
  assign n15337 = n15335 | n15336 ;
  assign n15339 = ( x87 & ~n15338 ) | ( x87 & n15337 ) | ( ~n15338 & n15337 ) ;
  assign n15340 = ( n1741 & ~n15339 ) | ( n1741 & n9153 ) | ( ~n15339 & n9153 ) ;
  assign n15341 = ~n9153 & n15340 ;
  assign n15342 = ( x62 & n15339 ) | ( x62 & n15341 ) | ( n15339 & n15341 ) ;
  assign n15343 = ( x62 & ~n15341 ) | ( x62 & n15339 ) | ( ~n15341 & n15339 ) ;
  assign n15344 = ( n15341 & ~n15342 ) | ( n15341 & n15343 ) | ( ~n15342 & n15343 ) ;
  assign n15345 = x85 &  n10104 ;
  assign n15346 = ( x86 & ~n9760 ) | ( x86 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n15347 = n15345 | n15346 ;
  assign n15349 = ( n15334 & n15344 ) | ( n15334 & n15347 ) | ( n15344 & n15347 ) ;
  assign n15348 = ( n15344 & ~n15334 ) | ( n15344 & n15347 ) | ( ~n15334 & n15347 ) ;
  assign n15350 = ( n15334 & ~n15349 ) | ( n15334 & n15348 ) | ( ~n15349 & n15348 ) ;
  assign n15351 = ( n15169 & ~n15333 ) | ( n15169 & n15350 ) | ( ~n15333 & n15350 ) ;
  assign n15352 = ( n15169 & ~n15350 ) | ( n15169 & n15333 ) | ( ~n15350 & n15333 ) ;
  assign n15353 = ( n15351 & ~n15169 ) | ( n15351 & n15352 ) | ( ~n15169 & n15352 ) ;
  assign n15354 = ( n14977 & ~n15171 ) | ( n14977 & n15151 ) | ( ~n15171 & n15151 ) ;
  assign n15358 = x93 &  n7731 ;
  assign n15355 = ( x95 & ~n7538 ) | ( x95 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n15356 = x94 &  n7533 ;
  assign n15357 = n15355 | n15356 ;
  assign n15359 = ( x93 & ~n15358 ) | ( x93 & n15357 ) | ( ~n15358 & n15357 ) ;
  assign n15360 = ( n2547 & ~n7541 ) | ( n2547 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n15361 = n15359 | n15360 ;
  assign n15362 = ( x56 & ~n15361 ) | ( x56 & 1'b0 ) | ( ~n15361 & 1'b0 ) ;
  assign n15363 = ~x56 & n15361 ;
  assign n15364 = n15362 | n15363 ;
  assign n15365 = ( n15353 & ~n15354 ) | ( n15353 & n15364 ) | ( ~n15354 & n15364 ) ;
  assign n15366 = ( n15353 & ~n15364 ) | ( n15353 & n15354 ) | ( ~n15364 & n15354 ) ;
  assign n15367 = ( n15365 & ~n15353 ) | ( n15365 & n15366 ) | ( ~n15353 & n15366 ) ;
  assign n15371 = x96 &  n6982 ;
  assign n15368 = ( x98 & ~n6727 ) | ( x98 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n15369 = x97 &  n6722 ;
  assign n15370 = n15368 | n15369 ;
  assign n15372 = ( x96 & ~n15371 ) | ( x96 & n15370 ) | ( ~n15371 & n15370 ) ;
  assign n15373 = ( n3170 & ~n6730 ) | ( n3170 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n15374 = n15372 | n15373 ;
  assign n15375 = ( x53 & ~n15374 ) | ( x53 & 1'b0 ) | ( ~n15374 & 1'b0 ) ;
  assign n15376 = ~x53 & n15374 ;
  assign n15377 = n15375 | n15376 ;
  assign n15379 = ( n15176 & n15367 ) | ( n15176 & n15377 ) | ( n15367 & n15377 ) ;
  assign n15378 = ( n15367 & ~n15176 ) | ( n15367 & n15377 ) | ( ~n15176 & n15377 ) ;
  assign n15380 = ( n15176 & ~n15379 ) | ( n15176 & n15378 ) | ( ~n15379 & n15378 ) ;
  assign n15384 = x99 &  n6288 ;
  assign n15381 = ( x101 & ~n6032 ) | ( x101 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n15382 = x100 &  n6027 ;
  assign n15383 = n15381 | n15382 ;
  assign n15385 = ( x99 & ~n15384 ) | ( x99 & n15383 ) | ( ~n15384 & n15383 ) ;
  assign n15386 = n3694 | n6035 ;
  assign n15387 = ~n15385 & n15386 ;
  assign n15388 = x50 &  n15387 ;
  assign n15389 = x50 | n15387 ;
  assign n15390 = ~n15388 & n15389 ;
  assign n15392 = ( n15180 & n15380 ) | ( n15180 & n15390 ) | ( n15380 & n15390 ) ;
  assign n15391 = ( n15380 & ~n15180 ) | ( n15380 & n15390 ) | ( ~n15180 & n15390 ) ;
  assign n15393 = ( n15180 & ~n15392 ) | ( n15180 & n15391 ) | ( ~n15392 & n15391 ) ;
  assign n15394 = ( n15313 & n15323 ) | ( n15313 & n15393 ) | ( n15323 & n15393 ) ;
  assign n15395 = ( n15323 & ~n15313 ) | ( n15323 & n15393 ) | ( ~n15313 & n15393 ) ;
  assign n15396 = ( n15313 & ~n15394 ) | ( n15313 & n15395 ) | ( ~n15394 & n15395 ) ;
  assign n15397 = ( n15197 & n15312 ) | ( n15197 & n15396 ) | ( n15312 & n15396 ) ;
  assign n15398 = ( n15312 & ~n15197 ) | ( n15312 & n15396 ) | ( ~n15197 & n15396 ) ;
  assign n15399 = ( n15197 & ~n15397 ) | ( n15197 & n15398 ) | ( ~n15397 & n15398 ) ;
  assign n15410 = ( n15200 & ~n15409 ) | ( n15200 & n15399 ) | ( ~n15409 & n15399 ) ;
  assign n15411 = ( n15200 & ~n15399 ) | ( n15200 & n15409 ) | ( ~n15399 & n15409 ) ;
  assign n15412 = ( n15410 & ~n15200 ) | ( n15410 & n15411 ) | ( ~n15200 & n15411 ) ;
  assign n15416 = x111 &  n3756 ;
  assign n15413 = ( x113 & ~n3602 ) | ( x113 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n15414 = x112 &  n3597 ;
  assign n15415 = n15413 | n15414 ;
  assign n15417 = ( x111 & ~n15416 ) | ( x111 & n15415 ) | ( ~n15416 & n15415 ) ;
  assign n15418 = n3605 | n6169 ;
  assign n15419 = ~n15417 & n15418 ;
  assign n15420 = x38 &  n15419 ;
  assign n15421 = x38 | n15419 ;
  assign n15422 = ~n15420 & n15421 ;
  assign n15423 = ( n15203 & n15412 ) | ( n15203 & n15422 ) | ( n15412 & n15422 ) ;
  assign n15424 = ( n15412 & ~n15203 ) | ( n15412 & n15422 ) | ( ~n15203 & n15422 ) ;
  assign n15425 = ( n15203 & ~n15423 ) | ( n15203 & n15424 ) | ( ~n15423 & n15424 ) ;
  assign n15429 = x114 &  n3214 ;
  assign n15426 = ( x116 & ~n3087 ) | ( x116 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n15427 = x115 &  n3082 ;
  assign n15428 = n15426 | n15427 ;
  assign n15430 = ( x114 & ~n15429 ) | ( x114 & n15428 ) | ( ~n15429 & n15428 ) ;
  assign n15431 = n3090 | n6885 ;
  assign n15432 = ~n15430 & n15431 ;
  assign n15433 = x35 &  n15432 ;
  assign n15434 = x35 | n15432 ;
  assign n15435 = ~n15433 & n15434 ;
  assign n15437 = ( n15207 & n15425 ) | ( n15207 & n15435 ) | ( n15425 & n15435 ) ;
  assign n15436 = ( n15425 & ~n15207 ) | ( n15425 & n15435 ) | ( ~n15207 & n15435 ) ;
  assign n15438 = ( n15207 & ~n15437 ) | ( n15207 & n15436 ) | ( ~n15437 & n15436 ) ;
  assign n15279 = ( n15209 & ~n15042 ) | ( n15209 & n15219 ) | ( ~n15042 & n15219 ) ;
  assign n15283 = x117 &  n2718 ;
  assign n15280 = ( x119 & ~n2642 ) | ( x119 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n15281 = x118 &  n2637 ;
  assign n15282 = n15280 | n15281 ;
  assign n15284 = ( x117 & ~n15283 ) | ( x117 & n15282 ) | ( ~n15283 & n15282 ) ;
  assign n15285 = ~n2645 & n7648 ;
  assign n15286 = n15284 | n15285 ;
  assign n15287 = ( x32 & n15279 ) | ( x32 & n15286 ) | ( n15279 & n15286 ) ;
  assign n15288 = ( x32 & ~n15279 ) | ( x32 & n15286 ) | ( ~n15279 & n15286 ) ;
  assign n15289 = ( n15279 & ~n15287 ) | ( n15279 & n15288 ) | ( ~n15287 & n15288 ) ;
  assign n15290 = ( x32 & ~n15080 ) | ( x32 & 1'b0 ) | ( ~n15080 & 1'b0 ) ;
  assign n15291 = n15223 | n15290 ;
  assign n15292 = ( n15081 & n15222 ) | ( n15081 & n15291 ) | ( n15222 & n15291 ) ;
  assign n15439 = ~n15289 & n15292 ;
  assign n15440 = n15289 | n15292 ;
  assign n15441 = ( n15439 & ~n15292 ) | ( n15439 & n15440 ) | ( ~n15292 & n15440 ) ;
  assign n15442 = ( n15302 & ~n15438 ) | ( n15302 & n15441 ) | ( ~n15438 & n15441 ) ;
  assign n15443 = ( n15438 & ~n15302 ) | ( n15438 & n15441 ) | ( ~n15302 & n15441 ) ;
  assign n15444 = ( n15442 & ~n15441 ) | ( n15442 & n15443 ) | ( ~n15441 & n15443 ) ;
  assign n15445 = n15278 &  n15444 ;
  assign n15446 = n15278 | n15444 ;
  assign n15447 = ~n15445 & n15446 ;
  assign n15448 = ( x126 & ~n1551 ) | ( x126 & 1'b0 ) | ( ~n1551 & 1'b0 ) ;
  assign n15449 = x127 &  n1446 ;
  assign n15450 = n15448 | n15449 ;
  assign n15451 = n1454 | n9960 ;
  assign n15452 = ( n15450 & ~n1454 ) | ( n15450 & n15451 ) | ( ~n1454 & n15451 ) ;
  assign n15453 = x23 | n15452 ;
  assign n15454 = ( x23 & ~n15452 ) | ( x23 & 1'b0 ) | ( ~n15452 & 1'b0 ) ;
  assign n15455 = ( n15453 & ~x23 ) | ( n15453 & n15454 ) | ( ~x23 & n15454 ) ;
  assign n15456 = ( n15267 & ~n15447 ) | ( n15267 & n15455 ) | ( ~n15447 & n15455 ) ;
  assign n15457 = ( n15267 & ~n15455 ) | ( n15267 & n15447 ) | ( ~n15455 & n15447 ) ;
  assign n15458 = ( n15456 & ~n15267 ) | ( n15456 & n15457 ) | ( ~n15267 & n15457 ) ;
  assign n15459 = ( n15063 & ~n15061 ) | ( n15063 & n15260 ) | ( ~n15061 & n15260 ) ;
  assign n15460 = ( n15264 & n15458 ) | ( n15264 & n15459 ) | ( n15458 & n15459 ) ;
  assign n15461 = ( n15458 & ~n15264 ) | ( n15458 & n15459 ) | ( ~n15264 & n15459 ) ;
  assign n15462 = ( n15264 & ~n15460 ) | ( n15264 & n15461 ) | ( ~n15460 & n15461 ) ;
  assign n15463 = ( n15267 & n15447 ) | ( n15267 & n15455 ) | ( n15447 & n15455 ) ;
  assign n15464 = ( n15264 & ~n15458 ) | ( n15264 & n15459 ) | ( ~n15458 & n15459 ) ;
  assign n15465 = ( x127 & ~n1551 ) | ( x127 & 1'b0 ) | ( ~n1551 & 1'b0 ) ;
  assign n15466 = n1454 | n10258 ;
  assign n15467 = ~n15465 & n15466 ;
  assign n15468 = ~x23 & n15467 ;
  assign n15469 = ( x23 & ~n15467 ) | ( x23 & 1'b0 ) | ( ~n15467 & 1'b0 ) ;
  assign n15470 = n15468 | n15469 ;
  assign n15471 = x26 &  n15274 ;
  assign n15472 = ( n15276 & ~n15471 ) | ( n15276 & n15445 ) | ( ~n15471 & n15445 ) ;
  assign n15473 = n15289 &  n15438 ;
  assign n15474 = n15289 | n15438 ;
  assign n15475 = ~n15473 & n15474 ;
  assign n15476 = ( n15292 & ~n15302 ) | ( n15292 & n15475 ) | ( ~n15302 & n15475 ) ;
  assign n15480 = x124 &  n1894 ;
  assign n15477 = ( x126 & ~n1816 ) | ( x126 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n15478 = x125 &  n1811 ;
  assign n15479 = n15477 | n15478 ;
  assign n15481 = ( x124 & ~n15480 ) | ( x124 & n15479 ) | ( ~n15480 & n15479 ) ;
  assign n15482 = n1819 | n9349 ;
  assign n15483 = ~n15481 & n15482 ;
  assign n15484 = x26 &  n15483 ;
  assign n15485 = x26 | n15483 ;
  assign n15486 = ~n15484 & n15485 ;
  assign n15488 = x32 &  n15286 ;
  assign n15487 = ~x32 & n15286 ;
  assign n15489 = ( x32 & ~n15488 ) | ( x32 & n15487 ) | ( ~n15488 & n15487 ) ;
  assign n15490 = ( n15279 & ~n15438 ) | ( n15279 & n15489 ) | ( ~n15438 & n15489 ) ;
  assign n15494 = x121 &  n2312 ;
  assign n15491 = ( x123 & ~n2195 ) | ( x123 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n15492 = x122 &  n2190 ;
  assign n15493 = n15491 | n15492 ;
  assign n15495 = ( x121 & ~n15494 ) | ( x121 & n15493 ) | ( ~n15494 & n15493 ) ;
  assign n15496 = ~n2198 & n8472 ;
  assign n15497 = n15495 | n15496 ;
  assign n15498 = ( x29 & ~n15497 ) | ( x29 & 1'b0 ) | ( ~n15497 & 1'b0 ) ;
  assign n15499 = ~x29 & n15497 ;
  assign n15500 = n15498 | n15499 ;
  assign n15501 = ( n15207 & ~n15435 ) | ( n15207 & n15425 ) | ( ~n15435 & n15425 ) ;
  assign n15505 = x118 &  n2718 ;
  assign n15502 = ( x120 & ~n2642 ) | ( x120 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n15503 = x119 &  n2637 ;
  assign n15504 = n15502 | n15503 ;
  assign n15506 = ( x118 & ~n15505 ) | ( x118 & n15504 ) | ( ~n15505 & n15504 ) ;
  assign n15507 = ~n2645 & n9364 ;
  assign n15508 = n15506 | n15507 ;
  assign n15509 = ( x32 & ~n15508 ) | ( x32 & 1'b0 ) | ( ~n15508 & 1'b0 ) ;
  assign n15510 = ~x32 & n15508 ;
  assign n15511 = n15509 | n15510 ;
  assign n15512 = ( n15203 & ~n15412 ) | ( n15203 & n15422 ) | ( ~n15412 & n15422 ) ;
  assign n15516 = x115 &  n3214 ;
  assign n15513 = ( x117 & ~n3087 ) | ( x117 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n15514 = x116 &  n3082 ;
  assign n15515 = n15513 | n15514 ;
  assign n15517 = ( x115 & ~n15516 ) | ( x115 & n15515 ) | ( ~n15516 & n15515 ) ;
  assign n15518 = n3090 | n7136 ;
  assign n15519 = ~n15517 & n15518 ;
  assign n15520 = x35 &  n15519 ;
  assign n15521 = x35 | n15519 ;
  assign n15522 = ~n15520 & n15521 ;
  assign n15523 = ( n15399 & ~n15200 ) | ( n15399 & n15409 ) | ( ~n15200 & n15409 ) ;
  assign n15527 = x106 &  n4934 ;
  assign n15524 = ( x108 & ~n4725 ) | ( x108 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n15525 = x107 &  n4720 ;
  assign n15526 = n15524 | n15525 ;
  assign n15528 = ( x106 & ~n15527 ) | ( x106 & n15526 ) | ( ~n15527 & n15526 ) ;
  assign n15529 = n4728 | n5055 ;
  assign n15530 = ~n15528 & n15529 ;
  assign n15531 = x44 &  n15530 ;
  assign n15532 = x44 | n15530 ;
  assign n15533 = ~n15531 & n15532 ;
  assign n15534 = ( n15180 & ~n15390 ) | ( n15180 & n15380 ) | ( ~n15390 & n15380 ) ;
  assign n15535 = ( n15354 & ~n15353 ) | ( n15354 & n15364 ) | ( ~n15353 & n15364 ) ;
  assign n15539 = x97 &  n6982 ;
  assign n15536 = ( x99 & ~n6727 ) | ( x99 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n15537 = x98 &  n6722 ;
  assign n15538 = n15536 | n15537 ;
  assign n15540 = ( x97 & ~n15539 ) | ( x97 & n15538 ) | ( ~n15539 & n15538 ) ;
  assign n15541 = ( n3338 & ~n6730 ) | ( n3338 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n15542 = n15540 | n15541 ;
  assign n15543 = ( x53 & ~n15542 ) | ( x53 & 1'b0 ) | ( ~n15542 & 1'b0 ) ;
  assign n15544 = ~x53 & n15542 ;
  assign n15545 = n15543 | n15544 ;
  assign n15546 = x86 &  n10104 ;
  assign n15547 = ( x87 & ~n9760 ) | ( x87 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n15548 = n15546 | n15547 ;
  assign n15552 = x88 &  n9457 ;
  assign n15549 = ( x90 & ~n9150 ) | ( x90 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n15550 = x89 &  n9145 ;
  assign n15551 = n15549 | n15550 ;
  assign n15553 = ( x88 & ~n15552 ) | ( x88 & n15551 ) | ( ~n15552 & n15551 ) ;
  assign n15554 = ( n1976 & ~n15553 ) | ( n1976 & n9153 ) | ( ~n15553 & n9153 ) ;
  assign n15555 = ~n9153 & n15554 ;
  assign n15556 = ( x62 & n15553 ) | ( x62 & n15555 ) | ( n15553 & n15555 ) ;
  assign n15557 = ( x62 & ~n15555 ) | ( x62 & n15553 ) | ( ~n15555 & n15553 ) ;
  assign n15558 = ( n15555 & ~n15556 ) | ( n15555 & n15557 ) | ( ~n15556 & n15557 ) ;
  assign n15559 = ( n15548 & ~n15347 ) | ( n15548 & n15558 ) | ( ~n15347 & n15558 ) ;
  assign n15560 = ( n15347 & ~n15558 ) | ( n15347 & n15548 ) | ( ~n15558 & n15548 ) ;
  assign n15561 = ( n15559 & ~n15548 ) | ( n15559 & n15560 ) | ( ~n15548 & n15560 ) ;
  assign n15562 = ( n15334 & ~n15347 ) | ( n15334 & n15344 ) | ( ~n15347 & n15344 ) ;
  assign n15566 = x91 &  n8558 ;
  assign n15563 = ( x93 & ~n8314 ) | ( x93 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n15564 = x92 &  n8309 ;
  assign n15565 = n15563 | n15564 ;
  assign n15567 = ( x91 & ~n15566 ) | ( x91 & n15565 ) | ( ~n15566 & n15565 ) ;
  assign n15568 = n2264 | n8317 ;
  assign n15569 = ~n15567 & n15568 ;
  assign n15570 = x59 &  n15569 ;
  assign n15571 = x59 | n15569 ;
  assign n15572 = ~n15570 & n15571 ;
  assign n15574 = ( n15561 & n15562 ) | ( n15561 & n15572 ) | ( n15562 & n15572 ) ;
  assign n15573 = ( n15562 & ~n15561 ) | ( n15562 & n15572 ) | ( ~n15561 & n15572 ) ;
  assign n15575 = ( n15561 & ~n15574 ) | ( n15561 & n15573 ) | ( ~n15574 & n15573 ) ;
  assign n15579 = x94 &  n7731 ;
  assign n15576 = ( x96 & ~n7538 ) | ( x96 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n15577 = x95 &  n7533 ;
  assign n15578 = n15576 | n15577 ;
  assign n15580 = ( x94 & ~n15579 ) | ( x94 & n15578 ) | ( ~n15579 & n15578 ) ;
  assign n15581 = ( n2836 & ~n7541 ) | ( n2836 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n15582 = n15580 | n15581 ;
  assign n15583 = ( x56 & ~n15582 ) | ( x56 & 1'b0 ) | ( ~n15582 & 1'b0 ) ;
  assign n15584 = ~x56 & n15582 ;
  assign n15585 = n15583 | n15584 ;
  assign n15586 = ( n15352 & ~n15575 ) | ( n15352 & n15585 ) | ( ~n15575 & n15585 ) ;
  assign n15587 = ( n15352 & ~n15585 ) | ( n15352 & n15575 ) | ( ~n15585 & n15575 ) ;
  assign n15588 = ( n15586 & ~n15352 ) | ( n15586 & n15587 ) | ( ~n15352 & n15587 ) ;
  assign n15590 = ( n15535 & n15545 ) | ( n15535 & n15588 ) | ( n15545 & n15588 ) ;
  assign n15589 = ( n15545 & ~n15535 ) | ( n15545 & n15588 ) | ( ~n15535 & n15588 ) ;
  assign n15591 = ( n15535 & ~n15590 ) | ( n15535 & n15589 ) | ( ~n15590 & n15589 ) ;
  assign n15592 = ( n15176 & ~n15377 ) | ( n15176 & n15367 ) | ( ~n15377 & n15367 ) ;
  assign n15596 = x100 &  n6288 ;
  assign n15593 = ( x102 & ~n6032 ) | ( x102 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n15594 = x101 &  n6027 ;
  assign n15595 = n15593 | n15594 ;
  assign n15597 = ( x100 & ~n15596 ) | ( x100 & n15595 ) | ( ~n15596 & n15595 ) ;
  assign n15598 = n3872 | n6035 ;
  assign n15599 = ~n15597 & n15598 ;
  assign n15600 = x50 &  n15599 ;
  assign n15601 = x50 | n15599 ;
  assign n15602 = ~n15600 & n15601 ;
  assign n15603 = ( n15591 & ~n15592 ) | ( n15591 & n15602 ) | ( ~n15592 & n15602 ) ;
  assign n15604 = ( n15591 & ~n15602 ) | ( n15591 & n15592 ) | ( ~n15602 & n15592 ) ;
  assign n15605 = ( n15603 & ~n15591 ) | ( n15603 & n15604 ) | ( ~n15591 & n15604 ) ;
  assign n15609 = x103 &  n5586 ;
  assign n15606 = ( x105 & ~n5389 ) | ( x105 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n15607 = x104 &  n5384 ;
  assign n15608 = n15606 | n15607 ;
  assign n15610 = ( x103 & ~n15609 ) | ( x103 & n15608 ) | ( ~n15609 & n15608 ) ;
  assign n15611 = ( n4442 & ~n5392 ) | ( n4442 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n15612 = n15610 | n15611 ;
  assign n15613 = ( x47 & ~n15612 ) | ( x47 & 1'b0 ) | ( ~n15612 & 1'b0 ) ;
  assign n15614 = ~x47 & n15612 ;
  assign n15615 = n15613 | n15614 ;
  assign n15616 = ( n15534 & ~n15605 ) | ( n15534 & n15615 ) | ( ~n15605 & n15615 ) ;
  assign n15617 = ( n15534 & ~n15615 ) | ( n15534 & n15605 ) | ( ~n15615 & n15605 ) ;
  assign n15618 = ( n15616 & ~n15534 ) | ( n15616 & n15617 ) | ( ~n15534 & n15617 ) ;
  assign n15620 = ( n15395 & n15533 ) | ( n15395 & n15618 ) | ( n15533 & n15618 ) ;
  assign n15619 = ( n15533 & ~n15395 ) | ( n15533 & n15618 ) | ( ~n15395 & n15618 ) ;
  assign n15621 = ( n15395 & ~n15620 ) | ( n15395 & n15619 ) | ( ~n15620 & n15619 ) ;
  assign n15625 = x109 &  n4344 ;
  assign n15622 = ( x111 & ~n4143 ) | ( x111 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n15623 = x110 &  n4138 ;
  assign n15624 = n15622 | n15623 ;
  assign n15626 = ( x109 & ~n15625 ) | ( x109 & n15624 ) | ( ~n15625 & n15624 ) ;
  assign n15627 = n4146 | n5711 ;
  assign n15628 = ~n15626 & n15627 ;
  assign n15629 = x41 &  n15628 ;
  assign n15630 = x41 | n15628 ;
  assign n15631 = ~n15629 & n15630 ;
  assign n15632 = ( n15398 & n15621 ) | ( n15398 & n15631 ) | ( n15621 & n15631 ) ;
  assign n15633 = ( n15398 & ~n15621 ) | ( n15398 & n15631 ) | ( ~n15621 & n15631 ) ;
  assign n15634 = ( n15621 & ~n15632 ) | ( n15621 & n15633 ) | ( ~n15632 & n15633 ) ;
  assign n15638 = x112 &  n3756 ;
  assign n15635 = ( x114 & ~n3602 ) | ( x114 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n15636 = x113 &  n3597 ;
  assign n15637 = n15635 | n15636 ;
  assign n15639 = ( x112 & ~n15638 ) | ( x112 & n15637 ) | ( ~n15638 & n15637 ) ;
  assign n15640 = n3605 | n6185 ;
  assign n15641 = ~n15639 & n15640 ;
  assign n15642 = x38 &  n15641 ;
  assign n15643 = x38 | n15641 ;
  assign n15644 = ~n15642 & n15643 ;
  assign n15645 = ( n15523 & ~n15634 ) | ( n15523 & n15644 ) | ( ~n15634 & n15644 ) ;
  assign n15646 = ( n15523 & ~n15644 ) | ( n15523 & n15634 ) | ( ~n15644 & n15634 ) ;
  assign n15647 = ( n15645 & ~n15523 ) | ( n15645 & n15646 ) | ( ~n15523 & n15646 ) ;
  assign n15649 = ( n15512 & n15522 ) | ( n15512 & n15647 ) | ( n15522 & n15647 ) ;
  assign n15648 = ( n15522 & ~n15512 ) | ( n15522 & n15647 ) | ( ~n15512 & n15647 ) ;
  assign n15650 = ( n15512 & ~n15649 ) | ( n15512 & n15648 ) | ( ~n15649 & n15648 ) ;
  assign n15652 = ( n15501 & n15511 ) | ( n15501 & n15650 ) | ( n15511 & n15650 ) ;
  assign n15651 = ( n15511 & ~n15501 ) | ( n15511 & n15650 ) | ( ~n15501 & n15650 ) ;
  assign n15653 = ( n15501 & ~n15652 ) | ( n15501 & n15651 ) | ( ~n15652 & n15651 ) ;
  assign n15655 = ( n15490 & n15500 ) | ( n15490 & n15653 ) | ( n15500 & n15653 ) ;
  assign n15654 = ( n15500 & ~n15490 ) | ( n15500 & n15653 ) | ( ~n15490 & n15653 ) ;
  assign n15656 = ( n15490 & ~n15655 ) | ( n15490 & n15654 ) | ( ~n15655 & n15654 ) ;
  assign n15657 = ( n15476 & ~n15486 ) | ( n15476 & n15656 ) | ( ~n15486 & n15656 ) ;
  assign n15658 = ( n15476 & ~n15656 ) | ( n15476 & n15486 ) | ( ~n15656 & n15486 ) ;
  assign n15659 = ( n15657 & ~n15476 ) | ( n15657 & n15658 ) | ( ~n15476 & n15658 ) ;
  assign n15660 = ( n15470 & n15472 ) | ( n15470 & n15659 ) | ( n15472 & n15659 ) ;
  assign n15661 = ( n15472 & ~n15470 ) | ( n15472 & n15659 ) | ( ~n15470 & n15659 ) ;
  assign n15662 = ( n15470 & ~n15660 ) | ( n15470 & n15661 ) | ( ~n15660 & n15661 ) ;
  assign n15663 = ( n15463 & n15464 ) | ( n15463 & n15662 ) | ( n15464 & n15662 ) ;
  assign n15664 = ( n15464 & ~n15463 ) | ( n15464 & n15662 ) | ( ~n15463 & n15662 ) ;
  assign n15665 = ( n15463 & ~n15663 ) | ( n15463 & n15664 ) | ( ~n15663 & n15664 ) ;
  assign n15666 = ( n15470 & ~n15472 ) | ( n15470 & n15659 ) | ( ~n15472 & n15659 ) ;
  assign n15667 = ( n15463 & ~n15464 ) | ( n15463 & n15662 ) | ( ~n15464 & n15662 ) ;
  assign n15671 = x125 &  n1894 ;
  assign n15668 = ( x127 & ~n1816 ) | ( x127 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n15669 = x126 &  n1811 ;
  assign n15670 = n15668 | n15669 ;
  assign n15672 = ( x125 & ~n15671 ) | ( x125 & n15670 ) | ( ~n15671 & n15670 ) ;
  assign n15673 = n1819 | n9941 ;
  assign n15674 = ~n15672 & n15673 ;
  assign n15675 = x26 &  n15674 ;
  assign n15676 = x26 | n15674 ;
  assign n15677 = ~n15675 & n15676 ;
  assign n15678 = ( n15476 & n15486 ) | ( n15476 & n15656 ) | ( n15486 & n15656 ) ;
  assign n15679 = ( n15490 & ~n15653 ) | ( n15490 & n15500 ) | ( ~n15653 & n15500 ) ;
  assign n15687 = ( n15501 & ~n15650 ) | ( n15501 & n15511 ) | ( ~n15650 & n15511 ) ;
  assign n15691 = x110 &  n4344 ;
  assign n15688 = ( x112 & ~n4143 ) | ( x112 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n15689 = x111 &  n4138 ;
  assign n15690 = n15688 | n15689 ;
  assign n15692 = ( x110 & ~n15691 ) | ( x110 & n15690 ) | ( ~n15691 & n15690 ) ;
  assign n15693 = ~n4146 & n5727 ;
  assign n15694 = n15692 | n15693 ;
  assign n15695 = ( x41 & ~n15694 ) | ( x41 & 1'b0 ) | ( ~n15694 & 1'b0 ) ;
  assign n15696 = ~x41 & n15694 ;
  assign n15697 = n15695 | n15696 ;
  assign n15701 = x101 &  n6288 ;
  assign n15698 = ( x103 & ~n6032 ) | ( x103 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n15699 = x102 &  n6027 ;
  assign n15700 = n15698 | n15699 ;
  assign n15702 = ( x101 & ~n15701 ) | ( x101 & n15700 ) | ( ~n15701 & n15700 ) ;
  assign n15703 = n4056 | n6035 ;
  assign n15704 = ~n15702 & n15703 ;
  assign n15705 = x50 &  n15704 ;
  assign n15706 = x50 | n15704 ;
  assign n15707 = ~n15705 & n15706 ;
  assign n15711 = x95 &  n7731 ;
  assign n15708 = ( x97 & ~n7538 ) | ( x97 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n15709 = x96 &  n7533 ;
  assign n15710 = n15708 | n15709 ;
  assign n15712 = ( x95 & ~n15711 ) | ( x95 & n15710 ) | ( ~n15711 & n15710 ) ;
  assign n15713 = ( n2999 & ~n7541 ) | ( n2999 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n15714 = n15712 | n15713 ;
  assign n15715 = ( x56 & ~n15714 ) | ( x56 & 1'b0 ) | ( ~n15714 & 1'b0 ) ;
  assign n15716 = ~x56 & n15714 ;
  assign n15717 = n15715 | n15716 ;
  assign n15718 = x87 &  n10104 ;
  assign n15719 = ( x88 & ~n9760 ) | ( x88 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n15720 = n15718 | n15719 ;
  assign n15721 = ( x23 & n15548 ) | ( x23 & n15720 ) | ( n15548 & n15720 ) ;
  assign n15722 = ( x23 & ~n15548 ) | ( x23 & n15720 ) | ( ~n15548 & n15720 ) ;
  assign n15723 = ( n15548 & ~n15721 ) | ( n15548 & n15722 ) | ( ~n15721 & n15722 ) ;
  assign n15724 = ( n15347 & ~n15548 ) | ( n15347 & n15558 ) | ( ~n15548 & n15558 ) ;
  assign n15728 = x89 &  n9457 ;
  assign n15725 = ( x91 & ~n9150 ) | ( x91 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n15726 = x90 &  n9145 ;
  assign n15727 = n15725 | n15726 ;
  assign n15729 = ( x89 & ~n15728 ) | ( x89 & n15727 ) | ( ~n15728 & n15727 ) ;
  assign n15730 = ( n2108 & ~n9153 ) | ( n2108 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n15731 = n15729 | n15730 ;
  assign n15732 = ( x62 & ~n15731 ) | ( x62 & 1'b0 ) | ( ~n15731 & 1'b0 ) ;
  assign n15733 = ~x62 & n15731 ;
  assign n15734 = n15732 | n15733 ;
  assign n15735 = ( n15723 & ~n15724 ) | ( n15723 & n15734 ) | ( ~n15724 & n15734 ) ;
  assign n15736 = ( n15723 & ~n15734 ) | ( n15723 & n15724 ) | ( ~n15734 & n15724 ) ;
  assign n15737 = ( n15735 & ~n15723 ) | ( n15735 & n15736 ) | ( ~n15723 & n15736 ) ;
  assign n15738 = ( n15561 & ~n15562 ) | ( n15561 & n15572 ) | ( ~n15562 & n15572 ) ;
  assign n15742 = x92 &  n8558 ;
  assign n15739 = ( x94 & ~n8314 ) | ( x94 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n15740 = x93 &  n8309 ;
  assign n15741 = n15739 | n15740 ;
  assign n15743 = ( x92 & ~n15742 ) | ( x92 & n15741 ) | ( ~n15742 & n15741 ) ;
  assign n15744 = ( n2401 & ~n8317 ) | ( n2401 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n15745 = n15743 | n15744 ;
  assign n15746 = ( x59 & ~n15745 ) | ( x59 & 1'b0 ) | ( ~n15745 & 1'b0 ) ;
  assign n15747 = ~x59 & n15745 ;
  assign n15748 = n15746 | n15747 ;
  assign n15750 = ( n15737 & n15738 ) | ( n15737 & n15748 ) | ( n15738 & n15748 ) ;
  assign n15749 = ( n15738 & ~n15737 ) | ( n15738 & n15748 ) | ( ~n15737 & n15748 ) ;
  assign n15751 = ( n15737 & ~n15750 ) | ( n15737 & n15749 ) | ( ~n15750 & n15749 ) ;
  assign n15752 = ( n15352 & n15575 ) | ( n15352 & n15585 ) | ( n15575 & n15585 ) ;
  assign n15753 = ( n15717 & n15751 ) | ( n15717 & n15752 ) | ( n15751 & n15752 ) ;
  assign n15754 = ( n15751 & ~n15717 ) | ( n15751 & n15752 ) | ( ~n15717 & n15752 ) ;
  assign n15755 = ( n15717 & ~n15753 ) | ( n15717 & n15754 ) | ( ~n15753 & n15754 ) ;
  assign n15759 = x98 &  n6982 ;
  assign n15756 = ( x100 & ~n6727 ) | ( x100 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n15757 = x99 &  n6722 ;
  assign n15758 = n15756 | n15757 ;
  assign n15760 = ( x98 & ~n15759 ) | ( x98 & n15758 ) | ( ~n15759 & n15758 ) ;
  assign n15761 = n3354 | n6730 ;
  assign n15762 = ~n15760 & n15761 ;
  assign n15763 = x53 &  n15762 ;
  assign n15764 = x53 | n15762 ;
  assign n15765 = ~n15763 & n15764 ;
  assign n15767 = ( n15590 & n15755 ) | ( n15590 & n15765 ) | ( n15755 & n15765 ) ;
  assign n15766 = ( n15590 & ~n15755 ) | ( n15590 & n15765 ) | ( ~n15755 & n15765 ) ;
  assign n15768 = ( n15755 & ~n15767 ) | ( n15755 & n15766 ) | ( ~n15767 & n15766 ) ;
  assign n15769 = ( n15592 & ~n15591 ) | ( n15592 & n15602 ) | ( ~n15591 & n15602 ) ;
  assign n15770 = ( n15707 & n15768 ) | ( n15707 & n15769 ) | ( n15768 & n15769 ) ;
  assign n15771 = ( n15768 & ~n15707 ) | ( n15768 & n15769 ) | ( ~n15707 & n15769 ) ;
  assign n15772 = ( n15707 & ~n15770 ) | ( n15707 & n15771 ) | ( ~n15770 & n15771 ) ;
  assign n15773 = ( n15534 & n15605 ) | ( n15534 & n15615 ) | ( n15605 & n15615 ) ;
  assign n15777 = x104 &  n5586 ;
  assign n15774 = ( x106 & ~n5389 ) | ( x106 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n15775 = x105 &  n5384 ;
  assign n15776 = n15774 | n15775 ;
  assign n15778 = ( x104 & ~n15777 ) | ( x104 & n15776 ) | ( ~n15777 & n15776 ) ;
  assign n15779 = ( n4458 & ~n5392 ) | ( n4458 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n15780 = n15778 | n15779 ;
  assign n15781 = ( x47 & ~n15780 ) | ( x47 & 1'b0 ) | ( ~n15780 & 1'b0 ) ;
  assign n15782 = ~x47 & n15780 ;
  assign n15783 = n15781 | n15782 ;
  assign n15784 = ( n15772 & ~n15773 ) | ( n15772 & n15783 ) | ( ~n15773 & n15783 ) ;
  assign n15785 = ( n15772 & ~n15783 ) | ( n15772 & n15773 ) | ( ~n15783 & n15773 ) ;
  assign n15786 = ( n15784 & ~n15772 ) | ( n15784 & n15785 ) | ( ~n15772 & n15785 ) ;
  assign n15787 = ( n15395 & ~n15618 ) | ( n15395 & n15533 ) | ( ~n15618 & n15533 ) ;
  assign n15791 = x107 &  n4934 ;
  assign n15788 = ( x109 & ~n4725 ) | ( x109 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n15789 = x108 &  n4720 ;
  assign n15790 = n15788 | n15789 ;
  assign n15792 = ( x107 & ~n15791 ) | ( x107 & n15790 ) | ( ~n15791 & n15790 ) ;
  assign n15793 = ~n4728 & n5267 ;
  assign n15794 = n15792 | n15793 ;
  assign n15795 = ( x44 & ~n15794 ) | ( x44 & 1'b0 ) | ( ~n15794 & 1'b0 ) ;
  assign n15796 = ~x44 & n15794 ;
  assign n15797 = n15795 | n15796 ;
  assign n15799 = ( n15786 & n15787 ) | ( n15786 & n15797 ) | ( n15787 & n15797 ) ;
  assign n15798 = ( n15787 & ~n15786 ) | ( n15787 & n15797 ) | ( ~n15786 & n15797 ) ;
  assign n15800 = ( n15786 & ~n15799 ) | ( n15786 & n15798 ) | ( ~n15799 & n15798 ) ;
  assign n15801 = ( n15398 & ~n15631 ) | ( n15398 & n15621 ) | ( ~n15631 & n15621 ) ;
  assign n15802 = ( n15697 & n15800 ) | ( n15697 & n15801 ) | ( n15800 & n15801 ) ;
  assign n15803 = ( n15800 & ~n15697 ) | ( n15800 & n15801 ) | ( ~n15697 & n15801 ) ;
  assign n15804 = ( n15697 & ~n15802 ) | ( n15697 & n15803 ) | ( ~n15802 & n15803 ) ;
  assign n15805 = ( n15523 & n15634 ) | ( n15523 & n15644 ) | ( n15634 & n15644 ) ;
  assign n15809 = x113 &  n3756 ;
  assign n15806 = ( x115 & ~n3602 ) | ( x115 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n15807 = x114 &  n3597 ;
  assign n15808 = n15806 | n15807 ;
  assign n15810 = ( x113 & ~n15809 ) | ( x113 & n15808 ) | ( ~n15809 & n15808 ) ;
  assign n15811 = ~n3605 & n6420 ;
  assign n15812 = n15810 | n15811 ;
  assign n15813 = ( x38 & ~n15812 ) | ( x38 & 1'b0 ) | ( ~n15812 & 1'b0 ) ;
  assign n15814 = ~x38 & n15812 ;
  assign n15815 = n15813 | n15814 ;
  assign n15817 = ( n15804 & n15805 ) | ( n15804 & n15815 ) | ( n15805 & n15815 ) ;
  assign n15816 = ( n15805 & ~n15804 ) | ( n15805 & n15815 ) | ( ~n15804 & n15815 ) ;
  assign n15818 = ( n15804 & ~n15817 ) | ( n15804 & n15816 ) | ( ~n15817 & n15816 ) ;
  assign n15822 = x116 &  n3214 ;
  assign n15819 = ( x118 & ~n3087 ) | ( x118 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n15820 = x117 &  n3082 ;
  assign n15821 = n15819 | n15820 ;
  assign n15823 = ( x116 & ~n15822 ) | ( x116 & n15821 ) | ( ~n15822 & n15821 ) ;
  assign n15824 = n3090 | n7152 ;
  assign n15825 = ~n15823 & n15824 ;
  assign n15826 = x35 &  n15825 ;
  assign n15827 = x35 | n15825 ;
  assign n15828 = ~n15826 & n15827 ;
  assign n15829 = ( n15818 & ~n15649 ) | ( n15818 & n15828 ) | ( ~n15649 & n15828 ) ;
  assign n15830 = ( n15649 & ~n15828 ) | ( n15649 & n15818 ) | ( ~n15828 & n15818 ) ;
  assign n15831 = ( n15829 & ~n15818 ) | ( n15829 & n15830 ) | ( ~n15818 & n15830 ) ;
  assign n15683 = x119 &  n2718 ;
  assign n15680 = ( x121 & ~n2642 ) | ( x121 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n15681 = x120 &  n2637 ;
  assign n15682 = n15680 | n15681 ;
  assign n15684 = ( x119 & ~n15683 ) | ( x119 & n15682 ) | ( ~n15683 & n15682 ) ;
  assign n15685 = ~n2645 & n8176 ;
  assign n15686 = n15684 | n15685 ;
  assign n15832 = x32 | n15686 ;
  assign n15833 = ~x32 & n15686 ;
  assign n15834 = ( n15832 & ~n15686 ) | ( n15832 & n15833 ) | ( ~n15686 & n15833 ) ;
  assign n15835 = ( n15687 & ~n15831 ) | ( n15687 & n15834 ) | ( ~n15831 & n15834 ) ;
  assign n15836 = ( n15831 & ~n15687 ) | ( n15831 & n15834 ) | ( ~n15687 & n15834 ) ;
  assign n15837 = ( n15835 & ~n15834 ) | ( n15835 & n15836 ) | ( ~n15834 & n15836 ) ;
  assign n15841 = x122 &  n2312 ;
  assign n15838 = ( x124 & ~n2195 ) | ( x124 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n15839 = x123 &  n2190 ;
  assign n15840 = n15838 | n15839 ;
  assign n15842 = ( x122 & ~n15841 ) | ( x122 & n15840 ) | ( ~n15841 & n15840 ) ;
  assign n15843 = ~n2198 & n8755 ;
  assign n15844 = n15842 | n15843 ;
  assign n15845 = ( x29 & ~n15844 ) | ( x29 & 1'b0 ) | ( ~n15844 & 1'b0 ) ;
  assign n15846 = ~x29 & n15844 ;
  assign n15847 = n15845 | n15846 ;
  assign n15848 = ( n15679 & n15837 ) | ( n15679 & n15847 ) | ( n15837 & n15847 ) ;
  assign n15849 = ( n15837 & ~n15679 ) | ( n15837 & n15847 ) | ( ~n15679 & n15847 ) ;
  assign n15850 = ( n15679 & ~n15848 ) | ( n15679 & n15849 ) | ( ~n15848 & n15849 ) ;
  assign n15851 = ( n15677 & ~n15678 ) | ( n15677 & n15850 ) | ( ~n15678 & n15850 ) ;
  assign n15852 = ( n15677 & ~n15850 ) | ( n15677 & n15678 ) | ( ~n15850 & n15678 ) ;
  assign n15853 = ( n15851 & ~n15677 ) | ( n15851 & n15852 ) | ( ~n15677 & n15852 ) ;
  assign n15854 = ( n15666 & n15667 ) | ( n15666 & n15853 ) | ( n15667 & n15853 ) ;
  assign n15855 = ( n15667 & ~n15666 ) | ( n15667 & n15853 ) | ( ~n15666 & n15853 ) ;
  assign n15856 = ( n15666 & ~n15854 ) | ( n15666 & n15855 ) | ( ~n15854 & n15855 ) ;
  assign n15857 = ( n15677 & n15678 ) | ( n15677 & n15850 ) | ( n15678 & n15850 ) ;
  assign n15858 = ( n15666 & ~n15667 ) | ( n15666 & n15853 ) | ( ~n15667 & n15853 ) ;
  assign n15859 = ( n15679 & ~n15837 ) | ( n15679 & n15847 ) | ( ~n15837 & n15847 ) ;
  assign n15860 = ( x32 & ~n15686 ) | ( x32 & 1'b0 ) | ( ~n15686 & 1'b0 ) ;
  assign n15861 = n15833 | n15860 ;
  assign n15862 = ( n15687 & ~n15831 ) | ( n15687 & n15861 ) | ( ~n15831 & n15861 ) ;
  assign n15866 = x123 &  n2312 ;
  assign n15863 = ( x125 & ~n2195 ) | ( x125 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n15864 = x124 &  n2190 ;
  assign n15865 = n15863 | n15864 ;
  assign n15867 = ( x123 & ~n15866 ) | ( x123 & n15865 ) | ( ~n15866 & n15865 ) ;
  assign n15868 = ~n2198 & n9324 ;
  assign n15869 = n15867 | n15868 ;
  assign n15871 = x29 &  n15869 ;
  assign n15870 = ~x29 & n15869 ;
  assign n15872 = ( x29 & ~n15871 ) | ( x29 & n15870 ) | ( ~n15871 & n15870 ) ;
  assign n15876 = x120 &  n2718 ;
  assign n15873 = ( x122 & ~n2642 ) | ( x122 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n15874 = x121 &  n2637 ;
  assign n15875 = n15873 | n15874 ;
  assign n15877 = ( x120 & ~n15876 ) | ( x120 & n15875 ) | ( ~n15876 & n15875 ) ;
  assign n15878 = ( n2645 & n9987 ) | ( n2645 & n15877 ) | ( n9987 & n15877 ) ;
  assign n15879 = ( n9987 & ~n15878 ) | ( n9987 & 1'b0 ) | ( ~n15878 & 1'b0 ) ;
  assign n15880 = ( x32 & n15877 ) | ( x32 & n15879 ) | ( n15877 & n15879 ) ;
  assign n15881 = ( x32 & ~n15879 ) | ( x32 & n15877 ) | ( ~n15879 & n15877 ) ;
  assign n15882 = ( n15879 & ~n15880 ) | ( n15879 & n15881 ) | ( ~n15880 & n15881 ) ;
  assign n15883 = ( n15649 & n15818 ) | ( n15649 & n15828 ) | ( n15818 & n15828 ) ;
  assign n15884 = ( n15786 & ~n15797 ) | ( n15786 & n15787 ) | ( ~n15797 & n15787 ) ;
  assign n15885 = ( n15773 & ~n15772 ) | ( n15773 & n15783 ) | ( ~n15772 & n15783 ) ;
  assign n15974 = x108 &  n4934 ;
  assign n15971 = ( x110 & ~n4725 ) | ( x110 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n15972 = x109 &  n4720 ;
  assign n15973 = n15971 | n15972 ;
  assign n15975 = ( x108 & ~n15974 ) | ( x108 & n15973 ) | ( ~n15974 & n15973 ) ;
  assign n15976 = n4728 | n5283 ;
  assign n15977 = ~n15975 & n15976 ;
  assign n15978 = x44 &  n15977 ;
  assign n15979 = x44 | n15977 ;
  assign n15980 = ~n15978 & n15979 ;
  assign n15889 = x105 &  n5586 ;
  assign n15886 = ( x107 & ~n5389 ) | ( x107 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n15887 = x106 &  n5384 ;
  assign n15888 = n15886 | n15887 ;
  assign n15890 = ( x105 & ~n15889 ) | ( x105 & n15888 ) | ( ~n15889 & n15888 ) ;
  assign n15891 = ( n4848 & ~n5392 ) | ( n4848 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n15892 = n15890 | n15891 ;
  assign n15893 = ( x47 & ~n15892 ) | ( x47 & 1'b0 ) | ( ~n15892 & 1'b0 ) ;
  assign n15894 = ~x47 & n15892 ;
  assign n15895 = n15893 | n15894 ;
  assign n15896 = ( n15590 & ~n15765 ) | ( n15590 & n15755 ) | ( ~n15765 & n15755 ) ;
  assign n15900 = x102 &  n6288 ;
  assign n15897 = ( x104 & ~n6032 ) | ( x104 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n15898 = x103 &  n6027 ;
  assign n15899 = n15897 | n15898 ;
  assign n15901 = ( x102 & ~n15900 ) | ( x102 & n15899 ) | ( ~n15900 & n15899 ) ;
  assign n15902 = n4249 | n6035 ;
  assign n15903 = ~n15901 & n15902 ;
  assign n15904 = x50 &  n15903 ;
  assign n15905 = x50 | n15903 ;
  assign n15906 = ~n15904 & n15905 ;
  assign n15907 = ( n15737 & ~n15748 ) | ( n15737 & n15738 ) | ( ~n15748 & n15738 ) ;
  assign n15929 = x93 &  n8558 ;
  assign n15926 = ( x95 & ~n8314 ) | ( x95 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n15927 = x94 &  n8309 ;
  assign n15928 = n15926 | n15927 ;
  assign n15930 = ( x93 & ~n15929 ) | ( x93 & n15928 ) | ( ~n15929 & n15928 ) ;
  assign n15931 = ( n2547 & ~n8317 ) | ( n2547 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n15932 = n15930 | n15931 ;
  assign n15909 = ( n15548 & ~x23 ) | ( n15548 & n15720 ) | ( ~x23 & n15720 ) ;
  assign n15910 = x88 &  n10104 ;
  assign n15911 = ( x89 & ~n9760 ) | ( x89 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n15912 = n15910 | n15911 ;
  assign n15916 = x90 &  n9457 ;
  assign n15913 = ( x92 & ~n9150 ) | ( x92 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n15914 = x91 &  n9145 ;
  assign n15915 = n15913 | n15914 ;
  assign n15917 = ( x90 & ~n15916 ) | ( x90 & n15915 ) | ( ~n15916 & n15915 ) ;
  assign n15918 = ( n2248 & ~n15917 ) | ( n2248 & n9153 ) | ( ~n15917 & n9153 ) ;
  assign n15919 = ~n9153 & n15918 ;
  assign n15920 = ( x62 & n15917 ) | ( x62 & n15919 ) | ( n15917 & n15919 ) ;
  assign n15921 = ( x62 & ~n15919 ) | ( x62 & n15917 ) | ( ~n15919 & n15917 ) ;
  assign n15922 = ( n15919 & ~n15920 ) | ( n15919 & n15921 ) | ( ~n15920 & n15921 ) ;
  assign n15923 = ( n15909 & ~n15912 ) | ( n15909 & n15922 ) | ( ~n15912 & n15922 ) ;
  assign n15924 = ( n15909 & ~n15922 ) | ( n15909 & n15912 ) | ( ~n15922 & n15912 ) ;
  assign n15925 = ( n15923 & ~n15909 ) | ( n15923 & n15924 ) | ( ~n15909 & n15924 ) ;
  assign n15908 = ( n15724 & ~n15723 ) | ( n15724 & n15734 ) | ( ~n15723 & n15734 ) ;
  assign n15933 = ~x59 & n15908 ;
  assign n15934 = x59 | n15908 ;
  assign n15935 = ( n15933 & ~n15908 ) | ( n15933 & n15934 ) | ( ~n15908 & n15934 ) ;
  assign n15936 = ( n15932 & ~n15925 ) | ( n15932 & n15935 ) | ( ~n15925 & n15935 ) ;
  assign n15937 = ( n15925 & ~n15932 ) | ( n15925 & n15935 ) | ( ~n15932 & n15935 ) ;
  assign n15938 = ( n15936 & ~n15935 ) | ( n15936 & n15937 ) | ( ~n15935 & n15937 ) ;
  assign n15942 = x96 &  n7731 ;
  assign n15939 = ( x98 & ~n7538 ) | ( x98 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n15940 = x97 &  n7533 ;
  assign n15941 = n15939 | n15940 ;
  assign n15943 = ( x96 & ~n15942 ) | ( x96 & n15941 ) | ( ~n15942 & n15941 ) ;
  assign n15944 = ( n3170 & ~n7541 ) | ( n3170 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n15945 = n15943 | n15944 ;
  assign n15946 = ( x56 & ~n15945 ) | ( x56 & 1'b0 ) | ( ~n15945 & 1'b0 ) ;
  assign n15947 = ~x56 & n15945 ;
  assign n15948 = n15946 | n15947 ;
  assign n15950 = ( n15907 & n15938 ) | ( n15907 & n15948 ) | ( n15938 & n15948 ) ;
  assign n15949 = ( n15938 & ~n15907 ) | ( n15938 & n15948 ) | ( ~n15907 & n15948 ) ;
  assign n15951 = ( n15907 & ~n15950 ) | ( n15907 & n15949 ) | ( ~n15950 & n15949 ) ;
  assign n15955 = x99 &  n6982 ;
  assign n15952 = ( x101 & ~n6727 ) | ( x101 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n15953 = x100 &  n6722 ;
  assign n15954 = n15952 | n15953 ;
  assign n15956 = ( x99 & ~n15955 ) | ( x99 & n15954 ) | ( ~n15955 & n15954 ) ;
  assign n15957 = n3694 | n6730 ;
  assign n15958 = ~n15956 & n15957 ;
  assign n15959 = x53 &  n15958 ;
  assign n15960 = x53 | n15958 ;
  assign n15961 = ~n15959 & n15960 ;
  assign n15963 = ( n15753 & n15951 ) | ( n15753 & n15961 ) | ( n15951 & n15961 ) ;
  assign n15962 = ( n15951 & ~n15753 ) | ( n15951 & n15961 ) | ( ~n15753 & n15961 ) ;
  assign n15964 = ( n15753 & ~n15963 ) | ( n15753 & n15962 ) | ( ~n15963 & n15962 ) ;
  assign n15965 = ( n15896 & n15906 ) | ( n15896 & n15964 ) | ( n15906 & n15964 ) ;
  assign n15966 = ( n15906 & ~n15896 ) | ( n15906 & n15964 ) | ( ~n15896 & n15964 ) ;
  assign n15967 = ( n15896 & ~n15965 ) | ( n15896 & n15966 ) | ( ~n15965 & n15966 ) ;
  assign n15968 = ( n15770 & n15895 ) | ( n15770 & n15967 ) | ( n15895 & n15967 ) ;
  assign n15969 = ( n15895 & ~n15770 ) | ( n15895 & n15967 ) | ( ~n15770 & n15967 ) ;
  assign n15970 = ( n15770 & ~n15968 ) | ( n15770 & n15969 ) | ( ~n15968 & n15969 ) ;
  assign n15981 = ( n15885 & ~n15980 ) | ( n15885 & n15970 ) | ( ~n15980 & n15970 ) ;
  assign n15982 = ( n15885 & ~n15970 ) | ( n15885 & n15980 ) | ( ~n15970 & n15980 ) ;
  assign n15983 = ( n15981 & ~n15885 ) | ( n15981 & n15982 ) | ( ~n15885 & n15982 ) ;
  assign n15987 = x111 &  n4344 ;
  assign n15984 = ( x113 & ~n4143 ) | ( x113 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n15985 = x112 &  n4138 ;
  assign n15986 = n15984 | n15985 ;
  assign n15988 = ( x111 & ~n15987 ) | ( x111 & n15986 ) | ( ~n15987 & n15986 ) ;
  assign n15989 = n4146 | n6169 ;
  assign n15990 = ~n15988 & n15989 ;
  assign n15991 = x41 &  n15990 ;
  assign n15992 = x41 | n15990 ;
  assign n15993 = ~n15991 & n15992 ;
  assign n15994 = ( n15884 & n15983 ) | ( n15884 & n15993 ) | ( n15983 & n15993 ) ;
  assign n15995 = ( n15983 & ~n15884 ) | ( n15983 & n15993 ) | ( ~n15884 & n15993 ) ;
  assign n15996 = ( n15884 & ~n15994 ) | ( n15884 & n15995 ) | ( ~n15994 & n15995 ) ;
  assign n16000 = x114 &  n3756 ;
  assign n15997 = ( x116 & ~n3602 ) | ( x116 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n15998 = x115 &  n3597 ;
  assign n15999 = n15997 | n15998 ;
  assign n16001 = ( x114 & ~n16000 ) | ( x114 & n15999 ) | ( ~n16000 & n15999 ) ;
  assign n16002 = n3605 | n6885 ;
  assign n16003 = ~n16001 & n16002 ;
  assign n16004 = x38 &  n16003 ;
  assign n16005 = x38 | n16003 ;
  assign n16006 = ~n16004 & n16005 ;
  assign n16008 = ( n15802 & n15996 ) | ( n15802 & n16006 ) | ( n15996 & n16006 ) ;
  assign n16007 = ( n15996 & ~n15802 ) | ( n15996 & n16006 ) | ( ~n15802 & n16006 ) ;
  assign n16009 = ( n15802 & ~n16008 ) | ( n15802 & n16007 ) | ( ~n16008 & n16007 ) ;
  assign n16014 = x117 &  n3214 ;
  assign n16011 = ( x119 & ~n3087 ) | ( x119 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n16012 = x118 &  n3082 ;
  assign n16013 = n16011 | n16012 ;
  assign n16015 = ( x117 & ~n16014 ) | ( x117 & n16013 ) | ( ~n16014 & n16013 ) ;
  assign n16016 = ~n3090 & n7648 ;
  assign n16017 = n16015 | n16016 ;
  assign n16018 = ( x35 & ~n16017 ) | ( x35 & 1'b0 ) | ( ~n16017 & 1'b0 ) ;
  assign n16019 = ~x35 & n16017 ;
  assign n16020 = n16018 | n16019 ;
  assign n16010 = ( n15804 & ~n15805 ) | ( n15804 & n15815 ) | ( ~n15805 & n15815 ) ;
  assign n16021 = ( n16009 & ~n16020 ) | ( n16009 & n16010 ) | ( ~n16020 & n16010 ) ;
  assign n16022 = ( n16009 & ~n16010 ) | ( n16009 & n16020 ) | ( ~n16010 & n16020 ) ;
  assign n16023 = ( n16021 & ~n16009 ) | ( n16021 & n16022 ) | ( ~n16009 & n16022 ) ;
  assign n16024 = ( n15882 & n15883 ) | ( n15882 & n16023 ) | ( n15883 & n16023 ) ;
  assign n16025 = ( n15883 & ~n15882 ) | ( n15883 & n16023 ) | ( ~n15882 & n16023 ) ;
  assign n16026 = ( n15882 & ~n16024 ) | ( n15882 & n16025 ) | ( ~n16024 & n16025 ) ;
  assign n16028 = ( n15862 & n15872 ) | ( n15862 & n16026 ) | ( n15872 & n16026 ) ;
  assign n16027 = ( n15872 & ~n15862 ) | ( n15872 & n16026 ) | ( ~n15862 & n16026 ) ;
  assign n16029 = ( n15862 & ~n16028 ) | ( n15862 & n16027 ) | ( ~n16028 & n16027 ) ;
  assign n16030 = ( x126 & ~n1894 ) | ( x126 & 1'b0 ) | ( ~n1894 & 1'b0 ) ;
  assign n16031 = x127 &  n1811 ;
  assign n16032 = n16030 | n16031 ;
  assign n16033 = n1819 | n9960 ;
  assign n16034 = ( n16032 & ~n1819 ) | ( n16032 & n16033 ) | ( ~n1819 & n16033 ) ;
  assign n16035 = x26 | n16034 ;
  assign n16036 = ( x26 & ~n16034 ) | ( x26 & 1'b0 ) | ( ~n16034 & 1'b0 ) ;
  assign n16037 = ( n16035 & ~x26 ) | ( n16035 & n16036 ) | ( ~x26 & n16036 ) ;
  assign n16038 = ( n15859 & ~n16029 ) | ( n15859 & n16037 ) | ( ~n16029 & n16037 ) ;
  assign n16039 = ( n15859 & ~n16037 ) | ( n15859 & n16029 ) | ( ~n16037 & n16029 ) ;
  assign n16040 = ( n16038 & ~n15859 ) | ( n16038 & n16039 ) | ( ~n15859 & n16039 ) ;
  assign n16041 = ( n15857 & ~n15858 ) | ( n15857 & n16040 ) | ( ~n15858 & n16040 ) ;
  assign n16042 = ( n15857 & ~n16040 ) | ( n15857 & n15858 ) | ( ~n16040 & n15858 ) ;
  assign n16043 = ( n16041 & ~n15857 ) | ( n16041 & n16042 ) | ( ~n15857 & n16042 ) ;
  assign n16054 = x124 &  n2312 ;
  assign n16051 = ( x126 & ~n2195 ) | ( x126 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n16052 = x125 &  n2190 ;
  assign n16053 = n16051 | n16052 ;
  assign n16055 = ( x124 & ~n16054 ) | ( x124 & n16053 ) | ( ~n16054 & n16053 ) ;
  assign n16056 = n2198 | n9349 ;
  assign n16057 = ~n16055 & n16056 ;
  assign n16058 = x29 &  n16057 ;
  assign n16059 = x29 | n16057 ;
  assign n16060 = ~n16058 & n16059 ;
  assign n16061 = ( n16010 & ~n16009 ) | ( n16010 & n16020 ) | ( ~n16009 & n16020 ) ;
  assign n16065 = x121 &  n2718 ;
  assign n16062 = ( x123 & ~n2642 ) | ( x123 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n16063 = x122 &  n2637 ;
  assign n16064 = n16062 | n16063 ;
  assign n16066 = ( x121 & ~n16065 ) | ( x121 & n16064 ) | ( ~n16065 & n16064 ) ;
  assign n16067 = ~n2645 & n8472 ;
  assign n16068 = n16066 | n16067 ;
  assign n16070 = x32 &  n16068 ;
  assign n16069 = ~x32 & n16068 ;
  assign n16071 = ( x32 & ~n16070 ) | ( x32 & n16069 ) | ( ~n16070 & n16069 ) ;
  assign n16072 = ( n15802 & ~n16006 ) | ( n15802 & n15996 ) | ( ~n16006 & n15996 ) ;
  assign n16076 = x118 &  n3214 ;
  assign n16073 = ( x120 & ~n3087 ) | ( x120 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n16074 = x119 &  n3082 ;
  assign n16075 = n16073 | n16074 ;
  assign n16077 = ( x118 & ~n16076 ) | ( x118 & n16075 ) | ( ~n16076 & n16075 ) ;
  assign n16078 = ~n3090 & n9364 ;
  assign n16079 = n16077 | n16078 ;
  assign n16080 = ( x35 & ~n16079 ) | ( x35 & 1'b0 ) | ( ~n16079 & 1'b0 ) ;
  assign n16081 = ~x35 & n16079 ;
  assign n16082 = n16080 | n16081 ;
  assign n16083 = ( n15884 & ~n15983 ) | ( n15884 & n15993 ) | ( ~n15983 & n15993 ) ;
  assign n16087 = x115 &  n3756 ;
  assign n16084 = ( x117 & ~n3602 ) | ( x117 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n16085 = x116 &  n3597 ;
  assign n16086 = n16084 | n16085 ;
  assign n16088 = ( x115 & ~n16087 ) | ( x115 & n16086 ) | ( ~n16087 & n16086 ) ;
  assign n16089 = n3605 | n7136 ;
  assign n16090 = ~n16088 & n16089 ;
  assign n16091 = x38 &  n16090 ;
  assign n16092 = x38 | n16090 ;
  assign n16093 = ~n16091 & n16092 ;
  assign n16094 = ( n15970 & ~n15885 ) | ( n15970 & n15980 ) | ( ~n15885 & n15980 ) ;
  assign n16098 = x106 &  n5586 ;
  assign n16095 = ( x108 & ~n5389 ) | ( x108 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n16096 = x107 &  n5384 ;
  assign n16097 = n16095 | n16096 ;
  assign n16099 = ( x106 & ~n16098 ) | ( x106 & n16097 ) | ( ~n16098 & n16097 ) ;
  assign n16100 = n5055 | n5392 ;
  assign n16101 = ~n16099 & n16100 ;
  assign n16102 = x47 &  n16101 ;
  assign n16103 = x47 | n16101 ;
  assign n16104 = ~n16102 & n16103 ;
  assign n16105 = ( n15753 & ~n15961 ) | ( n15753 & n15951 ) | ( ~n15961 & n15951 ) ;
  assign n16106 = ( x59 & ~n15932 ) | ( x59 & 1'b0 ) | ( ~n15932 & 1'b0 ) ;
  assign n16107 = ~x59 & n15932 ;
  assign n16108 = n16106 | n16107 ;
  assign n16109 = ( n15908 & ~n15925 ) | ( n15908 & n16108 ) | ( ~n15925 & n16108 ) ;
  assign n16113 = x97 &  n7731 ;
  assign n16110 = ( x99 & ~n7538 ) | ( x99 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n16111 = x98 &  n7533 ;
  assign n16112 = n16110 | n16111 ;
  assign n16114 = ( x97 & ~n16113 ) | ( x97 & n16112 ) | ( ~n16113 & n16112 ) ;
  assign n16115 = ( n3338 & ~n7541 ) | ( n3338 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n16116 = n16114 | n16115 ;
  assign n16117 = ( x56 & ~n16116 ) | ( x56 & 1'b0 ) | ( ~n16116 & 1'b0 ) ;
  assign n16118 = ~x56 & n16116 ;
  assign n16119 = n16117 | n16118 ;
  assign n16123 = x94 &  n8558 ;
  assign n16120 = ( x96 & ~n8314 ) | ( x96 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n16121 = x95 &  n8309 ;
  assign n16122 = n16120 | n16121 ;
  assign n16124 = ( x94 & ~n16123 ) | ( x94 & n16122 ) | ( ~n16123 & n16122 ) ;
  assign n16125 = ( n2836 & ~n8317 ) | ( n2836 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n16126 = n16124 | n16125 ;
  assign n16127 = ( x59 & ~n16126 ) | ( x59 & 1'b0 ) | ( ~n16126 & 1'b0 ) ;
  assign n16128 = ~x59 & n16126 ;
  assign n16129 = n16127 | n16128 ;
  assign n16130 = x89 &  n10104 ;
  assign n16131 = ( x90 & ~n9760 ) | ( x90 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n16132 = n16130 | n16131 ;
  assign n16133 = ( n15912 & ~n16132 ) | ( n15912 & 1'b0 ) | ( ~n16132 & 1'b0 ) ;
  assign n16134 = ~n15912 & n16132 ;
  assign n16135 = n16133 | n16134 ;
  assign n16139 = x91 &  n9457 ;
  assign n16136 = ( x93 & ~n9150 ) | ( x93 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n16137 = x92 &  n9145 ;
  assign n16138 = n16136 | n16137 ;
  assign n16140 = ( x91 & ~n16139 ) | ( x91 & n16138 ) | ( ~n16139 & n16138 ) ;
  assign n16141 = ~n2264 & n9153 ;
  assign n16142 = ( n2264 & ~n16140 ) | ( n2264 & n16141 ) | ( ~n16140 & n16141 ) ;
  assign n16143 = ( x62 & n16135 ) | ( x62 & n16142 ) | ( n16135 & n16142 ) ;
  assign n16144 = ( x62 & ~n16135 ) | ( x62 & n16142 ) | ( ~n16135 & n16142 ) ;
  assign n16145 = ( n16135 & ~n16143 ) | ( n16135 & n16144 ) | ( ~n16143 & n16144 ) ;
  assign n16147 = ( n15923 & n16129 ) | ( n15923 & n16145 ) | ( n16129 & n16145 ) ;
  assign n16146 = ( n16129 & ~n15923 ) | ( n16129 & n16145 ) | ( ~n15923 & n16145 ) ;
  assign n16148 = ( n15923 & ~n16147 ) | ( n15923 & n16146 ) | ( ~n16147 & n16146 ) ;
  assign n16150 = ( n16109 & n16119 ) | ( n16109 & n16148 ) | ( n16119 & n16148 ) ;
  assign n16149 = ( n16119 & ~n16109 ) | ( n16119 & n16148 ) | ( ~n16109 & n16148 ) ;
  assign n16151 = ( n16109 & ~n16150 ) | ( n16109 & n16149 ) | ( ~n16150 & n16149 ) ;
  assign n16152 = ( n15907 & ~n15948 ) | ( n15907 & n15938 ) | ( ~n15948 & n15938 ) ;
  assign n16156 = x100 &  n6982 ;
  assign n16153 = ( x102 & ~n6727 ) | ( x102 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n16154 = x101 &  n6722 ;
  assign n16155 = n16153 | n16154 ;
  assign n16157 = ( x100 & ~n16156 ) | ( x100 & n16155 ) | ( ~n16156 & n16155 ) ;
  assign n16158 = n3872 | n6730 ;
  assign n16159 = ~n16157 & n16158 ;
  assign n16160 = x53 &  n16159 ;
  assign n16161 = x53 | n16159 ;
  assign n16162 = ~n16160 & n16161 ;
  assign n16163 = ( n16151 & ~n16152 ) | ( n16151 & n16162 ) | ( ~n16152 & n16162 ) ;
  assign n16164 = ( n16151 & ~n16162 ) | ( n16151 & n16152 ) | ( ~n16162 & n16152 ) ;
  assign n16165 = ( n16163 & ~n16151 ) | ( n16163 & n16164 ) | ( ~n16151 & n16164 ) ;
  assign n16169 = x103 &  n6288 ;
  assign n16166 = ( x105 & ~n6032 ) | ( x105 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n16167 = x104 &  n6027 ;
  assign n16168 = n16166 | n16167 ;
  assign n16170 = ( x103 & ~n16169 ) | ( x103 & n16168 ) | ( ~n16169 & n16168 ) ;
  assign n16171 = ( n4442 & ~n6035 ) | ( n4442 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n16172 = n16170 | n16171 ;
  assign n16173 = ( x50 & ~n16172 ) | ( x50 & 1'b0 ) | ( ~n16172 & 1'b0 ) ;
  assign n16174 = ~x50 & n16172 ;
  assign n16175 = n16173 | n16174 ;
  assign n16176 = ( n16105 & ~n16165 ) | ( n16105 & n16175 ) | ( ~n16165 & n16175 ) ;
  assign n16177 = ( n16105 & ~n16175 ) | ( n16105 & n16165 ) | ( ~n16175 & n16165 ) ;
  assign n16178 = ( n16176 & ~n16105 ) | ( n16176 & n16177 ) | ( ~n16105 & n16177 ) ;
  assign n16180 = ( n15966 & n16104 ) | ( n15966 & n16178 ) | ( n16104 & n16178 ) ;
  assign n16179 = ( n16104 & ~n15966 ) | ( n16104 & n16178 ) | ( ~n15966 & n16178 ) ;
  assign n16181 = ( n15966 & ~n16180 ) | ( n15966 & n16179 ) | ( ~n16180 & n16179 ) ;
  assign n16185 = x109 &  n4934 ;
  assign n16182 = ( x111 & ~n4725 ) | ( x111 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n16183 = x110 &  n4720 ;
  assign n16184 = n16182 | n16183 ;
  assign n16186 = ( x109 & ~n16185 ) | ( x109 & n16184 ) | ( ~n16185 & n16184 ) ;
  assign n16187 = n4728 | n5711 ;
  assign n16188 = ~n16186 & n16187 ;
  assign n16189 = x44 &  n16188 ;
  assign n16190 = x44 | n16188 ;
  assign n16191 = ~n16189 & n16190 ;
  assign n16192 = ( n15969 & n16181 ) | ( n15969 & n16191 ) | ( n16181 & n16191 ) ;
  assign n16193 = ( n15969 & ~n16181 ) | ( n15969 & n16191 ) | ( ~n16181 & n16191 ) ;
  assign n16194 = ( n16181 & ~n16192 ) | ( n16181 & n16193 ) | ( ~n16192 & n16193 ) ;
  assign n16198 = x112 &  n4344 ;
  assign n16195 = ( x114 & ~n4143 ) | ( x114 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n16196 = x113 &  n4138 ;
  assign n16197 = n16195 | n16196 ;
  assign n16199 = ( x112 & ~n16198 ) | ( x112 & n16197 ) | ( ~n16198 & n16197 ) ;
  assign n16200 = n4146 | n6185 ;
  assign n16201 = ~n16199 & n16200 ;
  assign n16202 = x41 &  n16201 ;
  assign n16203 = x41 | n16201 ;
  assign n16204 = ~n16202 & n16203 ;
  assign n16205 = ( n16094 & ~n16194 ) | ( n16094 & n16204 ) | ( ~n16194 & n16204 ) ;
  assign n16206 = ( n16094 & ~n16204 ) | ( n16094 & n16194 ) | ( ~n16204 & n16194 ) ;
  assign n16207 = ( n16205 & ~n16094 ) | ( n16205 & n16206 ) | ( ~n16094 & n16206 ) ;
  assign n16209 = ( n16083 & n16093 ) | ( n16083 & n16207 ) | ( n16093 & n16207 ) ;
  assign n16208 = ( n16093 & ~n16083 ) | ( n16093 & n16207 ) | ( ~n16083 & n16207 ) ;
  assign n16210 = ( n16083 & ~n16209 ) | ( n16083 & n16208 ) | ( ~n16209 & n16208 ) ;
  assign n16211 = ( n16072 & ~n16082 ) | ( n16072 & n16210 ) | ( ~n16082 & n16210 ) ;
  assign n16212 = ( n16072 & ~n16210 ) | ( n16072 & n16082 ) | ( ~n16210 & n16082 ) ;
  assign n16213 = ( n16211 & ~n16072 ) | ( n16211 & n16212 ) | ( ~n16072 & n16212 ) ;
  assign n16215 = ( n16061 & n16071 ) | ( n16061 & n16213 ) | ( n16071 & n16213 ) ;
  assign n16214 = ( n16071 & ~n16061 ) | ( n16071 & n16213 ) | ( ~n16061 & n16213 ) ;
  assign n16216 = ( n16061 & ~n16215 ) | ( n16061 & n16214 ) | ( ~n16215 & n16214 ) ;
  assign n16217 = ( n16025 & ~n16060 ) | ( n16025 & n16216 ) | ( ~n16060 & n16216 ) ;
  assign n16218 = ( n16025 & ~n16216 ) | ( n16025 & n16060 ) | ( ~n16216 & n16060 ) ;
  assign n16219 = ( n16217 & ~n16025 ) | ( n16217 & n16218 ) | ( ~n16025 & n16218 ) ;
  assign n16045 = ( x127 & ~n1894 ) | ( x127 & 1'b0 ) | ( ~n1894 & 1'b0 ) ;
  assign n16046 = n1819 | n10258 ;
  assign n16047 = ~n16045 & n16046 ;
  assign n16048 = ~x26 & n16047 ;
  assign n16049 = ( x26 & ~n16047 ) | ( x26 & 1'b0 ) | ( ~n16047 & 1'b0 ) ;
  assign n16050 = n16048 | n16049 ;
  assign n16220 = ( n16028 & ~n16219 ) | ( n16028 & n16050 ) | ( ~n16219 & n16050 ) ;
  assign n16221 = ( n16050 & ~n16028 ) | ( n16050 & n16219 ) | ( ~n16028 & n16219 ) ;
  assign n16222 = ( n16220 & ~n16050 ) | ( n16220 & n16221 ) | ( ~n16050 & n16221 ) ;
  assign n16044 = ( n15859 & n16029 ) | ( n15859 & n16037 ) | ( n16029 & n16037 ) ;
  assign n16223 = ( n16042 & ~n16222 ) | ( n16042 & n16044 ) | ( ~n16222 & n16044 ) ;
  assign n16224 = ( n16044 & ~n16042 ) | ( n16044 & n16222 ) | ( ~n16042 & n16222 ) ;
  assign n16225 = ( n16223 & ~n16044 ) | ( n16223 & n16224 ) | ( ~n16044 & n16224 ) ;
  assign n16229 = x125 &  n2312 ;
  assign n16226 = ( x127 & ~n2195 ) | ( x127 & 1'b0 ) | ( ~n2195 & 1'b0 ) ;
  assign n16227 = x126 &  n2190 ;
  assign n16228 = n16226 | n16227 ;
  assign n16230 = ( x125 & ~n16229 ) | ( x125 & n16228 ) | ( ~n16229 & n16228 ) ;
  assign n16231 = n2198 | n9941 ;
  assign n16232 = ~n16230 & n16231 ;
  assign n16233 = x29 &  n16232 ;
  assign n16234 = x29 | n16232 ;
  assign n16235 = ~n16233 & n16234 ;
  assign n16236 = ( n16025 & n16060 ) | ( n16025 & n16216 ) | ( n16060 & n16216 ) ;
  assign n16240 = x122 &  n2718 ;
  assign n16237 = ( x124 & ~n2642 ) | ( x124 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n16238 = x123 &  n2637 ;
  assign n16239 = n16237 | n16238 ;
  assign n16241 = ( x122 & ~n16240 ) | ( x122 & n16239 ) | ( ~n16240 & n16239 ) ;
  assign n16242 = ~n2645 & n8755 ;
  assign n16243 = n16241 | n16242 ;
  assign n16244 = ( x32 & ~n16243 ) | ( x32 & 1'b0 ) | ( ~n16243 & 1'b0 ) ;
  assign n16245 = ~x32 & n16243 ;
  assign n16246 = n16244 | n16245 ;
  assign n16381 = x119 &  n3214 ;
  assign n16378 = ( x121 & ~n3087 ) | ( x121 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n16379 = x120 &  n3082 ;
  assign n16380 = n16378 | n16379 ;
  assign n16382 = ( x119 & ~n16381 ) | ( x119 & n16380 ) | ( ~n16381 & n16380 ) ;
  assign n16383 = ~n3090 & n8176 ;
  assign n16384 = n16382 | n16383 ;
  assign n16250 = x110 &  n4934 ;
  assign n16247 = ( x112 & ~n4725 ) | ( x112 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n16248 = x111 &  n4720 ;
  assign n16249 = n16247 | n16248 ;
  assign n16251 = ( x110 & ~n16250 ) | ( x110 & n16249 ) | ( ~n16250 & n16249 ) ;
  assign n16252 = ~n4728 & n5727 ;
  assign n16253 = n16251 | n16252 ;
  assign n16254 = ( x44 & ~n16253 ) | ( x44 & 1'b0 ) | ( ~n16253 & 1'b0 ) ;
  assign n16255 = ~x44 & n16253 ;
  assign n16256 = n16254 | n16255 ;
  assign n16260 = x101 &  n6982 ;
  assign n16257 = ( x103 & ~n6727 ) | ( x103 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n16258 = x102 &  n6722 ;
  assign n16259 = n16257 | n16258 ;
  assign n16261 = ( x101 & ~n16260 ) | ( x101 & n16259 ) | ( ~n16260 & n16259 ) ;
  assign n16262 = n4056 | n6730 ;
  assign n16263 = ~n16261 & n16262 ;
  assign n16264 = x53 &  n16263 ;
  assign n16265 = x53 | n16263 ;
  assign n16266 = ~n16264 & n16265 ;
  assign n16270 = x98 &  n7731 ;
  assign n16267 = ( x100 & ~n7538 ) | ( x100 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n16268 = x99 &  n7533 ;
  assign n16269 = n16267 | n16268 ;
  assign n16271 = ( x98 & ~n16270 ) | ( x98 & n16269 ) | ( ~n16270 & n16269 ) ;
  assign n16272 = n3354 | n7541 ;
  assign n16273 = ~n16271 & n16272 ;
  assign n16274 = x56 &  n16273 ;
  assign n16275 = x56 | n16273 ;
  assign n16276 = ~n16274 & n16275 ;
  assign n16280 = x95 &  n8558 ;
  assign n16277 = ( x97 & ~n8314 ) | ( x97 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n16278 = x96 &  n8309 ;
  assign n16279 = n16277 | n16278 ;
  assign n16281 = ( x95 & ~n16280 ) | ( x95 & n16279 ) | ( ~n16280 & n16279 ) ;
  assign n16282 = ( n2999 & ~n8317 ) | ( n2999 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n16283 = n16281 | n16282 ;
  assign n16284 = ( x59 & ~n16283 ) | ( x59 & 1'b0 ) | ( ~n16283 & 1'b0 ) ;
  assign n16285 = ~x59 & n16283 ;
  assign n16286 = n16284 | n16285 ;
  assign n16287 = x90 &  n10104 ;
  assign n16288 = ( x91 & ~n9760 ) | ( x91 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n16289 = n16287 | n16288 ;
  assign n16290 = ( x26 & n16132 ) | ( x26 & n16289 ) | ( n16132 & n16289 ) ;
  assign n16291 = ( x26 & ~n16132 ) | ( x26 & n16289 ) | ( ~n16132 & n16289 ) ;
  assign n16292 = ( n16132 & ~n16290 ) | ( n16132 & n16291 ) | ( ~n16290 & n16291 ) ;
  assign n16293 = ~x62 & n16142 ;
  assign n16294 = ( x62 & ~n16142 ) | ( x62 & n16135 ) | ( ~n16142 & n16135 ) ;
  assign n16295 = ( n16293 & ~n16133 ) | ( n16293 & n16294 ) | ( ~n16133 & n16294 ) ;
  assign n16299 = x92 &  n9457 ;
  assign n16296 = ( x94 & ~n9150 ) | ( x94 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n16297 = x93 &  n9145 ;
  assign n16298 = n16296 | n16297 ;
  assign n16300 = ( x92 & ~n16299 ) | ( x92 & n16298 ) | ( ~n16299 & n16298 ) ;
  assign n16301 = ( n2401 & ~n9153 ) | ( n2401 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n16302 = n16300 | n16301 ;
  assign n16303 = ( x62 & ~n16302 ) | ( x62 & 1'b0 ) | ( ~n16302 & 1'b0 ) ;
  assign n16304 = ~x62 & n16302 ;
  assign n16305 = n16303 | n16304 ;
  assign n16306 = ( n16292 & n16295 ) | ( n16292 & n16305 ) | ( n16295 & n16305 ) ;
  assign n16307 = ( n16295 & ~n16292 ) | ( n16295 & n16305 ) | ( ~n16292 & n16305 ) ;
  assign n16308 = ( n16292 & ~n16306 ) | ( n16292 & n16307 ) | ( ~n16306 & n16307 ) ;
  assign n16309 = ( n16147 & ~n16286 ) | ( n16147 & n16308 ) | ( ~n16286 & n16308 ) ;
  assign n16310 = ( n16147 & ~n16308 ) | ( n16147 & n16286 ) | ( ~n16308 & n16286 ) ;
  assign n16311 = ( n16309 & ~n16147 ) | ( n16309 & n16310 ) | ( ~n16147 & n16310 ) ;
  assign n16313 = ( n16150 & n16276 ) | ( n16150 & n16311 ) | ( n16276 & n16311 ) ;
  assign n16312 = ( n16150 & ~n16276 ) | ( n16150 & n16311 ) | ( ~n16276 & n16311 ) ;
  assign n16314 = ( n16276 & ~n16313 ) | ( n16276 & n16312 ) | ( ~n16313 & n16312 ) ;
  assign n16315 = ( n16152 & ~n16151 ) | ( n16152 & n16162 ) | ( ~n16151 & n16162 ) ;
  assign n16316 = ( n16266 & n16314 ) | ( n16266 & n16315 ) | ( n16314 & n16315 ) ;
  assign n16317 = ( n16314 & ~n16266 ) | ( n16314 & n16315 ) | ( ~n16266 & n16315 ) ;
  assign n16318 = ( n16266 & ~n16316 ) | ( n16266 & n16317 ) | ( ~n16316 & n16317 ) ;
  assign n16319 = ( n16105 & n16165 ) | ( n16105 & n16175 ) | ( n16165 & n16175 ) ;
  assign n16323 = x104 &  n6288 ;
  assign n16320 = ( x106 & ~n6032 ) | ( x106 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n16321 = x105 &  n6027 ;
  assign n16322 = n16320 | n16321 ;
  assign n16324 = ( x104 & ~n16323 ) | ( x104 & n16322 ) | ( ~n16323 & n16322 ) ;
  assign n16325 = ( n4458 & ~n6035 ) | ( n4458 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n16326 = n16324 | n16325 ;
  assign n16327 = ( x50 & ~n16326 ) | ( x50 & 1'b0 ) | ( ~n16326 & 1'b0 ) ;
  assign n16328 = ~x50 & n16326 ;
  assign n16329 = n16327 | n16328 ;
  assign n16330 = ( n16318 & ~n16319 ) | ( n16318 & n16329 ) | ( ~n16319 & n16329 ) ;
  assign n16331 = ( n16318 & ~n16329 ) | ( n16318 & n16319 ) | ( ~n16329 & n16319 ) ;
  assign n16332 = ( n16330 & ~n16318 ) | ( n16330 & n16331 ) | ( ~n16318 & n16331 ) ;
  assign n16333 = ( n15966 & ~n16178 ) | ( n15966 & n16104 ) | ( ~n16178 & n16104 ) ;
  assign n16337 = x107 &  n5586 ;
  assign n16334 = ( x109 & ~n5389 ) | ( x109 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n16335 = x108 &  n5384 ;
  assign n16336 = n16334 | n16335 ;
  assign n16338 = ( x107 & ~n16337 ) | ( x107 & n16336 ) | ( ~n16337 & n16336 ) ;
  assign n16339 = ( n5267 & ~n5392 ) | ( n5267 & 1'b0 ) | ( ~n5392 & 1'b0 ) ;
  assign n16340 = n16338 | n16339 ;
  assign n16341 = ( x47 & ~n16340 ) | ( x47 & 1'b0 ) | ( ~n16340 & 1'b0 ) ;
  assign n16342 = ~x47 & n16340 ;
  assign n16343 = n16341 | n16342 ;
  assign n16345 = ( n16332 & n16333 ) | ( n16332 & n16343 ) | ( n16333 & n16343 ) ;
  assign n16344 = ( n16333 & ~n16332 ) | ( n16333 & n16343 ) | ( ~n16332 & n16343 ) ;
  assign n16346 = ( n16332 & ~n16345 ) | ( n16332 & n16344 ) | ( ~n16345 & n16344 ) ;
  assign n16347 = ( n15969 & ~n16191 ) | ( n15969 & n16181 ) | ( ~n16191 & n16181 ) ;
  assign n16348 = ( n16256 & n16346 ) | ( n16256 & n16347 ) | ( n16346 & n16347 ) ;
  assign n16349 = ( n16346 & ~n16256 ) | ( n16346 & n16347 ) | ( ~n16256 & n16347 ) ;
  assign n16350 = ( n16256 & ~n16348 ) | ( n16256 & n16349 ) | ( ~n16348 & n16349 ) ;
  assign n16351 = ( n16094 & n16194 ) | ( n16094 & n16204 ) | ( n16194 & n16204 ) ;
  assign n16355 = x113 &  n4344 ;
  assign n16352 = ( x115 & ~n4143 ) | ( x115 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n16353 = x114 &  n4138 ;
  assign n16354 = n16352 | n16353 ;
  assign n16356 = ( x113 & ~n16355 ) | ( x113 & n16354 ) | ( ~n16355 & n16354 ) ;
  assign n16357 = ~n4146 & n6420 ;
  assign n16358 = n16356 | n16357 ;
  assign n16359 = ( x41 & ~n16358 ) | ( x41 & 1'b0 ) | ( ~n16358 & 1'b0 ) ;
  assign n16360 = ~x41 & n16358 ;
  assign n16361 = n16359 | n16360 ;
  assign n16363 = ( n16350 & n16351 ) | ( n16350 & n16361 ) | ( n16351 & n16361 ) ;
  assign n16362 = ( n16351 & ~n16350 ) | ( n16351 & n16361 ) | ( ~n16350 & n16361 ) ;
  assign n16364 = ( n16350 & ~n16363 ) | ( n16350 & n16362 ) | ( ~n16363 & n16362 ) ;
  assign n16368 = x116 &  n3756 ;
  assign n16365 = ( x118 & ~n3602 ) | ( x118 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n16366 = x117 &  n3597 ;
  assign n16367 = n16365 | n16366 ;
  assign n16369 = ( x116 & ~n16368 ) | ( x116 & n16367 ) | ( ~n16368 & n16367 ) ;
  assign n16370 = n3605 | n7152 ;
  assign n16371 = ~n16369 & n16370 ;
  assign n16372 = x38 &  n16371 ;
  assign n16373 = x38 | n16371 ;
  assign n16374 = ~n16372 & n16373 ;
  assign n16375 = ( n16364 & ~n16209 ) | ( n16364 & n16374 ) | ( ~n16209 & n16374 ) ;
  assign n16376 = ( n16209 & ~n16374 ) | ( n16209 & n16364 ) | ( ~n16374 & n16364 ) ;
  assign n16377 = ( n16375 & ~n16364 ) | ( n16375 & n16376 ) | ( ~n16364 & n16376 ) ;
  assign n16385 = ( x35 & n16377 ) | ( x35 & n16384 ) | ( n16377 & n16384 ) ;
  assign n16386 = ( x35 & ~n16384 ) | ( x35 & n16377 ) | ( ~n16384 & n16377 ) ;
  assign n16387 = ( n16384 & ~n16385 ) | ( n16384 & n16386 ) | ( ~n16385 & n16386 ) ;
  assign n16388 = ~n16212 & n16387 ;
  assign n16389 = ( n16212 & ~n16387 ) | ( n16212 & 1'b0 ) | ( ~n16387 & 1'b0 ) ;
  assign n16390 = n16388 | n16389 ;
  assign n16391 = ( n16061 & ~n16213 ) | ( n16061 & n16071 ) | ( ~n16213 & n16071 ) ;
  assign n16392 = ( n16246 & ~n16390 ) | ( n16246 & n16391 ) | ( ~n16390 & n16391 ) ;
  assign n16393 = ( n16246 & ~n16391 ) | ( n16246 & n16390 ) | ( ~n16391 & n16390 ) ;
  assign n16394 = ( n16392 & ~n16246 ) | ( n16392 & n16393 ) | ( ~n16246 & n16393 ) ;
  assign n16395 = ( n16235 & ~n16236 ) | ( n16235 & n16394 ) | ( ~n16236 & n16394 ) ;
  assign n16396 = ( n16235 & ~n16394 ) | ( n16235 & n16236 ) | ( ~n16394 & n16236 ) ;
  assign n16397 = ( n16395 & ~n16235 ) | ( n16395 & n16396 ) | ( ~n16235 & n16396 ) ;
  assign n16398 = ( n16221 & n16224 ) | ( n16221 & n16397 ) | ( n16224 & n16397 ) ;
  assign n16399 = ( n16221 & ~n16397 ) | ( n16221 & n16224 ) | ( ~n16397 & n16224 ) ;
  assign n16400 = ( n16397 & ~n16398 ) | ( n16397 & n16399 ) | ( ~n16398 & n16399 ) ;
  assign n16401 = ( n16235 & n16236 ) | ( n16235 & n16394 ) | ( n16236 & n16394 ) ;
  assign n16409 = ( x35 & ~n16384 ) | ( x35 & 1'b0 ) | ( ~n16384 & 1'b0 ) ;
  assign n16410 = ~x35 & n16384 ;
  assign n16411 = n16409 | n16410 ;
  assign n16412 = ( n16212 & ~n16377 ) | ( n16212 & n16411 ) | ( ~n16377 & n16411 ) ;
  assign n16405 = x123 &  n2718 ;
  assign n16402 = ( x125 & ~n2642 ) | ( x125 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n16403 = x124 &  n2637 ;
  assign n16404 = n16402 | n16403 ;
  assign n16406 = ( x123 & ~n16405 ) | ( x123 & n16404 ) | ( ~n16405 & n16404 ) ;
  assign n16407 = ~n2645 & n9324 ;
  assign n16408 = n16406 | n16407 ;
  assign n16413 = ( x32 & n16408 ) | ( x32 & n16412 ) | ( n16408 & n16412 ) ;
  assign n16414 = ( x32 & ~n16412 ) | ( x32 & n16408 ) | ( ~n16412 & n16408 ) ;
  assign n16415 = ( n16412 & ~n16413 ) | ( n16412 & n16414 ) | ( ~n16413 & n16414 ) ;
  assign n16416 = ( n16209 & n16364 ) | ( n16209 & n16374 ) | ( n16364 & n16374 ) ;
  assign n16427 = ( n16332 & ~n16343 ) | ( n16332 & n16333 ) | ( ~n16343 & n16333 ) ;
  assign n16428 = ( n16319 & ~n16318 ) | ( n16319 & n16329 ) | ( ~n16318 & n16329 ) ;
  assign n16503 = x108 &  n5586 ;
  assign n16500 = ( x110 & ~n5389 ) | ( x110 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n16501 = x109 &  n5384 ;
  assign n16502 = n16500 | n16501 ;
  assign n16504 = ( x108 & ~n16503 ) | ( x108 & n16502 ) | ( ~n16503 & n16502 ) ;
  assign n16505 = n5283 | n5392 ;
  assign n16506 = ~n16504 & n16505 ;
  assign n16507 = x47 &  n16506 ;
  assign n16508 = x47 | n16506 ;
  assign n16509 = ~n16507 & n16508 ;
  assign n16432 = x105 &  n6288 ;
  assign n16429 = ( x107 & ~n6032 ) | ( x107 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n16430 = x106 &  n6027 ;
  assign n16431 = n16429 | n16430 ;
  assign n16433 = ( x105 & ~n16432 ) | ( x105 & n16431 ) | ( ~n16432 & n16431 ) ;
  assign n16434 = ( n4848 & ~n6035 ) | ( n4848 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n16435 = n16433 | n16434 ;
  assign n16436 = ( x50 & ~n16435 ) | ( x50 & 1'b0 ) | ( ~n16435 & 1'b0 ) ;
  assign n16437 = ~x50 & n16435 ;
  assign n16438 = n16436 | n16437 ;
  assign n16449 = ( n16147 & n16286 ) | ( n16147 & n16308 ) | ( n16286 & n16308 ) ;
  assign n16453 = x96 &  n8558 ;
  assign n16450 = ( x98 & ~n8314 ) | ( x98 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n16451 = x97 &  n8309 ;
  assign n16452 = n16450 | n16451 ;
  assign n16454 = ( x96 & ~n16453 ) | ( x96 & n16452 ) | ( ~n16453 & n16452 ) ;
  assign n16455 = ( n3170 & ~n8317 ) | ( n3170 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n16456 = n16454 | n16455 ;
  assign n16475 = x59 | n16456 ;
  assign n16476 = ~x59 & n16456 ;
  assign n16477 = ( n16475 & ~n16456 ) | ( n16475 & n16476 ) | ( ~n16456 & n16476 ) ;
  assign n16457 = ( n16132 & ~x26 ) | ( n16132 & n16289 ) | ( ~x26 & n16289 ) ;
  assign n16458 = x91 &  n10104 ;
  assign n16459 = ( x92 & ~n9760 ) | ( x92 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n16460 = n16458 | n16459 ;
  assign n16464 = x93 &  n9457 ;
  assign n16461 = ( x95 & ~n9150 ) | ( x95 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n16462 = x94 &  n9145 ;
  assign n16463 = n16461 | n16462 ;
  assign n16465 = ( x93 & ~n16464 ) | ( x93 & n16463 ) | ( ~n16464 & n16463 ) ;
  assign n16466 = ( n2547 & ~n9153 ) | ( n2547 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n16467 = n16465 | n16466 ;
  assign n16468 = ( x62 & ~n16467 ) | ( x62 & 1'b0 ) | ( ~n16467 & 1'b0 ) ;
  assign n16469 = ~x62 & n16467 ;
  assign n16470 = n16468 | n16469 ;
  assign n16471 = ( n16457 & ~n16460 ) | ( n16457 & n16470 ) | ( ~n16460 & n16470 ) ;
  assign n16472 = ( n16457 & ~n16470 ) | ( n16457 & n16460 ) | ( ~n16470 & n16460 ) ;
  assign n16473 = ( n16471 & ~n16457 ) | ( n16471 & n16472 ) | ( ~n16457 & n16472 ) ;
  assign n16474 = ( n16292 & ~n16305 ) | ( n16292 & n16295 ) | ( ~n16305 & n16295 ) ;
  assign n16479 = ( n16473 & n16474 ) | ( n16473 & n16477 ) | ( n16474 & n16477 ) ;
  assign n16478 = ( n16473 & ~n16477 ) | ( n16473 & n16474 ) | ( ~n16477 & n16474 ) ;
  assign n16480 = ( n16477 & ~n16479 ) | ( n16477 & n16478 ) | ( ~n16479 & n16478 ) ;
  assign n16484 = x99 &  n7731 ;
  assign n16481 = ( x101 & ~n7538 ) | ( x101 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n16482 = x100 &  n7533 ;
  assign n16483 = n16481 | n16482 ;
  assign n16485 = ( x99 & ~n16484 ) | ( x99 & n16483 ) | ( ~n16484 & n16483 ) ;
  assign n16486 = n3694 | n7541 ;
  assign n16487 = ~n16485 & n16486 ;
  assign n16488 = x56 &  n16487 ;
  assign n16489 = x56 | n16487 ;
  assign n16490 = ~n16488 & n16489 ;
  assign n16492 = ( n16449 & n16480 ) | ( n16449 & n16490 ) | ( n16480 & n16490 ) ;
  assign n16491 = ( n16480 & ~n16449 ) | ( n16480 & n16490 ) | ( ~n16449 & n16490 ) ;
  assign n16493 = ( n16449 & ~n16492 ) | ( n16449 & n16491 ) | ( ~n16492 & n16491 ) ;
  assign n16442 = x102 &  n6982 ;
  assign n16439 = ( x104 & ~n6727 ) | ( x104 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n16440 = x103 &  n6722 ;
  assign n16441 = n16439 | n16440 ;
  assign n16443 = ( x102 & ~n16442 ) | ( x102 & n16441 ) | ( ~n16442 & n16441 ) ;
  assign n16444 = n4249 | n6730 ;
  assign n16445 = ~n16443 & n16444 ;
  assign n16446 = x53 &  n16445 ;
  assign n16447 = x53 | n16445 ;
  assign n16448 = ~n16446 & n16447 ;
  assign n16494 = ( n16312 & ~n16493 ) | ( n16312 & n16448 ) | ( ~n16493 & n16448 ) ;
  assign n16495 = ( n16312 & ~n16448 ) | ( n16312 & n16493 ) | ( ~n16448 & n16493 ) ;
  assign n16496 = ( n16494 & ~n16312 ) | ( n16494 & n16495 ) | ( ~n16312 & n16495 ) ;
  assign n16497 = ( n16316 & n16438 ) | ( n16316 & n16496 ) | ( n16438 & n16496 ) ;
  assign n16498 = ( n16438 & ~n16316 ) | ( n16438 & n16496 ) | ( ~n16316 & n16496 ) ;
  assign n16499 = ( n16316 & ~n16497 ) | ( n16316 & n16498 ) | ( ~n16497 & n16498 ) ;
  assign n16510 = ( n16428 & ~n16509 ) | ( n16428 & n16499 ) | ( ~n16509 & n16499 ) ;
  assign n16511 = ( n16428 & ~n16499 ) | ( n16428 & n16509 ) | ( ~n16499 & n16509 ) ;
  assign n16512 = ( n16510 & ~n16428 ) | ( n16510 & n16511 ) | ( ~n16428 & n16511 ) ;
  assign n16516 = x111 &  n4934 ;
  assign n16513 = ( x113 & ~n4725 ) | ( x113 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n16514 = x112 &  n4720 ;
  assign n16515 = n16513 | n16514 ;
  assign n16517 = ( x111 & ~n16516 ) | ( x111 & n16515 ) | ( ~n16516 & n16515 ) ;
  assign n16518 = n4728 | n6169 ;
  assign n16519 = ~n16517 & n16518 ;
  assign n16520 = x44 &  n16519 ;
  assign n16521 = x44 | n16519 ;
  assign n16522 = ~n16520 & n16521 ;
  assign n16523 = ( n16427 & n16512 ) | ( n16427 & n16522 ) | ( n16512 & n16522 ) ;
  assign n16524 = ( n16512 & ~n16427 ) | ( n16512 & n16522 ) | ( ~n16427 & n16522 ) ;
  assign n16525 = ( n16427 & ~n16523 ) | ( n16427 & n16524 ) | ( ~n16523 & n16524 ) ;
  assign n16529 = x114 &  n4344 ;
  assign n16526 = ( x116 & ~n4143 ) | ( x116 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n16527 = x115 &  n4138 ;
  assign n16528 = n16526 | n16527 ;
  assign n16530 = ( x114 & ~n16529 ) | ( x114 & n16528 ) | ( ~n16529 & n16528 ) ;
  assign n16531 = n4146 | n6885 ;
  assign n16532 = ~n16530 & n16531 ;
  assign n16533 = x41 &  n16532 ;
  assign n16534 = x41 | n16532 ;
  assign n16535 = ~n16533 & n16534 ;
  assign n16537 = ( n16348 & n16525 ) | ( n16348 & n16535 ) | ( n16525 & n16535 ) ;
  assign n16536 = ( n16525 & ~n16348 ) | ( n16525 & n16535 ) | ( ~n16348 & n16535 ) ;
  assign n16538 = ( n16348 & ~n16537 ) | ( n16348 & n16536 ) | ( ~n16537 & n16536 ) ;
  assign n16543 = x117 &  n3756 ;
  assign n16540 = ( x119 & ~n3602 ) | ( x119 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n16541 = x118 &  n3597 ;
  assign n16542 = n16540 | n16541 ;
  assign n16544 = ( x117 & ~n16543 ) | ( x117 & n16542 ) | ( ~n16543 & n16542 ) ;
  assign n16545 = ~n3605 & n7648 ;
  assign n16546 = n16544 | n16545 ;
  assign n16547 = ( x38 & ~n16546 ) | ( x38 & 1'b0 ) | ( ~n16546 & 1'b0 ) ;
  assign n16548 = ~x38 & n16546 ;
  assign n16549 = n16547 | n16548 ;
  assign n16539 = ( n16350 & ~n16351 ) | ( n16350 & n16361 ) | ( ~n16351 & n16361 ) ;
  assign n16550 = ( n16538 & ~n16549 ) | ( n16538 & n16539 ) | ( ~n16549 & n16539 ) ;
  assign n16551 = ( n16538 & ~n16539 ) | ( n16538 & n16549 ) | ( ~n16539 & n16549 ) ;
  assign n16552 = ( n16550 & ~n16538 ) | ( n16550 & n16551 ) | ( ~n16538 & n16551 ) ;
  assign n16420 = x120 &  n3214 ;
  assign n16417 = ( x122 & ~n3087 ) | ( x122 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n16418 = x121 &  n3082 ;
  assign n16419 = n16417 | n16418 ;
  assign n16421 = ( x120 & ~n16420 ) | ( x120 & n16419 ) | ( ~n16420 & n16419 ) ;
  assign n16422 = ~n3090 & n9987 ;
  assign n16423 = n16421 | n16422 ;
  assign n16424 = ( x35 & ~n16423 ) | ( x35 & 1'b0 ) | ( ~n16423 & 1'b0 ) ;
  assign n16425 = ~x35 & n16423 ;
  assign n16426 = n16424 | n16425 ;
  assign n16553 = ( n16416 & ~n16552 ) | ( n16416 & n16426 ) | ( ~n16552 & n16426 ) ;
  assign n16554 = ( n16416 & ~n16426 ) | ( n16416 & n16552 ) | ( ~n16426 & n16552 ) ;
  assign n16555 = ( n16553 & ~n16416 ) | ( n16553 & n16554 ) | ( ~n16416 & n16554 ) ;
  assign n16556 = n16415 &  n16555 ;
  assign n16557 = n16415 | n16555 ;
  assign n16558 = ~n16556 & n16557 ;
  assign n16559 = ( x126 & ~n2312 ) | ( x126 & 1'b0 ) | ( ~n2312 & 1'b0 ) ;
  assign n16560 = x127 &  n2190 ;
  assign n16561 = n16559 | n16560 ;
  assign n16562 = n2198 | n9960 ;
  assign n16563 = ( n16561 & ~n2198 ) | ( n16561 & n16562 ) | ( ~n2198 & n16562 ) ;
  assign n16564 = x29 | n16563 ;
  assign n16565 = ( x29 & ~n16563 ) | ( x29 & 1'b0 ) | ( ~n16563 & 1'b0 ) ;
  assign n16566 = ( n16564 & ~x29 ) | ( n16564 & n16565 ) | ( ~x29 & n16565 ) ;
  assign n16567 = ( n16392 & ~n16558 ) | ( n16392 & n16566 ) | ( ~n16558 & n16566 ) ;
  assign n16568 = ( n16392 & ~n16566 ) | ( n16392 & n16558 ) | ( ~n16566 & n16558 ) ;
  assign n16569 = ( n16567 & ~n16392 ) | ( n16567 & n16568 ) | ( ~n16392 & n16568 ) ;
  assign n16570 = ( n16221 & ~n16224 ) | ( n16221 & n16397 ) | ( ~n16224 & n16397 ) ;
  assign n16571 = ( n16401 & n16569 ) | ( n16401 & n16570 ) | ( n16569 & n16570 ) ;
  assign n16572 = ( n16569 & ~n16401 ) | ( n16569 & n16570 ) | ( ~n16401 & n16570 ) ;
  assign n16573 = ( n16401 & ~n16571 ) | ( n16401 & n16572 ) | ( ~n16571 & n16572 ) ;
  assign n16574 = ( n16392 & n16558 ) | ( n16392 & n16566 ) | ( n16558 & n16566 ) ;
  assign n16575 = ( n16401 & ~n16569 ) | ( n16401 & n16570 ) | ( ~n16569 & n16570 ) ;
  assign n16576 = ( x127 & ~n2312 ) | ( x127 & 1'b0 ) | ( ~n2312 & 1'b0 ) ;
  assign n16577 = n2198 | n10258 ;
  assign n16578 = ~n16576 & n16577 ;
  assign n16579 = ~x29 & n16578 ;
  assign n16580 = ( x29 & ~n16578 ) | ( x29 & 1'b0 ) | ( ~n16578 & 1'b0 ) ;
  assign n16581 = n16579 | n16580 ;
  assign n16582 = ( x32 & ~n16408 ) | ( x32 & 1'b0 ) | ( ~n16408 & 1'b0 ) ;
  assign n16583 = ~x32 & n16408 ;
  assign n16584 = n16582 | n16583 ;
  assign n16585 = ( n16412 & n16555 ) | ( n16412 & n16584 ) | ( n16555 & n16584 ) ;
  assign n16589 = x124 &  n2718 ;
  assign n16586 = ( x126 & ~n2642 ) | ( x126 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n16587 = x125 &  n2637 ;
  assign n16588 = n16586 | n16587 ;
  assign n16590 = ( x124 & ~n16589 ) | ( x124 & n16588 ) | ( ~n16589 & n16588 ) ;
  assign n16591 = n2645 | n9349 ;
  assign n16592 = ~n16590 & n16591 ;
  assign n16593 = x32 &  n16592 ;
  assign n16594 = x32 | n16592 ;
  assign n16595 = ~n16593 & n16594 ;
  assign n16596 = ( n16348 & ~n16535 ) | ( n16348 & n16525 ) | ( ~n16535 & n16525 ) ;
  assign n16600 = x118 &  n3756 ;
  assign n16597 = ( x120 & ~n3602 ) | ( x120 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n16598 = x119 &  n3597 ;
  assign n16599 = n16597 | n16598 ;
  assign n16601 = ( x118 & ~n16600 ) | ( x118 & n16599 ) | ( ~n16600 & n16599 ) ;
  assign n16602 = ~n3605 & n9364 ;
  assign n16603 = n16601 | n16602 ;
  assign n16604 = ( x38 & ~n16603 ) | ( x38 & 1'b0 ) | ( ~n16603 & 1'b0 ) ;
  assign n16605 = ~x38 & n16603 ;
  assign n16606 = n16604 | n16605 ;
  assign n16607 = ( n16427 & ~n16512 ) | ( n16427 & n16522 ) | ( ~n16512 & n16522 ) ;
  assign n16611 = x115 &  n4344 ;
  assign n16608 = ( x117 & ~n4143 ) | ( x117 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n16609 = x116 &  n4138 ;
  assign n16610 = n16608 | n16609 ;
  assign n16612 = ( x115 & ~n16611 ) | ( x115 & n16610 ) | ( ~n16611 & n16610 ) ;
  assign n16613 = n4146 | n7136 ;
  assign n16614 = ~n16612 & n16613 ;
  assign n16615 = x41 &  n16614 ;
  assign n16616 = x41 | n16614 ;
  assign n16617 = ~n16615 & n16616 ;
  assign n16618 = ( n16499 & ~n16428 ) | ( n16499 & n16509 ) | ( ~n16428 & n16509 ) ;
  assign n16619 = ( n16448 & ~n16312 ) | ( n16448 & n16493 ) | ( ~n16312 & n16493 ) ;
  assign n16623 = x106 &  n6288 ;
  assign n16620 = ( x108 & ~n6032 ) | ( x108 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n16621 = x107 &  n6027 ;
  assign n16622 = n16620 | n16621 ;
  assign n16624 = ( x106 & ~n16623 ) | ( x106 & n16622 ) | ( ~n16623 & n16622 ) ;
  assign n16625 = n5055 | n6035 ;
  assign n16626 = ~n16624 & n16625 ;
  assign n16627 = x50 &  n16626 ;
  assign n16628 = x50 | n16626 ;
  assign n16629 = ~n16627 & n16628 ;
  assign n16630 = ( n16449 & ~n16490 ) | ( n16449 & n16480 ) | ( ~n16490 & n16480 ) ;
  assign n16631 = x92 &  n10104 ;
  assign n16632 = ( x93 & ~n9760 ) | ( x93 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n16633 = n16631 | n16632 ;
  assign n16634 = ( n16460 & n16471 ) | ( n16460 & n16633 ) | ( n16471 & n16633 ) ;
  assign n16635 = ( n16460 & ~n16471 ) | ( n16460 & n16633 ) | ( ~n16471 & n16633 ) ;
  assign n16636 = ( n16471 & ~n16634 ) | ( n16471 & n16635 ) | ( ~n16634 & n16635 ) ;
  assign n16650 = x94 &  n9457 ;
  assign n16647 = ( x96 & ~n9150 ) | ( x96 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n16648 = x95 &  n9145 ;
  assign n16649 = n16647 | n16648 ;
  assign n16651 = ( x94 & ~n16650 ) | ( x94 & n16649 ) | ( ~n16650 & n16649 ) ;
  assign n16652 = ( n2836 & ~n9153 ) | ( n2836 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n16653 = n16651 | n16652 ;
  assign n16654 = ( x62 & ~n16653 ) | ( x62 & 1'b0 ) | ( ~n16653 & 1'b0 ) ;
  assign n16655 = ~x62 & n16653 ;
  assign n16656 = n16654 | n16655 ;
  assign n16640 = x97 &  n8558 ;
  assign n16637 = ( x99 & ~n8314 ) | ( x99 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n16638 = x98 &  n8309 ;
  assign n16639 = n16637 | n16638 ;
  assign n16641 = ( x97 & ~n16640 ) | ( x97 & n16639 ) | ( ~n16640 & n16639 ) ;
  assign n16642 = ( n3338 & ~n8317 ) | ( n3338 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n16643 = n16641 | n16642 ;
  assign n16644 = ( x59 & ~n16643 ) | ( x59 & 1'b0 ) | ( ~n16643 & 1'b0 ) ;
  assign n16645 = ~x59 & n16643 ;
  assign n16646 = n16644 | n16645 ;
  assign n16657 = ( n16636 & ~n16656 ) | ( n16636 & n16646 ) | ( ~n16656 & n16646 ) ;
  assign n16658 = ( n16636 & ~n16646 ) | ( n16636 & n16656 ) | ( ~n16646 & n16656 ) ;
  assign n16659 = ( n16657 & ~n16636 ) | ( n16657 & n16658 ) | ( ~n16636 & n16658 ) ;
  assign n16666 = x100 &  n7731 ;
  assign n16663 = ( x102 & ~n7538 ) | ( x102 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n16664 = x101 &  n7533 ;
  assign n16665 = n16663 | n16664 ;
  assign n16667 = ( x100 & ~n16666 ) | ( x100 & n16665 ) | ( ~n16666 & n16665 ) ;
  assign n16668 = n3872 | n7541 ;
  assign n16669 = ~n16667 & n16668 ;
  assign n16670 = x56 &  n16669 ;
  assign n16671 = x56 | n16669 ;
  assign n16672 = ~n16670 & n16671 ;
  assign n16660 = ( x59 & ~n16456 ) | ( x59 & 1'b0 ) | ( ~n16456 & 1'b0 ) ;
  assign n16661 = n16476 | n16660 ;
  assign n16662 = ( n16473 & ~n16661 ) | ( n16473 & n16474 ) | ( ~n16661 & n16474 ) ;
  assign n16673 = ( n16659 & ~n16672 ) | ( n16659 & n16662 ) | ( ~n16672 & n16662 ) ;
  assign n16674 = ( n16659 & ~n16662 ) | ( n16659 & n16672 ) | ( ~n16662 & n16672 ) ;
  assign n16675 = ( n16673 & ~n16659 ) | ( n16673 & n16674 ) | ( ~n16659 & n16674 ) ;
  assign n16679 = x103 &  n6982 ;
  assign n16676 = ( x105 & ~n6727 ) | ( x105 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n16677 = x104 &  n6722 ;
  assign n16678 = n16676 | n16677 ;
  assign n16680 = ( x103 & ~n16679 ) | ( x103 & n16678 ) | ( ~n16679 & n16678 ) ;
  assign n16681 = ( n4442 & ~n6730 ) | ( n4442 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n16682 = n16680 | n16681 ;
  assign n16683 = ( x53 & ~n16682 ) | ( x53 & 1'b0 ) | ( ~n16682 & 1'b0 ) ;
  assign n16684 = ~x53 & n16682 ;
  assign n16685 = n16683 | n16684 ;
  assign n16686 = ( n16630 & n16675 ) | ( n16630 & n16685 ) | ( n16675 & n16685 ) ;
  assign n16687 = ( n16675 & ~n16630 ) | ( n16675 & n16685 ) | ( ~n16630 & n16685 ) ;
  assign n16688 = ( n16630 & ~n16686 ) | ( n16630 & n16687 ) | ( ~n16686 & n16687 ) ;
  assign n16689 = ( n16619 & ~n16629 ) | ( n16619 & n16688 ) | ( ~n16629 & n16688 ) ;
  assign n16690 = ( n16619 & ~n16688 ) | ( n16619 & n16629 ) | ( ~n16688 & n16629 ) ;
  assign n16691 = ( n16689 & ~n16619 ) | ( n16689 & n16690 ) | ( ~n16619 & n16690 ) ;
  assign n16695 = x109 &  n5586 ;
  assign n16692 = ( x111 & ~n5389 ) | ( x111 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n16693 = x110 &  n5384 ;
  assign n16694 = n16692 | n16693 ;
  assign n16696 = ( x109 & ~n16695 ) | ( x109 & n16694 ) | ( ~n16695 & n16694 ) ;
  assign n16697 = n5392 | n5711 ;
  assign n16698 = ~n16696 & n16697 ;
  assign n16699 = x47 &  n16698 ;
  assign n16700 = x47 | n16698 ;
  assign n16701 = ~n16699 & n16700 ;
  assign n16703 = ( n16498 & n16691 ) | ( n16498 & n16701 ) | ( n16691 & n16701 ) ;
  assign n16702 = ( n16498 & ~n16691 ) | ( n16498 & n16701 ) | ( ~n16691 & n16701 ) ;
  assign n16704 = ( n16691 & ~n16703 ) | ( n16691 & n16702 ) | ( ~n16703 & n16702 ) ;
  assign n16708 = x112 &  n4934 ;
  assign n16705 = ( x114 & ~n4725 ) | ( x114 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n16706 = x113 &  n4720 ;
  assign n16707 = n16705 | n16706 ;
  assign n16709 = ( x112 & ~n16708 ) | ( x112 & n16707 ) | ( ~n16708 & n16707 ) ;
  assign n16710 = n4728 | n6185 ;
  assign n16711 = ~n16709 & n16710 ;
  assign n16712 = x44 &  n16711 ;
  assign n16713 = x44 | n16711 ;
  assign n16714 = ~n16712 & n16713 ;
  assign n16715 = ( n16618 & n16704 ) | ( n16618 & n16714 ) | ( n16704 & n16714 ) ;
  assign n16716 = ( n16704 & ~n16618 ) | ( n16704 & n16714 ) | ( ~n16618 & n16714 ) ;
  assign n16717 = ( n16618 & ~n16715 ) | ( n16618 & n16716 ) | ( ~n16715 & n16716 ) ;
  assign n16718 = ( n16607 & ~n16617 ) | ( n16607 & n16717 ) | ( ~n16617 & n16717 ) ;
  assign n16719 = ( n16607 & ~n16717 ) | ( n16607 & n16617 ) | ( ~n16717 & n16617 ) ;
  assign n16720 = ( n16718 & ~n16607 ) | ( n16718 & n16719 ) | ( ~n16607 & n16719 ) ;
  assign n16722 = ( n16596 & n16606 ) | ( n16596 & n16720 ) | ( n16606 & n16720 ) ;
  assign n16721 = ( n16606 & ~n16596 ) | ( n16606 & n16720 ) | ( ~n16596 & n16720 ) ;
  assign n16723 = ( n16596 & ~n16722 ) | ( n16596 & n16721 ) | ( ~n16722 & n16721 ) ;
  assign n16728 = x121 &  n3214 ;
  assign n16725 = ( x123 & ~n3087 ) | ( x123 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n16726 = x122 &  n3082 ;
  assign n16727 = n16725 | n16726 ;
  assign n16729 = ( x121 & ~n16728 ) | ( x121 & n16727 ) | ( ~n16728 & n16727 ) ;
  assign n16730 = ~n3090 & n8472 ;
  assign n16731 = n16729 | n16730 ;
  assign n16732 = ( x35 & ~n16731 ) | ( x35 & 1'b0 ) | ( ~n16731 & 1'b0 ) ;
  assign n16733 = ~x35 & n16731 ;
  assign n16734 = n16732 | n16733 ;
  assign n16724 = ( n16539 & ~n16538 ) | ( n16539 & n16549 ) | ( ~n16538 & n16549 ) ;
  assign n16735 = ( n16723 & ~n16734 ) | ( n16723 & n16724 ) | ( ~n16734 & n16724 ) ;
  assign n16736 = ( n16723 & ~n16724 ) | ( n16723 & n16734 ) | ( ~n16724 & n16734 ) ;
  assign n16737 = ( n16735 & ~n16723 ) | ( n16735 & n16736 ) | ( ~n16723 & n16736 ) ;
  assign n16739 = ( n16554 & n16595 ) | ( n16554 & n16737 ) | ( n16595 & n16737 ) ;
  assign n16738 = ( n16595 & ~n16554 ) | ( n16595 & n16737 ) | ( ~n16554 & n16737 ) ;
  assign n16740 = ( n16554 & ~n16739 ) | ( n16554 & n16738 ) | ( ~n16739 & n16738 ) ;
  assign n16741 = ( n16581 & n16585 ) | ( n16581 & n16740 ) | ( n16585 & n16740 ) ;
  assign n16742 = ( n16585 & ~n16581 ) | ( n16585 & n16740 ) | ( ~n16581 & n16740 ) ;
  assign n16743 = ( n16581 & ~n16741 ) | ( n16581 & n16742 ) | ( ~n16741 & n16742 ) ;
  assign n16744 = ( n16574 & n16575 ) | ( n16574 & n16743 ) | ( n16575 & n16743 ) ;
  assign n16745 = ( n16575 & ~n16574 ) | ( n16575 & n16743 ) | ( ~n16574 & n16743 ) ;
  assign n16746 = ( n16574 & ~n16744 ) | ( n16574 & n16745 ) | ( ~n16744 & n16745 ) ;
  assign n16747 = ( n16554 & ~n16737 ) | ( n16554 & n16595 ) | ( ~n16737 & n16595 ) ;
  assign n16748 = ( n16723 & n16724 ) | ( n16723 & n16734 ) | ( n16724 & n16734 ) ;
  assign n16869 = x119 &  n3756 ;
  assign n16866 = ( x121 & ~n3602 ) | ( x121 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n16867 = x120 &  n3597 ;
  assign n16868 = n16866 | n16867 ;
  assign n16870 = ( x119 & ~n16869 ) | ( x119 & n16868 ) | ( ~n16869 & n16868 ) ;
  assign n16871 = ~n3605 & n8176 ;
  assign n16872 = n16870 | n16871 ;
  assign n16752 = x110 &  n5586 ;
  assign n16749 = ( x112 & ~n5389 ) | ( x112 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n16750 = x111 &  n5384 ;
  assign n16751 = n16749 | n16750 ;
  assign n16753 = ( x110 & ~n16752 ) | ( x110 & n16751 ) | ( ~n16752 & n16751 ) ;
  assign n16754 = ~n5392 & n5727 ;
  assign n16755 = n16753 | n16754 ;
  assign n16756 = ( x47 & ~n16755 ) | ( x47 & 1'b0 ) | ( ~n16755 & 1'b0 ) ;
  assign n16757 = ~x47 & n16755 ;
  assign n16758 = n16756 | n16757 ;
  assign n16759 = x93 &  n10104 ;
  assign n16760 = ( x94 & ~n9760 ) | ( x94 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n16761 = n16759 | n16760 ;
  assign n16762 = ( x29 & n16633 ) | ( x29 & n16761 ) | ( n16633 & n16761 ) ;
  assign n16763 = ( x29 & ~n16633 ) | ( x29 & n16761 ) | ( ~n16633 & n16761 ) ;
  assign n16764 = ( n16633 & ~n16762 ) | ( n16633 & n16763 ) | ( ~n16762 & n16763 ) ;
  assign n16769 = x95 &  n9457 ;
  assign n16766 = ( x97 & ~n9150 ) | ( x97 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n16767 = x96 &  n9145 ;
  assign n16768 = n16766 | n16767 ;
  assign n16770 = ( x95 & ~n16769 ) | ( x95 & n16768 ) | ( ~n16769 & n16768 ) ;
  assign n16771 = ( n2999 & ~n9153 ) | ( n2999 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n16772 = n16770 | n16771 ;
  assign n16773 = ( x62 & ~n16772 ) | ( x62 & 1'b0 ) | ( ~n16772 & 1'b0 ) ;
  assign n16774 = ~x62 & n16772 ;
  assign n16775 = n16773 | n16774 ;
  assign n16765 = ( n16460 & ~n16633 ) | ( n16460 & n16471 ) | ( ~n16633 & n16471 ) ;
  assign n16776 = ( n16764 & ~n16775 ) | ( n16764 & n16765 ) | ( ~n16775 & n16765 ) ;
  assign n16777 = ( n16764 & ~n16765 ) | ( n16764 & n16775 ) | ( ~n16765 & n16775 ) ;
  assign n16778 = ( n16776 & ~n16764 ) | ( n16776 & n16777 ) | ( ~n16764 & n16777 ) ;
  assign n16779 = ( n16646 & ~n16636 ) | ( n16646 & n16656 ) | ( ~n16636 & n16656 ) ;
  assign n16783 = x98 &  n8558 ;
  assign n16780 = ( x100 & ~n8314 ) | ( x100 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n16781 = x99 &  n8309 ;
  assign n16782 = n16780 | n16781 ;
  assign n16784 = ( x98 & ~n16783 ) | ( x98 & n16782 ) | ( ~n16783 & n16782 ) ;
  assign n16785 = n3354 | n8317 ;
  assign n16786 = ~n16784 & n16785 ;
  assign n16787 = x59 &  n16786 ;
  assign n16788 = x59 | n16786 ;
  assign n16789 = ~n16787 & n16788 ;
  assign n16790 = ( n16778 & n16779 ) | ( n16778 & n16789 ) | ( n16779 & n16789 ) ;
  assign n16791 = ( n16779 & ~n16778 ) | ( n16779 & n16789 ) | ( ~n16778 & n16789 ) ;
  assign n16792 = ( n16778 & ~n16790 ) | ( n16778 & n16791 ) | ( ~n16790 & n16791 ) ;
  assign n16796 = x101 &  n7731 ;
  assign n16793 = ( x103 & ~n7538 ) | ( x103 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n16794 = x102 &  n7533 ;
  assign n16795 = n16793 | n16794 ;
  assign n16797 = ( x101 & ~n16796 ) | ( x101 & n16795 ) | ( ~n16796 & n16795 ) ;
  assign n16798 = n4056 | n7541 ;
  assign n16799 = ~n16797 & n16798 ;
  assign n16800 = x56 &  n16799 ;
  assign n16801 = x56 | n16799 ;
  assign n16802 = ~n16800 & n16801 ;
  assign n16803 = ( n16659 & n16662 ) | ( n16659 & n16672 ) | ( n16662 & n16672 ) ;
  assign n16804 = ( n16792 & ~n16802 ) | ( n16792 & n16803 ) | ( ~n16802 & n16803 ) ;
  assign n16805 = ( n16792 & ~n16803 ) | ( n16792 & n16802 ) | ( ~n16803 & n16802 ) ;
  assign n16806 = ( n16804 & ~n16792 ) | ( n16804 & n16805 ) | ( ~n16792 & n16805 ) ;
  assign n16811 = x104 &  n6982 ;
  assign n16808 = ( x106 & ~n6727 ) | ( x106 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n16809 = x105 &  n6722 ;
  assign n16810 = n16808 | n16809 ;
  assign n16812 = ( x104 & ~n16811 ) | ( x104 & n16810 ) | ( ~n16811 & n16810 ) ;
  assign n16813 = ( n4458 & ~n6730 ) | ( n4458 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n16814 = n16812 | n16813 ;
  assign n16815 = ( x53 & ~n16814 ) | ( x53 & 1'b0 ) | ( ~n16814 & 1'b0 ) ;
  assign n16816 = ~x53 & n16814 ;
  assign n16817 = n16815 | n16816 ;
  assign n16807 = ( n16630 & ~n16675 ) | ( n16630 & n16685 ) | ( ~n16675 & n16685 ) ;
  assign n16818 = ( n16806 & ~n16817 ) | ( n16806 & n16807 ) | ( ~n16817 & n16807 ) ;
  assign n16819 = ( n16806 & ~n16807 ) | ( n16806 & n16817 ) | ( ~n16807 & n16817 ) ;
  assign n16820 = ( n16818 & ~n16806 ) | ( n16818 & n16819 ) | ( ~n16806 & n16819 ) ;
  assign n16821 = ( n16619 & n16629 ) | ( n16619 & n16688 ) | ( n16629 & n16688 ) ;
  assign n16825 = x107 &  n6288 ;
  assign n16822 = ( x109 & ~n6032 ) | ( x109 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n16823 = x108 &  n6027 ;
  assign n16824 = n16822 | n16823 ;
  assign n16826 = ( x107 & ~n16825 ) | ( x107 & n16824 ) | ( ~n16825 & n16824 ) ;
  assign n16827 = ( n5267 & ~n6035 ) | ( n5267 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n16828 = n16826 | n16827 ;
  assign n16829 = ( x50 & ~n16828 ) | ( x50 & 1'b0 ) | ( ~n16828 & 1'b0 ) ;
  assign n16830 = ~x50 & n16828 ;
  assign n16831 = n16829 | n16830 ;
  assign n16832 = ( n16820 & n16821 ) | ( n16820 & n16831 ) | ( n16821 & n16831 ) ;
  assign n16833 = ( n16821 & ~n16820 ) | ( n16821 & n16831 ) | ( ~n16820 & n16831 ) ;
  assign n16834 = ( n16820 & ~n16832 ) | ( n16820 & n16833 ) | ( ~n16832 & n16833 ) ;
  assign n16835 = ( n16691 & ~n16498 ) | ( n16691 & n16701 ) | ( ~n16498 & n16701 ) ;
  assign n16837 = ( n16758 & n16834 ) | ( n16758 & n16835 ) | ( n16834 & n16835 ) ;
  assign n16836 = ( n16834 & ~n16758 ) | ( n16834 & n16835 ) | ( ~n16758 & n16835 ) ;
  assign n16838 = ( n16758 & ~n16837 ) | ( n16758 & n16836 ) | ( ~n16837 & n16836 ) ;
  assign n16839 = ( n16618 & ~n16704 ) | ( n16618 & n16714 ) | ( ~n16704 & n16714 ) ;
  assign n16843 = x113 &  n4934 ;
  assign n16840 = ( x115 & ~n4725 ) | ( x115 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n16841 = x114 &  n4720 ;
  assign n16842 = n16840 | n16841 ;
  assign n16844 = ( x113 & ~n16843 ) | ( x113 & n16842 ) | ( ~n16843 & n16842 ) ;
  assign n16845 = ~n4728 & n6420 ;
  assign n16846 = n16844 | n16845 ;
  assign n16847 = ( x44 & ~n16846 ) | ( x44 & 1'b0 ) | ( ~n16846 & 1'b0 ) ;
  assign n16848 = ~x44 & n16846 ;
  assign n16849 = n16847 | n16848 ;
  assign n16851 = ( n16838 & n16839 ) | ( n16838 & n16849 ) | ( n16839 & n16849 ) ;
  assign n16850 = ( n16839 & ~n16838 ) | ( n16839 & n16849 ) | ( ~n16838 & n16849 ) ;
  assign n16852 = ( n16838 & ~n16851 ) | ( n16838 & n16850 ) | ( ~n16851 & n16850 ) ;
  assign n16856 = x116 &  n4344 ;
  assign n16853 = ( x118 & ~n4143 ) | ( x118 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n16854 = x117 &  n4138 ;
  assign n16855 = n16853 | n16854 ;
  assign n16857 = ( x116 & ~n16856 ) | ( x116 & n16855 ) | ( ~n16856 & n16855 ) ;
  assign n16858 = n4146 | n7152 ;
  assign n16859 = ~n16857 & n16858 ;
  assign n16860 = x41 &  n16859 ;
  assign n16861 = x41 | n16859 ;
  assign n16862 = ~n16860 & n16861 ;
  assign n16863 = ( n16852 & ~n16719 ) | ( n16852 & n16862 ) | ( ~n16719 & n16862 ) ;
  assign n16864 = ( n16719 & ~n16862 ) | ( n16719 & n16852 ) | ( ~n16862 & n16852 ) ;
  assign n16865 = ( n16863 & ~n16852 ) | ( n16863 & n16864 ) | ( ~n16852 & n16864 ) ;
  assign n16873 = ( x38 & n16865 ) | ( x38 & n16872 ) | ( n16865 & n16872 ) ;
  assign n16874 = ( x38 & ~n16872 ) | ( x38 & n16865 ) | ( ~n16872 & n16865 ) ;
  assign n16875 = ( n16872 & ~n16873 ) | ( n16872 & n16874 ) | ( ~n16873 & n16874 ) ;
  assign n16876 = ~n16722 & n16875 ;
  assign n16877 = ( n16722 & ~n16875 ) | ( n16722 & 1'b0 ) | ( ~n16875 & 1'b0 ) ;
  assign n16878 = n16876 | n16877 ;
  assign n16882 = x122 &  n3214 ;
  assign n16879 = ( x124 & ~n3087 ) | ( x124 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n16880 = x123 &  n3082 ;
  assign n16881 = n16879 | n16880 ;
  assign n16883 = ( x122 & ~n16882 ) | ( x122 & n16881 ) | ( ~n16882 & n16881 ) ;
  assign n16884 = ~n3090 & n8755 ;
  assign n16885 = n16883 | n16884 ;
  assign n16886 = ( n16878 & ~x35 ) | ( n16878 & n16885 ) | ( ~x35 & n16885 ) ;
  assign n16887 = ( x35 & ~n16878 ) | ( x35 & n16885 ) | ( ~n16878 & n16885 ) ;
  assign n16888 = ( n16886 & ~n16885 ) | ( n16886 & n16887 ) | ( ~n16885 & n16887 ) ;
  assign n16889 = n16748 &  n16888 ;
  assign n16890 = n16748 | n16888 ;
  assign n16891 = ~n16889 & n16890 ;
  assign n16895 = x125 &  n2718 ;
  assign n16892 = ( x127 & ~n2642 ) | ( x127 & 1'b0 ) | ( ~n2642 & 1'b0 ) ;
  assign n16893 = x126 &  n2637 ;
  assign n16894 = n16892 | n16893 ;
  assign n16896 = ( x125 & ~n16895 ) | ( x125 & n16894 ) | ( ~n16895 & n16894 ) ;
  assign n16897 = n2645 | n9941 ;
  assign n16898 = ~n16896 & n16897 ;
  assign n16899 = x32 &  n16898 ;
  assign n16900 = x32 | n16898 ;
  assign n16901 = ~n16899 & n16900 ;
  assign n16902 = ( n16747 & n16891 ) | ( n16747 & n16901 ) | ( n16891 & n16901 ) ;
  assign n16903 = ( n16891 & ~n16747 ) | ( n16891 & n16901 ) | ( ~n16747 & n16901 ) ;
  assign n16904 = ( n16747 & ~n16902 ) | ( n16747 & n16903 ) | ( ~n16902 & n16903 ) ;
  assign n16905 = ( n16742 & n16745 ) | ( n16742 & n16904 ) | ( n16745 & n16904 ) ;
  assign n16906 = ( n16745 & ~n16742 ) | ( n16745 & n16904 ) | ( ~n16742 & n16904 ) ;
  assign n16907 = ( n16742 & ~n16905 ) | ( n16742 & n16906 ) | ( ~n16905 & n16906 ) ;
  assign n16908 = ~x35 & n16885 ;
  assign n16909 = ( x35 & ~n16885 ) | ( x35 & 1'b0 ) | ( ~n16885 & 1'b0 ) ;
  assign n16910 = n16908 | n16909 ;
  assign n16911 = ( n16748 & ~n16878 ) | ( n16748 & n16910 ) | ( ~n16878 & n16910 ) ;
  assign n17040 = x38 | n16872 ;
  assign n17041 = ( n16877 & ~n16873 ) | ( n16877 & n17040 ) | ( ~n16873 & n17040 ) ;
  assign n16912 = ( n16719 & n16852 ) | ( n16719 & n16862 ) | ( n16852 & n16862 ) ;
  assign n16923 = ( n16820 & ~n16821 ) | ( n16820 & n16831 ) | ( ~n16821 & n16831 ) ;
  assign n16924 = ( n16806 & n16807 ) | ( n16806 & n16817 ) | ( n16807 & n16817 ) ;
  assign n16987 = x108 &  n6288 ;
  assign n16984 = ( x110 & ~n6032 ) | ( x110 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n16985 = x109 &  n6027 ;
  assign n16986 = n16984 | n16985 ;
  assign n16988 = ( x108 & ~n16987 ) | ( x108 & n16986 ) | ( ~n16987 & n16986 ) ;
  assign n16989 = n5283 | n6035 ;
  assign n16990 = ~n16988 & n16989 ;
  assign n16991 = x50 &  n16990 ;
  assign n16992 = x50 | n16990 ;
  assign n16993 = ~n16991 & n16992 ;
  assign n16925 = ( n16802 & ~n16792 ) | ( n16802 & n16803 ) | ( ~n16792 & n16803 ) ;
  assign n16929 = x105 &  n6982 ;
  assign n16926 = ( x107 & ~n6727 ) | ( x107 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n16927 = x106 &  n6722 ;
  assign n16928 = n16926 | n16927 ;
  assign n16930 = ( x105 & ~n16929 ) | ( x105 & n16928 ) | ( ~n16929 & n16928 ) ;
  assign n16931 = ( n4848 & ~n6730 ) | ( n4848 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n16932 = n16930 | n16931 ;
  assign n16933 = ( x53 & ~n16932 ) | ( x53 & 1'b0 ) | ( ~n16932 & 1'b0 ) ;
  assign n16934 = ~x53 & n16932 ;
  assign n16935 = n16933 | n16934 ;
  assign n16936 = ( n16778 & ~n16779 ) | ( n16778 & n16789 ) | ( ~n16779 & n16789 ) ;
  assign n16940 = x102 &  n7731 ;
  assign n16937 = ( x104 & ~n7538 ) | ( x104 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n16938 = x103 &  n7533 ;
  assign n16939 = n16937 | n16938 ;
  assign n16941 = ( x102 & ~n16940 ) | ( x102 & n16939 ) | ( ~n16940 & n16939 ) ;
  assign n16942 = n4249 | n7541 ;
  assign n16943 = ~n16941 & n16942 ;
  assign n16944 = x56 &  n16943 ;
  assign n16945 = x56 | n16943 ;
  assign n16946 = ~n16944 & n16945 ;
  assign n16947 = ( n16765 & ~n16764 ) | ( n16765 & n16775 ) | ( ~n16764 & n16775 ) ;
  assign n16951 = x99 &  n8558 ;
  assign n16948 = ( x101 & ~n8314 ) | ( x101 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n16949 = x100 &  n8309 ;
  assign n16950 = n16948 | n16949 ;
  assign n16952 = ( x99 & ~n16951 ) | ( x99 & n16950 ) | ( ~n16951 & n16950 ) ;
  assign n16953 = n3694 | n8317 ;
  assign n16954 = ~n16952 & n16953 ;
  assign n16955 = x59 &  n16954 ;
  assign n16956 = x59 | n16954 ;
  assign n16957 = ~n16955 & n16956 ;
  assign n16958 = ( n16633 & ~x29 ) | ( n16633 & n16761 ) | ( ~x29 & n16761 ) ;
  assign n16959 = x94 &  n10104 ;
  assign n16960 = ( x95 & ~n9760 ) | ( x95 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n16961 = n16959 | n16960 ;
  assign n16965 = x96 &  n9457 ;
  assign n16962 = ( x98 & ~n9150 ) | ( x98 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n16963 = x97 &  n9145 ;
  assign n16964 = n16962 | n16963 ;
  assign n16966 = ( x96 & ~n16965 ) | ( x96 & n16964 ) | ( ~n16965 & n16964 ) ;
  assign n16967 = ( n3170 & ~n9153 ) | ( n3170 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n16968 = n16966 | n16967 ;
  assign n16969 = ( x62 & ~n16968 ) | ( x62 & 1'b0 ) | ( ~n16968 & 1'b0 ) ;
  assign n16970 = ~x62 & n16968 ;
  assign n16971 = n16969 | n16970 ;
  assign n16972 = ( n16958 & ~n16961 ) | ( n16958 & n16971 ) | ( ~n16961 & n16971 ) ;
  assign n16973 = ( n16958 & ~n16971 ) | ( n16958 & n16961 ) | ( ~n16971 & n16961 ) ;
  assign n16974 = ( n16972 & ~n16958 ) | ( n16972 & n16973 ) | ( ~n16958 & n16973 ) ;
  assign n16975 = ( n16947 & n16957 ) | ( n16947 & n16974 ) | ( n16957 & n16974 ) ;
  assign n16976 = ( n16957 & ~n16947 ) | ( n16957 & n16974 ) | ( ~n16947 & n16974 ) ;
  assign n16977 = ( n16947 & ~n16975 ) | ( n16947 & n16976 ) | ( ~n16975 & n16976 ) ;
  assign n16978 = ( n16936 & ~n16946 ) | ( n16936 & n16977 ) | ( ~n16946 & n16977 ) ;
  assign n16979 = ( n16936 & ~n16977 ) | ( n16936 & n16946 ) | ( ~n16977 & n16946 ) ;
  assign n16980 = ( n16978 & ~n16936 ) | ( n16978 & n16979 ) | ( ~n16936 & n16979 ) ;
  assign n16981 = ( n16925 & n16935 ) | ( n16925 & n16980 ) | ( n16935 & n16980 ) ;
  assign n16982 = ( n16935 & ~n16925 ) | ( n16935 & n16980 ) | ( ~n16925 & n16980 ) ;
  assign n16983 = ( n16925 & ~n16981 ) | ( n16925 & n16982 ) | ( ~n16981 & n16982 ) ;
  assign n16994 = ( n16924 & ~n16993 ) | ( n16924 & n16983 ) | ( ~n16993 & n16983 ) ;
  assign n16995 = ( n16924 & ~n16983 ) | ( n16924 & n16993 ) | ( ~n16983 & n16993 ) ;
  assign n16996 = ( n16994 & ~n16924 ) | ( n16994 & n16995 ) | ( ~n16924 & n16995 ) ;
  assign n17000 = x111 &  n5586 ;
  assign n16997 = ( x113 & ~n5389 ) | ( x113 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n16998 = x112 &  n5384 ;
  assign n16999 = n16997 | n16998 ;
  assign n17001 = ( x111 & ~n17000 ) | ( x111 & n16999 ) | ( ~n17000 & n16999 ) ;
  assign n17002 = n5392 | n6169 ;
  assign n17003 = ~n17001 & n17002 ;
  assign n17004 = x47 &  n17003 ;
  assign n17005 = x47 | n17003 ;
  assign n17006 = ~n17004 & n17005 ;
  assign n17008 = ( n16923 & n16996 ) | ( n16923 & n17006 ) | ( n16996 & n17006 ) ;
  assign n17007 = ( n16996 & ~n16923 ) | ( n16996 & n17006 ) | ( ~n16923 & n17006 ) ;
  assign n17009 = ( n16923 & ~n17008 ) | ( n16923 & n17007 ) | ( ~n17008 & n17007 ) ;
  assign n17013 = x114 &  n4934 ;
  assign n17010 = ( x116 & ~n4725 ) | ( x116 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n17011 = x115 &  n4720 ;
  assign n17012 = n17010 | n17011 ;
  assign n17014 = ( x114 & ~n17013 ) | ( x114 & n17012 ) | ( ~n17013 & n17012 ) ;
  assign n17015 = n4728 | n6885 ;
  assign n17016 = ~n17014 & n17015 ;
  assign n17017 = x44 &  n17016 ;
  assign n17018 = x44 | n17016 ;
  assign n17019 = ~n17017 & n17018 ;
  assign n17020 = ( n16836 & ~n17009 ) | ( n16836 & n17019 ) | ( ~n17009 & n17019 ) ;
  assign n17021 = ( n16836 & ~n17019 ) | ( n16836 & n17009 ) | ( ~n17019 & n17009 ) ;
  assign n17022 = ( n17020 & ~n16836 ) | ( n17020 & n17021 ) | ( ~n16836 & n17021 ) ;
  assign n17027 = x117 &  n4344 ;
  assign n17024 = ( x119 & ~n4143 ) | ( x119 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n17025 = x118 &  n4138 ;
  assign n17026 = n17024 | n17025 ;
  assign n17028 = ( x117 & ~n17027 ) | ( x117 & n17026 ) | ( ~n17027 & n17026 ) ;
  assign n17029 = ~n4146 & n7648 ;
  assign n17030 = n17028 | n17029 ;
  assign n17031 = ( x41 & ~n17030 ) | ( x41 & 1'b0 ) | ( ~n17030 & 1'b0 ) ;
  assign n17032 = ~x41 & n17030 ;
  assign n17033 = n17031 | n17032 ;
  assign n17023 = ( n16838 & ~n16839 ) | ( n16838 & n16849 ) | ( ~n16839 & n16849 ) ;
  assign n17034 = ( n17022 & ~n17033 ) | ( n17022 & n17023 ) | ( ~n17033 & n17023 ) ;
  assign n17035 = ( n17022 & ~n17023 ) | ( n17022 & n17033 ) | ( ~n17023 & n17033 ) ;
  assign n17036 = ( n17034 & ~n17022 ) | ( n17034 & n17035 ) | ( ~n17022 & n17035 ) ;
  assign n16916 = x120 &  n3756 ;
  assign n16913 = ( x122 & ~n3602 ) | ( x122 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n16914 = x121 &  n3597 ;
  assign n16915 = n16913 | n16914 ;
  assign n16917 = ( x120 & ~n16916 ) | ( x120 & n16915 ) | ( ~n16916 & n16915 ) ;
  assign n16918 = ~n3605 & n9987 ;
  assign n16919 = n16917 | n16918 ;
  assign n16920 = ( x38 & ~n16919 ) | ( x38 & 1'b0 ) | ( ~n16919 & 1'b0 ) ;
  assign n16921 = ~x38 & n16919 ;
  assign n16922 = n16920 | n16921 ;
  assign n17037 = ( n16912 & ~n17036 ) | ( n16912 & n16922 ) | ( ~n17036 & n16922 ) ;
  assign n17038 = ( n16912 & ~n16922 ) | ( n16912 & n17036 ) | ( ~n16922 & n17036 ) ;
  assign n17039 = ( n17037 & ~n16912 ) | ( n17037 & n17038 ) | ( ~n16912 & n17038 ) ;
  assign n17045 = x123 &  n3214 ;
  assign n17042 = ( x125 & ~n3087 ) | ( x125 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n17043 = x124 &  n3082 ;
  assign n17044 = n17042 | n17043 ;
  assign n17046 = ( x123 & ~n17045 ) | ( x123 & n17044 ) | ( ~n17045 & n17044 ) ;
  assign n17047 = ~n3090 & n9324 ;
  assign n17048 = n17046 | n17047 ;
  assign n17049 = ( x35 & ~n17048 ) | ( x35 & 1'b0 ) | ( ~n17048 & 1'b0 ) ;
  assign n17050 = ~x35 & n17048 ;
  assign n17051 = n17049 | n17050 ;
  assign n17053 = ( n17039 & n17041 ) | ( n17039 & n17051 ) | ( n17041 & n17051 ) ;
  assign n17052 = ( n17039 & ~n17041 ) | ( n17039 & n17051 ) | ( ~n17041 & n17051 ) ;
  assign n17054 = ( n17041 & ~n17053 ) | ( n17041 & n17052 ) | ( ~n17053 & n17052 ) ;
  assign n17055 = ( x126 & ~n2718 ) | ( x126 & 1'b0 ) | ( ~n2718 & 1'b0 ) ;
  assign n17056 = x127 &  n2637 ;
  assign n17057 = n17055 | n17056 ;
  assign n17058 = n2645 | n9960 ;
  assign n17059 = ( n17057 & ~n2645 ) | ( n17057 & n17058 ) | ( ~n2645 & n17058 ) ;
  assign n17060 = x32 | n17059 ;
  assign n17061 = ( x32 & ~n17059 ) | ( x32 & 1'b0 ) | ( ~n17059 & 1'b0 ) ;
  assign n17062 = ( n17060 & ~x32 ) | ( n17060 & n17061 ) | ( ~x32 & n17061 ) ;
  assign n17063 = ( n16911 & ~n17054 ) | ( n16911 & n17062 ) | ( ~n17054 & n17062 ) ;
  assign n17064 = ( n16911 & ~n17062 ) | ( n16911 & n17054 ) | ( ~n17062 & n17054 ) ;
  assign n17065 = ( n17063 & ~n16911 ) | ( n17063 & n17064 ) | ( ~n16911 & n17064 ) ;
  assign n17066 = ( n16902 & n16906 ) | ( n16902 & n17065 ) | ( n16906 & n17065 ) ;
  assign n17067 = ( n16906 & ~n16902 ) | ( n16906 & n17065 ) | ( ~n16902 & n17065 ) ;
  assign n17068 = ( n16902 & ~n17066 ) | ( n16902 & n17067 ) | ( ~n17066 & n17067 ) ;
  assign n17069 = ( n16911 & n17054 ) | ( n16911 & n17062 ) | ( n17054 & n17062 ) ;
  assign n17077 = ( n16836 & n17009 ) | ( n16836 & n17019 ) | ( n17009 & n17019 ) ;
  assign n17088 = ( n16923 & ~n17006 ) | ( n16923 & n16996 ) | ( ~n17006 & n16996 ) ;
  assign n17099 = ( n16983 & ~n16924 ) | ( n16983 & n16993 ) | ( ~n16924 & n16993 ) ;
  assign n17103 = x106 &  n6982 ;
  assign n17100 = ( x108 & ~n6727 ) | ( x108 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n17101 = x107 &  n6722 ;
  assign n17102 = n17100 | n17101 ;
  assign n17104 = ( x106 & ~n17103 ) | ( x106 & n17102 ) | ( ~n17103 & n17102 ) ;
  assign n17105 = n5055 | n6730 ;
  assign n17106 = ~n17104 & n17105 ;
  assign n17107 = x53 &  n17106 ;
  assign n17108 = x53 | n17106 ;
  assign n17109 = ~n17107 & n17108 ;
  assign n17123 = x97 &  n9457 ;
  assign n17120 = ( x99 & ~n9150 ) | ( x99 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n17121 = x98 &  n9145 ;
  assign n17122 = n17120 | n17121 ;
  assign n17124 = ( x97 & ~n17123 ) | ( x97 & n17122 ) | ( ~n17123 & n17122 ) ;
  assign n17125 = ( n3338 & ~n9153 ) | ( n3338 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n17126 = n17124 | n17125 ;
  assign n17127 = ( x62 & ~n17126 ) | ( x62 & 1'b0 ) | ( ~n17126 & 1'b0 ) ;
  assign n17128 = ~x62 & n17126 ;
  assign n17129 = n17127 | n17128 ;
  assign n17139 = x100 &  n8558 ;
  assign n17136 = ( x102 & ~n8314 ) | ( x102 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n17137 = x101 &  n8309 ;
  assign n17138 = n17136 | n17137 ;
  assign n17140 = ( x100 & ~n17139 ) | ( x100 & n17138 ) | ( ~n17139 & n17138 ) ;
  assign n17141 = n3872 | n8317 ;
  assign n17142 = ~n17140 & n17141 ;
  assign n17143 = x59 &  n17142 ;
  assign n17144 = x59 | n17142 ;
  assign n17145 = ~n17143 & n17144 ;
  assign n17130 = x95 &  n10104 ;
  assign n17131 = ( x96 & ~n9760 ) | ( x96 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n17132 = n17130 | n17131 ;
  assign n17133 = ( n16961 & n16972 ) | ( n16961 & n17132 ) | ( n16972 & n17132 ) ;
  assign n17134 = ( n16961 & ~n16972 ) | ( n16961 & n17132 ) | ( ~n16972 & n17132 ) ;
  assign n17135 = ( n16972 & ~n17133 ) | ( n16972 & n17134 ) | ( ~n17133 & n17134 ) ;
  assign n17146 = ( n17129 & ~n17145 ) | ( n17129 & n17135 ) | ( ~n17145 & n17135 ) ;
  assign n17147 = ( n17129 & ~n17135 ) | ( n17129 & n17145 ) | ( ~n17135 & n17145 ) ;
  assign n17148 = ( n17146 & ~n17129 ) | ( n17146 & n17147 ) | ( ~n17129 & n17147 ) ;
  assign n17113 = x103 &  n7731 ;
  assign n17110 = ( x105 & ~n7538 ) | ( x105 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n17111 = x104 &  n7533 ;
  assign n17112 = n17110 | n17111 ;
  assign n17114 = ( x103 & ~n17113 ) | ( x103 & n17112 ) | ( ~n17113 & n17112 ) ;
  assign n17115 = ( n4442 & ~n7541 ) | ( n4442 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n17116 = n17114 | n17115 ;
  assign n17117 = ( x56 & ~n17116 ) | ( x56 & 1'b0 ) | ( ~n17116 & 1'b0 ) ;
  assign n17118 = ~x56 & n17116 ;
  assign n17119 = n17117 | n17118 ;
  assign n17149 = ( n16976 & ~n17148 ) | ( n16976 & n17119 ) | ( ~n17148 & n17119 ) ;
  assign n17150 = ( n16976 & ~n17119 ) | ( n16976 & n17148 ) | ( ~n17119 & n17148 ) ;
  assign n17151 = ( n17149 & ~n16976 ) | ( n17149 & n17150 ) | ( ~n16976 & n17150 ) ;
  assign n17153 = ( n16979 & n17109 ) | ( n16979 & n17151 ) | ( n17109 & n17151 ) ;
  assign n17152 = ( n17109 & ~n16979 ) | ( n17109 & n17151 ) | ( ~n16979 & n17151 ) ;
  assign n17154 = ( n16979 & ~n17153 ) | ( n16979 & n17152 ) | ( ~n17153 & n17152 ) ;
  assign n17158 = x109 &  n6288 ;
  assign n17155 = ( x111 & ~n6032 ) | ( x111 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n17156 = x110 &  n6027 ;
  assign n17157 = n17155 | n17156 ;
  assign n17159 = ( x109 & ~n17158 ) | ( x109 & n17157 ) | ( ~n17158 & n17157 ) ;
  assign n17160 = n5711 | n6035 ;
  assign n17161 = ~n17159 & n17160 ;
  assign n17162 = x50 &  n17161 ;
  assign n17163 = x50 | n17161 ;
  assign n17164 = ~n17162 & n17163 ;
  assign n17166 = ( n16982 & n17154 ) | ( n16982 & n17164 ) | ( n17154 & n17164 ) ;
  assign n17165 = ( n16982 & ~n17154 ) | ( n16982 & n17164 ) | ( ~n17154 & n17164 ) ;
  assign n17167 = ( n17154 & ~n17166 ) | ( n17154 & n17165 ) | ( ~n17166 & n17165 ) ;
  assign n17171 = x112 &  n5586 ;
  assign n17168 = ( x114 & ~n5389 ) | ( x114 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n17169 = x113 &  n5384 ;
  assign n17170 = n17168 | n17169 ;
  assign n17172 = ( x112 & ~n17171 ) | ( x112 & n17170 ) | ( ~n17171 & n17170 ) ;
  assign n17173 = n5392 | n6185 ;
  assign n17174 = ~n17172 & n17173 ;
  assign n17175 = x47 &  n17174 ;
  assign n17176 = x47 | n17174 ;
  assign n17177 = ~n17175 & n17176 ;
  assign n17178 = ( n17099 & n17167 ) | ( n17099 & n17177 ) | ( n17167 & n17177 ) ;
  assign n17179 = ( n17167 & ~n17099 ) | ( n17167 & n17177 ) | ( ~n17099 & n17177 ) ;
  assign n17180 = ( n17099 & ~n17178 ) | ( n17099 & n17179 ) | ( ~n17178 & n17179 ) ;
  assign n17092 = x115 &  n4934 ;
  assign n17089 = ( x117 & ~n4725 ) | ( x117 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n17090 = x116 &  n4720 ;
  assign n17091 = n17089 | n17090 ;
  assign n17093 = ( x115 & ~n17092 ) | ( x115 & n17091 ) | ( ~n17092 & n17091 ) ;
  assign n17094 = n4728 | n7136 ;
  assign n17095 = ~n17093 & n17094 ;
  assign n17096 = x44 &  n17095 ;
  assign n17097 = x44 | n17095 ;
  assign n17098 = ~n17096 & n17097 ;
  assign n17181 = ( n17088 & ~n17180 ) | ( n17088 & n17098 ) | ( ~n17180 & n17098 ) ;
  assign n17182 = ( n17088 & ~n17098 ) | ( n17088 & n17180 ) | ( ~n17098 & n17180 ) ;
  assign n17183 = ( n17181 & ~n17088 ) | ( n17181 & n17182 ) | ( ~n17088 & n17182 ) ;
  assign n17081 = x118 &  n4344 ;
  assign n17078 = ( x120 & ~n4143 ) | ( x120 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n17079 = x119 &  n4138 ;
  assign n17080 = n17078 | n17079 ;
  assign n17082 = ( x118 & ~n17081 ) | ( x118 & n17080 ) | ( ~n17081 & n17080 ) ;
  assign n17083 = ~n4146 & n9364 ;
  assign n17084 = n17082 | n17083 ;
  assign n17085 = ( x41 & ~n17084 ) | ( x41 & 1'b0 ) | ( ~n17084 & 1'b0 ) ;
  assign n17086 = ~x41 & n17084 ;
  assign n17087 = n17085 | n17086 ;
  assign n17184 = ( n17077 & ~n17183 ) | ( n17077 & n17087 ) | ( ~n17183 & n17087 ) ;
  assign n17185 = ( n17077 & ~n17087 ) | ( n17077 & n17183 ) | ( ~n17087 & n17183 ) ;
  assign n17186 = ( n17184 & ~n17077 ) | ( n17184 & n17185 ) | ( ~n17077 & n17185 ) ;
  assign n17191 = x121 &  n3756 ;
  assign n17188 = ( x123 & ~n3602 ) | ( x123 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n17189 = x122 &  n3597 ;
  assign n17190 = n17188 | n17189 ;
  assign n17192 = ( x121 & ~n17191 ) | ( x121 & n17190 ) | ( ~n17191 & n17190 ) ;
  assign n17193 = ~n3605 & n8472 ;
  assign n17194 = n17192 | n17193 ;
  assign n17195 = ( x38 & ~n17194 ) | ( x38 & 1'b0 ) | ( ~n17194 & 1'b0 ) ;
  assign n17196 = ~x38 & n17194 ;
  assign n17197 = n17195 | n17196 ;
  assign n17187 = ( n17023 & ~n17022 ) | ( n17023 & n17033 ) | ( ~n17022 & n17033 ) ;
  assign n17198 = ( n17186 & ~n17197 ) | ( n17186 & n17187 ) | ( ~n17197 & n17187 ) ;
  assign n17199 = ( n17186 & ~n17187 ) | ( n17186 & n17197 ) | ( ~n17187 & n17197 ) ;
  assign n17200 = ( n17198 & ~n17186 ) | ( n17198 & n17199 ) | ( ~n17186 & n17199 ) ;
  assign n17204 = x124 &  n3214 ;
  assign n17201 = ( x126 & ~n3087 ) | ( x126 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n17202 = x125 &  n3082 ;
  assign n17203 = n17201 | n17202 ;
  assign n17205 = ( x124 & ~n17204 ) | ( x124 & n17203 ) | ( ~n17204 & n17203 ) ;
  assign n17206 = n3090 | n9349 ;
  assign n17207 = ~n17205 & n17206 ;
  assign n17208 = x35 &  n17207 ;
  assign n17209 = x35 | n17207 ;
  assign n17210 = ~n17208 & n17209 ;
  assign n17211 = ( n17038 & n17200 ) | ( n17038 & n17210 ) | ( n17200 & n17210 ) ;
  assign n17212 = ( n17200 & ~n17038 ) | ( n17200 & n17210 ) | ( ~n17038 & n17210 ) ;
  assign n17213 = ( n17038 & ~n17211 ) | ( n17038 & n17212 ) | ( ~n17211 & n17212 ) ;
  assign n17071 = ( x127 & ~n2718 ) | ( x127 & 1'b0 ) | ( ~n2718 & 1'b0 ) ;
  assign n17072 = n2645 | n10258 ;
  assign n17073 = ~n17071 & n17072 ;
  assign n17074 = ~x32 & n17073 ;
  assign n17075 = ( x32 & ~n17073 ) | ( x32 & 1'b0 ) | ( ~n17073 & 1'b0 ) ;
  assign n17076 = n17074 | n17075 ;
  assign n17214 = ( n17053 & ~n17213 ) | ( n17053 & n17076 ) | ( ~n17213 & n17076 ) ;
  assign n17215 = ( n17076 & ~n17053 ) | ( n17076 & n17213 ) | ( ~n17053 & n17213 ) ;
  assign n17216 = ( n17214 & ~n17076 ) | ( n17214 & n17215 ) | ( ~n17076 & n17215 ) ;
  assign n17070 = ( n16902 & ~n17065 ) | ( n16902 & n16906 ) | ( ~n17065 & n16906 ) ;
  assign n17217 = ( n17069 & ~n17216 ) | ( n17069 & n17070 ) | ( ~n17216 & n17070 ) ;
  assign n17218 = ( n17069 & ~n17070 ) | ( n17069 & n17216 ) | ( ~n17070 & n17216 ) ;
  assign n17219 = ( n17217 & ~n17069 ) | ( n17217 & n17218 ) | ( ~n17069 & n17218 ) ;
  assign n17220 = ( n17053 & ~n17076 ) | ( n17053 & n17213 ) | ( ~n17076 & n17213 ) ;
  assign n17221 = ( n17070 & ~n17069 ) | ( n17070 & n17216 ) | ( ~n17069 & n17216 ) ;
  assign n17222 = ( n17038 & ~n17200 ) | ( n17038 & n17210 ) | ( ~n17200 & n17210 ) ;
  assign n17223 = ( n17186 & n17187 ) | ( n17186 & n17197 ) | ( n17187 & n17197 ) ;
  assign n17227 = x110 &  n6288 ;
  assign n17224 = ( x112 & ~n6032 ) | ( x112 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n17225 = x111 &  n6027 ;
  assign n17226 = n17224 | n17225 ;
  assign n17228 = ( x110 & ~n17227 ) | ( x110 & n17226 ) | ( ~n17227 & n17226 ) ;
  assign n17229 = ( n5727 & ~n6035 ) | ( n5727 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n17230 = n17228 | n17229 ;
  assign n17231 = ( x50 & ~n17230 ) | ( x50 & 1'b0 ) | ( ~n17230 & 1'b0 ) ;
  assign n17232 = ~x50 & n17230 ;
  assign n17233 = n17231 | n17232 ;
  assign n17237 = x107 &  n6982 ;
  assign n17234 = ( x109 & ~n6727 ) | ( x109 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n17235 = x108 &  n6722 ;
  assign n17236 = n17234 | n17235 ;
  assign n17238 = ( x107 & ~n17237 ) | ( x107 & n17236 ) | ( ~n17237 & n17236 ) ;
  assign n17239 = ( n5267 & ~n6730 ) | ( n5267 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n17240 = n17238 | n17239 ;
  assign n17241 = ( x53 & ~n17240 ) | ( x53 & 1'b0 ) | ( ~n17240 & 1'b0 ) ;
  assign n17242 = ~x53 & n17240 ;
  assign n17243 = n17241 | n17242 ;
  assign n17244 = x96 &  n10104 ;
  assign n17245 = ( x97 & ~n9760 ) | ( x97 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n17246 = n17244 | n17245 ;
  assign n17247 = ( x32 & n17132 ) | ( x32 & n17246 ) | ( n17132 & n17246 ) ;
  assign n17248 = ( x32 & ~n17132 ) | ( x32 & n17246 ) | ( ~n17132 & n17246 ) ;
  assign n17249 = ( n17132 & ~n17247 ) | ( n17132 & n17248 ) | ( ~n17247 & n17248 ) ;
  assign n17250 = ( n16961 & ~n17132 ) | ( n16961 & n16972 ) | ( ~n17132 & n16972 ) ;
  assign n17254 = x98 &  n9457 ;
  assign n17251 = ( x100 & ~n9150 ) | ( x100 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n17252 = x99 &  n9145 ;
  assign n17253 = n17251 | n17252 ;
  assign n17255 = ( x98 & ~n17254 ) | ( x98 & n17253 ) | ( ~n17254 & n17253 ) ;
  assign n17256 = n3354 | n9153 ;
  assign n17257 = ~n17255 & n17256 ;
  assign n17258 = x62 &  n17257 ;
  assign n17259 = x62 | n17257 ;
  assign n17260 = ~n17258 & n17259 ;
  assign n17261 = ( n17249 & n17250 ) | ( n17249 & n17260 ) | ( n17250 & n17260 ) ;
  assign n17262 = ( n17250 & ~n17249 ) | ( n17250 & n17260 ) | ( ~n17249 & n17260 ) ;
  assign n17263 = ( n17249 & ~n17261 ) | ( n17249 & n17262 ) | ( ~n17261 & n17262 ) ;
  assign n17268 = x101 &  n8558 ;
  assign n17265 = ( x103 & ~n8314 ) | ( x103 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n17266 = x102 &  n8309 ;
  assign n17267 = n17265 | n17266 ;
  assign n17269 = ( x101 & ~n17268 ) | ( x101 & n17267 ) | ( ~n17268 & n17267 ) ;
  assign n17270 = n4056 | n8317 ;
  assign n17271 = ~n17269 & n17270 ;
  assign n17272 = x59 &  n17271 ;
  assign n17273 = x59 | n17271 ;
  assign n17274 = ~n17272 & n17273 ;
  assign n17264 = ( n17135 & ~n17129 ) | ( n17135 & n17145 ) | ( ~n17129 & n17145 ) ;
  assign n17275 = ( n17263 & ~n17274 ) | ( n17263 & n17264 ) | ( ~n17274 & n17264 ) ;
  assign n17276 = ( n17263 & ~n17264 ) | ( n17263 & n17274 ) | ( ~n17264 & n17274 ) ;
  assign n17277 = ( n17275 & ~n17263 ) | ( n17275 & n17276 ) | ( ~n17263 & n17276 ) ;
  assign n17288 = ( n17119 & ~n16976 ) | ( n17119 & n17148 ) | ( ~n16976 & n17148 ) ;
  assign n17281 = x104 &  n7731 ;
  assign n17278 = ( x106 & ~n7538 ) | ( x106 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n17279 = x105 &  n7533 ;
  assign n17280 = n17278 | n17279 ;
  assign n17282 = ( x104 & ~n17281 ) | ( x104 & n17280 ) | ( ~n17281 & n17280 ) ;
  assign n17283 = ( n4458 & ~n7541 ) | ( n4458 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n17284 = n17282 | n17283 ;
  assign n17285 = ( x56 & ~n17284 ) | ( x56 & 1'b0 ) | ( ~n17284 & 1'b0 ) ;
  assign n17286 = ~x56 & n17284 ;
  assign n17287 = n17285 | n17286 ;
  assign n17289 = ( n17277 & ~n17288 ) | ( n17277 & n17287 ) | ( ~n17288 & n17287 ) ;
  assign n17290 = ( n17277 & ~n17287 ) | ( n17277 & n17288 ) | ( ~n17287 & n17288 ) ;
  assign n17291 = ( n17289 & ~n17277 ) | ( n17289 & n17290 ) | ( ~n17277 & n17290 ) ;
  assign n17292 = ( n17243 & ~n17153 ) | ( n17243 & n17291 ) | ( ~n17153 & n17291 ) ;
  assign n17293 = ( n17153 & ~n17291 ) | ( n17153 & n17243 ) | ( ~n17291 & n17243 ) ;
  assign n17294 = ( n17292 & ~n17243 ) | ( n17292 & n17293 ) | ( ~n17243 & n17293 ) ;
  assign n17295 = ( n17154 & ~n16982 ) | ( n17154 & n17164 ) | ( ~n16982 & n17164 ) ;
  assign n17297 = ( n17233 & n17294 ) | ( n17233 & n17295 ) | ( n17294 & n17295 ) ;
  assign n17296 = ( n17294 & ~n17233 ) | ( n17294 & n17295 ) | ( ~n17233 & n17295 ) ;
  assign n17298 = ( n17233 & ~n17297 ) | ( n17233 & n17296 ) | ( ~n17297 & n17296 ) ;
  assign n17299 = ( n17099 & ~n17167 ) | ( n17099 & n17177 ) | ( ~n17167 & n17177 ) ;
  assign n17303 = x113 &  n5586 ;
  assign n17300 = ( x115 & ~n5389 ) | ( x115 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n17301 = x114 &  n5384 ;
  assign n17302 = n17300 | n17301 ;
  assign n17304 = ( x113 & ~n17303 ) | ( x113 & n17302 ) | ( ~n17303 & n17302 ) ;
  assign n17305 = ~n5392 & n6420 ;
  assign n17306 = n17304 | n17305 ;
  assign n17307 = ( x47 & ~n17306 ) | ( x47 & 1'b0 ) | ( ~n17306 & 1'b0 ) ;
  assign n17308 = ~x47 & n17306 ;
  assign n17309 = n17307 | n17308 ;
  assign n17311 = ( n17298 & n17299 ) | ( n17298 & n17309 ) | ( n17299 & n17309 ) ;
  assign n17310 = ( n17299 & ~n17298 ) | ( n17299 & n17309 ) | ( ~n17298 & n17309 ) ;
  assign n17312 = ( n17298 & ~n17311 ) | ( n17298 & n17310 ) | ( ~n17311 & n17310 ) ;
  assign n17316 = x116 &  n4934 ;
  assign n17313 = ( x118 & ~n4725 ) | ( x118 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n17314 = x117 &  n4720 ;
  assign n17315 = n17313 | n17314 ;
  assign n17317 = ( x116 & ~n17316 ) | ( x116 & n17315 ) | ( ~n17316 & n17315 ) ;
  assign n17318 = n4728 | n7152 ;
  assign n17319 = ~n17317 & n17318 ;
  assign n17320 = x44 &  n17319 ;
  assign n17321 = x44 | n17319 ;
  assign n17322 = ~n17320 & n17321 ;
  assign n17323 = ( n17182 & n17312 ) | ( n17182 & n17322 ) | ( n17312 & n17322 ) ;
  assign n17324 = ( n17182 & ~n17312 ) | ( n17182 & n17322 ) | ( ~n17312 & n17322 ) ;
  assign n17325 = ( n17312 & ~n17323 ) | ( n17312 & n17324 ) | ( ~n17323 & n17324 ) ;
  assign n17329 = x119 &  n4344 ;
  assign n17326 = ( x121 & ~n4143 ) | ( x121 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n17327 = x120 &  n4138 ;
  assign n17328 = n17326 | n17327 ;
  assign n17330 = ( x119 & ~n17329 ) | ( x119 & n17328 ) | ( ~n17329 & n17328 ) ;
  assign n17331 = ~n4146 & n8176 ;
  assign n17332 = n17330 | n17331 ;
  assign n17333 = ( x41 & ~n17325 ) | ( x41 & n17332 ) | ( ~n17325 & n17332 ) ;
  assign n17334 = ( n17325 & ~x41 ) | ( n17325 & n17332 ) | ( ~x41 & n17332 ) ;
  assign n17335 = ( n17333 & ~n17332 ) | ( n17333 & n17334 ) | ( ~n17332 & n17334 ) ;
  assign n17336 = ( n17185 & ~n17335 ) | ( n17185 & 1'b0 ) | ( ~n17335 & 1'b0 ) ;
  assign n17337 = ~n17185 & n17335 ;
  assign n17338 = n17336 | n17337 ;
  assign n17342 = x122 &  n3756 ;
  assign n17339 = ( x124 & ~n3602 ) | ( x124 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n17340 = x123 &  n3597 ;
  assign n17341 = n17339 | n17340 ;
  assign n17343 = ( x122 & ~n17342 ) | ( x122 & n17341 ) | ( ~n17342 & n17341 ) ;
  assign n17344 = ~n3605 & n8755 ;
  assign n17345 = n17343 | n17344 ;
  assign n17346 = ( n17338 & ~x38 ) | ( n17338 & n17345 ) | ( ~x38 & n17345 ) ;
  assign n17347 = ( x38 & ~n17338 ) | ( x38 & n17345 ) | ( ~n17338 & n17345 ) ;
  assign n17348 = ( n17346 & ~n17345 ) | ( n17346 & n17347 ) | ( ~n17345 & n17347 ) ;
  assign n17349 = n17223 &  n17348 ;
  assign n17350 = n17223 | n17348 ;
  assign n17351 = ~n17349 & n17350 ;
  assign n17355 = x125 &  n3214 ;
  assign n17352 = ( x127 & ~n3087 ) | ( x127 & 1'b0 ) | ( ~n3087 & 1'b0 ) ;
  assign n17353 = x126 &  n3082 ;
  assign n17354 = n17352 | n17353 ;
  assign n17356 = ( x125 & ~n17355 ) | ( x125 & n17354 ) | ( ~n17355 & n17354 ) ;
  assign n17357 = n3090 | n9941 ;
  assign n17358 = ~n17356 & n17357 ;
  assign n17359 = x35 &  n17358 ;
  assign n17360 = x35 | n17358 ;
  assign n17361 = ~n17359 & n17360 ;
  assign n17362 = ( n17222 & n17351 ) | ( n17222 & n17361 ) | ( n17351 & n17361 ) ;
  assign n17363 = ( n17351 & ~n17222 ) | ( n17351 & n17361 ) | ( ~n17222 & n17361 ) ;
  assign n17364 = ( n17222 & ~n17362 ) | ( n17222 & n17363 ) | ( ~n17362 & n17363 ) ;
  assign n17365 = ( n17220 & n17221 ) | ( n17220 & n17364 ) | ( n17221 & n17364 ) ;
  assign n17366 = ( n17221 & ~n17220 ) | ( n17221 & n17364 ) | ( ~n17220 & n17364 ) ;
  assign n17367 = ( n17220 & ~n17365 ) | ( n17220 & n17366 ) | ( ~n17365 & n17366 ) ;
  assign n17496 = ~x38 & n17345 ;
  assign n17497 = ( x38 & ~n17345 ) | ( x38 & 1'b0 ) | ( ~n17345 & 1'b0 ) ;
  assign n17498 = n17496 | n17497 ;
  assign n17499 = ( n17223 & ~n17338 ) | ( n17223 & n17498 ) | ( ~n17338 & n17498 ) ;
  assign n17500 = ( x126 & ~n3214 ) | ( x126 & 1'b0 ) | ( ~n3214 & 1'b0 ) ;
  assign n17501 = x127 &  n3082 ;
  assign n17502 = n17500 | n17501 ;
  assign n17503 = n3090 | n9960 ;
  assign n17504 = ( n17502 & ~n3090 ) | ( n17502 & n17503 ) | ( ~n3090 & n17503 ) ;
  assign n17508 = ( n17499 & ~x35 ) | ( n17499 & n17504 ) | ( ~x35 & n17504 ) ;
  assign n17509 = ( x35 & ~n17504 ) | ( x35 & n17499 ) | ( ~n17504 & n17499 ) ;
  assign n17510 = ( n17508 & ~n17499 ) | ( n17508 & n17509 ) | ( ~n17499 & n17509 ) ;
  assign n17368 = ( n17312 & ~n17182 ) | ( n17312 & n17322 ) | ( ~n17182 & n17322 ) ;
  assign n17379 = ( n17277 & n17287 ) | ( n17277 & n17288 ) | ( n17287 & n17288 ) ;
  assign n17428 = x108 &  n6982 ;
  assign n17425 = ( x110 & ~n6727 ) | ( x110 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n17426 = x109 &  n6722 ;
  assign n17427 = n17425 | n17426 ;
  assign n17429 = ( x108 & ~n17428 ) | ( x108 & n17427 ) | ( ~n17428 & n17427 ) ;
  assign n17430 = n5283 | n6730 ;
  assign n17431 = ~n17429 & n17430 ;
  assign n17432 = x53 &  n17431 ;
  assign n17433 = x53 | n17431 ;
  assign n17434 = ~n17432 & n17433 ;
  assign n17380 = ( n17264 & ~n17263 ) | ( n17264 & n17274 ) | ( ~n17263 & n17274 ) ;
  assign n17384 = x105 &  n7731 ;
  assign n17381 = ( x107 & ~n7538 ) | ( x107 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n17382 = x106 &  n7533 ;
  assign n17383 = n17381 | n17382 ;
  assign n17385 = ( x105 & ~n17384 ) | ( x105 & n17383 ) | ( ~n17384 & n17383 ) ;
  assign n17386 = ( n4848 & ~n7541 ) | ( n4848 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n17387 = n17385 | n17386 ;
  assign n17388 = ( x56 & ~n17387 ) | ( x56 & 1'b0 ) | ( ~n17387 & 1'b0 ) ;
  assign n17389 = ~x56 & n17387 ;
  assign n17390 = n17388 | n17389 ;
  assign n17391 = ( n17249 & ~n17250 ) | ( n17249 & n17260 ) | ( ~n17250 & n17260 ) ;
  assign n17395 = x102 &  n8558 ;
  assign n17392 = ( x104 & ~n8314 ) | ( x104 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n17393 = x103 &  n8309 ;
  assign n17394 = n17392 | n17393 ;
  assign n17396 = ( x102 & ~n17395 ) | ( x102 & n17394 ) | ( ~n17395 & n17394 ) ;
  assign n17397 = n4249 | n8317 ;
  assign n17398 = ~n17396 & n17397 ;
  assign n17399 = x59 &  n17398 ;
  assign n17400 = x59 | n17398 ;
  assign n17401 = ~n17399 & n17400 ;
  assign n17402 = ( n17132 & ~x32 ) | ( n17132 & n17246 ) | ( ~x32 & n17246 ) ;
  assign n17403 = x97 &  n10104 ;
  assign n17404 = ( x98 & ~n9760 ) | ( x98 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n17405 = n17403 | n17404 ;
  assign n17409 = x99 &  n9457 ;
  assign n17406 = ( x101 & ~n9150 ) | ( x101 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n17407 = x100 &  n9145 ;
  assign n17408 = n17406 | n17407 ;
  assign n17410 = ( x99 & ~n17409 ) | ( x99 & n17408 ) | ( ~n17409 & n17408 ) ;
  assign n17411 = n3694 | n9153 ;
  assign n17412 = ~n17410 & n17411 ;
  assign n17413 = x62 &  n17412 ;
  assign n17414 = x62 | n17412 ;
  assign n17415 = ~n17413 & n17414 ;
  assign n17417 = ( n17402 & n17405 ) | ( n17402 & n17415 ) | ( n17405 & n17415 ) ;
  assign n17416 = ( n17405 & ~n17402 ) | ( n17405 & n17415 ) | ( ~n17402 & n17415 ) ;
  assign n17418 = ( n17402 & ~n17417 ) | ( n17402 & n17416 ) | ( ~n17417 & n17416 ) ;
  assign n17419 = ( n17391 & ~n17401 ) | ( n17391 & n17418 ) | ( ~n17401 & n17418 ) ;
  assign n17420 = ( n17391 & ~n17418 ) | ( n17391 & n17401 ) | ( ~n17418 & n17401 ) ;
  assign n17421 = ( n17419 & ~n17391 ) | ( n17419 & n17420 ) | ( ~n17391 & n17420 ) ;
  assign n17422 = ( n17380 & n17390 ) | ( n17380 & n17421 ) | ( n17390 & n17421 ) ;
  assign n17423 = ( n17390 & ~n17380 ) | ( n17390 & n17421 ) | ( ~n17380 & n17421 ) ;
  assign n17424 = ( n17380 & ~n17422 ) | ( n17380 & n17423 ) | ( ~n17422 & n17423 ) ;
  assign n17435 = ( n17379 & ~n17434 ) | ( n17379 & n17424 ) | ( ~n17434 & n17424 ) ;
  assign n17436 = ( n17379 & ~n17424 ) | ( n17379 & n17434 ) | ( ~n17424 & n17434 ) ;
  assign n17437 = ( n17435 & ~n17379 ) | ( n17435 & n17436 ) | ( ~n17379 & n17436 ) ;
  assign n17441 = x111 &  n6288 ;
  assign n17438 = ( x113 & ~n6032 ) | ( x113 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n17439 = x112 &  n6027 ;
  assign n17440 = n17438 | n17439 ;
  assign n17442 = ( x111 & ~n17441 ) | ( x111 & n17440 ) | ( ~n17441 & n17440 ) ;
  assign n17443 = n6035 | n6169 ;
  assign n17444 = ~n17442 & n17443 ;
  assign n17445 = x50 &  n17444 ;
  assign n17446 = x50 | n17444 ;
  assign n17447 = ~n17445 & n17446 ;
  assign n17449 = ( n17292 & n17437 ) | ( n17292 & n17447 ) | ( n17437 & n17447 ) ;
  assign n17448 = ( n17437 & ~n17292 ) | ( n17437 & n17447 ) | ( ~n17292 & n17447 ) ;
  assign n17450 = ( n17292 & ~n17449 ) | ( n17292 & n17448 ) | ( ~n17449 & n17448 ) ;
  assign n17454 = x114 &  n5586 ;
  assign n17451 = ( x116 & ~n5389 ) | ( x116 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n17452 = x115 &  n5384 ;
  assign n17453 = n17451 | n17452 ;
  assign n17455 = ( x114 & ~n17454 ) | ( x114 & n17453 ) | ( ~n17454 & n17453 ) ;
  assign n17456 = n5392 | n6885 ;
  assign n17457 = ~n17455 & n17456 ;
  assign n17458 = x47 &  n17457 ;
  assign n17459 = x47 | n17457 ;
  assign n17460 = ~n17458 & n17459 ;
  assign n17461 = ( n17296 & ~n17450 ) | ( n17296 & n17460 ) | ( ~n17450 & n17460 ) ;
  assign n17462 = ( n17296 & ~n17460 ) | ( n17296 & n17450 ) | ( ~n17460 & n17450 ) ;
  assign n17463 = ( n17461 & ~n17296 ) | ( n17461 & n17462 ) | ( ~n17296 & n17462 ) ;
  assign n17468 = x117 &  n4934 ;
  assign n17465 = ( x119 & ~n4725 ) | ( x119 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n17466 = x118 &  n4720 ;
  assign n17467 = n17465 | n17466 ;
  assign n17469 = ( x117 & ~n17468 ) | ( x117 & n17467 ) | ( ~n17468 & n17467 ) ;
  assign n17470 = ~n4728 & n7648 ;
  assign n17471 = n17469 | n17470 ;
  assign n17472 = ( x44 & ~n17471 ) | ( x44 & 1'b0 ) | ( ~n17471 & 1'b0 ) ;
  assign n17473 = ~x44 & n17471 ;
  assign n17474 = n17472 | n17473 ;
  assign n17464 = ( n17298 & ~n17299 ) | ( n17298 & n17309 ) | ( ~n17299 & n17309 ) ;
  assign n17475 = ( n17463 & ~n17474 ) | ( n17463 & n17464 ) | ( ~n17474 & n17464 ) ;
  assign n17476 = ( n17463 & ~n17464 ) | ( n17463 & n17474 ) | ( ~n17464 & n17474 ) ;
  assign n17477 = ( n17475 & ~n17463 ) | ( n17475 & n17476 ) | ( ~n17463 & n17476 ) ;
  assign n17372 = x120 &  n4344 ;
  assign n17369 = ( x122 & ~n4143 ) | ( x122 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n17370 = x121 &  n4138 ;
  assign n17371 = n17369 | n17370 ;
  assign n17373 = ( x120 & ~n17372 ) | ( x120 & n17371 ) | ( ~n17372 & n17371 ) ;
  assign n17374 = ~n4146 & n9987 ;
  assign n17375 = n17373 | n17374 ;
  assign n17376 = ( x41 & ~n17375 ) | ( x41 & 1'b0 ) | ( ~n17375 & 1'b0 ) ;
  assign n17377 = ~x41 & n17375 ;
  assign n17378 = n17376 | n17377 ;
  assign n17478 = ( n17368 & ~n17477 ) | ( n17368 & n17378 ) | ( ~n17477 & n17378 ) ;
  assign n17479 = ( n17368 & ~n17378 ) | ( n17368 & n17477 ) | ( ~n17378 & n17477 ) ;
  assign n17480 = ( n17478 & ~n17368 ) | ( n17478 & n17479 ) | ( ~n17368 & n17479 ) ;
  assign n17481 = x41 | n17332 ;
  assign n17482 = ( n17337 & ~n17333 ) | ( n17337 & n17481 ) | ( ~n17333 & n17481 ) ;
  assign n17483 = n17480 &  n17482 ;
  assign n17484 = ~n17480 & n17482 ;
  assign n17485 = ( n17480 & ~n17483 ) | ( n17480 & n17484 ) | ( ~n17483 & n17484 ) ;
  assign n17489 = x123 &  n3756 ;
  assign n17486 = ( x125 & ~n3602 ) | ( x125 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n17487 = x124 &  n3597 ;
  assign n17488 = n17486 | n17487 ;
  assign n17490 = ( x123 & ~n17489 ) | ( x123 & n17488 ) | ( ~n17489 & n17488 ) ;
  assign n17491 = ~n3605 & n9324 ;
  assign n17492 = n17490 | n17491 ;
  assign n17493 = ( x38 & ~n17492 ) | ( x38 & 1'b0 ) | ( ~n17492 & 1'b0 ) ;
  assign n17494 = ~x38 & n17492 ;
  assign n17495 = n17493 | n17494 ;
  assign n17511 = ( n17485 & n17495 ) | ( n17485 & n17510 ) | ( n17495 & n17510 ) ;
  assign n17512 = ( n17485 & ~n17510 ) | ( n17485 & n17495 ) | ( ~n17510 & n17495 ) ;
  assign n17513 = ( n17510 & ~n17511 ) | ( n17510 & n17512 ) | ( ~n17511 & n17512 ) ;
  assign n17514 = ( n17362 & n17366 ) | ( n17362 & n17513 ) | ( n17366 & n17513 ) ;
  assign n17515 = ( n17366 & ~n17362 ) | ( n17366 & n17513 ) | ( ~n17362 & n17513 ) ;
  assign n17516 = ( n17362 & ~n17514 ) | ( n17362 & n17515 ) | ( ~n17514 & n17515 ) ;
  assign n17505 = x35 | n17504 ;
  assign n17506 = ( x35 & ~n17504 ) | ( x35 & 1'b0 ) | ( ~n17504 & 1'b0 ) ;
  assign n17507 = ( n17505 & ~x35 ) | ( n17505 & n17506 ) | ( ~x35 & n17506 ) ;
  assign n17517 = n17485 &  n17495 ;
  assign n17518 = n17485 | n17495 ;
  assign n17519 = ~n17517 & n17518 ;
  assign n17520 = ( n17499 & n17507 ) | ( n17499 & n17519 ) | ( n17507 & n17519 ) ;
  assign n17522 = ( x127 & ~n3214 ) | ( x127 & 1'b0 ) | ( ~n3214 & 1'b0 ) ;
  assign n17523 = n3090 | n10258 ;
  assign n17524 = ~n17522 & n17523 ;
  assign n17525 = ~x35 & n17524 ;
  assign n17526 = ( x35 & ~n17524 ) | ( x35 & 1'b0 ) | ( ~n17524 & 1'b0 ) ;
  assign n17527 = n17525 | n17526 ;
  assign n17529 = ( n17296 & n17450 ) | ( n17296 & n17460 ) | ( n17450 & n17460 ) ;
  assign n17540 = ( n17292 & ~n17447 ) | ( n17292 & n17437 ) | ( ~n17447 & n17437 ) ;
  assign n17551 = ( n17424 & ~n17379 ) | ( n17424 & n17434 ) | ( ~n17379 & n17434 ) ;
  assign n17555 = x106 &  n7731 ;
  assign n17552 = ( x108 & ~n7538 ) | ( x108 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n17553 = x107 &  n7533 ;
  assign n17554 = n17552 | n17553 ;
  assign n17556 = ( x106 & ~n17555 ) | ( x106 & n17554 ) | ( ~n17555 & n17554 ) ;
  assign n17557 = n5055 | n7541 ;
  assign n17558 = ~n17556 & n17557 ;
  assign n17559 = x56 &  n17558 ;
  assign n17560 = x56 | n17558 ;
  assign n17561 = ~n17559 & n17560 ;
  assign n17565 = x100 &  n9457 ;
  assign n17562 = ( x102 & ~n9150 ) | ( x102 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n17563 = x101 &  n9145 ;
  assign n17564 = n17562 | n17563 ;
  assign n17566 = ( x100 & ~n17565 ) | ( x100 & n17564 ) | ( ~n17565 & n17564 ) ;
  assign n17567 = n3872 | n9153 ;
  assign n17568 = ~n17566 & n17567 ;
  assign n17569 = x62 &  n17568 ;
  assign n17570 = x62 | n17568 ;
  assign n17571 = ~n17569 & n17570 ;
  assign n17581 = x103 &  n8558 ;
  assign n17578 = ( x105 & ~n8314 ) | ( x105 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n17579 = x104 &  n8309 ;
  assign n17580 = n17578 | n17579 ;
  assign n17582 = ( x103 & ~n17581 ) | ( x103 & n17580 ) | ( ~n17581 & n17580 ) ;
  assign n17583 = ( n4442 & ~n8317 ) | ( n4442 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n17584 = n17582 | n17583 ;
  assign n17585 = ( x59 & ~n17584 ) | ( x59 & 1'b0 ) | ( ~n17584 & 1'b0 ) ;
  assign n17586 = ~x59 & n17584 ;
  assign n17587 = n17585 | n17586 ;
  assign n17572 = x98 &  n10104 ;
  assign n17573 = ( x99 & ~n9760 ) | ( x99 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n17574 = n17572 | n17573 ;
  assign n17576 = ( n17405 & n17416 ) | ( n17405 & n17574 ) | ( n17416 & n17574 ) ;
  assign n17575 = ( n17405 & ~n17416 ) | ( n17405 & n17574 ) | ( ~n17416 & n17574 ) ;
  assign n17577 = ( n17416 & ~n17576 ) | ( n17416 & n17575 ) | ( ~n17576 & n17575 ) ;
  assign n17588 = ( n17571 & ~n17587 ) | ( n17571 & n17577 ) | ( ~n17587 & n17577 ) ;
  assign n17589 = ( n17571 & ~n17577 ) | ( n17571 & n17587 ) | ( ~n17577 & n17587 ) ;
  assign n17590 = ( n17588 & ~n17571 ) | ( n17588 & n17589 ) | ( ~n17571 & n17589 ) ;
  assign n17591 = ( n17420 & ~n17561 ) | ( n17420 & n17590 ) | ( ~n17561 & n17590 ) ;
  assign n17592 = ( n17420 & ~n17590 ) | ( n17420 & n17561 ) | ( ~n17590 & n17561 ) ;
  assign n17593 = ( n17591 & ~n17420 ) | ( n17591 & n17592 ) | ( ~n17420 & n17592 ) ;
  assign n17597 = x109 &  n6982 ;
  assign n17594 = ( x111 & ~n6727 ) | ( x111 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n17595 = x110 &  n6722 ;
  assign n17596 = n17594 | n17595 ;
  assign n17598 = ( x109 & ~n17597 ) | ( x109 & n17596 ) | ( ~n17597 & n17596 ) ;
  assign n17599 = n5711 | n6730 ;
  assign n17600 = ~n17598 & n17599 ;
  assign n17601 = x53 &  n17600 ;
  assign n17602 = x53 | n17600 ;
  assign n17603 = ~n17601 & n17602 ;
  assign n17605 = ( n17423 & n17593 ) | ( n17423 & n17603 ) | ( n17593 & n17603 ) ;
  assign n17604 = ( n17423 & ~n17593 ) | ( n17423 & n17603 ) | ( ~n17593 & n17603 ) ;
  assign n17606 = ( n17593 & ~n17605 ) | ( n17593 & n17604 ) | ( ~n17605 & n17604 ) ;
  assign n17610 = x112 &  n6288 ;
  assign n17607 = ( x114 & ~n6032 ) | ( x114 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n17608 = x113 &  n6027 ;
  assign n17609 = n17607 | n17608 ;
  assign n17611 = ( x112 & ~n17610 ) | ( x112 & n17609 ) | ( ~n17610 & n17609 ) ;
  assign n17612 = n6035 | n6185 ;
  assign n17613 = ~n17611 & n17612 ;
  assign n17614 = x50 &  n17613 ;
  assign n17615 = x50 | n17613 ;
  assign n17616 = ~n17614 & n17615 ;
  assign n17617 = ( n17551 & n17606 ) | ( n17551 & n17616 ) | ( n17606 & n17616 ) ;
  assign n17618 = ( n17606 & ~n17551 ) | ( n17606 & n17616 ) | ( ~n17551 & n17616 ) ;
  assign n17619 = ( n17551 & ~n17617 ) | ( n17551 & n17618 ) | ( ~n17617 & n17618 ) ;
  assign n17544 = x115 &  n5586 ;
  assign n17541 = ( x117 & ~n5389 ) | ( x117 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n17542 = x116 &  n5384 ;
  assign n17543 = n17541 | n17542 ;
  assign n17545 = ( x115 & ~n17544 ) | ( x115 & n17543 ) | ( ~n17544 & n17543 ) ;
  assign n17546 = n5392 | n7136 ;
  assign n17547 = ~n17545 & n17546 ;
  assign n17548 = x47 &  n17547 ;
  assign n17549 = x47 | n17547 ;
  assign n17550 = ~n17548 & n17549 ;
  assign n17620 = ( n17540 & ~n17619 ) | ( n17540 & n17550 ) | ( ~n17619 & n17550 ) ;
  assign n17621 = ( n17540 & ~n17550 ) | ( n17540 & n17619 ) | ( ~n17550 & n17619 ) ;
  assign n17622 = ( n17620 & ~n17540 ) | ( n17620 & n17621 ) | ( ~n17540 & n17621 ) ;
  assign n17533 = x118 &  n4934 ;
  assign n17530 = ( x120 & ~n4725 ) | ( x120 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n17531 = x119 &  n4720 ;
  assign n17532 = n17530 | n17531 ;
  assign n17534 = ( x118 & ~n17533 ) | ( x118 & n17532 ) | ( ~n17533 & n17532 ) ;
  assign n17535 = ~n4728 & n9364 ;
  assign n17536 = n17534 | n17535 ;
  assign n17537 = ( x44 & ~n17536 ) | ( x44 & 1'b0 ) | ( ~n17536 & 1'b0 ) ;
  assign n17538 = ~x44 & n17536 ;
  assign n17539 = n17537 | n17538 ;
  assign n17623 = ( n17529 & ~n17622 ) | ( n17529 & n17539 ) | ( ~n17622 & n17539 ) ;
  assign n17624 = ( n17529 & ~n17539 ) | ( n17529 & n17622 ) | ( ~n17539 & n17622 ) ;
  assign n17625 = ( n17623 & ~n17529 ) | ( n17623 & n17624 ) | ( ~n17529 & n17624 ) ;
  assign n17630 = x121 &  n4344 ;
  assign n17627 = ( x123 & ~n4143 ) | ( x123 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n17628 = x122 &  n4138 ;
  assign n17629 = n17627 | n17628 ;
  assign n17631 = ( x121 & ~n17630 ) | ( x121 & n17629 ) | ( ~n17630 & n17629 ) ;
  assign n17632 = ~n4146 & n8472 ;
  assign n17633 = n17631 | n17632 ;
  assign n17634 = ( x41 & ~n17633 ) | ( x41 & 1'b0 ) | ( ~n17633 & 1'b0 ) ;
  assign n17635 = ~x41 & n17633 ;
  assign n17636 = n17634 | n17635 ;
  assign n17626 = ( n17464 & ~n17463 ) | ( n17464 & n17474 ) | ( ~n17463 & n17474 ) ;
  assign n17637 = ( n17625 & ~n17636 ) | ( n17625 & n17626 ) | ( ~n17636 & n17626 ) ;
  assign n17638 = ( n17625 & ~n17626 ) | ( n17625 & n17636 ) | ( ~n17626 & n17636 ) ;
  assign n17639 = ( n17637 & ~n17625 ) | ( n17637 & n17638 ) | ( ~n17625 & n17638 ) ;
  assign n17643 = x124 &  n3756 ;
  assign n17640 = ( x126 & ~n3602 ) | ( x126 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n17641 = x125 &  n3597 ;
  assign n17642 = n17640 | n17641 ;
  assign n17644 = ( x124 & ~n17643 ) | ( x124 & n17642 ) | ( ~n17643 & n17642 ) ;
  assign n17645 = n3605 | n9349 ;
  assign n17646 = ~n17644 & n17645 ;
  assign n17647 = x38 &  n17646 ;
  assign n17648 = x38 | n17646 ;
  assign n17649 = ~n17647 & n17648 ;
  assign n17650 = ( n17479 & n17639 ) | ( n17479 & n17649 ) | ( n17639 & n17649 ) ;
  assign n17651 = ( n17639 & ~n17479 ) | ( n17639 & n17649 ) | ( ~n17479 & n17649 ) ;
  assign n17652 = ( n17479 & ~n17650 ) | ( n17479 & n17651 ) | ( ~n17650 & n17651 ) ;
  assign n17528 = ( n17480 & n17482 ) | ( n17480 & n17495 ) | ( n17482 & n17495 ) ;
  assign n17653 = ( n17527 & ~n17652 ) | ( n17527 & n17528 ) | ( ~n17652 & n17528 ) ;
  assign n17654 = ( n17527 & ~n17528 ) | ( n17527 & n17652 ) | ( ~n17528 & n17652 ) ;
  assign n17655 = ( n17653 & ~n17527 ) | ( n17653 & n17654 ) | ( ~n17527 & n17654 ) ;
  assign n17521 = ( n17362 & ~n17513 ) | ( n17362 & n17366 ) | ( ~n17513 & n17366 ) ;
  assign n17656 = ( n17520 & ~n17655 ) | ( n17520 & n17521 ) | ( ~n17655 & n17521 ) ;
  assign n17657 = ( n17520 & ~n17521 ) | ( n17520 & n17655 ) | ( ~n17521 & n17655 ) ;
  assign n17658 = ( n17656 & ~n17520 ) | ( n17656 & n17657 ) | ( ~n17520 & n17657 ) ;
  assign n17662 = x125 &  n3756 ;
  assign n17659 = ( x127 & ~n3602 ) | ( x127 & 1'b0 ) | ( ~n3602 & 1'b0 ) ;
  assign n17660 = x126 &  n3597 ;
  assign n17661 = n17659 | n17660 ;
  assign n17663 = ( x125 & ~n17662 ) | ( x125 & n17661 ) | ( ~n17662 & n17661 ) ;
  assign n17664 = n3605 | n9941 ;
  assign n17665 = ~n17663 & n17664 ;
  assign n17666 = x38 &  n17665 ;
  assign n17667 = x38 | n17665 ;
  assign n17668 = ~n17666 & n17667 ;
  assign n17672 = x122 &  n4344 ;
  assign n17669 = ( x124 & ~n4143 ) | ( x124 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n17670 = x123 &  n4138 ;
  assign n17671 = n17669 | n17670 ;
  assign n17673 = ( x122 & ~n17672 ) | ( x122 & n17671 ) | ( ~n17672 & n17671 ) ;
  assign n17674 = ~n4146 & n8755 ;
  assign n17675 = n17673 | n17674 ;
  assign n17676 = ( x41 & ~n17675 ) | ( x41 & 1'b0 ) | ( ~n17675 & 1'b0 ) ;
  assign n17677 = ~x41 & n17675 ;
  assign n17678 = n17676 | n17677 ;
  assign n17682 = x119 &  n4934 ;
  assign n17679 = ( x121 & ~n4725 ) | ( x121 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n17680 = x120 &  n4720 ;
  assign n17681 = n17679 | n17680 ;
  assign n17683 = ( x119 & ~n17682 ) | ( x119 & n17681 ) | ( ~n17682 & n17681 ) ;
  assign n17684 = ~n4728 & n8176 ;
  assign n17685 = n17683 | n17684 ;
  assign n17686 = ( x44 & ~n17685 ) | ( x44 & 1'b0 ) | ( ~n17685 & 1'b0 ) ;
  assign n17687 = ~x44 & n17685 ;
  assign n17688 = n17686 | n17687 ;
  assign n17692 = x116 &  n5586 ;
  assign n17689 = ( x118 & ~n5389 ) | ( x118 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n17690 = x117 &  n5384 ;
  assign n17691 = n17689 | n17690 ;
  assign n17693 = ( x116 & ~n17692 ) | ( x116 & n17691 ) | ( ~n17692 & n17691 ) ;
  assign n17694 = n5392 | n7152 ;
  assign n17695 = ~n17693 & n17694 ;
  assign n17696 = x47 &  n17695 ;
  assign n17697 = x47 | n17695 ;
  assign n17698 = ~n17696 & n17697 ;
  assign n17702 = x110 &  n6982 ;
  assign n17699 = ( x112 & ~n6727 ) | ( x112 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n17700 = x111 &  n6722 ;
  assign n17701 = n17699 | n17700 ;
  assign n17703 = ( x110 & ~n17702 ) | ( x110 & n17701 ) | ( ~n17702 & n17701 ) ;
  assign n17704 = ( n5727 & ~n6730 ) | ( n5727 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n17705 = n17703 | n17704 ;
  assign n17706 = ( x53 & ~n17705 ) | ( x53 & 1'b0 ) | ( ~n17705 & 1'b0 ) ;
  assign n17707 = ~x53 & n17705 ;
  assign n17708 = n17706 | n17707 ;
  assign n17757 = ( n17593 & ~n17423 ) | ( n17593 & n17603 ) | ( ~n17423 & n17603 ) ;
  assign n17712 = x107 &  n7731 ;
  assign n17709 = ( x109 & ~n7538 ) | ( x109 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n17710 = x108 &  n7533 ;
  assign n17711 = n17709 | n17710 ;
  assign n17713 = ( x107 & ~n17712 ) | ( x107 & n17711 ) | ( ~n17712 & n17711 ) ;
  assign n17714 = ( n5267 & ~n7541 ) | ( n5267 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n17715 = n17713 | n17714 ;
  assign n17716 = ( x56 & ~n17715 ) | ( x56 & 1'b0 ) | ( ~n17715 & 1'b0 ) ;
  assign n17717 = ~x56 & n17715 ;
  assign n17718 = n17716 | n17717 ;
  assign n17753 = ( n17420 & n17561 ) | ( n17420 & n17590 ) | ( n17561 & n17590 ) ;
  assign n17722 = x104 &  n8558 ;
  assign n17719 = ( x106 & ~n8314 ) | ( x106 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n17720 = x105 &  n8309 ;
  assign n17721 = n17719 | n17720 ;
  assign n17723 = ( x104 & ~n17722 ) | ( x104 & n17721 ) | ( ~n17722 & n17721 ) ;
  assign n17724 = ( n4458 & ~n8317 ) | ( n4458 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n17725 = n17723 | n17724 ;
  assign n17726 = ( x59 & ~n17725 ) | ( x59 & 1'b0 ) | ( ~n17725 & 1'b0 ) ;
  assign n17727 = ~x59 & n17725 ;
  assign n17728 = n17726 | n17727 ;
  assign n17729 = x99 &  n10104 ;
  assign n17730 = ( x100 & ~n9760 ) | ( x100 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n17731 = n17729 | n17730 ;
  assign n17732 = ( x35 & n17574 ) | ( x35 & n17731 ) | ( n17574 & n17731 ) ;
  assign n17733 = ( x35 & ~n17574 ) | ( x35 & n17731 ) | ( ~n17574 & n17731 ) ;
  assign n17734 = ( n17574 & ~n17732 ) | ( n17574 & n17733 ) | ( ~n17732 & n17733 ) ;
  assign n17739 = x101 &  n9457 ;
  assign n17736 = ( x103 & ~n9150 ) | ( x103 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n17737 = x102 &  n9145 ;
  assign n17738 = n17736 | n17737 ;
  assign n17740 = ( x101 & ~n17739 ) | ( x101 & n17738 ) | ( ~n17739 & n17738 ) ;
  assign n17741 = n4056 | n9153 ;
  assign n17742 = ~n17740 & n17741 ;
  assign n17743 = x62 &  n17742 ;
  assign n17744 = x62 | n17742 ;
  assign n17745 = ~n17743 & n17744 ;
  assign n17735 = ( n17416 & ~n17405 ) | ( n17416 & n17574 ) | ( ~n17405 & n17574 ) ;
  assign n17746 = ( n17734 & ~n17745 ) | ( n17734 & n17735 ) | ( ~n17745 & n17735 ) ;
  assign n17747 = ( n17734 & ~n17735 ) | ( n17734 & n17745 ) | ( ~n17735 & n17745 ) ;
  assign n17748 = ( n17746 & ~n17734 ) | ( n17746 & n17747 ) | ( ~n17734 & n17747 ) ;
  assign n17749 = ( n17577 & ~n17571 ) | ( n17577 & n17587 ) | ( ~n17571 & n17587 ) ;
  assign n17750 = ( n17728 & ~n17748 ) | ( n17728 & n17749 ) | ( ~n17748 & n17749 ) ;
  assign n17751 = ( n17728 & ~n17749 ) | ( n17728 & n17748 ) | ( ~n17749 & n17748 ) ;
  assign n17752 = ( n17750 & ~n17728 ) | ( n17750 & n17751 ) | ( ~n17728 & n17751 ) ;
  assign n17754 = ( n17718 & ~n17753 ) | ( n17718 & n17752 ) | ( ~n17753 & n17752 ) ;
  assign n17755 = ( n17718 & ~n17752 ) | ( n17718 & n17753 ) | ( ~n17752 & n17753 ) ;
  assign n17756 = ( n17754 & ~n17718 ) | ( n17754 & n17755 ) | ( ~n17718 & n17755 ) ;
  assign n17758 = ( n17708 & ~n17757 ) | ( n17708 & n17756 ) | ( ~n17757 & n17756 ) ;
  assign n17759 = ( n17708 & ~n17756 ) | ( n17708 & n17757 ) | ( ~n17756 & n17757 ) ;
  assign n17760 = ( n17758 & ~n17708 ) | ( n17758 & n17759 ) | ( ~n17708 & n17759 ) ;
  assign n17761 = ( n17551 & ~n17606 ) | ( n17551 & n17616 ) | ( ~n17606 & n17616 ) ;
  assign n17765 = x113 &  n6288 ;
  assign n17762 = ( x115 & ~n6032 ) | ( x115 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n17763 = x114 &  n6027 ;
  assign n17764 = n17762 | n17763 ;
  assign n17766 = ( x113 & ~n17765 ) | ( x113 & n17764 ) | ( ~n17765 & n17764 ) ;
  assign n17767 = ~n6035 & n6420 ;
  assign n17768 = n17766 | n17767 ;
  assign n17769 = ( x50 & ~n17768 ) | ( x50 & 1'b0 ) | ( ~n17768 & 1'b0 ) ;
  assign n17770 = ~x50 & n17768 ;
  assign n17771 = n17769 | n17770 ;
  assign n17772 = ( n17760 & n17761 ) | ( n17760 & n17771 ) | ( n17761 & n17771 ) ;
  assign n17773 = ( n17761 & ~n17760 ) | ( n17761 & n17771 ) | ( ~n17760 & n17771 ) ;
  assign n17774 = ( n17760 & ~n17772 ) | ( n17760 & n17773 ) | ( ~n17772 & n17773 ) ;
  assign n17775 = ( n17621 & n17698 ) | ( n17621 & n17774 ) | ( n17698 & n17774 ) ;
  assign n17776 = ( n17621 & ~n17698 ) | ( n17621 & n17774 ) | ( ~n17698 & n17774 ) ;
  assign n17777 = ( n17698 & ~n17775 ) | ( n17698 & n17776 ) | ( ~n17775 & n17776 ) ;
  assign n17779 = ( n17624 & n17688 ) | ( n17624 & n17777 ) | ( n17688 & n17777 ) ;
  assign n17778 = ( n17624 & ~n17688 ) | ( n17624 & n17777 ) | ( ~n17688 & n17777 ) ;
  assign n17780 = ( n17688 & ~n17779 ) | ( n17688 & n17778 ) | ( ~n17779 & n17778 ) ;
  assign n17781 = ( n17625 & n17626 ) | ( n17625 & n17636 ) | ( n17626 & n17636 ) ;
  assign n17782 = ( n17678 & n17780 ) | ( n17678 & n17781 ) | ( n17780 & n17781 ) ;
  assign n17783 = ( n17780 & ~n17678 ) | ( n17780 & n17781 ) | ( ~n17678 & n17781 ) ;
  assign n17784 = ( n17678 & ~n17782 ) | ( n17678 & n17783 ) | ( ~n17782 & n17783 ) ;
  assign n17785 = ( n17479 & ~n17639 ) | ( n17479 & n17649 ) | ( ~n17639 & n17649 ) ;
  assign n17786 = ( n17668 & ~n17784 ) | ( n17668 & n17785 ) | ( ~n17784 & n17785 ) ;
  assign n17787 = ( n17668 & ~n17785 ) | ( n17668 & n17784 ) | ( ~n17785 & n17784 ) ;
  assign n17788 = ( n17786 & ~n17668 ) | ( n17786 & n17787 ) | ( ~n17668 & n17787 ) ;
  assign n17789 = ( n17521 & ~n17520 ) | ( n17521 & n17655 ) | ( ~n17520 & n17655 ) ;
  assign n17790 = ( n17528 & ~n17527 ) | ( n17528 & n17652 ) | ( ~n17527 & n17652 ) ;
  assign n17792 = ( n17788 & n17789 ) | ( n17788 & n17790 ) | ( n17789 & n17790 ) ;
  assign n17791 = ( n17789 & ~n17788 ) | ( n17789 & n17790 ) | ( ~n17788 & n17790 ) ;
  assign n17793 = ( n17788 & ~n17792 ) | ( n17788 & n17791 ) | ( ~n17792 & n17791 ) ;
  assign n17794 = ( n17760 & ~n17771 ) | ( n17760 & n17761 ) | ( ~n17771 & n17761 ) ;
  assign n17795 = ( n17752 & ~n17718 ) | ( n17752 & n17753 ) | ( ~n17718 & n17753 ) ;
  assign n17830 = x108 &  n7731 ;
  assign n17827 = ( x110 & ~n7538 ) | ( x110 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n17828 = x109 &  n7533 ;
  assign n17829 = n17827 | n17828 ;
  assign n17831 = ( x108 & ~n17830 ) | ( x108 & n17829 ) | ( ~n17830 & n17829 ) ;
  assign n17832 = n5283 | n7541 ;
  assign n17833 = ~n17831 & n17832 ;
  assign n17834 = x56 &  n17833 ;
  assign n17835 = x56 | n17833 ;
  assign n17836 = ~n17834 & n17835 ;
  assign n17807 = x100 &  n10104 ;
  assign n17808 = ( x101 & ~n9760 ) | ( x101 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n17809 = n17807 | n17808 ;
  assign n17796 = ( n17574 & ~x35 ) | ( n17574 & n17731 ) | ( ~x35 & n17731 ) ;
  assign n17800 = x102 &  n9457 ;
  assign n17797 = ( x104 & ~n9150 ) | ( x104 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n17798 = x103 &  n9145 ;
  assign n17799 = n17797 | n17798 ;
  assign n17801 = ( x102 & ~n17800 ) | ( x102 & n17799 ) | ( ~n17800 & n17799 ) ;
  assign n17802 = n4249 | n9153 ;
  assign n17803 = ~n17801 & n17802 ;
  assign n17804 = x62 &  n17803 ;
  assign n17805 = x62 | n17803 ;
  assign n17806 = ~n17804 & n17805 ;
  assign n17810 = ( n17796 & n17806 ) | ( n17796 & n17809 ) | ( n17806 & n17809 ) ;
  assign n17811 = ( n17796 & ~n17809 ) | ( n17796 & n17806 ) | ( ~n17809 & n17806 ) ;
  assign n17812 = ( n17809 & ~n17810 ) | ( n17809 & n17811 ) | ( ~n17810 & n17811 ) ;
  assign n17813 = ( n17734 & n17735 ) | ( n17734 & n17745 ) | ( n17735 & n17745 ) ;
  assign n17814 = ~n17812 & n17813 ;
  assign n17815 = ( n17812 & ~n17813 ) | ( n17812 & 1'b0 ) | ( ~n17813 & 1'b0 ) ;
  assign n17816 = n17814 | n17815 ;
  assign n17820 = x105 &  n8558 ;
  assign n17817 = ( x107 & ~n8314 ) | ( x107 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n17818 = x106 &  n8309 ;
  assign n17819 = n17817 | n17818 ;
  assign n17821 = ( x105 & ~n17820 ) | ( x105 & n17819 ) | ( ~n17820 & n17819 ) ;
  assign n17822 = ( n4848 & ~n8317 ) | ( n4848 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n17823 = n17821 | n17822 ;
  assign n17824 = ( n17816 & ~x59 ) | ( n17816 & n17823 ) | ( ~x59 & n17823 ) ;
  assign n17825 = ( x59 & ~n17816 ) | ( x59 & n17823 ) | ( ~n17816 & n17823 ) ;
  assign n17826 = ( n17824 & ~n17823 ) | ( n17824 & n17825 ) | ( ~n17823 & n17825 ) ;
  assign n17837 = ( n17750 & ~n17836 ) | ( n17750 & n17826 ) | ( ~n17836 & n17826 ) ;
  assign n17838 = ( n17750 & ~n17826 ) | ( n17750 & n17836 ) | ( ~n17826 & n17836 ) ;
  assign n17839 = ( n17837 & ~n17750 ) | ( n17837 & n17838 ) | ( ~n17750 & n17838 ) ;
  assign n17843 = x111 &  n6982 ;
  assign n17840 = ( x113 & ~n6727 ) | ( x113 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n17841 = x112 &  n6722 ;
  assign n17842 = n17840 | n17841 ;
  assign n17844 = ( x111 & ~n17843 ) | ( x111 & n17842 ) | ( ~n17843 & n17842 ) ;
  assign n17845 = n6169 | n6730 ;
  assign n17846 = ~n17844 & n17845 ;
  assign n17847 = x53 &  n17846 ;
  assign n17848 = x53 | n17846 ;
  assign n17849 = ~n17847 & n17848 ;
  assign n17850 = ( n17795 & n17839 ) | ( n17795 & n17849 ) | ( n17839 & n17849 ) ;
  assign n17851 = ( n17839 & ~n17795 ) | ( n17839 & n17849 ) | ( ~n17795 & n17849 ) ;
  assign n17852 = ( n17795 & ~n17850 ) | ( n17795 & n17851 ) | ( ~n17850 & n17851 ) ;
  assign n17856 = x114 &  n6288 ;
  assign n17853 = ( x116 & ~n6032 ) | ( x116 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n17854 = x115 &  n6027 ;
  assign n17855 = n17853 | n17854 ;
  assign n17857 = ( x114 & ~n17856 ) | ( x114 & n17855 ) | ( ~n17856 & n17855 ) ;
  assign n17858 = n6035 | n6885 ;
  assign n17859 = ~n17857 & n17858 ;
  assign n17860 = x50 &  n17859 ;
  assign n17861 = x50 | n17859 ;
  assign n17862 = ~n17860 & n17861 ;
  assign n17864 = ( n17758 & n17852 ) | ( n17758 & n17862 ) | ( n17852 & n17862 ) ;
  assign n17863 = ( n17852 & ~n17758 ) | ( n17852 & n17862 ) | ( ~n17758 & n17862 ) ;
  assign n17865 = ( n17758 & ~n17864 ) | ( n17758 & n17863 ) | ( ~n17864 & n17863 ) ;
  assign n17869 = x117 &  n5586 ;
  assign n17866 = ( x119 & ~n5389 ) | ( x119 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n17867 = x118 &  n5384 ;
  assign n17868 = n17866 | n17867 ;
  assign n17870 = ( x117 & ~n17869 ) | ( x117 & n17868 ) | ( ~n17869 & n17868 ) ;
  assign n17871 = ~n5392 & n7648 ;
  assign n17872 = n17870 | n17871 ;
  assign n17874 = x47 &  n17872 ;
  assign n17873 = ~x47 & n17872 ;
  assign n17875 = ( x47 & ~n17874 ) | ( x47 & n17873 ) | ( ~n17874 & n17873 ) ;
  assign n17877 = ( n17794 & n17865 ) | ( n17794 & n17875 ) | ( n17865 & n17875 ) ;
  assign n17876 = ( n17865 & ~n17794 ) | ( n17865 & n17875 ) | ( ~n17794 & n17875 ) ;
  assign n17878 = ( n17794 & ~n17877 ) | ( n17794 & n17876 ) | ( ~n17877 & n17876 ) ;
  assign n17882 = x120 &  n4934 ;
  assign n17879 = ( x122 & ~n4725 ) | ( x122 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n17880 = x121 &  n4720 ;
  assign n17881 = n17879 | n17880 ;
  assign n17883 = ( x120 & ~n17882 ) | ( x120 & n17881 ) | ( ~n17882 & n17881 ) ;
  assign n17884 = ~n4728 & n9987 ;
  assign n17885 = n17883 | n17884 ;
  assign n17886 = ( x44 & ~n17885 ) | ( x44 & 1'b0 ) | ( ~n17885 & 1'b0 ) ;
  assign n17887 = ~x44 & n17885 ;
  assign n17888 = n17886 | n17887 ;
  assign n17889 = ( n17776 & ~n17878 ) | ( n17776 & n17888 ) | ( ~n17878 & n17888 ) ;
  assign n17890 = ( n17776 & ~n17888 ) | ( n17776 & n17878 ) | ( ~n17888 & n17878 ) ;
  assign n17891 = ( n17889 & ~n17776 ) | ( n17889 & n17890 ) | ( ~n17776 & n17890 ) ;
  assign n17892 = n17778 | n17891 ;
  assign n17893 = n17778 &  n17891 ;
  assign n17894 = ( n17892 & ~n17893 ) | ( n17892 & 1'b0 ) | ( ~n17893 & 1'b0 ) ;
  assign n17895 = ( x126 & ~n3756 ) | ( x126 & 1'b0 ) | ( ~n3756 & 1'b0 ) ;
  assign n17896 = x127 &  n3597 ;
  assign n17897 = n17895 | n17896 ;
  assign n17898 = n3605 | n9960 ;
  assign n17899 = ( n17897 & ~n3605 ) | ( n17897 & n17898 ) | ( ~n3605 & n17898 ) ;
  assign n17903 = ( n17782 & ~x38 ) | ( n17782 & n17899 ) | ( ~x38 & n17899 ) ;
  assign n17904 = ( x38 & ~n17899 ) | ( x38 & n17782 ) | ( ~n17899 & n17782 ) ;
  assign n17905 = ( n17903 & ~n17782 ) | ( n17903 & n17904 ) | ( ~n17782 & n17904 ) ;
  assign n17909 = x123 &  n4344 ;
  assign n17906 = ( x125 & ~n4143 ) | ( x125 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n17907 = x124 &  n4138 ;
  assign n17908 = n17906 | n17907 ;
  assign n17910 = ( x123 & ~n17909 ) | ( x123 & n17908 ) | ( ~n17909 & n17908 ) ;
  assign n17911 = ~n4146 & n9324 ;
  assign n17912 = n17910 | n17911 ;
  assign n17913 = ( x41 & ~n17912 ) | ( x41 & 1'b0 ) | ( ~n17912 & 1'b0 ) ;
  assign n17914 = ~x41 & n17912 ;
  assign n17915 = n17913 | n17914 ;
  assign n17916 = ( n17894 & ~n17905 ) | ( n17894 & n17915 ) | ( ~n17905 & n17915 ) ;
  assign n17917 = ( n17894 & ~n17915 ) | ( n17894 & n17905 ) | ( ~n17915 & n17905 ) ;
  assign n17918 = ( n17916 & ~n17894 ) | ( n17916 & n17917 ) | ( ~n17894 & n17917 ) ;
  assign n17919 = ( n17788 & ~n17789 ) | ( n17788 & n17790 ) | ( ~n17789 & n17790 ) ;
  assign n17921 = ( n17786 & n17918 ) | ( n17786 & n17919 ) | ( n17918 & n17919 ) ;
  assign n17920 = ( n17918 & ~n17786 ) | ( n17918 & n17919 ) | ( ~n17786 & n17919 ) ;
  assign n17922 = ( n17786 & ~n17921 ) | ( n17786 & n17920 ) | ( ~n17921 & n17920 ) ;
  assign n17923 = ~n17894 & n17915 ;
  assign n17924 = ( n17894 & ~n17915 ) | ( n17894 & 1'b0 ) | ( ~n17915 & 1'b0 ) ;
  assign n17925 = n17923 | n17924 ;
  assign n17900 = x38 | n17899 ;
  assign n17901 = ( x38 & ~n17899 ) | ( x38 & 1'b0 ) | ( ~n17899 & 1'b0 ) ;
  assign n17902 = ( n17900 & ~x38 ) | ( n17900 & n17901 ) | ( ~x38 & n17901 ) ;
  assign n17926 = ( n17782 & ~n17925 ) | ( n17782 & n17902 ) | ( ~n17925 & n17902 ) ;
  assign n17928 = ( x127 & ~n3756 ) | ( x127 & 1'b0 ) | ( ~n3756 & 1'b0 ) ;
  assign n17929 = n3605 | n10258 ;
  assign n17930 = ~n17928 & n17929 ;
  assign n17931 = ~x38 & n17930 ;
  assign n17932 = ( x38 & ~n17930 ) | ( x38 & 1'b0 ) | ( ~n17930 & 1'b0 ) ;
  assign n17933 = n17931 | n17932 ;
  assign n17935 = ( n17776 & n17878 ) | ( n17776 & n17888 ) | ( n17878 & n17888 ) ;
  assign n18041 = x124 &  n4344 ;
  assign n18038 = ( x126 & ~n4143 ) | ( x126 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n18039 = x125 &  n4138 ;
  assign n18040 = n18038 | n18039 ;
  assign n18042 = ( x124 & ~n18041 ) | ( x124 & n18040 ) | ( ~n18041 & n18040 ) ;
  assign n18043 = n4146 | n9349 ;
  assign n18044 = ~n18042 & n18043 ;
  assign n18045 = x41 &  n18044 ;
  assign n18046 = x41 | n18044 ;
  assign n18047 = ~n18045 & n18046 ;
  assign n17936 = ( n17758 & ~n17862 ) | ( n17758 & n17852 ) | ( ~n17862 & n17852 ) ;
  assign n17940 = x118 &  n5586 ;
  assign n17937 = ( x120 & ~n5389 ) | ( x120 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n17938 = x119 &  n5384 ;
  assign n17939 = n17937 | n17938 ;
  assign n17941 = ( x118 & ~n17940 ) | ( x118 & n17939 ) | ( ~n17940 & n17939 ) ;
  assign n17942 = ~n5392 & n9364 ;
  assign n17943 = n17941 | n17942 ;
  assign n17944 = ( x47 & ~n17943 ) | ( x47 & 1'b0 ) | ( ~n17943 & 1'b0 ) ;
  assign n17945 = ~x47 & n17943 ;
  assign n17946 = n17944 | n17945 ;
  assign n17947 = ( n17795 & ~n17839 ) | ( n17795 & n17849 ) | ( ~n17839 & n17849 ) ;
  assign n17951 = x115 &  n6288 ;
  assign n17948 = ( x117 & ~n6032 ) | ( x117 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n17949 = x116 &  n6027 ;
  assign n17950 = n17948 | n17949 ;
  assign n17952 = ( x115 & ~n17951 ) | ( x115 & n17950 ) | ( ~n17951 & n17950 ) ;
  assign n17953 = n6035 | n7136 ;
  assign n17954 = ~n17952 & n17953 ;
  assign n17955 = x50 &  n17954 ;
  assign n17956 = x50 | n17954 ;
  assign n17957 = ~n17955 & n17956 ;
  assign n17958 = ( n17826 & ~n17750 ) | ( n17826 & n17836 ) | ( ~n17750 & n17836 ) ;
  assign n17960 = ( x59 & n17814 ) | ( x59 & n17823 ) | ( n17814 & n17823 ) ;
  assign n17959 = x59 | n17823 ;
  assign n17961 = ( n17815 & ~n17960 ) | ( n17815 & n17959 ) | ( ~n17960 & n17959 ) ;
  assign n17995 = x109 &  n7731 ;
  assign n17992 = ( x111 & ~n7538 ) | ( x111 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n17993 = x110 &  n7533 ;
  assign n17994 = n17992 | n17993 ;
  assign n17996 = ( x109 & ~n17995 ) | ( x109 & n17994 ) | ( ~n17995 & n17994 ) ;
  assign n17997 = n5711 | n7541 ;
  assign n17998 = ~n17996 & n17997 ;
  assign n17999 = x56 &  n17998 ;
  assign n18000 = x56 | n17998 ;
  assign n18001 = ~n17999 & n18000 ;
  assign n17965 = x103 &  n9457 ;
  assign n17962 = ( x105 & ~n9150 ) | ( x105 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n17963 = x104 &  n9145 ;
  assign n17964 = n17962 | n17963 ;
  assign n17966 = ( x103 & ~n17965 ) | ( x103 & n17964 ) | ( ~n17965 & n17964 ) ;
  assign n17967 = ( n4442 & ~n9153 ) | ( n4442 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n17968 = n17966 | n17967 ;
  assign n17969 = ( x62 & ~n17968 ) | ( x62 & 1'b0 ) | ( ~n17968 & 1'b0 ) ;
  assign n17970 = ~x62 & n17968 ;
  assign n17971 = n17969 | n17970 ;
  assign n17973 = x101 &  n10104 ;
  assign n17974 = ( x102 & ~n9760 ) | ( x102 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n17975 = n17973 | n17974 ;
  assign n17972 = ( n17806 & ~n17796 ) | ( n17806 & n17809 ) | ( ~n17796 & n17809 ) ;
  assign n17976 = ( n17809 & ~n17975 ) | ( n17809 & n17972 ) | ( ~n17975 & n17972 ) ;
  assign n17977 = ( n17972 & ~n17809 ) | ( n17972 & n17975 ) | ( ~n17809 & n17975 ) ;
  assign n17978 = ( n17976 & ~n17972 ) | ( n17976 & n17977 ) | ( ~n17972 & n17977 ) ;
  assign n17982 = x106 &  n8558 ;
  assign n17979 = ( x108 & ~n8314 ) | ( x108 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n17980 = x107 &  n8309 ;
  assign n17981 = n17979 | n17980 ;
  assign n17983 = ( x106 & ~n17982 ) | ( x106 & n17981 ) | ( ~n17982 & n17981 ) ;
  assign n17984 = n5055 | n8317 ;
  assign n17985 = ~n17983 & n17984 ;
  assign n17986 = x59 &  n17985 ;
  assign n17987 = x59 | n17985 ;
  assign n17988 = ~n17986 & n17987 ;
  assign n17990 = ( n17971 & n17978 ) | ( n17971 & n17988 ) | ( n17978 & n17988 ) ;
  assign n17989 = ( n17978 & ~n17971 ) | ( n17978 & n17988 ) | ( ~n17971 & n17988 ) ;
  assign n17991 = ( n17971 & ~n17990 ) | ( n17971 & n17989 ) | ( ~n17990 & n17989 ) ;
  assign n18002 = ( n17961 & ~n18001 ) | ( n17961 & n17991 ) | ( ~n18001 & n17991 ) ;
  assign n18003 = ( n17961 & ~n17991 ) | ( n17961 & n18001 ) | ( ~n17991 & n18001 ) ;
  assign n18004 = ( n18002 & ~n17961 ) | ( n18002 & n18003 ) | ( ~n17961 & n18003 ) ;
  assign n18008 = x112 &  n6982 ;
  assign n18005 = ( x114 & ~n6727 ) | ( x114 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n18006 = x113 &  n6722 ;
  assign n18007 = n18005 | n18006 ;
  assign n18009 = ( x112 & ~n18008 ) | ( x112 & n18007 ) | ( ~n18008 & n18007 ) ;
  assign n18010 = n6185 | n6730 ;
  assign n18011 = ~n18009 & n18010 ;
  assign n18012 = x53 &  n18011 ;
  assign n18013 = x53 | n18011 ;
  assign n18014 = ~n18012 & n18013 ;
  assign n18015 = ( n17958 & n18004 ) | ( n17958 & n18014 ) | ( n18004 & n18014 ) ;
  assign n18016 = ( n18004 & ~n17958 ) | ( n18004 & n18014 ) | ( ~n17958 & n18014 ) ;
  assign n18017 = ( n17958 & ~n18015 ) | ( n17958 & n18016 ) | ( ~n18015 & n18016 ) ;
  assign n18018 = ( n17947 & ~n17957 ) | ( n17947 & n18017 ) | ( ~n17957 & n18017 ) ;
  assign n18019 = ( n17947 & ~n18017 ) | ( n17947 & n17957 ) | ( ~n18017 & n17957 ) ;
  assign n18020 = ( n18018 & ~n17947 ) | ( n18018 & n18019 ) | ( ~n17947 & n18019 ) ;
  assign n18022 = ( n17936 & n17946 ) | ( n17936 & n18020 ) | ( n17946 & n18020 ) ;
  assign n18021 = ( n17946 & ~n17936 ) | ( n17946 & n18020 ) | ( ~n17936 & n18020 ) ;
  assign n18023 = ( n17936 & ~n18022 ) | ( n17936 & n18021 ) | ( ~n18022 & n18021 ) ;
  assign n18024 = ( n17794 & ~n17875 ) | ( n17794 & n17865 ) | ( ~n17875 & n17865 ) ;
  assign n18028 = x121 &  n4934 ;
  assign n18025 = ( x123 & ~n4725 ) | ( x123 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n18026 = x122 &  n4720 ;
  assign n18027 = n18025 | n18026 ;
  assign n18029 = ( x121 & ~n18028 ) | ( x121 & n18027 ) | ( ~n18028 & n18027 ) ;
  assign n18030 = ~n4728 & n8472 ;
  assign n18031 = n18029 | n18030 ;
  assign n18032 = ( x44 & ~n18031 ) | ( x44 & 1'b0 ) | ( ~n18031 & 1'b0 ) ;
  assign n18033 = ~x44 & n18031 ;
  assign n18034 = n18032 | n18033 ;
  assign n18036 = ( n18023 & n18024 ) | ( n18023 & n18034 ) | ( n18024 & n18034 ) ;
  assign n18035 = ( n18024 & ~n18023 ) | ( n18024 & n18034 ) | ( ~n18023 & n18034 ) ;
  assign n18037 = ( n18023 & ~n18036 ) | ( n18023 & n18035 ) | ( ~n18036 & n18035 ) ;
  assign n18048 = ( n17935 & ~n18047 ) | ( n17935 & n18037 ) | ( ~n18047 & n18037 ) ;
  assign n18049 = ( n17935 & ~n18037 ) | ( n17935 & n18047 ) | ( ~n18037 & n18047 ) ;
  assign n18050 = ( n18048 & ~n17935 ) | ( n18048 & n18049 ) | ( ~n17935 & n18049 ) ;
  assign n17934 = ( n17891 & ~n17778 ) | ( n17891 & n17915 ) | ( ~n17778 & n17915 ) ;
  assign n18051 = ( n17933 & ~n18050 ) | ( n17933 & n17934 ) | ( ~n18050 & n17934 ) ;
  assign n18052 = ( n17933 & ~n17934 ) | ( n17933 & n18050 ) | ( ~n17934 & n18050 ) ;
  assign n18053 = ( n18051 & ~n17933 ) | ( n18051 & n18052 ) | ( ~n17933 & n18052 ) ;
  assign n17927 = ( n17786 & ~n17919 ) | ( n17786 & n17918 ) | ( ~n17919 & n17918 ) ;
  assign n18054 = ( n17926 & ~n18053 ) | ( n17926 & n17927 ) | ( ~n18053 & n17927 ) ;
  assign n18055 = ( n17926 & ~n17927 ) | ( n17926 & n18053 ) | ( ~n17927 & n18053 ) ;
  assign n18056 = ( n18054 & ~n17926 ) | ( n18054 & n18055 ) | ( ~n17926 & n18055 ) ;
  assign n18060 = x125 &  n4344 ;
  assign n18057 = ( x127 & ~n4143 ) | ( x127 & 1'b0 ) | ( ~n4143 & 1'b0 ) ;
  assign n18058 = x126 &  n4138 ;
  assign n18059 = n18057 | n18058 ;
  assign n18061 = ( x125 & ~n18060 ) | ( x125 & n18059 ) | ( ~n18060 & n18059 ) ;
  assign n18062 = n4146 | n9941 ;
  assign n18063 = ~n18061 & n18062 ;
  assign n18064 = x41 &  n18063 ;
  assign n18065 = x41 | n18063 ;
  assign n18066 = ~n18064 & n18065 ;
  assign n18070 = x122 &  n4934 ;
  assign n18067 = ( x124 & ~n4725 ) | ( x124 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n18068 = x123 &  n4720 ;
  assign n18069 = n18067 | n18068 ;
  assign n18071 = ( x122 & ~n18070 ) | ( x122 & n18069 ) | ( ~n18070 & n18069 ) ;
  assign n18072 = ~n4728 & n8755 ;
  assign n18073 = n18071 | n18072 ;
  assign n18074 = ( x44 & ~n18073 ) | ( x44 & 1'b0 ) | ( ~n18073 & 1'b0 ) ;
  assign n18075 = ~x44 & n18073 ;
  assign n18076 = n18074 | n18075 ;
  assign n18080 = x119 &  n5586 ;
  assign n18077 = ( x121 & ~n5389 ) | ( x121 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n18078 = x120 &  n5384 ;
  assign n18079 = n18077 | n18078 ;
  assign n18081 = ( x119 & ~n18080 ) | ( x119 & n18079 ) | ( ~n18080 & n18079 ) ;
  assign n18082 = ~n5392 & n8176 ;
  assign n18083 = n18081 | n18082 ;
  assign n18084 = ( x47 & ~n18083 ) | ( x47 & 1'b0 ) | ( ~n18083 & 1'b0 ) ;
  assign n18085 = ~x47 & n18083 ;
  assign n18086 = n18084 | n18085 ;
  assign n18090 = x116 &  n6288 ;
  assign n18087 = ( x118 & ~n6032 ) | ( x118 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n18088 = x117 &  n6027 ;
  assign n18089 = n18087 | n18088 ;
  assign n18091 = ( x116 & ~n18090 ) | ( x116 & n18089 ) | ( ~n18090 & n18089 ) ;
  assign n18092 = n6035 | n7152 ;
  assign n18093 = ~n18091 & n18092 ;
  assign n18094 = x50 &  n18093 ;
  assign n18095 = x50 | n18093 ;
  assign n18096 = ~n18094 & n18095 ;
  assign n18100 = x110 &  n7731 ;
  assign n18097 = ( x112 & ~n7538 ) | ( x112 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n18098 = x111 &  n7533 ;
  assign n18099 = n18097 | n18098 ;
  assign n18101 = ( x110 & ~n18100 ) | ( x110 & n18099 ) | ( ~n18100 & n18099 ) ;
  assign n18102 = ( n5727 & ~n7541 ) | ( n5727 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n18103 = n18101 | n18102 ;
  assign n18104 = ( x56 & ~n18103 ) | ( x56 & 1'b0 ) | ( ~n18103 & 1'b0 ) ;
  assign n18105 = ~x56 & n18103 ;
  assign n18106 = n18104 | n18105 ;
  assign n18110 = x107 &  n8558 ;
  assign n18107 = ( x109 & ~n8314 ) | ( x109 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n18108 = x108 &  n8309 ;
  assign n18109 = n18107 | n18108 ;
  assign n18111 = ( x107 & ~n18110 ) | ( x107 & n18109 ) | ( ~n18110 & n18109 ) ;
  assign n18112 = ( n5267 & ~n8317 ) | ( n5267 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n18113 = n18111 | n18112 ;
  assign n18114 = ( x59 & ~n18113 ) | ( x59 & 1'b0 ) | ( ~n18113 & 1'b0 ) ;
  assign n18115 = ~x59 & n18113 ;
  assign n18116 = n18114 | n18115 ;
  assign n18117 = x102 &  n10104 ;
  assign n18118 = ( x103 & ~n9760 ) | ( x103 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n18119 = n18117 | n18118 ;
  assign n18120 = ( x38 & n17809 ) | ( x38 & n18119 ) | ( n17809 & n18119 ) ;
  assign n18121 = ( x38 & ~n17809 ) | ( x38 & n18119 ) | ( ~n17809 & n18119 ) ;
  assign n18122 = ( n17809 & ~n18120 ) | ( n17809 & n18121 ) | ( ~n18120 & n18121 ) ;
  assign n18126 = x104 &  n9457 ;
  assign n18123 = ( x106 & ~n9150 ) | ( x106 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n18124 = x105 &  n9145 ;
  assign n18125 = n18123 | n18124 ;
  assign n18127 = ( x104 & ~n18126 ) | ( x104 & n18125 ) | ( ~n18126 & n18125 ) ;
  assign n18128 = ( n4458 & ~n9153 ) | ( n4458 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n18129 = n18127 | n18128 ;
  assign n18130 = ( x62 & ~n18129 ) | ( x62 & 1'b0 ) | ( ~n18129 & 1'b0 ) ;
  assign n18131 = ~x62 & n18129 ;
  assign n18132 = n18130 | n18131 ;
  assign n18133 = ( n17976 & n18122 ) | ( n17976 & n18132 ) | ( n18122 & n18132 ) ;
  assign n18134 = ( n17976 & ~n18122 ) | ( n17976 & n18132 ) | ( ~n18122 & n18132 ) ;
  assign n18135 = ( n18122 & ~n18133 ) | ( n18122 & n18134 ) | ( ~n18133 & n18134 ) ;
  assign n18136 = ( n17971 & ~n17988 ) | ( n17971 & n17978 ) | ( ~n17988 & n17978 ) ;
  assign n18137 = ( n18116 & ~n18135 ) | ( n18116 & n18136 ) | ( ~n18135 & n18136 ) ;
  assign n18138 = ( n18116 & ~n18136 ) | ( n18116 & n18135 ) | ( ~n18136 & n18135 ) ;
  assign n18139 = ( n18137 & ~n18116 ) | ( n18137 & n18138 ) | ( ~n18116 & n18138 ) ;
  assign n18140 = ( n17991 & ~n17961 ) | ( n17991 & n18001 ) | ( ~n17961 & n18001 ) ;
  assign n18142 = ( n18106 & n18139 ) | ( n18106 & n18140 ) | ( n18139 & n18140 ) ;
  assign n18141 = ( n18139 & ~n18106 ) | ( n18139 & n18140 ) | ( ~n18106 & n18140 ) ;
  assign n18143 = ( n18106 & ~n18142 ) | ( n18106 & n18141 ) | ( ~n18142 & n18141 ) ;
  assign n18144 = ( n17958 & ~n18004 ) | ( n17958 & n18014 ) | ( ~n18004 & n18014 ) ;
  assign n18148 = x113 &  n6982 ;
  assign n18145 = ( x115 & ~n6727 ) | ( x115 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n18146 = x114 &  n6722 ;
  assign n18147 = n18145 | n18146 ;
  assign n18149 = ( x113 & ~n18148 ) | ( x113 & n18147 ) | ( ~n18148 & n18147 ) ;
  assign n18150 = ( n6420 & ~n6730 ) | ( n6420 & 1'b0 ) | ( ~n6730 & 1'b0 ) ;
  assign n18151 = n18149 | n18150 ;
  assign n18152 = ( x53 & ~n18151 ) | ( x53 & 1'b0 ) | ( ~n18151 & 1'b0 ) ;
  assign n18153 = ~x53 & n18151 ;
  assign n18154 = n18152 | n18153 ;
  assign n18155 = ( n18143 & n18144 ) | ( n18143 & n18154 ) | ( n18144 & n18154 ) ;
  assign n18156 = ( n18144 & ~n18143 ) | ( n18144 & n18154 ) | ( ~n18143 & n18154 ) ;
  assign n18157 = ( n18143 & ~n18155 ) | ( n18143 & n18156 ) | ( ~n18155 & n18156 ) ;
  assign n18158 = ( n18096 & ~n18019 ) | ( n18096 & n18157 ) | ( ~n18019 & n18157 ) ;
  assign n18159 = ( n18019 & ~n18157 ) | ( n18019 & n18096 ) | ( ~n18157 & n18096 ) ;
  assign n18160 = ( n18158 & ~n18096 ) | ( n18158 & n18159 ) | ( ~n18096 & n18159 ) ;
  assign n18161 = ( n18022 & n18086 ) | ( n18022 & n18160 ) | ( n18086 & n18160 ) ;
  assign n18162 = ( n18022 & ~n18086 ) | ( n18022 & n18160 ) | ( ~n18086 & n18160 ) ;
  assign n18163 = ( n18086 & ~n18161 ) | ( n18086 & n18162 ) | ( ~n18161 & n18162 ) ;
  assign n18164 = ( n18023 & ~n18024 ) | ( n18023 & n18034 ) | ( ~n18024 & n18034 ) ;
  assign n18165 = ( n18076 & n18163 ) | ( n18076 & n18164 ) | ( n18163 & n18164 ) ;
  assign n18166 = ( n18163 & ~n18076 ) | ( n18163 & n18164 ) | ( ~n18076 & n18164 ) ;
  assign n18167 = ( n18076 & ~n18165 ) | ( n18076 & n18166 ) | ( ~n18165 & n18166 ) ;
  assign n18168 = ( n18037 & ~n17935 ) | ( n18037 & n18047 ) | ( ~n17935 & n18047 ) ;
  assign n18169 = ( n18066 & ~n18167 ) | ( n18066 & n18168 ) | ( ~n18167 & n18168 ) ;
  assign n18170 = ( n18066 & ~n18168 ) | ( n18066 & n18167 ) | ( ~n18168 & n18167 ) ;
  assign n18171 = ( n18169 & ~n18066 ) | ( n18169 & n18170 ) | ( ~n18066 & n18170 ) ;
  assign n18172 = ( n17927 & ~n17926 ) | ( n17927 & n18053 ) | ( ~n17926 & n18053 ) ;
  assign n18173 = ( n17934 & ~n17933 ) | ( n17934 & n18050 ) | ( ~n17933 & n18050 ) ;
  assign n18175 = ( n18171 & n18172 ) | ( n18171 & n18173 ) | ( n18172 & n18173 ) ;
  assign n18174 = ( n18172 & ~n18171 ) | ( n18172 & n18173 ) | ( ~n18171 & n18173 ) ;
  assign n18176 = ( n18171 & ~n18175 ) | ( n18171 & n18174 ) | ( ~n18175 & n18174 ) ;
  assign n18253 = x120 &  n5586 ;
  assign n18250 = ( x122 & ~n5389 ) | ( x122 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n18251 = x121 &  n5384 ;
  assign n18252 = n18250 | n18251 ;
  assign n18254 = ( x120 & ~n18253 ) | ( x120 & n18252 ) | ( ~n18253 & n18252 ) ;
  assign n18255 = ~n5392 & n9987 ;
  assign n18256 = n18254 | n18255 ;
  assign n18257 = ( x47 & ~n18256 ) | ( x47 & 1'b0 ) | ( ~n18256 & 1'b0 ) ;
  assign n18258 = ~x47 & n18256 ;
  assign n18259 = n18257 | n18258 ;
  assign n18177 = ( n18143 & ~n18154 ) | ( n18143 & n18144 ) | ( ~n18154 & n18144 ) ;
  assign n18178 = ( n18106 & ~n18140 ) | ( n18106 & n18139 ) | ( ~n18140 & n18139 ) ;
  assign n18179 = ( n18116 & n18135 ) | ( n18116 & n18136 ) | ( n18135 & n18136 ) ;
  assign n18214 = x111 &  n7731 ;
  assign n18211 = ( x113 & ~n7538 ) | ( x113 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n18212 = x112 &  n7533 ;
  assign n18213 = n18211 | n18212 ;
  assign n18215 = ( x111 & ~n18214 ) | ( x111 & n18213 ) | ( ~n18214 & n18213 ) ;
  assign n18216 = n6169 | n7541 ;
  assign n18217 = ~n18215 & n18216 ;
  assign n18218 = x56 &  n18217 ;
  assign n18219 = x56 | n18217 ;
  assign n18220 = ~n18218 & n18219 ;
  assign n18180 = ( n17809 & ~x38 ) | ( n17809 & n18119 ) | ( ~x38 & n18119 ) ;
  assign n18181 = x103 &  n10104 ;
  assign n18182 = ( x104 & ~n9760 ) | ( x104 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n18183 = n18181 | n18182 ;
  assign n18187 = x105 &  n9457 ;
  assign n18184 = ( x107 & ~n9150 ) | ( x107 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n18185 = x106 &  n9145 ;
  assign n18186 = n18184 | n18185 ;
  assign n18188 = ( x105 & ~n18187 ) | ( x105 & n18186 ) | ( ~n18187 & n18186 ) ;
  assign n18189 = ( n4848 & ~n18188 ) | ( n4848 & n9153 ) | ( ~n18188 & n9153 ) ;
  assign n18190 = ~n9153 & n18189 ;
  assign n18191 = ( x62 & n18188 ) | ( x62 & n18190 ) | ( n18188 & n18190 ) ;
  assign n18192 = ( x62 & ~n18190 ) | ( x62 & n18188 ) | ( ~n18190 & n18188 ) ;
  assign n18193 = ( n18190 & ~n18191 ) | ( n18190 & n18192 ) | ( ~n18191 & n18192 ) ;
  assign n18194 = ( n18180 & ~n18183 ) | ( n18180 & n18193 ) | ( ~n18183 & n18193 ) ;
  assign n18195 = ( n18180 & ~n18193 ) | ( n18180 & n18183 ) | ( ~n18193 & n18183 ) ;
  assign n18196 = ( n18194 & ~n18180 ) | ( n18194 & n18195 ) | ( ~n18180 & n18195 ) ;
  assign n18201 = x108 &  n8558 ;
  assign n18198 = ( x110 & ~n8314 ) | ( x110 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n18199 = x109 &  n8309 ;
  assign n18200 = n18198 | n18199 ;
  assign n18202 = ( x108 & ~n18201 ) | ( x108 & n18200 ) | ( ~n18201 & n18200 ) ;
  assign n18203 = n5283 | n8317 ;
  assign n18204 = ~n18202 & n18203 ;
  assign n18205 = x59 &  n18204 ;
  assign n18206 = x59 | n18204 ;
  assign n18207 = ~n18205 & n18206 ;
  assign n18197 = ( n17976 & ~n18132 ) | ( n17976 & n18122 ) | ( ~n18132 & n18122 ) ;
  assign n18208 = ( n18196 & ~n18207 ) | ( n18196 & n18197 ) | ( ~n18207 & n18197 ) ;
  assign n18209 = ( n18196 & ~n18197 ) | ( n18196 & n18207 ) | ( ~n18197 & n18207 ) ;
  assign n18210 = ( n18208 & ~n18196 ) | ( n18208 & n18209 ) | ( ~n18196 & n18209 ) ;
  assign n18221 = ( n18179 & ~n18220 ) | ( n18179 & n18210 ) | ( ~n18220 & n18210 ) ;
  assign n18222 = ( n18179 & ~n18210 ) | ( n18179 & n18220 ) | ( ~n18210 & n18220 ) ;
  assign n18223 = ( n18221 & ~n18179 ) | ( n18221 & n18222 ) | ( ~n18179 & n18222 ) ;
  assign n18227 = x114 &  n6982 ;
  assign n18224 = ( x116 & ~n6727 ) | ( x116 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n18225 = x115 &  n6722 ;
  assign n18226 = n18224 | n18225 ;
  assign n18228 = ( x114 & ~n18227 ) | ( x114 & n18226 ) | ( ~n18227 & n18226 ) ;
  assign n18229 = n6730 | n6885 ;
  assign n18230 = ~n18228 & n18229 ;
  assign n18231 = x53 &  n18230 ;
  assign n18232 = x53 | n18230 ;
  assign n18233 = ~n18231 & n18232 ;
  assign n18235 = ( n18178 & n18223 ) | ( n18178 & n18233 ) | ( n18223 & n18233 ) ;
  assign n18234 = ( n18223 & ~n18178 ) | ( n18223 & n18233 ) | ( ~n18178 & n18233 ) ;
  assign n18236 = ( n18178 & ~n18235 ) | ( n18178 & n18234 ) | ( ~n18235 & n18234 ) ;
  assign n18240 = x117 &  n6288 ;
  assign n18237 = ( x119 & ~n6032 ) | ( x119 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n18238 = x118 &  n6027 ;
  assign n18239 = n18237 | n18238 ;
  assign n18241 = ( x117 & ~n18240 ) | ( x117 & n18239 ) | ( ~n18240 & n18239 ) ;
  assign n18242 = ~n6035 & n7648 ;
  assign n18243 = n18241 | n18242 ;
  assign n18245 = x50 &  n18243 ;
  assign n18244 = ~x50 & n18243 ;
  assign n18246 = ( x50 & ~n18245 ) | ( x50 & n18244 ) | ( ~n18245 & n18244 ) ;
  assign n18248 = ( n18177 & n18236 ) | ( n18177 & n18246 ) | ( n18236 & n18246 ) ;
  assign n18247 = ( n18236 & ~n18177 ) | ( n18236 & n18246 ) | ( ~n18177 & n18246 ) ;
  assign n18249 = ( n18177 & ~n18248 ) | ( n18177 & n18247 ) | ( ~n18248 & n18247 ) ;
  assign n18260 = ( n18159 & ~n18259 ) | ( n18159 & n18249 ) | ( ~n18259 & n18249 ) ;
  assign n18261 = ( n18159 & ~n18249 ) | ( n18159 & n18259 ) | ( ~n18249 & n18259 ) ;
  assign n18262 = ( n18260 & ~n18159 ) | ( n18260 & n18261 ) | ( ~n18159 & n18261 ) ;
  assign n18263 = n18161 &  n18262 ;
  assign n18264 = n18161 | n18262 ;
  assign n18265 = ~n18263 & n18264 ;
  assign n18266 = ( x126 & ~n4344 ) | ( x126 & 1'b0 ) | ( ~n4344 & 1'b0 ) ;
  assign n18267 = x127 &  n4138 ;
  assign n18268 = n18266 | n18267 ;
  assign n18269 = n4146 | n9960 ;
  assign n18270 = ( n18268 & ~n4146 ) | ( n18268 & n18269 ) | ( ~n4146 & n18269 ) ;
  assign n18274 = ( n18165 & ~x41 ) | ( n18165 & n18270 ) | ( ~x41 & n18270 ) ;
  assign n18275 = ( x41 & ~n18270 ) | ( x41 & n18165 ) | ( ~n18270 & n18165 ) ;
  assign n18276 = ( n18274 & ~n18165 ) | ( n18274 & n18275 ) | ( ~n18165 & n18275 ) ;
  assign n18280 = x123 &  n4934 ;
  assign n18277 = ( x125 & ~n4725 ) | ( x125 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n18278 = x124 &  n4720 ;
  assign n18279 = n18277 | n18278 ;
  assign n18281 = ( x123 & ~n18280 ) | ( x123 & n18279 ) | ( ~n18280 & n18279 ) ;
  assign n18282 = ~n4728 & n9324 ;
  assign n18283 = n18281 | n18282 ;
  assign n18284 = ( x44 & ~n18283 ) | ( x44 & 1'b0 ) | ( ~n18283 & 1'b0 ) ;
  assign n18285 = ~x44 & n18283 ;
  assign n18286 = n18284 | n18285 ;
  assign n18287 = ( n18265 & ~n18276 ) | ( n18265 & n18286 ) | ( ~n18276 & n18286 ) ;
  assign n18288 = ( n18265 & ~n18286 ) | ( n18265 & n18276 ) | ( ~n18286 & n18276 ) ;
  assign n18289 = ( n18287 & ~n18265 ) | ( n18287 & n18288 ) | ( ~n18265 & n18288 ) ;
  assign n18290 = ( n18171 & ~n18172 ) | ( n18171 & n18173 ) | ( ~n18172 & n18173 ) ;
  assign n18292 = ( n18169 & n18289 ) | ( n18169 & n18290 ) | ( n18289 & n18290 ) ;
  assign n18291 = ( n18289 & ~n18169 ) | ( n18289 & n18290 ) | ( ~n18169 & n18290 ) ;
  assign n18293 = ( n18169 & ~n18292 ) | ( n18169 & n18291 ) | ( ~n18292 & n18291 ) ;
  assign n18294 = ~n18265 & n18286 ;
  assign n18295 = ( n18265 & ~n18286 ) | ( n18265 & 1'b0 ) | ( ~n18286 & 1'b0 ) ;
  assign n18296 = n18294 | n18295 ;
  assign n18271 = x41 | n18270 ;
  assign n18272 = ( x41 & ~n18270 ) | ( x41 & 1'b0 ) | ( ~n18270 & 1'b0 ) ;
  assign n18273 = ( n18271 & ~x41 ) | ( n18271 & n18272 ) | ( ~x41 & n18272 ) ;
  assign n18297 = ( n18165 & ~n18296 ) | ( n18165 & n18273 ) | ( ~n18296 & n18273 ) ;
  assign n18298 = ( n18169 & ~n18290 ) | ( n18169 & n18289 ) | ( ~n18290 & n18289 ) ;
  assign n18299 = ( x127 & ~n4344 ) | ( x127 & 1'b0 ) | ( ~n4344 & 1'b0 ) ;
  assign n18300 = n4146 | n10258 ;
  assign n18301 = ~n18299 & n18300 ;
  assign n18302 = ~x41 & n18301 ;
  assign n18303 = ( x41 & ~n18301 ) | ( x41 & 1'b0 ) | ( ~n18301 & 1'b0 ) ;
  assign n18304 = n18302 | n18303 ;
  assign n18305 = ( n18161 & ~n18262 ) | ( n18161 & n18286 ) | ( ~n18262 & n18286 ) ;
  assign n18306 = ( n18249 & ~n18159 ) | ( n18249 & n18259 ) | ( ~n18159 & n18259 ) ;
  assign n18307 = ( n18177 & ~n18246 ) | ( n18177 & n18236 ) | ( ~n18246 & n18236 ) ;
  assign n18318 = ( n18178 & ~n18233 ) | ( n18178 & n18223 ) | ( ~n18233 & n18223 ) ;
  assign n18322 = x118 &  n6288 ;
  assign n18319 = ( x120 & ~n6032 ) | ( x120 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n18320 = x119 &  n6027 ;
  assign n18321 = n18319 | n18320 ;
  assign n18323 = ( x118 & ~n18322 ) | ( x118 & n18321 ) | ( ~n18322 & n18321 ) ;
  assign n18324 = ~n6035 & n9364 ;
  assign n18325 = n18323 | n18324 ;
  assign n18326 = ( x50 & ~n18325 ) | ( x50 & 1'b0 ) | ( ~n18325 & 1'b0 ) ;
  assign n18327 = ~x50 & n18325 ;
  assign n18328 = n18326 | n18327 ;
  assign n18329 = ( n18210 & ~n18179 ) | ( n18210 & n18220 ) | ( ~n18179 & n18220 ) ;
  assign n18333 = x115 &  n6982 ;
  assign n18330 = ( x117 & ~n6727 ) | ( x117 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n18331 = x116 &  n6722 ;
  assign n18332 = n18330 | n18331 ;
  assign n18334 = ( x115 & ~n18333 ) | ( x115 & n18332 ) | ( ~n18333 & n18332 ) ;
  assign n18335 = n6730 | n7136 ;
  assign n18336 = ~n18334 & n18335 ;
  assign n18337 = x53 &  n18336 ;
  assign n18338 = x53 | n18336 ;
  assign n18339 = ~n18337 & n18338 ;
  assign n18343 = x106 &  n9457 ;
  assign n18340 = ( x108 & ~n9150 ) | ( x108 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n18341 = x107 &  n9145 ;
  assign n18342 = n18340 | n18341 ;
  assign n18344 = ( x106 & ~n18343 ) | ( x106 & n18342 ) | ( ~n18343 & n18342 ) ;
  assign n18345 = n5055 | n9153 ;
  assign n18346 = ~n18344 & n18345 ;
  assign n18347 = x62 &  n18346 ;
  assign n18348 = x62 | n18346 ;
  assign n18349 = ~n18347 & n18348 ;
  assign n18350 = x104 &  n10104 ;
  assign n18351 = ( x105 & ~n9760 ) | ( x105 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n18352 = n18350 | n18351 ;
  assign n18353 = ( n18194 & ~n18183 ) | ( n18194 & n18352 ) | ( ~n18183 & n18352 ) ;
  assign n18354 = ( n18183 & ~n18352 ) | ( n18183 & n18194 ) | ( ~n18352 & n18194 ) ;
  assign n18355 = ( n18353 & ~n18194 ) | ( n18353 & n18354 ) | ( ~n18194 & n18354 ) ;
  assign n18359 = x109 &  n8558 ;
  assign n18356 = ( x111 & ~n8314 ) | ( x111 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n18357 = x110 &  n8309 ;
  assign n18358 = n18356 | n18357 ;
  assign n18360 = ( x109 & ~n18359 ) | ( x109 & n18358 ) | ( ~n18359 & n18358 ) ;
  assign n18361 = n5711 | n8317 ;
  assign n18362 = ~n18360 & n18361 ;
  assign n18363 = x59 &  n18362 ;
  assign n18364 = x59 | n18362 ;
  assign n18365 = ~n18363 & n18364 ;
  assign n18366 = ( n18349 & ~n18355 ) | ( n18349 & n18365 ) | ( ~n18355 & n18365 ) ;
  assign n18367 = ( n18349 & ~n18365 ) | ( n18349 & n18355 ) | ( ~n18365 & n18355 ) ;
  assign n18368 = ( n18366 & ~n18349 ) | ( n18366 & n18367 ) | ( ~n18349 & n18367 ) ;
  assign n18373 = x112 &  n7731 ;
  assign n18370 = ( x114 & ~n7538 ) | ( x114 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n18371 = x113 &  n7533 ;
  assign n18372 = n18370 | n18371 ;
  assign n18374 = ( x112 & ~n18373 ) | ( x112 & n18372 ) | ( ~n18373 & n18372 ) ;
  assign n18375 = n6185 | n7541 ;
  assign n18376 = ~n18374 & n18375 ;
  assign n18377 = x56 &  n18376 ;
  assign n18378 = x56 | n18376 ;
  assign n18379 = ~n18377 & n18378 ;
  assign n18369 = ( n18196 & n18197 ) | ( n18196 & n18207 ) | ( n18197 & n18207 ) ;
  assign n18380 = ( n18368 & ~n18379 ) | ( n18368 & n18369 ) | ( ~n18379 & n18369 ) ;
  assign n18381 = ( n18368 & ~n18369 ) | ( n18368 & n18379 ) | ( ~n18369 & n18379 ) ;
  assign n18382 = ( n18380 & ~n18368 ) | ( n18380 & n18381 ) | ( ~n18368 & n18381 ) ;
  assign n18384 = ( n18329 & n18339 ) | ( n18329 & n18382 ) | ( n18339 & n18382 ) ;
  assign n18383 = ( n18339 & ~n18329 ) | ( n18339 & n18382 ) | ( ~n18329 & n18382 ) ;
  assign n18385 = ( n18329 & ~n18384 ) | ( n18329 & n18383 ) | ( ~n18384 & n18383 ) ;
  assign n18386 = ( n18318 & ~n18328 ) | ( n18318 & n18385 ) | ( ~n18328 & n18385 ) ;
  assign n18387 = ( n18318 & ~n18385 ) | ( n18318 & n18328 ) | ( ~n18385 & n18328 ) ;
  assign n18388 = ( n18386 & ~n18318 ) | ( n18386 & n18387 ) | ( ~n18318 & n18387 ) ;
  assign n18311 = x121 &  n5586 ;
  assign n18308 = ( x123 & ~n5389 ) | ( x123 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n18309 = x122 &  n5384 ;
  assign n18310 = n18308 | n18309 ;
  assign n18312 = ( x121 & ~n18311 ) | ( x121 & n18310 ) | ( ~n18311 & n18310 ) ;
  assign n18313 = ~n5392 & n8472 ;
  assign n18314 = n18312 | n18313 ;
  assign n18315 = ( x47 & ~n18314 ) | ( x47 & 1'b0 ) | ( ~n18314 & 1'b0 ) ;
  assign n18316 = ~x47 & n18314 ;
  assign n18317 = n18315 | n18316 ;
  assign n18389 = ( n18307 & ~n18388 ) | ( n18307 & n18317 ) | ( ~n18388 & n18317 ) ;
  assign n18390 = ( n18307 & ~n18317 ) | ( n18307 & n18388 ) | ( ~n18317 & n18388 ) ;
  assign n18391 = ( n18389 & ~n18307 ) | ( n18389 & n18390 ) | ( ~n18307 & n18390 ) ;
  assign n18395 = x124 &  n4934 ;
  assign n18392 = ( x126 & ~n4725 ) | ( x126 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n18393 = x125 &  n4720 ;
  assign n18394 = n18392 | n18393 ;
  assign n18396 = ( x124 & ~n18395 ) | ( x124 & n18394 ) | ( ~n18395 & n18394 ) ;
  assign n18397 = n4728 | n9349 ;
  assign n18398 = ~n18396 & n18397 ;
  assign n18399 = x44 &  n18398 ;
  assign n18400 = x44 | n18398 ;
  assign n18401 = ~n18399 & n18400 ;
  assign n18403 = ( n18306 & n18391 ) | ( n18306 & n18401 ) | ( n18391 & n18401 ) ;
  assign n18402 = ( n18391 & ~n18306 ) | ( n18391 & n18401 ) | ( ~n18306 & n18401 ) ;
  assign n18404 = ( n18306 & ~n18403 ) | ( n18306 & n18402 ) | ( ~n18403 & n18402 ) ;
  assign n18405 = ( n18304 & n18305 ) | ( n18304 & n18404 ) | ( n18305 & n18404 ) ;
  assign n18406 = ( n18305 & ~n18304 ) | ( n18305 & n18404 ) | ( ~n18304 & n18404 ) ;
  assign n18407 = ( n18304 & ~n18405 ) | ( n18304 & n18406 ) | ( ~n18405 & n18406 ) ;
  assign n18408 = ( n18297 & n18298 ) | ( n18297 & n18407 ) | ( n18298 & n18407 ) ;
  assign n18409 = ( n18298 & ~n18297 ) | ( n18298 & n18407 ) | ( ~n18297 & n18407 ) ;
  assign n18410 = ( n18297 & ~n18408 ) | ( n18297 & n18409 ) | ( ~n18408 & n18409 ) ;
  assign n18414 = x125 &  n4934 ;
  assign n18411 = ( x127 & ~n4725 ) | ( x127 & 1'b0 ) | ( ~n4725 & 1'b0 ) ;
  assign n18412 = x126 &  n4720 ;
  assign n18413 = n18411 | n18412 ;
  assign n18415 = ( x125 & ~n18414 ) | ( x125 & n18413 ) | ( ~n18414 & n18413 ) ;
  assign n18416 = n4728 | n9941 ;
  assign n18417 = ~n18415 & n18416 ;
  assign n18418 = x44 &  n18417 ;
  assign n18419 = x44 | n18417 ;
  assign n18420 = ~n18418 & n18419 ;
  assign n18424 = x119 &  n6288 ;
  assign n18421 = ( x121 & ~n6032 ) | ( x121 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n18422 = x120 &  n6027 ;
  assign n18423 = n18421 | n18422 ;
  assign n18425 = ( x119 & ~n18424 ) | ( x119 & n18423 ) | ( ~n18424 & n18423 ) ;
  assign n18426 = ~n6035 & n8176 ;
  assign n18427 = n18425 | n18426 ;
  assign n18428 = ( x50 & ~n18427 ) | ( x50 & 1'b0 ) | ( ~n18427 & 1'b0 ) ;
  assign n18429 = ~x50 & n18427 ;
  assign n18430 = n18428 | n18429 ;
  assign n18434 = x113 &  n7731 ;
  assign n18431 = ( x115 & ~n7538 ) | ( x115 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n18432 = x114 &  n7533 ;
  assign n18433 = n18431 | n18432 ;
  assign n18435 = ( x113 & ~n18434 ) | ( x113 & n18433 ) | ( ~n18434 & n18433 ) ;
  assign n18436 = ( n6420 & ~n7541 ) | ( n6420 & 1'b0 ) | ( ~n7541 & 1'b0 ) ;
  assign n18437 = n18435 | n18436 ;
  assign n18438 = ( x56 & ~n18437 ) | ( x56 & 1'b0 ) | ( ~n18437 & 1'b0 ) ;
  assign n18439 = ~x56 & n18437 ;
  assign n18440 = n18438 | n18439 ;
  assign n18445 = x110 &  n8558 ;
  assign n18442 = ( x112 & ~n8314 ) | ( x112 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n18443 = x111 &  n8309 ;
  assign n18444 = n18442 | n18443 ;
  assign n18446 = ( x110 & ~n18445 ) | ( x110 & n18444 ) | ( ~n18445 & n18444 ) ;
  assign n18447 = ( n5727 & ~n8317 ) | ( n5727 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n18448 = n18446 | n18447 ;
  assign n18449 = ( x59 & ~n18448 ) | ( x59 & 1'b0 ) | ( ~n18448 & 1'b0 ) ;
  assign n18450 = ~x59 & n18448 ;
  assign n18451 = n18449 | n18450 ;
  assign n18452 = x105 &  n10104 ;
  assign n18453 = ( x106 & ~n9760 ) | ( x106 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n18454 = n18452 | n18453 ;
  assign n18455 = ( x41 & n18183 ) | ( x41 & n18454 ) | ( n18183 & n18454 ) ;
  assign n18456 = ( x41 & ~n18183 ) | ( x41 & n18454 ) | ( ~n18183 & n18454 ) ;
  assign n18457 = ( n18183 & ~n18455 ) | ( n18183 & n18456 ) | ( ~n18455 & n18456 ) ;
  assign n18461 = x107 &  n9457 ;
  assign n18458 = ( x109 & ~n9150 ) | ( x109 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n18459 = x108 &  n9145 ;
  assign n18460 = n18458 | n18459 ;
  assign n18462 = ( x107 & ~n18461 ) | ( x107 & n18460 ) | ( ~n18461 & n18460 ) ;
  assign n18463 = ( n5267 & ~n9153 ) | ( n5267 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n18464 = n18462 | n18463 ;
  assign n18465 = ( x62 & ~n18464 ) | ( x62 & 1'b0 ) | ( ~n18464 & 1'b0 ) ;
  assign n18466 = ~x62 & n18464 ;
  assign n18467 = n18465 | n18466 ;
  assign n18468 = ( n18353 & ~n18457 ) | ( n18353 & n18467 ) | ( ~n18457 & n18467 ) ;
  assign n18469 = ( n18457 & ~n18353 ) | ( n18457 & n18467 ) | ( ~n18353 & n18467 ) ;
  assign n18470 = ( n18468 & ~n18467 ) | ( n18468 & n18469 ) | ( ~n18467 & n18469 ) ;
  assign n18471 = ( n18349 & n18355 ) | ( n18349 & n18365 ) | ( n18355 & n18365 ) ;
  assign n18473 = ( n18451 & n18470 ) | ( n18451 & n18471 ) | ( n18470 & n18471 ) ;
  assign n18472 = ( n18470 & ~n18451 ) | ( n18470 & n18471 ) | ( ~n18451 & n18471 ) ;
  assign n18474 = ( n18451 & ~n18473 ) | ( n18451 & n18472 ) | ( ~n18473 & n18472 ) ;
  assign n18441 = ( n18368 & n18369 ) | ( n18368 & n18379 ) | ( n18369 & n18379 ) ;
  assign n18475 = ( n18440 & ~n18474 ) | ( n18440 & n18441 ) | ( ~n18474 & n18441 ) ;
  assign n18476 = ( n18440 & ~n18441 ) | ( n18440 & n18474 ) | ( ~n18441 & n18474 ) ;
  assign n18477 = ( n18475 & ~n18440 ) | ( n18475 & n18476 ) | ( ~n18440 & n18476 ) ;
  assign n18481 = x116 &  n6982 ;
  assign n18478 = ( x118 & ~n6727 ) | ( x118 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n18479 = x117 &  n6722 ;
  assign n18480 = n18478 | n18479 ;
  assign n18482 = ( x116 & ~n18481 ) | ( x116 & n18480 ) | ( ~n18481 & n18480 ) ;
  assign n18483 = n6730 | n7152 ;
  assign n18484 = ~n18482 & n18483 ;
  assign n18485 = x53 &  n18484 ;
  assign n18486 = x53 | n18484 ;
  assign n18487 = ~n18485 & n18486 ;
  assign n18488 = ( n18477 & ~n18384 ) | ( n18477 & n18487 ) | ( ~n18384 & n18487 ) ;
  assign n18489 = ( n18384 & ~n18487 ) | ( n18384 & n18477 ) | ( ~n18487 & n18477 ) ;
  assign n18490 = ( n18488 & ~n18477 ) | ( n18488 & n18489 ) | ( ~n18477 & n18489 ) ;
  assign n18491 = ( n18430 & ~n18387 ) | ( n18430 & n18490 ) | ( ~n18387 & n18490 ) ;
  assign n18492 = ( n18387 & ~n18490 ) | ( n18387 & n18430 ) | ( ~n18490 & n18430 ) ;
  assign n18493 = ( n18491 & ~n18430 ) | ( n18491 & n18492 ) | ( ~n18430 & n18492 ) ;
  assign n18497 = x122 &  n5586 ;
  assign n18494 = ( x124 & ~n5389 ) | ( x124 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n18495 = x123 &  n5384 ;
  assign n18496 = n18494 | n18495 ;
  assign n18498 = ( x122 & ~n18497 ) | ( x122 & n18496 ) | ( ~n18497 & n18496 ) ;
  assign n18499 = ~n5392 & n8755 ;
  assign n18500 = n18498 | n18499 ;
  assign n18501 = ( x47 & ~n18500 ) | ( x47 & 1'b0 ) | ( ~n18500 & 1'b0 ) ;
  assign n18502 = ~x47 & n18500 ;
  assign n18503 = n18501 | n18502 ;
  assign n18505 = ( n18390 & n18493 ) | ( n18390 & n18503 ) | ( n18493 & n18503 ) ;
  assign n18504 = ( n18390 & ~n18493 ) | ( n18390 & n18503 ) | ( ~n18493 & n18503 ) ;
  assign n18506 = ( n18493 & ~n18505 ) | ( n18493 & n18504 ) | ( ~n18505 & n18504 ) ;
  assign n18507 = ( n18306 & ~n18401 ) | ( n18306 & n18391 ) | ( ~n18401 & n18391 ) ;
  assign n18509 = ( n18420 & n18506 ) | ( n18420 & n18507 ) | ( n18506 & n18507 ) ;
  assign n18508 = ( n18506 & ~n18420 ) | ( n18506 & n18507 ) | ( ~n18420 & n18507 ) ;
  assign n18510 = ( n18420 & ~n18509 ) | ( n18420 & n18508 ) | ( ~n18509 & n18508 ) ;
  assign n18511 = ( n18297 & ~n18298 ) | ( n18297 & n18407 ) | ( ~n18298 & n18407 ) ;
  assign n18512 = ( n18304 & ~n18305 ) | ( n18304 & n18404 ) | ( ~n18305 & n18404 ) ;
  assign n18514 = ( n18510 & n18511 ) | ( n18510 & n18512 ) | ( n18511 & n18512 ) ;
  assign n18513 = ( n18511 & ~n18510 ) | ( n18511 & n18512 ) | ( ~n18510 & n18512 ) ;
  assign n18515 = ( n18510 & ~n18514 ) | ( n18510 & n18513 ) | ( ~n18514 & n18513 ) ;
  assign n18611 = ( n18510 & ~n18511 ) | ( n18510 & n18512 ) | ( ~n18511 & n18512 ) ;
  assign n18516 = ( x126 & ~n4934 ) | ( x126 & 1'b0 ) | ( ~n4934 & 1'b0 ) ;
  assign n18517 = x127 &  n4720 ;
  assign n18518 = n18516 | n18517 ;
  assign n18519 = n4728 | n9960 ;
  assign n18520 = ( n18518 & ~n4728 ) | ( n18518 & n18519 ) | ( ~n4728 & n18519 ) ;
  assign n18521 = x44 | n18520 ;
  assign n18522 = ( x44 & ~n18520 ) | ( x44 & 1'b0 ) | ( ~n18520 & 1'b0 ) ;
  assign n18523 = ( n18521 & ~x44 ) | ( n18521 & n18522 ) | ( ~x44 & n18522 ) ;
  assign n18524 = ( n18390 & ~n18503 ) | ( n18390 & n18493 ) | ( ~n18503 & n18493 ) ;
  assign n18528 = x123 &  n5586 ;
  assign n18525 = ( x125 & ~n5389 ) | ( x125 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n18526 = x124 &  n5384 ;
  assign n18527 = n18525 | n18526 ;
  assign n18529 = ( x123 & ~n18528 ) | ( x123 & n18527 ) | ( ~n18528 & n18527 ) ;
  assign n18530 = ~n5392 & n9324 ;
  assign n18531 = n18529 | n18530 ;
  assign n18532 = ( x47 & ~n18531 ) | ( x47 & 1'b0 ) | ( ~n18531 & 1'b0 ) ;
  assign n18533 = ~x47 & n18531 ;
  assign n18534 = n18532 | n18533 ;
  assign n18535 = ( n18183 & ~x41 ) | ( n18183 & n18454 ) | ( ~x41 & n18454 ) ;
  assign n18536 = x106 &  n10104 ;
  assign n18537 = ( x107 & ~n9760 ) | ( x107 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n18538 = n18536 | n18537 ;
  assign n18542 = x108 &  n9457 ;
  assign n18539 = ( x110 & ~n9150 ) | ( x110 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n18540 = x109 &  n9145 ;
  assign n18541 = n18539 | n18540 ;
  assign n18543 = ( x108 & ~n18542 ) | ( x108 & n18541 ) | ( ~n18542 & n18541 ) ;
  assign n18544 = ( n5283 & ~n9153 ) | ( n5283 & n18543 ) | ( ~n9153 & n18543 ) ;
  assign n18545 = n9153 | n18544 ;
  assign n18547 = ( x62 & n18543 ) | ( x62 & n18545 ) | ( n18543 & n18545 ) ;
  assign n18546 = ( x62 & ~n18545 ) | ( x62 & n18543 ) | ( ~n18545 & n18543 ) ;
  assign n18548 = ( n18545 & ~n18547 ) | ( n18545 & n18546 ) | ( ~n18547 & n18546 ) ;
  assign n18550 = ( n18535 & n18538 ) | ( n18535 & n18548 ) | ( n18538 & n18548 ) ;
  assign n18549 = ( n18538 & ~n18535 ) | ( n18538 & n18548 ) | ( ~n18535 & n18548 ) ;
  assign n18551 = ( n18535 & ~n18550 ) | ( n18535 & n18549 ) | ( ~n18550 & n18549 ) ;
  assign n18555 = x111 &  n8558 ;
  assign n18552 = ( x113 & ~n8314 ) | ( x113 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n18553 = x112 &  n8309 ;
  assign n18554 = n18552 | n18553 ;
  assign n18556 = ( x111 & ~n18555 ) | ( x111 & n18554 ) | ( ~n18555 & n18554 ) ;
  assign n18557 = n6169 | n8317 ;
  assign n18558 = ~n18556 & n18557 ;
  assign n18559 = x59 &  n18558 ;
  assign n18560 = x59 | n18558 ;
  assign n18561 = ~n18559 & n18560 ;
  assign n18562 = ( n18468 & n18551 ) | ( n18468 & n18561 ) | ( n18551 & n18561 ) ;
  assign n18563 = ( n18468 & ~n18551 ) | ( n18468 & n18561 ) | ( ~n18551 & n18561 ) ;
  assign n18564 = ( n18551 & ~n18562 ) | ( n18551 & n18563 ) | ( ~n18562 & n18563 ) ;
  assign n18568 = x114 &  n7731 ;
  assign n18565 = ( x116 & ~n7538 ) | ( x116 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n18566 = x115 &  n7533 ;
  assign n18567 = n18565 | n18566 ;
  assign n18569 = ( x114 & ~n18568 ) | ( x114 & n18567 ) | ( ~n18568 & n18567 ) ;
  assign n18570 = n6885 | n7541 ;
  assign n18571 = ~n18569 & n18570 ;
  assign n18572 = x56 &  n18571 ;
  assign n18573 = x56 | n18571 ;
  assign n18574 = ~n18572 & n18573 ;
  assign n18575 = ( n18472 & ~n18564 ) | ( n18472 & n18574 ) | ( ~n18564 & n18574 ) ;
  assign n18576 = ( n18472 & ~n18574 ) | ( n18472 & n18564 ) | ( ~n18574 & n18564 ) ;
  assign n18577 = ( n18575 & ~n18472 ) | ( n18575 & n18576 ) | ( ~n18472 & n18576 ) ;
  assign n18581 = x117 &  n6982 ;
  assign n18578 = ( x119 & ~n6727 ) | ( x119 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n18579 = x118 &  n6722 ;
  assign n18580 = n18578 | n18579 ;
  assign n18582 = ( x117 & ~n18581 ) | ( x117 & n18580 ) | ( ~n18581 & n18580 ) ;
  assign n18583 = ~n6730 & n7648 ;
  assign n18584 = n18582 | n18583 ;
  assign n18585 = ( x53 & ~n18584 ) | ( x53 & 1'b0 ) | ( ~n18584 & 1'b0 ) ;
  assign n18586 = ~x53 & n18584 ;
  assign n18587 = n18585 | n18586 ;
  assign n18588 = ( n18476 & n18577 ) | ( n18476 & n18587 ) | ( n18577 & n18587 ) ;
  assign n18589 = ( n18577 & ~n18476 ) | ( n18577 & n18587 ) | ( ~n18476 & n18587 ) ;
  assign n18590 = ( n18476 & ~n18588 ) | ( n18476 & n18589 ) | ( ~n18588 & n18589 ) ;
  assign n18591 = ( n18384 & n18477 ) | ( n18384 & n18487 ) | ( n18477 & n18487 ) ;
  assign n18595 = x120 &  n6288 ;
  assign n18592 = ( x122 & ~n6032 ) | ( x122 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n18593 = x121 &  n6027 ;
  assign n18594 = n18592 | n18593 ;
  assign n18596 = ( x120 & ~n18595 ) | ( x120 & n18594 ) | ( ~n18595 & n18594 ) ;
  assign n18597 = ~n6035 & n9987 ;
  assign n18598 = n18596 | n18597 ;
  assign n18599 = ( x50 & ~n18598 ) | ( x50 & 1'b0 ) | ( ~n18598 & 1'b0 ) ;
  assign n18600 = ~x50 & n18598 ;
  assign n18601 = n18599 | n18600 ;
  assign n18603 = ( n18590 & n18591 ) | ( n18590 & n18601 ) | ( n18591 & n18601 ) ;
  assign n18602 = ( n18591 & ~n18590 ) | ( n18591 & n18601 ) | ( ~n18590 & n18601 ) ;
  assign n18604 = ( n18590 & ~n18603 ) | ( n18590 & n18602 ) | ( ~n18603 & n18602 ) ;
  assign n18606 = ( n18492 & n18534 ) | ( n18492 & n18604 ) | ( n18534 & n18604 ) ;
  assign n18605 = ( n18534 & ~n18492 ) | ( n18534 & n18604 ) | ( ~n18492 & n18604 ) ;
  assign n18607 = ( n18492 & ~n18606 ) | ( n18492 & n18605 ) | ( ~n18606 & n18605 ) ;
  assign n18608 = ( n18523 & n18524 ) | ( n18523 & n18607 ) | ( n18524 & n18607 ) ;
  assign n18609 = ( n18524 & ~n18523 ) | ( n18524 & n18607 ) | ( ~n18523 & n18607 ) ;
  assign n18610 = ( n18523 & ~n18608 ) | ( n18523 & n18609 ) | ( ~n18608 & n18609 ) ;
  assign n18612 = ( n18508 & ~n18611 ) | ( n18508 & n18610 ) | ( ~n18611 & n18610 ) ;
  assign n18613 = ( n18508 & ~n18610 ) | ( n18508 & n18611 ) | ( ~n18610 & n18611 ) ;
  assign n18614 = ( n18612 & ~n18508 ) | ( n18612 & n18613 ) | ( ~n18508 & n18613 ) ;
  assign n18615 = ( n18523 & ~n18524 ) | ( n18523 & n18607 ) | ( ~n18524 & n18607 ) ;
  assign n18623 = ( n18590 & ~n18601 ) | ( n18590 & n18591 ) | ( ~n18601 & n18591 ) ;
  assign n18624 = ( n18476 & ~n18577 ) | ( n18476 & n18587 ) | ( ~n18577 & n18587 ) ;
  assign n18628 = x121 &  n6288 ;
  assign n18625 = ( x123 & ~n6032 ) | ( x123 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n18626 = x122 &  n6027 ;
  assign n18627 = n18625 | n18626 ;
  assign n18629 = ( x121 & ~n18628 ) | ( x121 & n18627 ) | ( ~n18628 & n18627 ) ;
  assign n18630 = ~n6035 & n8472 ;
  assign n18631 = n18629 | n18630 ;
  assign n18632 = ( x50 & ~n18631 ) | ( x50 & 1'b0 ) | ( ~n18631 & 1'b0 ) ;
  assign n18633 = ~x50 & n18631 ;
  assign n18634 = n18632 | n18633 ;
  assign n18635 = ( n18472 & n18564 ) | ( n18472 & n18574 ) | ( n18564 & n18574 ) ;
  assign n18646 = ( n18468 & ~n18561 ) | ( n18468 & n18551 ) | ( ~n18561 & n18551 ) ;
  assign n18660 = x112 &  n8558 ;
  assign n18657 = ( x114 & ~n8314 ) | ( x114 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n18658 = x113 &  n8309 ;
  assign n18659 = n18657 | n18658 ;
  assign n18661 = ( x112 & ~n18660 ) | ( x112 & n18659 ) | ( ~n18660 & n18659 ) ;
  assign n18662 = n6185 | n8317 ;
  assign n18663 = ~n18661 & n18662 ;
  assign n18664 = x59 &  n18663 ;
  assign n18665 = x59 | n18663 ;
  assign n18666 = ~n18664 & n18665 ;
  assign n18667 = x107 &  n10104 ;
  assign n18668 = ( x108 & ~n9760 ) | ( x108 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n18669 = n18667 | n18668 ;
  assign n18673 = x109 &  n9457 ;
  assign n18670 = ( x111 & ~n9150 ) | ( x111 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n18671 = x110 &  n9145 ;
  assign n18672 = n18670 | n18671 ;
  assign n18674 = ( x109 & ~n18673 ) | ( x109 & n18672 ) | ( ~n18673 & n18672 ) ;
  assign n18675 = ( n5711 & ~n9153 ) | ( n5711 & n18674 ) | ( ~n9153 & n18674 ) ;
  assign n18676 = n9153 | n18675 ;
  assign n18678 = ( x62 & n18674 ) | ( x62 & n18676 ) | ( n18674 & n18676 ) ;
  assign n18677 = ( x62 & ~n18676 ) | ( x62 & n18674 ) | ( ~n18676 & n18674 ) ;
  assign n18679 = ( n18676 & ~n18678 ) | ( n18676 & n18677 ) | ( ~n18678 & n18677 ) ;
  assign n18681 = ( n18538 & n18669 ) | ( n18538 & n18679 ) | ( n18669 & n18679 ) ;
  assign n18680 = ( n18538 & ~n18669 ) | ( n18538 & n18679 ) | ( ~n18669 & n18679 ) ;
  assign n18682 = ( n18669 & ~n18681 ) | ( n18669 & n18680 ) | ( ~n18681 & n18680 ) ;
  assign n18683 = ( n18549 & ~n18666 ) | ( n18549 & n18682 ) | ( ~n18666 & n18682 ) ;
  assign n18684 = ( n18549 & ~n18682 ) | ( n18549 & n18666 ) | ( ~n18682 & n18666 ) ;
  assign n18685 = ( n18683 & ~n18549 ) | ( n18683 & n18684 ) | ( ~n18549 & n18684 ) ;
  assign n18650 = x115 &  n7731 ;
  assign n18647 = ( x117 & ~n7538 ) | ( x117 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n18648 = x116 &  n7533 ;
  assign n18649 = n18647 | n18648 ;
  assign n18651 = ( x115 & ~n18650 ) | ( x115 & n18649 ) | ( ~n18650 & n18649 ) ;
  assign n18652 = n7136 | n7541 ;
  assign n18653 = ~n18651 & n18652 ;
  assign n18654 = x56 &  n18653 ;
  assign n18655 = x56 | n18653 ;
  assign n18656 = ~n18654 & n18655 ;
  assign n18686 = ( n18646 & ~n18685 ) | ( n18646 & n18656 ) | ( ~n18685 & n18656 ) ;
  assign n18687 = ( n18646 & ~n18656 ) | ( n18646 & n18685 ) | ( ~n18656 & n18685 ) ;
  assign n18688 = ( n18686 & ~n18646 ) | ( n18686 & n18687 ) | ( ~n18646 & n18687 ) ;
  assign n18639 = x118 &  n6982 ;
  assign n18636 = ( x120 & ~n6727 ) | ( x120 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n18637 = x119 &  n6722 ;
  assign n18638 = n18636 | n18637 ;
  assign n18640 = ( x118 & ~n18639 ) | ( x118 & n18638 ) | ( ~n18639 & n18638 ) ;
  assign n18641 = ~n6730 & n9364 ;
  assign n18642 = n18640 | n18641 ;
  assign n18643 = ( x53 & ~n18642 ) | ( x53 & 1'b0 ) | ( ~n18642 & 1'b0 ) ;
  assign n18644 = ~x53 & n18642 ;
  assign n18645 = n18643 | n18644 ;
  assign n18689 = ( n18635 & ~n18688 ) | ( n18635 & n18645 ) | ( ~n18688 & n18645 ) ;
  assign n18690 = ( n18635 & ~n18645 ) | ( n18635 & n18688 ) | ( ~n18645 & n18688 ) ;
  assign n18691 = ( n18689 & ~n18635 ) | ( n18689 & n18690 ) | ( ~n18635 & n18690 ) ;
  assign n18693 = ( n18624 & n18634 ) | ( n18624 & n18691 ) | ( n18634 & n18691 ) ;
  assign n18692 = ( n18634 & ~n18624 ) | ( n18634 & n18691 ) | ( ~n18624 & n18691 ) ;
  assign n18694 = ( n18624 & ~n18693 ) | ( n18624 & n18692 ) | ( ~n18693 & n18692 ) ;
  assign n18698 = x124 &  n5586 ;
  assign n18695 = ( x126 & ~n5389 ) | ( x126 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n18696 = x125 &  n5384 ;
  assign n18697 = n18695 | n18696 ;
  assign n18699 = ( x124 & ~n18698 ) | ( x124 & n18697 ) | ( ~n18698 & n18697 ) ;
  assign n18700 = n5392 | n9349 ;
  assign n18701 = ~n18699 & n18700 ;
  assign n18702 = x47 &  n18701 ;
  assign n18703 = x47 | n18701 ;
  assign n18704 = ~n18702 & n18703 ;
  assign n18705 = ( n18623 & n18694 ) | ( n18623 & n18704 ) | ( n18694 & n18704 ) ;
  assign n18706 = ( n18694 & ~n18623 ) | ( n18694 & n18704 ) | ( ~n18623 & n18704 ) ;
  assign n18707 = ( n18623 & ~n18705 ) | ( n18623 & n18706 ) | ( ~n18705 & n18706 ) ;
  assign n18617 = ( x127 & ~n4934 ) | ( x127 & 1'b0 ) | ( ~n4934 & 1'b0 ) ;
  assign n18618 = n4728 | n10258 ;
  assign n18619 = ~n18617 & n18618 ;
  assign n18620 = ~x44 & n18619 ;
  assign n18621 = ( x44 & ~n18619 ) | ( x44 & 1'b0 ) | ( ~n18619 & 1'b0 ) ;
  assign n18622 = n18620 | n18621 ;
  assign n18708 = ( n18606 & ~n18707 ) | ( n18606 & n18622 ) | ( ~n18707 & n18622 ) ;
  assign n18709 = ( n18622 & ~n18606 ) | ( n18622 & n18707 ) | ( ~n18606 & n18707 ) ;
  assign n18710 = ( n18708 & ~n18622 ) | ( n18708 & n18709 ) | ( ~n18622 & n18709 ) ;
  assign n18616 = ( n18610 & ~n18508 ) | ( n18610 & n18611 ) | ( ~n18508 & n18611 ) ;
  assign n18711 = ( n18615 & ~n18710 ) | ( n18615 & n18616 ) | ( ~n18710 & n18616 ) ;
  assign n18712 = ( n18615 & ~n18616 ) | ( n18615 & n18710 ) | ( ~n18616 & n18710 ) ;
  assign n18713 = ( n18711 & ~n18615 ) | ( n18711 & n18712 ) | ( ~n18615 & n18712 ) ;
  assign n18717 = x122 &  n6288 ;
  assign n18714 = ( x124 & ~n6032 ) | ( x124 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n18715 = x123 &  n6027 ;
  assign n18716 = n18714 | n18715 ;
  assign n18718 = ( x122 & ~n18717 ) | ( x122 & n18716 ) | ( ~n18717 & n18716 ) ;
  assign n18719 = ~n6035 & n8755 ;
  assign n18720 = n18718 | n18719 ;
  assign n18721 = ( x50 & ~n18720 ) | ( x50 & 1'b0 ) | ( ~n18720 & 1'b0 ) ;
  assign n18722 = ~x50 & n18720 ;
  assign n18723 = n18721 | n18722 ;
  assign n18744 = x108 &  n10104 ;
  assign n18745 = ( x109 & ~n9760 ) | ( x109 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n18746 = n18744 | n18745 ;
  assign n18747 = ( x44 & n18538 ) | ( x44 & n18746 ) | ( n18538 & n18746 ) ;
  assign n18748 = ( x44 & ~n18538 ) | ( x44 & n18746 ) | ( ~n18538 & n18746 ) ;
  assign n18749 = ( n18538 & ~n18747 ) | ( n18538 & n18748 ) | ( ~n18747 & n18748 ) ;
  assign n18753 = x110 &  n9457 ;
  assign n18750 = ( x112 & ~n9150 ) | ( x112 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n18751 = x111 &  n9145 ;
  assign n18752 = n18750 | n18751 ;
  assign n18754 = ( x110 & ~n18753 ) | ( x110 & n18752 ) | ( ~n18753 & n18752 ) ;
  assign n18755 = ( n5727 & ~n9153 ) | ( n5727 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n18756 = n18754 | n18755 ;
  assign n18757 = ( x62 & ~n18756 ) | ( x62 & 1'b0 ) | ( ~n18756 & 1'b0 ) ;
  assign n18758 = ~x62 & n18756 ;
  assign n18759 = n18757 | n18758 ;
  assign n18761 = ( n18680 & n18749 ) | ( n18680 & n18759 ) | ( n18749 & n18759 ) ;
  assign n18760 = ( n18680 & ~n18749 ) | ( n18680 & n18759 ) | ( ~n18749 & n18759 ) ;
  assign n18762 = ( n18749 & ~n18761 ) | ( n18749 & n18760 ) | ( ~n18761 & n18760 ) ;
  assign n18766 = x113 &  n8558 ;
  assign n18763 = ( x115 & ~n8314 ) | ( x115 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n18764 = x114 &  n8309 ;
  assign n18765 = n18763 | n18764 ;
  assign n18767 = ( x113 & ~n18766 ) | ( x113 & n18765 ) | ( ~n18766 & n18765 ) ;
  assign n18768 = ( n6420 & ~n8317 ) | ( n6420 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n18769 = n18767 | n18768 ;
  assign n18770 = ( x59 & ~n18769 ) | ( x59 & 1'b0 ) | ( ~n18769 & 1'b0 ) ;
  assign n18771 = ~x59 & n18769 ;
  assign n18772 = n18770 | n18771 ;
  assign n18773 = ( n18684 & n18762 ) | ( n18684 & n18772 ) | ( n18762 & n18772 ) ;
  assign n18774 = ( n18684 & ~n18762 ) | ( n18684 & n18772 ) | ( ~n18762 & n18772 ) ;
  assign n18775 = ( n18762 & ~n18773 ) | ( n18762 & n18774 ) | ( ~n18773 & n18774 ) ;
  assign n18737 = x116 &  n7731 ;
  assign n18734 = ( x118 & ~n7538 ) | ( x118 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n18735 = x117 &  n7533 ;
  assign n18736 = n18734 | n18735 ;
  assign n18738 = ( x116 & ~n18737 ) | ( x116 & n18736 ) | ( ~n18737 & n18736 ) ;
  assign n18739 = n7152 | n7541 ;
  assign n18740 = ~n18738 & n18739 ;
  assign n18741 = x56 &  n18740 ;
  assign n18742 = x56 | n18740 ;
  assign n18743 = ~n18741 & n18742 ;
  assign n18776 = ( n18687 & ~n18775 ) | ( n18687 & n18743 ) | ( ~n18775 & n18743 ) ;
  assign n18777 = ( n18743 & ~n18687 ) | ( n18743 & n18775 ) | ( ~n18687 & n18775 ) ;
  assign n18778 = ( n18776 & ~n18743 ) | ( n18776 & n18777 ) | ( ~n18743 & n18777 ) ;
  assign n18727 = x119 &  n6982 ;
  assign n18724 = ( x121 & ~n6727 ) | ( x121 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n18725 = x120 &  n6722 ;
  assign n18726 = n18724 | n18725 ;
  assign n18728 = ( x119 & ~n18727 ) | ( x119 & n18726 ) | ( ~n18727 & n18726 ) ;
  assign n18729 = ~n6730 & n8176 ;
  assign n18730 = n18728 | n18729 ;
  assign n18731 = ( x53 & ~n18730 ) | ( x53 & 1'b0 ) | ( ~n18730 & 1'b0 ) ;
  assign n18732 = ~x53 & n18730 ;
  assign n18733 = n18731 | n18732 ;
  assign n18779 = ( n18690 & ~n18778 ) | ( n18690 & n18733 ) | ( ~n18778 & n18733 ) ;
  assign n18780 = ( n18733 & ~n18690 ) | ( n18733 & n18778 ) | ( ~n18690 & n18778 ) ;
  assign n18781 = ( n18779 & ~n18733 ) | ( n18779 & n18780 ) | ( ~n18733 & n18780 ) ;
  assign n18782 = ( n18723 & ~n18693 ) | ( n18723 & n18781 ) | ( ~n18693 & n18781 ) ;
  assign n18783 = ( n18693 & ~n18781 ) | ( n18693 & n18723 ) | ( ~n18781 & n18723 ) ;
  assign n18784 = ( n18782 & ~n18723 ) | ( n18782 & n18783 ) | ( ~n18723 & n18783 ) ;
  assign n18795 = ( n18623 & ~n18694 ) | ( n18623 & n18704 ) | ( ~n18694 & n18704 ) ;
  assign n18788 = x125 &  n5586 ;
  assign n18785 = ( x127 & ~n5389 ) | ( x127 & 1'b0 ) | ( ~n5389 & 1'b0 ) ;
  assign n18786 = x126 &  n5384 ;
  assign n18787 = n18785 | n18786 ;
  assign n18789 = ( x125 & ~n18788 ) | ( x125 & n18787 ) | ( ~n18788 & n18787 ) ;
  assign n18790 = n5392 | n9941 ;
  assign n18791 = ~n18789 & n18790 ;
  assign n18792 = x47 &  n18791 ;
  assign n18793 = x47 | n18791 ;
  assign n18794 = ~n18792 & n18793 ;
  assign n18796 = ( n18784 & ~n18795 ) | ( n18784 & n18794 ) | ( ~n18795 & n18794 ) ;
  assign n18797 = ( n18784 & ~n18794 ) | ( n18784 & n18795 ) | ( ~n18794 & n18795 ) ;
  assign n18798 = ( n18796 & ~n18784 ) | ( n18796 & n18797 ) | ( ~n18784 & n18797 ) ;
  assign n18799 = ( n18616 & ~n18615 ) | ( n18616 & n18710 ) | ( ~n18615 & n18710 ) ;
  assign n18800 = ( n18606 & ~n18622 ) | ( n18606 & n18707 ) | ( ~n18622 & n18707 ) ;
  assign n18801 = ( n18798 & n18799 ) | ( n18798 & n18800 ) | ( n18799 & n18800 ) ;
  assign n18802 = ( n18799 & ~n18798 ) | ( n18799 & n18800 ) | ( ~n18798 & n18800 ) ;
  assign n18803 = ( n18798 & ~n18801 ) | ( n18798 & n18802 ) | ( ~n18801 & n18802 ) ;
  assign n18804 = ( n18784 & n18794 ) | ( n18784 & n18795 ) | ( n18794 & n18795 ) ;
  assign n18805 = ( x126 & ~n5586 ) | ( x126 & 1'b0 ) | ( ~n5586 & 1'b0 ) ;
  assign n18806 = x127 &  n5384 ;
  assign n18807 = n18805 | n18806 ;
  assign n18808 = n5392 | n9960 ;
  assign n18809 = ( n18807 & ~n5392 ) | ( n18807 & n18808 ) | ( ~n5392 & n18808 ) ;
  assign n18810 = x47 | n18809 ;
  assign n18811 = ( x47 & ~n18809 ) | ( x47 & 1'b0 ) | ( ~n18809 & 1'b0 ) ;
  assign n18812 = ( n18810 & ~x47 ) | ( n18810 & n18811 ) | ( ~x47 & n18811 ) ;
  assign n18816 = x123 &  n6288 ;
  assign n18813 = ( x125 & ~n6032 ) | ( x125 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n18814 = x124 &  n6027 ;
  assign n18815 = n18813 | n18814 ;
  assign n18817 = ( x123 & ~n18816 ) | ( x123 & n18815 ) | ( ~n18816 & n18815 ) ;
  assign n18818 = ~n6035 & n9324 ;
  assign n18819 = n18817 | n18818 ;
  assign n18821 = x50 &  n18819 ;
  assign n18820 = ~x50 & n18819 ;
  assign n18822 = ( x50 & ~n18821 ) | ( x50 & n18820 ) | ( ~n18821 & n18820 ) ;
  assign n18823 = ( n18762 & ~n18684 ) | ( n18762 & n18772 ) | ( ~n18684 & n18772 ) ;
  assign n18827 = x117 &  n7731 ;
  assign n18824 = ( x119 & ~n7538 ) | ( x119 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n18825 = x118 &  n7533 ;
  assign n18826 = n18824 | n18825 ;
  assign n18828 = ( x117 & ~n18827 ) | ( x117 & n18826 ) | ( ~n18827 & n18826 ) ;
  assign n18829 = ~n7541 & n7648 ;
  assign n18830 = n18828 | n18829 ;
  assign n18831 = ( x56 & ~n18830 ) | ( x56 & 1'b0 ) | ( ~n18830 & 1'b0 ) ;
  assign n18832 = ~x56 & n18830 ;
  assign n18833 = n18831 | n18832 ;
  assign n18834 = ( n18680 & ~n18759 ) | ( n18680 & n18749 ) | ( ~n18759 & n18749 ) ;
  assign n18838 = x114 &  n8558 ;
  assign n18835 = ( x116 & ~n8314 ) | ( x116 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n18836 = x115 &  n8309 ;
  assign n18837 = n18835 | n18836 ;
  assign n18839 = ( x114 & ~n18838 ) | ( x114 & n18837 ) | ( ~n18838 & n18837 ) ;
  assign n18840 = n6885 | n8317 ;
  assign n18841 = ~n18839 & n18840 ;
  assign n18842 = x59 &  n18841 ;
  assign n18843 = x59 | n18841 ;
  assign n18844 = ~n18842 & n18843 ;
  assign n18845 = ( n18538 & ~x44 ) | ( n18538 & n18746 ) | ( ~x44 & n18746 ) ;
  assign n18846 = x109 &  n10104 ;
  assign n18847 = ( x110 & ~n9760 ) | ( x110 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n18848 = n18846 | n18847 ;
  assign n18852 = x111 &  n9457 ;
  assign n18849 = ( x113 & ~n9150 ) | ( x113 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n18850 = x112 &  n9145 ;
  assign n18851 = n18849 | n18850 ;
  assign n18853 = ( x111 & ~n18852 ) | ( x111 & n18851 ) | ( ~n18852 & n18851 ) ;
  assign n18854 = n6169 | n9153 ;
  assign n18855 = ~n18853 & n18854 ;
  assign n18856 = x62 &  n18855 ;
  assign n18857 = x62 | n18855 ;
  assign n18858 = ~n18856 & n18857 ;
  assign n18860 = ( n18845 & n18848 ) | ( n18845 & n18858 ) | ( n18848 & n18858 ) ;
  assign n18859 = ( n18848 & ~n18845 ) | ( n18848 & n18858 ) | ( ~n18845 & n18858 ) ;
  assign n18861 = ( n18845 & ~n18860 ) | ( n18845 & n18859 ) | ( ~n18860 & n18859 ) ;
  assign n18862 = ( n18834 & ~n18844 ) | ( n18834 & n18861 ) | ( ~n18844 & n18861 ) ;
  assign n18863 = ( n18834 & ~n18861 ) | ( n18834 & n18844 ) | ( ~n18861 & n18844 ) ;
  assign n18864 = ( n18862 & ~n18834 ) | ( n18862 & n18863 ) | ( ~n18834 & n18863 ) ;
  assign n18866 = ( n18823 & n18833 ) | ( n18823 & n18864 ) | ( n18833 & n18864 ) ;
  assign n18865 = ( n18833 & ~n18823 ) | ( n18833 & n18864 ) | ( ~n18823 & n18864 ) ;
  assign n18867 = ( n18823 & ~n18866 ) | ( n18823 & n18865 ) | ( ~n18866 & n18865 ) ;
  assign n18871 = x120 &  n6982 ;
  assign n18868 = ( x122 & ~n6727 ) | ( x122 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n18869 = x121 &  n6722 ;
  assign n18870 = n18868 | n18869 ;
  assign n18872 = ( x120 & ~n18871 ) | ( x120 & n18870 ) | ( ~n18871 & n18870 ) ;
  assign n18873 = ~n6730 & n9987 ;
  assign n18874 = n18872 | n18873 ;
  assign n18875 = ( x53 & ~n18874 ) | ( x53 & 1'b0 ) | ( ~n18874 & 1'b0 ) ;
  assign n18876 = ~x53 & n18874 ;
  assign n18877 = n18875 | n18876 ;
  assign n18878 = ( n18777 & n18867 ) | ( n18777 & n18877 ) | ( n18867 & n18877 ) ;
  assign n18879 = ( n18777 & ~n18867 ) | ( n18777 & n18877 ) | ( ~n18867 & n18877 ) ;
  assign n18880 = ( n18867 & ~n18878 ) | ( n18867 & n18879 ) | ( ~n18878 & n18879 ) ;
  assign n18881 = ( n18780 & ~n18822 ) | ( n18780 & n18880 ) | ( ~n18822 & n18880 ) ;
  assign n18882 = ( n18780 & ~n18880 ) | ( n18780 & n18822 ) | ( ~n18880 & n18822 ) ;
  assign n18883 = ( n18881 & ~n18780 ) | ( n18881 & n18882 ) | ( ~n18780 & n18882 ) ;
  assign n18885 = ( n18783 & n18812 ) | ( n18783 & n18883 ) | ( n18812 & n18883 ) ;
  assign n18884 = ( n18783 & ~n18812 ) | ( n18783 & n18883 ) | ( ~n18812 & n18883 ) ;
  assign n18886 = ( n18812 & ~n18885 ) | ( n18812 & n18884 ) | ( ~n18885 & n18884 ) ;
  assign n18887 = ( n18798 & ~n18800 ) | ( n18798 & n18799 ) | ( ~n18800 & n18799 ) ;
  assign n18888 = ( n18804 & ~n18886 ) | ( n18804 & n18887 ) | ( ~n18886 & n18887 ) ;
  assign n18889 = ( n18804 & ~n18887 ) | ( n18804 & n18886 ) | ( ~n18887 & n18886 ) ;
  assign n18890 = ( n18888 & ~n18804 ) | ( n18888 & n18889 ) | ( ~n18804 & n18889 ) ;
  assign n18891 = ( n18783 & ~n18883 ) | ( n18783 & n18812 ) | ( ~n18883 & n18812 ) ;
  assign n18970 = ( n18804 & n18886 ) | ( n18804 & n18887 ) | ( n18886 & n18887 ) ;
  assign n18892 = ( n18867 & ~n18777 ) | ( n18867 & n18877 ) | ( ~n18777 & n18877 ) ;
  assign n18951 = x124 &  n6288 ;
  assign n18948 = ( x126 & ~n6032 ) | ( x126 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n18949 = x125 &  n6027 ;
  assign n18950 = n18948 | n18949 ;
  assign n18952 = ( x124 & ~n18951 ) | ( x124 & n18950 ) | ( ~n18951 & n18950 ) ;
  assign n18953 = n6035 | n9349 ;
  assign n18954 = ~n18952 & n18953 ;
  assign n18955 = x50 &  n18954 ;
  assign n18956 = x50 | n18954 ;
  assign n18957 = ~n18955 & n18956 ;
  assign n18896 = x121 &  n6982 ;
  assign n18893 = ( x123 & ~n6727 ) | ( x123 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n18894 = x122 &  n6722 ;
  assign n18895 = n18893 | n18894 ;
  assign n18897 = ( x121 & ~n18896 ) | ( x121 & n18895 ) | ( ~n18896 & n18895 ) ;
  assign n18898 = ~n6730 & n8472 ;
  assign n18899 = n18897 | n18898 ;
  assign n18900 = ( x53 & ~n18899 ) | ( x53 & 1'b0 ) | ( ~n18899 & 1'b0 ) ;
  assign n18901 = ~x53 & n18899 ;
  assign n18902 = n18900 | n18901 ;
  assign n18906 = x118 &  n7731 ;
  assign n18903 = ( x120 & ~n7538 ) | ( x120 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n18904 = x119 &  n7533 ;
  assign n18905 = n18903 | n18904 ;
  assign n18907 = ( x118 & ~n18906 ) | ( x118 & n18905 ) | ( ~n18906 & n18905 ) ;
  assign n18908 = ~n7541 & n9364 ;
  assign n18909 = n18907 | n18908 ;
  assign n18910 = ( x56 & ~n18909 ) | ( x56 & 1'b0 ) | ( ~n18909 & 1'b0 ) ;
  assign n18911 = ~x56 & n18909 ;
  assign n18912 = n18910 | n18911 ;
  assign n18913 = x110 &  n10104 ;
  assign n18914 = ( x111 & ~n9760 ) | ( x111 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n18915 = n18913 | n18914 ;
  assign n18917 = ( n18848 & n18859 ) | ( n18848 & n18915 ) | ( n18859 & n18915 ) ;
  assign n18916 = ( n18848 & ~n18859 ) | ( n18848 & n18915 ) | ( ~n18859 & n18915 ) ;
  assign n18918 = ( n18859 & ~n18917 ) | ( n18859 & n18916 ) | ( ~n18917 & n18916 ) ;
  assign n18932 = x112 &  n9457 ;
  assign n18929 = ( x114 & ~n9150 ) | ( x114 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n18930 = x113 &  n9145 ;
  assign n18931 = n18929 | n18930 ;
  assign n18933 = ( x112 & ~n18932 ) | ( x112 & n18931 ) | ( ~n18932 & n18931 ) ;
  assign n18934 = n6185 | n9153 ;
  assign n18935 = ~n18933 & n18934 ;
  assign n18936 = x62 &  n18935 ;
  assign n18937 = x62 | n18935 ;
  assign n18938 = ~n18936 & n18937 ;
  assign n18922 = x115 &  n8558 ;
  assign n18919 = ( x117 & ~n8314 ) | ( x117 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n18920 = x116 &  n8309 ;
  assign n18921 = n18919 | n18920 ;
  assign n18923 = ( x115 & ~n18922 ) | ( x115 & n18921 ) | ( ~n18922 & n18921 ) ;
  assign n18924 = n7136 | n8317 ;
  assign n18925 = ~n18923 & n18924 ;
  assign n18926 = x59 &  n18925 ;
  assign n18927 = x59 | n18925 ;
  assign n18928 = ~n18926 & n18927 ;
  assign n18939 = ( n18918 & ~n18938 ) | ( n18918 & n18928 ) | ( ~n18938 & n18928 ) ;
  assign n18940 = ( n18918 & ~n18928 ) | ( n18918 & n18938 ) | ( ~n18928 & n18938 ) ;
  assign n18941 = ( n18939 & ~n18918 ) | ( n18939 & n18940 ) | ( ~n18918 & n18940 ) ;
  assign n18942 = ( n18863 & n18912 ) | ( n18863 & n18941 ) | ( n18912 & n18941 ) ;
  assign n18943 = ( n18912 & ~n18863 ) | ( n18912 & n18941 ) | ( ~n18863 & n18941 ) ;
  assign n18944 = ( n18863 & ~n18942 ) | ( n18863 & n18943 ) | ( ~n18942 & n18943 ) ;
  assign n18945 = ( n18866 & ~n18902 ) | ( n18866 & n18944 ) | ( ~n18902 & n18944 ) ;
  assign n18946 = ( n18866 & ~n18944 ) | ( n18866 & n18902 ) | ( ~n18944 & n18902 ) ;
  assign n18947 = ( n18945 & ~n18866 ) | ( n18945 & n18946 ) | ( ~n18866 & n18946 ) ;
  assign n18958 = ( n18892 & ~n18957 ) | ( n18892 & n18947 ) | ( ~n18957 & n18947 ) ;
  assign n18959 = ( n18892 & ~n18947 ) | ( n18892 & n18957 ) | ( ~n18947 & n18957 ) ;
  assign n18960 = ( n18958 & ~n18892 ) | ( n18958 & n18959 ) | ( ~n18892 & n18959 ) ;
  assign n18961 = ( x127 & ~n5586 ) | ( x127 & 1'b0 ) | ( ~n5586 & 1'b0 ) ;
  assign n18962 = ( n5392 & ~n10258 ) | ( n5392 & n18961 ) | ( ~n10258 & n18961 ) ;
  assign n18963 = n10258 | n18962 ;
  assign n18964 = ( x47 & ~n18961 ) | ( x47 & n18963 ) | ( ~n18961 & n18963 ) ;
  assign n18965 = ( n18961 & ~x47 ) | ( n18961 & n18963 ) | ( ~x47 & n18963 ) ;
  assign n18966 = ( n18964 & ~n18963 ) | ( n18964 & n18965 ) | ( ~n18963 & n18965 ) ;
  assign n18968 = ( n18882 & n18960 ) | ( n18882 & n18966 ) | ( n18960 & n18966 ) ;
  assign n18967 = ( n18960 & ~n18882 ) | ( n18960 & n18966 ) | ( ~n18882 & n18966 ) ;
  assign n18969 = ( n18882 & ~n18968 ) | ( n18882 & n18967 ) | ( ~n18968 & n18967 ) ;
  assign n18971 = ( n18891 & ~n18970 ) | ( n18891 & n18969 ) | ( ~n18970 & n18969 ) ;
  assign n18972 = ( n18891 & ~n18969 ) | ( n18891 & n18970 ) | ( ~n18969 & n18970 ) ;
  assign n18973 = ( n18971 & ~n18891 ) | ( n18971 & n18972 ) | ( ~n18891 & n18972 ) ;
  assign n18974 = ( n18882 & ~n18966 ) | ( n18882 & n18960 ) | ( ~n18966 & n18960 ) ;
  assign n19049 = ( n18969 & ~n18891 ) | ( n18969 & n18970 ) | ( ~n18891 & n18970 ) ;
  assign n18978 = x122 &  n6982 ;
  assign n18975 = ( x124 & ~n6727 ) | ( x124 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n18976 = x123 &  n6722 ;
  assign n18977 = n18975 | n18976 ;
  assign n18979 = ( x122 & ~n18978 ) | ( x122 & n18977 ) | ( ~n18978 & n18977 ) ;
  assign n18980 = ~n6730 & n8755 ;
  assign n18981 = n18979 | n18980 ;
  assign n18982 = ( x53 & ~n18981 ) | ( x53 & 1'b0 ) | ( ~n18981 & 1'b0 ) ;
  assign n18983 = ~x53 & n18981 ;
  assign n18984 = n18982 | n18983 ;
  assign n18988 = x119 &  n7731 ;
  assign n18985 = ( x121 & ~n7538 ) | ( x121 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n18986 = x120 &  n7533 ;
  assign n18987 = n18985 | n18986 ;
  assign n18989 = ( x119 & ~n18988 ) | ( x119 & n18987 ) | ( ~n18988 & n18987 ) ;
  assign n18990 = ~n7541 & n8176 ;
  assign n18991 = n18989 | n18990 ;
  assign n18992 = ( x56 & ~n18991 ) | ( x56 & 1'b0 ) | ( ~n18991 & 1'b0 ) ;
  assign n18993 = ~x56 & n18991 ;
  assign n18994 = n18992 | n18993 ;
  assign n18998 = x113 &  n9457 ;
  assign n18995 = ( x115 & ~n9150 ) | ( x115 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n18996 = x114 &  n9145 ;
  assign n18997 = n18995 | n18996 ;
  assign n18999 = ( x113 & ~n18998 ) | ( x113 & n18997 ) | ( ~n18998 & n18997 ) ;
  assign n19000 = ( n6420 & ~n9153 ) | ( n6420 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n19001 = n18999 | n19000 ;
  assign n19002 = ( x62 & ~n19001 ) | ( x62 & 1'b0 ) | ( ~n19001 & 1'b0 ) ;
  assign n19003 = ~x62 & n19001 ;
  assign n19004 = n19002 | n19003 ;
  assign n19005 = ( n18859 & ~n18848 ) | ( n18859 & n18915 ) | ( ~n18848 & n18915 ) ;
  assign n19006 = x111 &  n10104 ;
  assign n19007 = ( x112 & ~n9760 ) | ( x112 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n19008 = n19006 | n19007 ;
  assign n19009 = ( x47 & n18915 ) | ( x47 & n19008 ) | ( n18915 & n19008 ) ;
  assign n19010 = ( x47 & ~n18915 ) | ( x47 & n19008 ) | ( ~n18915 & n19008 ) ;
  assign n19011 = ( n18915 & ~n19009 ) | ( n18915 & n19010 ) | ( ~n19009 & n19010 ) ;
  assign n19012 = ( n19004 & n19005 ) | ( n19004 & n19011 ) | ( n19005 & n19011 ) ;
  assign n19013 = ( n19005 & ~n19004 ) | ( n19005 & n19011 ) | ( ~n19004 & n19011 ) ;
  assign n19014 = ( n19004 & ~n19012 ) | ( n19004 & n19013 ) | ( ~n19012 & n19013 ) ;
  assign n19019 = x116 &  n8558 ;
  assign n19016 = ( x118 & ~n8314 ) | ( x118 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n19017 = x117 &  n8309 ;
  assign n19018 = n19016 | n19017 ;
  assign n19020 = ( x116 & ~n19019 ) | ( x116 & n19018 ) | ( ~n19019 & n19018 ) ;
  assign n19021 = n7152 | n8317 ;
  assign n19022 = ~n19020 & n19021 ;
  assign n19023 = x59 &  n19022 ;
  assign n19024 = x59 | n19022 ;
  assign n19025 = ~n19023 & n19024 ;
  assign n19015 = ( n18928 & ~n18918 ) | ( n18928 & n18938 ) | ( ~n18918 & n18938 ) ;
  assign n19026 = ( n19014 & ~n19025 ) | ( n19014 & n19015 ) | ( ~n19025 & n19015 ) ;
  assign n19027 = ( n19014 & ~n19015 ) | ( n19014 & n19025 ) | ( ~n19015 & n19025 ) ;
  assign n19028 = ( n19026 & ~n19014 ) | ( n19026 & n19027 ) | ( ~n19014 & n19027 ) ;
  assign n19030 = ( n18943 & n18994 ) | ( n18943 & n19028 ) | ( n18994 & n19028 ) ;
  assign n19029 = ( n18943 & ~n18994 ) | ( n18943 & n19028 ) | ( ~n18994 & n19028 ) ;
  assign n19031 = ( n18994 & ~n19030 ) | ( n18994 & n19029 ) | ( ~n19030 & n19029 ) ;
  assign n19033 = ( n18946 & n18984 ) | ( n18946 & n19031 ) | ( n18984 & n19031 ) ;
  assign n19032 = ( n18946 & ~n18984 ) | ( n18946 & n19031 ) | ( ~n18984 & n19031 ) ;
  assign n19034 = ( n18984 & ~n19033 ) | ( n18984 & n19032 ) | ( ~n19033 & n19032 ) ;
  assign n19038 = x125 &  n6288 ;
  assign n19035 = ( x127 & ~n6032 ) | ( x127 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n19036 = x126 &  n6027 ;
  assign n19037 = n19035 | n19036 ;
  assign n19039 = ( x125 & ~n19038 ) | ( x125 & n19037 ) | ( ~n19038 & n19037 ) ;
  assign n19040 = n6035 | n9941 ;
  assign n19041 = ~n19039 & n19040 ;
  assign n19042 = x50 &  n19041 ;
  assign n19043 = x50 | n19041 ;
  assign n19044 = ~n19042 & n19043 ;
  assign n19045 = ( n18947 & ~n18892 ) | ( n18947 & n18957 ) | ( ~n18892 & n18957 ) ;
  assign n19046 = ( n19034 & ~n19044 ) | ( n19034 & n19045 ) | ( ~n19044 & n19045 ) ;
  assign n19047 = ( n19034 & ~n19045 ) | ( n19034 & n19044 ) | ( ~n19045 & n19044 ) ;
  assign n19048 = ( n19046 & ~n19034 ) | ( n19046 & n19047 ) | ( ~n19034 & n19047 ) ;
  assign n19050 = ( n18974 & ~n19049 ) | ( n18974 & n19048 ) | ( ~n19049 & n19048 ) ;
  assign n19051 = ( n18974 & ~n19048 ) | ( n18974 & n19049 ) | ( ~n19048 & n19049 ) ;
  assign n19052 = ( n19050 & ~n18974 ) | ( n19050 & n19051 ) | ( ~n18974 & n19051 ) ;
  assign n19053 = ( n19044 & ~n19034 ) | ( n19044 & n19045 ) | ( ~n19034 & n19045 ) ;
  assign n19057 = x123 &  n6982 ;
  assign n19054 = ( x125 & ~n6727 ) | ( x125 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n19055 = x124 &  n6722 ;
  assign n19056 = n19054 | n19055 ;
  assign n19058 = ( x123 & ~n19057 ) | ( x123 & n19056 ) | ( ~n19057 & n19056 ) ;
  assign n19059 = ~n6730 & n9324 ;
  assign n19060 = n19058 | n19059 ;
  assign n19061 = ( x53 & ~n19060 ) | ( x53 & 1'b0 ) | ( ~n19060 & 1'b0 ) ;
  assign n19062 = ~x53 & n19060 ;
  assign n19063 = n19061 | n19062 ;
  assign n19064 = ( n19015 & ~n19014 ) | ( n19015 & n19025 ) | ( ~n19014 & n19025 ) ;
  assign n19078 = x117 &  n8558 ;
  assign n19075 = ( x119 & ~n8314 ) | ( x119 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n19076 = x118 &  n8309 ;
  assign n19077 = n19075 | n19076 ;
  assign n19079 = ( x117 & ~n19078 ) | ( x117 & n19077 ) | ( ~n19078 & n19077 ) ;
  assign n19080 = ( n7648 & ~n8317 ) | ( n7648 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n19081 = n19079 | n19080 ;
  assign n19082 = ( x59 & ~n19081 ) | ( x59 & 1'b0 ) | ( ~n19081 & 1'b0 ) ;
  assign n19083 = ~x59 & n19081 ;
  assign n19084 = n19082 | n19083 ;
  assign n19085 = ( n18915 & ~x47 ) | ( n18915 & n19008 ) | ( ~x47 & n19008 ) ;
  assign n19086 = x112 &  n10104 ;
  assign n19087 = ( x113 & ~n9760 ) | ( x113 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n19088 = n19086 | n19087 ;
  assign n19092 = x114 &  n9457 ;
  assign n19089 = ( x116 & ~n9150 ) | ( x116 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n19090 = x115 &  n9145 ;
  assign n19091 = n19089 | n19090 ;
  assign n19093 = ( x114 & ~n19092 ) | ( x114 & n19091 ) | ( ~n19092 & n19091 ) ;
  assign n19094 = ( n6885 & ~n9153 ) | ( n6885 & n19093 ) | ( ~n9153 & n19093 ) ;
  assign n19095 = n9153 | n19094 ;
  assign n19097 = ( x62 & n19093 ) | ( x62 & n19095 ) | ( n19093 & n19095 ) ;
  assign n19096 = ( x62 & ~n19095 ) | ( x62 & n19093 ) | ( ~n19095 & n19093 ) ;
  assign n19098 = ( n19095 & ~n19097 ) | ( n19095 & n19096 ) | ( ~n19097 & n19096 ) ;
  assign n19100 = ( n19085 & n19088 ) | ( n19085 & n19098 ) | ( n19088 & n19098 ) ;
  assign n19099 = ( n19088 & ~n19085 ) | ( n19088 & n19098 ) | ( ~n19085 & n19098 ) ;
  assign n19101 = ( n19085 & ~n19100 ) | ( n19085 & n19099 ) | ( ~n19100 & n19099 ) ;
  assign n19102 = ( n19013 & n19084 ) | ( n19013 & n19101 ) | ( n19084 & n19101 ) ;
  assign n19103 = ( n19084 & ~n19013 ) | ( n19084 & n19101 ) | ( ~n19013 & n19101 ) ;
  assign n19104 = ( n19013 & ~n19102 ) | ( n19013 & n19103 ) | ( ~n19102 & n19103 ) ;
  assign n19068 = x120 &  n7731 ;
  assign n19065 = ( x122 & ~n7538 ) | ( x122 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n19066 = x121 &  n7533 ;
  assign n19067 = n19065 | n19066 ;
  assign n19069 = ( x120 & ~n19068 ) | ( x120 & n19067 ) | ( ~n19068 & n19067 ) ;
  assign n19070 = ~n7541 & n9987 ;
  assign n19071 = n19069 | n19070 ;
  assign n19072 = ( x56 & ~n19071 ) | ( x56 & 1'b0 ) | ( ~n19071 & 1'b0 ) ;
  assign n19073 = ~x56 & n19071 ;
  assign n19074 = n19072 | n19073 ;
  assign n19105 = ( n19064 & ~n19104 ) | ( n19064 & n19074 ) | ( ~n19104 & n19074 ) ;
  assign n19106 = ( n19064 & ~n19074 ) | ( n19064 & n19104 ) | ( ~n19074 & n19104 ) ;
  assign n19107 = ( n19105 & ~n19064 ) | ( n19105 & n19106 ) | ( ~n19064 & n19106 ) ;
  assign n19109 = ( n19030 & n19063 ) | ( n19030 & n19107 ) | ( n19063 & n19107 ) ;
  assign n19108 = ( n19063 & ~n19030 ) | ( n19063 & n19107 ) | ( ~n19030 & n19107 ) ;
  assign n19110 = ( n19030 & ~n19109 ) | ( n19030 & n19108 ) | ( ~n19109 & n19108 ) ;
  assign n19111 = ( x126 & ~n6288 ) | ( x126 & 1'b0 ) | ( ~n6288 & 1'b0 ) ;
  assign n19112 = x127 &  n6027 ;
  assign n19113 = n19111 | n19112 ;
  assign n19114 = n6035 | n9960 ;
  assign n19115 = ( n19113 & ~n6035 ) | ( n19113 & n19114 ) | ( ~n6035 & n19114 ) ;
  assign n19116 = x50 | n19033 ;
  assign n19117 = ~x50 & n19033 ;
  assign n19118 = ( n19116 & ~n19033 ) | ( n19116 & n19117 ) | ( ~n19033 & n19117 ) ;
  assign n19119 = ( n19110 & ~n19115 ) | ( n19110 & n19118 ) | ( ~n19115 & n19118 ) ;
  assign n19120 = ( n19115 & ~n19110 ) | ( n19115 & n19118 ) | ( ~n19110 & n19118 ) ;
  assign n19121 = ( n19119 & ~n19118 ) | ( n19119 & n19120 ) | ( ~n19118 & n19120 ) ;
  assign n19122 = ( n19053 & ~n19050 ) | ( n19053 & n19121 ) | ( ~n19050 & n19121 ) ;
  assign n19123 = ( n19050 & ~n19121 ) | ( n19050 & n19053 ) | ( ~n19121 & n19053 ) ;
  assign n19124 = ( n19122 & ~n19053 ) | ( n19122 & n19123 ) | ( ~n19053 & n19123 ) ;
  assign n19125 = x50 | n19115 ;
  assign n19126 = x50 &  n19115 ;
  assign n19127 = ( n19125 & ~n19126 ) | ( n19125 & 1'b0 ) | ( ~n19126 & 1'b0 ) ;
  assign n19128 = ( n19033 & n19110 ) | ( n19033 & n19127 ) | ( n19110 & n19127 ) ;
  assign n19184 = ( x127 & ~n6288 ) | ( x127 & 1'b0 ) | ( ~n6288 & 1'b0 ) ;
  assign n19185 = ( n6035 & ~n10258 ) | ( n6035 & n19184 ) | ( ~n10258 & n19184 ) ;
  assign n19186 = n10258 | n19185 ;
  assign n19187 = ( x50 & ~n19184 ) | ( x50 & n19186 ) | ( ~n19184 & n19186 ) ;
  assign n19188 = ( n19184 & ~x50 ) | ( n19184 & n19186 ) | ( ~x50 & n19186 ) ;
  assign n19189 = ( n19187 & ~n19186 ) | ( n19187 & n19188 ) | ( ~n19186 & n19188 ) ;
  assign n19132 = x121 &  n7731 ;
  assign n19129 = ( x123 & ~n7538 ) | ( x123 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n19130 = x122 &  n7533 ;
  assign n19131 = n19129 | n19130 ;
  assign n19133 = ( x121 & ~n19132 ) | ( x121 & n19131 ) | ( ~n19132 & n19131 ) ;
  assign n19134 = ~n7541 & n8472 ;
  assign n19135 = n19133 | n19134 ;
  assign n19136 = ( x56 & ~n19135 ) | ( x56 & 1'b0 ) | ( ~n19135 & 1'b0 ) ;
  assign n19137 = ~x56 & n19135 ;
  assign n19138 = n19136 | n19137 ;
  assign n19158 = x118 &  n8558 ;
  assign n19155 = ( x120 & ~n8314 ) | ( x120 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n19156 = x119 &  n8309 ;
  assign n19157 = n19155 | n19156 ;
  assign n19159 = ( x118 & ~n19158 ) | ( x118 & n19157 ) | ( ~n19158 & n19157 ) ;
  assign n19160 = ~n8317 & n9364 ;
  assign n19161 = n19159 | n19160 ;
  assign n19162 = ( x59 & ~n19161 ) | ( x59 & 1'b0 ) | ( ~n19161 & 1'b0 ) ;
  assign n19163 = ~x59 & n19161 ;
  assign n19164 = n19162 | n19163 ;
  assign n19149 = x113 &  n10104 ;
  assign n19150 = ( x114 & ~n9760 ) | ( x114 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n19151 = n19149 | n19150 ;
  assign n19142 = x115 &  n9457 ;
  assign n19139 = ( x117 & ~n9150 ) | ( x117 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n19140 = x116 &  n9145 ;
  assign n19141 = n19139 | n19140 ;
  assign n19143 = ( x115 & ~n19142 ) | ( x115 & n19141 ) | ( ~n19142 & n19141 ) ;
  assign n19144 = n7136 | n9153 ;
  assign n19145 = ~n19143 & n19144 ;
  assign n19146 = x62 &  n19145 ;
  assign n19147 = x62 | n19145 ;
  assign n19148 = ~n19146 & n19147 ;
  assign n19152 = ( n19088 & ~n19151 ) | ( n19088 & n19148 ) | ( ~n19151 & n19148 ) ;
  assign n19153 = ( n19148 & ~n19088 ) | ( n19148 & n19151 ) | ( ~n19088 & n19151 ) ;
  assign n19154 = ( n19152 & ~n19148 ) | ( n19152 & n19153 ) | ( ~n19148 & n19153 ) ;
  assign n19165 = ( n19099 & ~n19164 ) | ( n19099 & n19154 ) | ( ~n19164 & n19154 ) ;
  assign n19166 = ( n19099 & ~n19154 ) | ( n19099 & n19164 ) | ( ~n19154 & n19164 ) ;
  assign n19167 = ( n19165 & ~n19099 ) | ( n19165 & n19166 ) | ( ~n19099 & n19166 ) ;
  assign n19168 = ( n19103 & ~n19138 ) | ( n19103 & n19167 ) | ( ~n19138 & n19167 ) ;
  assign n19169 = ( n19103 & ~n19167 ) | ( n19103 & n19138 ) | ( ~n19167 & n19138 ) ;
  assign n19170 = ( n19168 & ~n19103 ) | ( n19168 & n19169 ) | ( ~n19103 & n19169 ) ;
  assign n19174 = x124 &  n6982 ;
  assign n19171 = ( x126 & ~n6727 ) | ( x126 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n19172 = x125 &  n6722 ;
  assign n19173 = n19171 | n19172 ;
  assign n19175 = ( x124 & ~n19174 ) | ( x124 & n19173 ) | ( ~n19174 & n19173 ) ;
  assign n19176 = n6730 | n9349 ;
  assign n19177 = ~n19175 & n19176 ;
  assign n19178 = x53 &  n19177 ;
  assign n19179 = x53 | n19177 ;
  assign n19180 = ~n19178 & n19179 ;
  assign n19181 = ( n19106 & ~n19170 ) | ( n19106 & n19180 ) | ( ~n19170 & n19180 ) ;
  assign n19182 = ( n19106 & ~n19180 ) | ( n19106 & n19170 ) | ( ~n19180 & n19170 ) ;
  assign n19183 = ( n19181 & ~n19106 ) | ( n19181 & n19182 ) | ( ~n19106 & n19182 ) ;
  assign n19190 = ( n19109 & ~n19189 ) | ( n19109 & n19183 ) | ( ~n19189 & n19183 ) ;
  assign n19191 = ( n19109 & ~n19183 ) | ( n19109 & n19189 ) | ( ~n19183 & n19189 ) ;
  assign n19192 = ( n19190 & ~n19109 ) | ( n19190 & n19191 ) | ( ~n19109 & n19191 ) ;
  assign n19193 = ( n19050 & ~n19053 ) | ( n19050 & n19121 ) | ( ~n19053 & n19121 ) ;
  assign n19194 = ( n19128 & ~n19192 ) | ( n19128 & n19193 ) | ( ~n19192 & n19193 ) ;
  assign n19195 = ( n19128 & ~n19193 ) | ( n19128 & n19192 ) | ( ~n19193 & n19192 ) ;
  assign n19196 = ( n19194 & ~n19128 ) | ( n19194 & n19195 ) | ( ~n19128 & n19195 ) ;
  assign n19197 = ( n19183 & ~n19109 ) | ( n19183 & n19189 ) | ( ~n19109 & n19189 ) ;
  assign n19258 = ( n19128 & n19192 ) | ( n19128 & n19193 ) | ( n19192 & n19193 ) ;
  assign n19201 = x125 &  n6982 ;
  assign n19198 = ( x127 & ~n6727 ) | ( x127 & 1'b0 ) | ( ~n6727 & 1'b0 ) ;
  assign n19199 = x126 &  n6722 ;
  assign n19200 = n19198 | n19199 ;
  assign n19202 = ( x125 & ~n19201 ) | ( x125 & n19200 ) | ( ~n19201 & n19200 ) ;
  assign n19203 = n6730 | n9941 ;
  assign n19204 = ~n19202 & n19203 ;
  assign n19205 = x53 &  n19204 ;
  assign n19206 = x53 | n19204 ;
  assign n19207 = ~n19205 & n19206 ;
  assign n19211 = x122 &  n7731 ;
  assign n19208 = ( x124 & ~n7538 ) | ( x124 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n19209 = x123 &  n7533 ;
  assign n19210 = n19208 | n19209 ;
  assign n19212 = ( x122 & ~n19211 ) | ( x122 & n19210 ) | ( ~n19211 & n19210 ) ;
  assign n19213 = ~n7541 & n8755 ;
  assign n19214 = n19212 | n19213 ;
  assign n19215 = ( x56 & ~n19214 ) | ( x56 & 1'b0 ) | ( ~n19214 & 1'b0 ) ;
  assign n19216 = ~x56 & n19214 ;
  assign n19217 = n19215 | n19216 ;
  assign n19221 = x119 &  n8558 ;
  assign n19218 = ( x121 & ~n8314 ) | ( x121 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n19219 = x120 &  n8309 ;
  assign n19220 = n19218 | n19219 ;
  assign n19222 = ( x119 & ~n19221 ) | ( x119 & n19220 ) | ( ~n19221 & n19220 ) ;
  assign n19223 = ( n8176 & ~n8317 ) | ( n8176 & 1'b0 ) | ( ~n8317 & 1'b0 ) ;
  assign n19224 = n19222 | n19223 ;
  assign n19225 = ( x59 & ~n19224 ) | ( x59 & 1'b0 ) | ( ~n19224 & 1'b0 ) ;
  assign n19226 = ~x59 & n19224 ;
  assign n19227 = n19225 | n19226 ;
  assign n19228 = ( n19154 & ~n19099 ) | ( n19154 & n19164 ) | ( ~n19099 & n19164 ) ;
  assign n19232 = x116 &  n9457 ;
  assign n19229 = ( x118 & ~n9150 ) | ( x118 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n19230 = x117 &  n9145 ;
  assign n19231 = n19229 | n19230 ;
  assign n19233 = ( x116 & ~n19232 ) | ( x116 & n19231 ) | ( ~n19232 & n19231 ) ;
  assign n19234 = n7152 | n9153 ;
  assign n19235 = ~n19233 & n19234 ;
  assign n19236 = x62 &  n19235 ;
  assign n19237 = x62 | n19235 ;
  assign n19238 = ~n19236 & n19237 ;
  assign n19239 = x114 &  n10104 ;
  assign n19240 = ( x115 & ~n9760 ) | ( x115 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n19241 = n19239 | n19240 ;
  assign n19242 = ( x50 & n19088 ) | ( x50 & n19241 ) | ( n19088 & n19241 ) ;
  assign n19243 = ( x50 & ~n19088 ) | ( x50 & n19241 ) | ( ~n19088 & n19241 ) ;
  assign n19244 = ( n19088 & ~n19242 ) | ( n19088 & n19243 ) | ( ~n19242 & n19243 ) ;
  assign n19246 = ( n19152 & n19238 ) | ( n19152 & n19244 ) | ( n19238 & n19244 ) ;
  assign n19245 = ( n19238 & ~n19152 ) | ( n19238 & n19244 ) | ( ~n19152 & n19244 ) ;
  assign n19247 = ( n19152 & ~n19246 ) | ( n19152 & n19245 ) | ( ~n19246 & n19245 ) ;
  assign n19248 = ( n19227 & ~n19228 ) | ( n19227 & n19247 ) | ( ~n19228 & n19247 ) ;
  assign n19249 = ( n19227 & ~n19247 ) | ( n19227 & n19228 ) | ( ~n19247 & n19228 ) ;
  assign n19250 = ( n19248 & ~n19227 ) | ( n19248 & n19249 ) | ( ~n19227 & n19249 ) ;
  assign n19251 = ( n19217 & ~n19169 ) | ( n19217 & n19250 ) | ( ~n19169 & n19250 ) ;
  assign n19252 = ( n19169 & ~n19250 ) | ( n19169 & n19217 ) | ( ~n19250 & n19217 ) ;
  assign n19253 = ( n19251 & ~n19217 ) | ( n19251 & n19252 ) | ( ~n19217 & n19252 ) ;
  assign n19254 = ( n19106 & n19170 ) | ( n19106 & n19180 ) | ( n19170 & n19180 ) ;
  assign n19255 = ( n19207 & n19253 ) | ( n19207 & n19254 ) | ( n19253 & n19254 ) ;
  assign n19256 = ( n19253 & ~n19207 ) | ( n19253 & n19254 ) | ( ~n19207 & n19254 ) ;
  assign n19257 = ( n19207 & ~n19255 ) | ( n19207 & n19256 ) | ( ~n19255 & n19256 ) ;
  assign n19259 = ( n19197 & ~n19258 ) | ( n19197 & n19257 ) | ( ~n19258 & n19257 ) ;
  assign n19260 = ( n19197 & ~n19257 ) | ( n19197 & n19258 ) | ( ~n19257 & n19258 ) ;
  assign n19261 = ( n19259 & ~n19197 ) | ( n19259 & n19260 ) | ( ~n19197 & n19260 ) ;
  assign n19265 = x123 &  n7731 ;
  assign n19262 = ( x125 & ~n7538 ) | ( x125 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n19263 = x124 &  n7533 ;
  assign n19264 = n19262 | n19263 ;
  assign n19266 = ( x123 & ~n19265 ) | ( x123 & n19264 ) | ( ~n19265 & n19264 ) ;
  assign n19267 = ~n7541 & n9324 ;
  assign n19268 = n19266 | n19267 ;
  assign n19269 = ( x56 & ~n19268 ) | ( x56 & 1'b0 ) | ( ~n19268 & 1'b0 ) ;
  assign n19270 = ~x56 & n19268 ;
  assign n19271 = n19269 | n19270 ;
  assign n19282 = ( n19088 & ~x50 ) | ( n19088 & n19241 ) | ( ~x50 & n19241 ) ;
  assign n19283 = x115 &  n10104 ;
  assign n19284 = ( x116 & ~n9760 ) | ( x116 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n19285 = n19283 | n19284 ;
  assign n19289 = x117 &  n9457 ;
  assign n19286 = ( x119 & ~n9150 ) | ( x119 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n19287 = x118 &  n9145 ;
  assign n19288 = n19286 | n19287 ;
  assign n19290 = ( x117 & ~n19289 ) | ( x117 & n19288 ) | ( ~n19289 & n19288 ) ;
  assign n19291 = ( n7648 & ~n9153 ) | ( n7648 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n19292 = n19290 | n19291 ;
  assign n19293 = ( x62 & ~n19292 ) | ( x62 & 1'b0 ) | ( ~n19292 & 1'b0 ) ;
  assign n19294 = ~x62 & n19292 ;
  assign n19295 = n19293 | n19294 ;
  assign n19296 = ( n19282 & ~n19285 ) | ( n19282 & n19295 ) | ( ~n19285 & n19295 ) ;
  assign n19297 = ( n19282 & ~n19295 ) | ( n19282 & n19285 ) | ( ~n19295 & n19285 ) ;
  assign n19298 = ( n19296 & ~n19282 ) | ( n19296 & n19297 ) | ( ~n19282 & n19297 ) ;
  assign n19275 = x120 &  n8558 ;
  assign n19272 = ( x122 & ~n8314 ) | ( x122 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n19273 = x121 &  n8309 ;
  assign n19274 = n19272 | n19273 ;
  assign n19276 = ( x120 & ~n19275 ) | ( x120 & n19274 ) | ( ~n19275 & n19274 ) ;
  assign n19277 = ~n8317 & n9987 ;
  assign n19278 = n19276 | n19277 ;
  assign n19279 = ( x59 & ~n19278 ) | ( x59 & 1'b0 ) | ( ~n19278 & 1'b0 ) ;
  assign n19280 = ~x59 & n19278 ;
  assign n19281 = n19279 | n19280 ;
  assign n19299 = ( n19246 & ~n19298 ) | ( n19246 & n19281 ) | ( ~n19298 & n19281 ) ;
  assign n19300 = ( n19246 & ~n19281 ) | ( n19246 & n19298 ) | ( ~n19281 & n19298 ) ;
  assign n19301 = ( n19299 & ~n19246 ) | ( n19299 & n19300 ) | ( ~n19246 & n19300 ) ;
  assign n19303 = ( n19249 & n19271 ) | ( n19249 & n19301 ) | ( n19271 & n19301 ) ;
  assign n19302 = ( n19271 & ~n19249 ) | ( n19271 & n19301 ) | ( ~n19249 & n19301 ) ;
  assign n19304 = ( n19249 & ~n19303 ) | ( n19249 & n19302 ) | ( ~n19303 & n19302 ) ;
  assign n19305 = ( x126 & ~n6982 ) | ( x126 & 1'b0 ) | ( ~n6982 & 1'b0 ) ;
  assign n19306 = x127 &  n6722 ;
  assign n19307 = n19305 | n19306 ;
  assign n19308 = n6730 | n9960 ;
  assign n19309 = ( n19307 & ~n6730 ) | ( n19307 & n19308 ) | ( ~n6730 & n19308 ) ;
  assign n19310 = x53 | n19252 ;
  assign n19311 = ~x53 & n19252 ;
  assign n19312 = ( n19310 & ~n19252 ) | ( n19310 & n19311 ) | ( ~n19252 & n19311 ) ;
  assign n19313 = ( n19304 & ~n19309 ) | ( n19304 & n19312 ) | ( ~n19309 & n19312 ) ;
  assign n19314 = ( n19309 & ~n19304 ) | ( n19309 & n19312 ) | ( ~n19304 & n19312 ) ;
  assign n19315 = ( n19313 & ~n19312 ) | ( n19313 & n19314 ) | ( ~n19312 & n19314 ) ;
  assign n19316 = ( n19255 & n19259 ) | ( n19255 & n19315 ) | ( n19259 & n19315 ) ;
  assign n19317 = ( n19259 & ~n19255 ) | ( n19259 & n19315 ) | ( ~n19255 & n19315 ) ;
  assign n19318 = ( n19255 & ~n19316 ) | ( n19255 & n19317 ) | ( ~n19316 & n19317 ) ;
  assign n19319 = x53 | n19309 ;
  assign n19320 = x53 &  n19309 ;
  assign n19321 = ( n19319 & ~n19320 ) | ( n19319 & 1'b0 ) | ( ~n19320 & 1'b0 ) ;
  assign n19322 = ( n19252 & n19304 ) | ( n19252 & n19321 ) | ( n19304 & n19321 ) ;
  assign n19365 = ( x127 & ~n6982 ) | ( x127 & 1'b0 ) | ( ~n6982 & 1'b0 ) ;
  assign n19366 = ( n6730 & ~n10258 ) | ( n6730 & n19365 ) | ( ~n10258 & n19365 ) ;
  assign n19367 = n10258 | n19366 ;
  assign n19368 = ( x53 & ~n19365 ) | ( x53 & n19367 ) | ( ~n19365 & n19367 ) ;
  assign n19369 = ( n19365 & ~x53 ) | ( n19365 & n19367 ) | ( ~x53 & n19367 ) ;
  assign n19370 = ( n19368 & ~n19367 ) | ( n19368 & n19369 ) | ( ~n19367 & n19369 ) ;
  assign n19355 = x124 &  n7731 ;
  assign n19352 = ( x126 & ~n7538 ) | ( x126 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n19353 = x125 &  n7533 ;
  assign n19354 = n19352 | n19353 ;
  assign n19356 = ( x124 & ~n19355 ) | ( x124 & n19354 ) | ( ~n19355 & n19354 ) ;
  assign n19357 = n7541 | n9349 ;
  assign n19358 = ~n19356 & n19357 ;
  assign n19359 = x56 &  n19358 ;
  assign n19360 = x56 | n19358 ;
  assign n19361 = ~n19359 & n19360 ;
  assign n19326 = x118 &  n9457 ;
  assign n19323 = ( x120 & ~n9150 ) | ( x120 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n19324 = x119 &  n9145 ;
  assign n19325 = n19323 | n19324 ;
  assign n19327 = ( x118 & ~n19326 ) | ( x118 & n19325 ) | ( ~n19326 & n19325 ) ;
  assign n19328 = ~n9153 & n9364 ;
  assign n19329 = n19327 | n19328 ;
  assign n19330 = ( x62 & ~n19329 ) | ( x62 & 1'b0 ) | ( ~n19329 & 1'b0 ) ;
  assign n19331 = ~x62 & n19329 ;
  assign n19332 = n19330 | n19331 ;
  assign n19333 = x116 &  n10104 ;
  assign n19334 = ( x117 & ~n9760 ) | ( x117 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n19335 = n19333 | n19334 ;
  assign n19336 = ( n19285 & n19296 ) | ( n19285 & n19335 ) | ( n19296 & n19335 ) ;
  assign n19337 = ( n19285 & ~n19296 ) | ( n19285 & n19335 ) | ( ~n19296 & n19335 ) ;
  assign n19338 = ( n19296 & ~n19336 ) | ( n19296 & n19337 ) | ( ~n19336 & n19337 ) ;
  assign n19342 = x121 &  n8558 ;
  assign n19339 = ( x123 & ~n8314 ) | ( x123 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n19340 = x122 &  n8309 ;
  assign n19341 = n19339 | n19340 ;
  assign n19343 = ( x121 & ~n19342 ) | ( x121 & n19341 ) | ( ~n19342 & n19341 ) ;
  assign n19344 = ~n8317 & n8472 ;
  assign n19345 = n19343 | n19344 ;
  assign n19346 = ( x59 & ~n19345 ) | ( x59 & 1'b0 ) | ( ~n19345 & 1'b0 ) ;
  assign n19347 = ~x59 & n19345 ;
  assign n19348 = n19346 | n19347 ;
  assign n19349 = ( n19332 & n19338 ) | ( n19332 & n19348 ) | ( n19338 & n19348 ) ;
  assign n19350 = ( n19338 & ~n19332 ) | ( n19338 & n19348 ) | ( ~n19332 & n19348 ) ;
  assign n19351 = ( n19332 & ~n19349 ) | ( n19332 & n19350 ) | ( ~n19349 & n19350 ) ;
  assign n19362 = ( n19300 & ~n19361 ) | ( n19300 & n19351 ) | ( ~n19361 & n19351 ) ;
  assign n19363 = ( n19351 & ~n19300 ) | ( n19351 & n19361 ) | ( ~n19300 & n19361 ) ;
  assign n19364 = ( n19362 & ~n19351 ) | ( n19362 & n19363 ) | ( ~n19351 & n19363 ) ;
  assign n19371 = ( n19303 & ~n19370 ) | ( n19303 & n19364 ) | ( ~n19370 & n19364 ) ;
  assign n19372 = ( n19303 & ~n19364 ) | ( n19303 & n19370 ) | ( ~n19364 & n19370 ) ;
  assign n19373 = ( n19371 & ~n19303 ) | ( n19371 & n19372 ) | ( ~n19303 & n19372 ) ;
  assign n19374 = ( n19255 & ~n19315 ) | ( n19255 & n19259 ) | ( ~n19315 & n19259 ) ;
  assign n19376 = ( n19322 & n19373 ) | ( n19322 & n19374 ) | ( n19373 & n19374 ) ;
  assign n19375 = ( n19373 & ~n19322 ) | ( n19373 & n19374 ) | ( ~n19322 & n19374 ) ;
  assign n19377 = ( n19322 & ~n19376 ) | ( n19322 & n19375 ) | ( ~n19376 & n19375 ) ;
  assign n19378 = ( n19364 & ~n19303 ) | ( n19364 & n19370 ) | ( ~n19303 & n19370 ) ;
  assign n19379 = ( n19322 & ~n19374 ) | ( n19322 & n19373 ) | ( ~n19374 & n19373 ) ;
  assign n19383 = x125 &  n7731 ;
  assign n19380 = ( x127 & ~n7538 ) | ( x127 & 1'b0 ) | ( ~n7538 & 1'b0 ) ;
  assign n19381 = x126 &  n7533 ;
  assign n19382 = n19380 | n19381 ;
  assign n19384 = ( x125 & ~n19383 ) | ( x125 & n19382 ) | ( ~n19383 & n19382 ) ;
  assign n19385 = n7541 | n9941 ;
  assign n19386 = ~n19384 & n19385 ;
  assign n19387 = x56 &  n19386 ;
  assign n19388 = x56 | n19386 ;
  assign n19389 = ~n19387 & n19388 ;
  assign n19390 = ( n19300 & n19351 ) | ( n19300 & n19361 ) | ( n19351 & n19361 ) ;
  assign n19394 = x122 &  n8558 ;
  assign n19391 = ( x124 & ~n8314 ) | ( x124 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n19392 = x123 &  n8309 ;
  assign n19393 = n19391 | n19392 ;
  assign n19395 = ( x122 & ~n19394 ) | ( x122 & n19393 ) | ( ~n19394 & n19393 ) ;
  assign n19396 = ~n8317 & n8755 ;
  assign n19397 = n19395 | n19396 ;
  assign n19399 = x59 &  n19397 ;
  assign n19398 = ~x59 & n19397 ;
  assign n19400 = ( x59 & ~n19399 ) | ( x59 & n19398 ) | ( ~n19399 & n19398 ) ;
  assign n19401 = ( n19332 & ~n19338 ) | ( n19332 & n19348 ) | ( ~n19338 & n19348 ) ;
  assign n19402 = x117 &  n10104 ;
  assign n19403 = ( x118 & ~n9760 ) | ( x118 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n19404 = n19402 | n19403 ;
  assign n19405 = ( x53 & n19335 ) | ( x53 & n19404 ) | ( n19335 & n19404 ) ;
  assign n19406 = ( x53 & ~n19335 ) | ( x53 & n19404 ) | ( ~n19335 & n19404 ) ;
  assign n19407 = ( n19335 & ~n19405 ) | ( n19335 & n19406 ) | ( ~n19405 & n19406 ) ;
  assign n19408 = ( n19285 & ~n19335 ) | ( n19285 & n19296 ) | ( ~n19335 & n19296 ) ;
  assign n19412 = x119 &  n9457 ;
  assign n19409 = ( x121 & ~n9150 ) | ( x121 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n19410 = x120 &  n9145 ;
  assign n19411 = n19409 | n19410 ;
  assign n19413 = ( x119 & ~n19412 ) | ( x119 & n19411 ) | ( ~n19412 & n19411 ) ;
  assign n19414 = ( n8176 & ~n9153 ) | ( n8176 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n19415 = n19413 | n19414 ;
  assign n19416 = ( x62 & ~n19415 ) | ( x62 & 1'b0 ) | ( ~n19415 & 1'b0 ) ;
  assign n19417 = ~x62 & n19415 ;
  assign n19418 = n19416 | n19417 ;
  assign n19419 = ( n19407 & ~n19408 ) | ( n19407 & n19418 ) | ( ~n19408 & n19418 ) ;
  assign n19420 = ( n19407 & ~n19418 ) | ( n19407 & n19408 ) | ( ~n19418 & n19408 ) ;
  assign n19421 = ( n19419 & ~n19407 ) | ( n19419 & n19420 ) | ( ~n19407 & n19420 ) ;
  assign n19422 = ( n19400 & ~n19401 ) | ( n19400 & n19421 ) | ( ~n19401 & n19421 ) ;
  assign n19423 = ( n19400 & ~n19421 ) | ( n19400 & n19401 ) | ( ~n19421 & n19401 ) ;
  assign n19424 = ( n19422 & ~n19400 ) | ( n19422 & n19423 ) | ( ~n19400 & n19423 ) ;
  assign n19425 = ( n19389 & ~n19390 ) | ( n19389 & n19424 ) | ( ~n19390 & n19424 ) ;
  assign n19426 = ( n19389 & ~n19424 ) | ( n19389 & n19390 ) | ( ~n19424 & n19390 ) ;
  assign n19427 = ( n19425 & ~n19389 ) | ( n19425 & n19426 ) | ( ~n19389 & n19426 ) ;
  assign n19428 = ( n19378 & n19379 ) | ( n19378 & n19427 ) | ( n19379 & n19427 ) ;
  assign n19429 = ( n19379 & ~n19378 ) | ( n19379 & n19427 ) | ( ~n19378 & n19427 ) ;
  assign n19430 = ( n19378 & ~n19428 ) | ( n19378 & n19429 ) | ( ~n19428 & n19429 ) ;
  assign n19431 = ( n19389 & n19390 ) | ( n19389 & n19424 ) | ( n19390 & n19424 ) ;
  assign n19432 = ( x126 & ~n7731 ) | ( x126 & 1'b0 ) | ( ~n7731 & 1'b0 ) ;
  assign n19433 = x127 &  n7533 ;
  assign n19434 = n19432 | n19433 ;
  assign n19435 = n7541 | n9960 ;
  assign n19436 = ( n19434 & ~n7541 ) | ( n19434 & n19435 ) | ( ~n7541 & n19435 ) ;
  assign n19438 = x56 &  n19436 ;
  assign n19437 = ~x56 & n19436 ;
  assign n19439 = ( x56 & ~n19438 ) | ( x56 & n19437 ) | ( ~n19438 & n19437 ) ;
  assign n19440 = ( n19408 & ~n19407 ) | ( n19408 & n19418 ) | ( ~n19407 & n19418 ) ;
  assign n19444 = x123 &  n8558 ;
  assign n19441 = ( x125 & ~n8314 ) | ( x125 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n19442 = x124 &  n8309 ;
  assign n19443 = n19441 | n19442 ;
  assign n19445 = ( x123 & ~n19444 ) | ( x123 & n19443 ) | ( ~n19444 & n19443 ) ;
  assign n19446 = ~n8317 & n9324 ;
  assign n19447 = n19445 | n19446 ;
  assign n19448 = ( x59 & ~n19447 ) | ( x59 & 1'b0 ) | ( ~n19447 & 1'b0 ) ;
  assign n19449 = ~x59 & n19447 ;
  assign n19450 = n19448 | n19449 ;
  assign n19451 = ( n19335 & ~x53 ) | ( n19335 & n19404 ) | ( ~x53 & n19404 ) ;
  assign n19452 = x118 &  n10104 ;
  assign n19453 = ( x119 & ~n9760 ) | ( x119 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n19454 = n19452 | n19453 ;
  assign n19458 = x120 &  n9457 ;
  assign n19455 = ( x122 & ~n9150 ) | ( x122 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n19456 = x121 &  n9145 ;
  assign n19457 = n19455 | n19456 ;
  assign n19459 = ( x120 & ~n19458 ) | ( x120 & n19457 ) | ( ~n19458 & n19457 ) ;
  assign n19460 = ( n9153 & ~n19459 ) | ( n9153 & n9987 ) | ( ~n19459 & n9987 ) ;
  assign n19461 = ~n9153 & n19460 ;
  assign n19462 = ( x62 & n19459 ) | ( x62 & n19461 ) | ( n19459 & n19461 ) ;
  assign n19463 = ( x62 & ~n19461 ) | ( x62 & n19459 ) | ( ~n19461 & n19459 ) ;
  assign n19464 = ( n19461 & ~n19462 ) | ( n19461 & n19463 ) | ( ~n19462 & n19463 ) ;
  assign n19465 = ( n19451 & ~n19454 ) | ( n19451 & n19464 ) | ( ~n19454 & n19464 ) ;
  assign n19466 = ( n19451 & ~n19464 ) | ( n19451 & n19454 ) | ( ~n19464 & n19454 ) ;
  assign n19467 = ( n19465 & ~n19451 ) | ( n19465 & n19466 ) | ( ~n19451 & n19466 ) ;
  assign n19468 = ( n19440 & ~n19450 ) | ( n19440 & n19467 ) | ( ~n19450 & n19467 ) ;
  assign n19469 = ( n19440 & ~n19467 ) | ( n19440 & n19450 ) | ( ~n19467 & n19450 ) ;
  assign n19470 = ( n19468 & ~n19440 ) | ( n19468 & n19469 ) | ( ~n19440 & n19469 ) ;
  assign n19471 = ( n19423 & ~n19439 ) | ( n19423 & n19470 ) | ( ~n19439 & n19470 ) ;
  assign n19472 = ( n19423 & ~n19470 ) | ( n19423 & n19439 ) | ( ~n19470 & n19439 ) ;
  assign n19473 = ( n19471 & ~n19423 ) | ( n19471 & n19472 ) | ( ~n19423 & n19472 ) ;
  assign n19474 = ( n19378 & ~n19379 ) | ( n19378 & n19427 ) | ( ~n19379 & n19427 ) ;
  assign n19475 = ( n19431 & ~n19473 ) | ( n19431 & n19474 ) | ( ~n19473 & n19474 ) ;
  assign n19476 = ( n19431 & ~n19474 ) | ( n19431 & n19473 ) | ( ~n19474 & n19473 ) ;
  assign n19477 = ( n19475 & ~n19431 ) | ( n19475 & n19476 ) | ( ~n19431 & n19476 ) ;
  assign n19516 = ( n19431 & n19473 ) | ( n19431 & n19474 ) | ( n19473 & n19474 ) ;
  assign n19497 = x124 &  n8558 ;
  assign n19494 = ( x126 & ~n8314 ) | ( x126 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n19495 = x125 &  n8309 ;
  assign n19496 = n19494 | n19495 ;
  assign n19498 = ( x124 & ~n19497 ) | ( x124 & n19496 ) | ( ~n19497 & n19496 ) ;
  assign n19499 = n8317 | n9349 ;
  assign n19500 = ~n19498 & n19499 ;
  assign n19501 = x59 &  n19500 ;
  assign n19502 = x59 | n19500 ;
  assign n19503 = ~n19501 & n19502 ;
  assign n19481 = x121 &  n9457 ;
  assign n19478 = ( x123 & ~n9150 ) | ( x123 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n19479 = x122 &  n9145 ;
  assign n19480 = n19478 | n19479 ;
  assign n19482 = ( x121 & ~n19481 ) | ( x121 & n19480 ) | ( ~n19481 & n19480 ) ;
  assign n19483 = ( n8472 & ~n9153 ) | ( n8472 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n19484 = n19482 | n19483 ;
  assign n19485 = ( x62 & ~n19484 ) | ( x62 & 1'b0 ) | ( ~n19484 & 1'b0 ) ;
  assign n19486 = ~x62 & n19484 ;
  assign n19487 = n19485 | n19486 ;
  assign n19488 = x119 &  n10104 ;
  assign n19489 = ( x120 & ~n9760 ) | ( x120 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n19490 = n19488 | n19489 ;
  assign n19491 = ( n19487 & ~n19454 ) | ( n19487 & n19490 ) | ( ~n19454 & n19490 ) ;
  assign n19492 = ( n19454 & ~n19490 ) | ( n19454 & n19487 ) | ( ~n19490 & n19487 ) ;
  assign n19493 = ( n19491 & ~n19487 ) | ( n19491 & n19492 ) | ( ~n19487 & n19492 ) ;
  assign n19504 = ( n19465 & ~n19503 ) | ( n19465 & n19493 ) | ( ~n19503 & n19493 ) ;
  assign n19505 = ( n19465 & ~n19493 ) | ( n19465 & n19503 ) | ( ~n19493 & n19503 ) ;
  assign n19506 = ( n19504 & ~n19465 ) | ( n19504 & n19505 ) | ( ~n19465 & n19505 ) ;
  assign n19507 = ( x127 & ~n7731 ) | ( x127 & 1'b0 ) | ( ~n7731 & 1'b0 ) ;
  assign n19508 = ( n7541 & ~n10258 ) | ( n7541 & n19507 ) | ( ~n10258 & n19507 ) ;
  assign n19509 = n10258 | n19508 ;
  assign n19510 = ( x56 & ~n19507 ) | ( x56 & n19509 ) | ( ~n19507 & n19509 ) ;
  assign n19511 = ( n19507 & ~x56 ) | ( n19507 & n19509 ) | ( ~x56 & n19509 ) ;
  assign n19512 = ( n19510 & ~n19509 ) | ( n19510 & n19511 ) | ( ~n19509 & n19511 ) ;
  assign n19514 = ( n19469 & n19506 ) | ( n19469 & n19512 ) | ( n19506 & n19512 ) ;
  assign n19513 = ( n19506 & ~n19469 ) | ( n19506 & n19512 ) | ( ~n19469 & n19512 ) ;
  assign n19515 = ( n19469 & ~n19514 ) | ( n19469 & n19513 ) | ( ~n19514 & n19513 ) ;
  assign n19517 = ( n19472 & ~n19516 ) | ( n19472 & n19515 ) | ( ~n19516 & n19515 ) ;
  assign n19518 = ( n19472 & ~n19515 ) | ( n19472 & n19516 ) | ( ~n19515 & n19516 ) ;
  assign n19519 = ( n19517 & ~n19472 ) | ( n19517 & n19518 ) | ( ~n19472 & n19518 ) ;
  assign n19520 = ( n19469 & ~n19512 ) | ( n19469 & n19506 ) | ( ~n19512 & n19506 ) ;
  assign n19554 = ( n19515 & ~n19472 ) | ( n19515 & n19516 ) | ( ~n19472 & n19516 ) ;
  assign n19521 = x120 &  n10104 ;
  assign n19522 = ( x121 & ~n9760 ) | ( x121 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n19523 = n19521 | n19522 ;
  assign n19524 = ( x56 & n19454 ) | ( x56 & n19523 ) | ( n19454 & n19523 ) ;
  assign n19525 = ( x56 & ~n19454 ) | ( x56 & n19523 ) | ( ~n19454 & n19523 ) ;
  assign n19526 = ( n19454 & ~n19524 ) | ( n19454 & n19525 ) | ( ~n19524 & n19525 ) ;
  assign n19527 = n19491 &  n19526 ;
  assign n19528 = n19491 | n19526 ;
  assign n19529 = ~n19527 & n19528 ;
  assign n19534 = x125 &  n8558 ;
  assign n19531 = ( x127 & ~n8314 ) | ( x127 & 1'b0 ) | ( ~n8314 & 1'b0 ) ;
  assign n19532 = x126 &  n8309 ;
  assign n19533 = n19531 | n19532 ;
  assign n19535 = ( x125 & ~n19534 ) | ( x125 & n19533 ) | ( ~n19534 & n19533 ) ;
  assign n19536 = n8317 | n9941 ;
  assign n19537 = ~n19535 & n19536 ;
  assign n19530 = ( n19493 & ~n19465 ) | ( n19493 & n19503 ) | ( ~n19465 & n19503 ) ;
  assign n19538 = ( x59 & ~n19537 ) | ( x59 & n19530 ) | ( ~n19537 & n19530 ) ;
  assign n19539 = ( x59 & ~n19530 ) | ( x59 & n19537 ) | ( ~n19530 & n19537 ) ;
  assign n19540 = ( n19538 & ~x59 ) | ( n19538 & n19539 ) | ( ~x59 & n19539 ) ;
  assign n19544 = x122 &  n9457 ;
  assign n19541 = ( x124 & ~n9150 ) | ( x124 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n19542 = x123 &  n9145 ;
  assign n19543 = n19541 | n19542 ;
  assign n19545 = ( x122 & ~n19544 ) | ( x122 & n19543 ) | ( ~n19544 & n19543 ) ;
  assign n19546 = ( n8755 & ~n9153 ) | ( n8755 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n19547 = n19545 | n19546 ;
  assign n19548 = ( x62 & ~n19547 ) | ( x62 & 1'b0 ) | ( ~n19547 & 1'b0 ) ;
  assign n19549 = ~x62 & n19547 ;
  assign n19550 = n19548 | n19549 ;
  assign n19551 = ( n19529 & ~n19540 ) | ( n19529 & n19550 ) | ( ~n19540 & n19550 ) ;
  assign n19552 = ( n19529 & ~n19550 ) | ( n19529 & n19540 ) | ( ~n19550 & n19540 ) ;
  assign n19553 = ( n19551 & ~n19529 ) | ( n19551 & n19552 ) | ( ~n19529 & n19552 ) ;
  assign n19555 = ( n19520 & ~n19554 ) | ( n19520 & n19553 ) | ( ~n19554 & n19553 ) ;
  assign n19556 = ( n19520 & ~n19553 ) | ( n19520 & n19554 ) | ( ~n19553 & n19554 ) ;
  assign n19557 = ( n19555 & ~n19520 ) | ( n19555 & n19556 ) | ( ~n19520 & n19556 ) ;
  assign n19558 = ( n19530 & ~x59 ) | ( n19530 & n19537 ) | ( ~x59 & n19537 ) ;
  assign n19559 = n19538 | n19558 ;
  assign n19561 = ( n19540 & ~n19529 ) | ( n19540 & n19550 ) | ( ~n19529 & n19550 ) ;
  assign n19560 = ~n19529 & n19550 ;
  assign n19562 = ( n19559 & ~n19561 ) | ( n19559 & n19560 ) | ( ~n19561 & n19560 ) ;
  assign n19563 = ( n19491 & ~n19526 ) | ( n19491 & n19550 ) | ( ~n19526 & n19550 ) ;
  assign n19586 = ~x59 & n19563 ;
  assign n19587 = x59 | n19563 ;
  assign n19588 = ( n19586 & ~n19563 ) | ( n19586 & n19587 ) | ( ~n19563 & n19587 ) ;
  assign n19564 = ( n19454 & ~x56 ) | ( n19454 & n19523 ) | ( ~x56 & n19523 ) ;
  assign n19565 = x121 &  n10104 ;
  assign n19566 = ( x122 & ~n9760 ) | ( x122 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n19567 = n19565 | n19566 ;
  assign n19571 = x123 &  n9457 ;
  assign n19568 = ( x125 & ~n9150 ) | ( x125 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n19569 = x124 &  n9145 ;
  assign n19570 = n19568 | n19569 ;
  assign n19572 = ( x123 & ~n19571 ) | ( x123 & n19570 ) | ( ~n19571 & n19570 ) ;
  assign n19573 = ( n9153 & n9324 ) | ( n9153 & n19572 ) | ( n9324 & n19572 ) ;
  assign n19574 = ( n9324 & ~n19573 ) | ( n9324 & 1'b0 ) | ( ~n19573 & 1'b0 ) ;
  assign n19575 = ( x62 & n19572 ) | ( x62 & n19574 ) | ( n19572 & n19574 ) ;
  assign n19576 = ( x62 & ~n19574 ) | ( x62 & n19572 ) | ( ~n19574 & n19572 ) ;
  assign n19577 = ( n19574 & ~n19575 ) | ( n19574 & n19576 ) | ( ~n19575 & n19576 ) ;
  assign n19578 = ( n19564 & ~n19567 ) | ( n19564 & n19577 ) | ( ~n19567 & n19577 ) ;
  assign n19579 = ( n19564 & ~n19577 ) | ( n19564 & n19567 ) | ( ~n19577 & n19567 ) ;
  assign n19580 = ( n19578 & ~n19564 ) | ( n19578 & n19579 ) | ( ~n19564 & n19579 ) ;
  assign n19581 = ( x126 & ~n8558 ) | ( x126 & 1'b0 ) | ( ~n8558 & 1'b0 ) ;
  assign n19582 = x127 &  n8309 ;
  assign n19583 = n19581 | n19582 ;
  assign n19584 = n8317 | n9960 ;
  assign n19585 = ( n19583 & ~n8317 ) | ( n19583 & n19584 ) | ( ~n8317 & n19584 ) ;
  assign n19589 = ( n19580 & n19585 ) | ( n19580 & n19588 ) | ( n19585 & n19588 ) ;
  assign n19590 = ( n19580 & ~n19588 ) | ( n19580 & n19585 ) | ( ~n19588 & n19585 ) ;
  assign n19591 = ( n19588 & ~n19589 ) | ( n19588 & n19590 ) | ( ~n19589 & n19590 ) ;
  assign n19592 = ( n19553 & ~n19520 ) | ( n19553 & n19554 ) | ( ~n19520 & n19554 ) ;
  assign n19593 = ( n19562 & ~n19591 ) | ( n19562 & n19592 ) | ( ~n19591 & n19592 ) ;
  assign n19594 = ( n19562 & ~n19592 ) | ( n19562 & n19591 ) | ( ~n19592 & n19591 ) ;
  assign n19595 = ( n19593 & ~n19562 ) | ( n19593 & n19594 ) | ( ~n19562 & n19594 ) ;
  assign n19596 = x59 | n19585 ;
  assign n19597 = x59 &  n19585 ;
  assign n19598 = ( n19596 & ~n19597 ) | ( n19596 & 1'b0 ) | ( ~n19597 & 1'b0 ) ;
  assign n19599 = ( n19563 & ~n19580 ) | ( n19563 & n19598 ) | ( ~n19580 & n19598 ) ;
  assign n19604 = x124 &  n9457 ;
  assign n19601 = ( x126 & ~n9150 ) | ( x126 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n19602 = x125 &  n9145 ;
  assign n19603 = n19601 | n19602 ;
  assign n19605 = ( x124 & ~n19604 ) | ( x124 & n19603 ) | ( ~n19604 & n19603 ) ;
  assign n19606 = n9153 | n9349 ;
  assign n19607 = ~n19605 & n19606 ;
  assign n19608 = x62 &  n19607 ;
  assign n19609 = x62 | n19607 ;
  assign n19610 = ~n19608 & n19609 ;
  assign n19611 = x122 &  n10104 ;
  assign n19612 = ( x123 & ~n9760 ) | ( x123 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n19613 = n19611 | n19612 ;
  assign n19614 = ( n19567 & n19578 ) | ( n19567 & n19613 ) | ( n19578 & n19613 ) ;
  assign n19615 = ( n19567 & ~n19578 ) | ( n19567 & n19613 ) | ( ~n19578 & n19613 ) ;
  assign n19616 = ( n19578 & ~n19614 ) | ( n19578 & n19615 ) | ( ~n19614 & n19615 ) ;
  assign n19617 = ( x127 & ~n8558 ) | ( x127 & 1'b0 ) | ( ~n8558 & 1'b0 ) ;
  assign n19618 = n8317 | n10258 ;
  assign n19619 = ~n19617 & n19618 ;
  assign n19620 = ~x59 & n19619 ;
  assign n19621 = ( x59 & ~n19619 ) | ( x59 & 1'b0 ) | ( ~n19619 & 1'b0 ) ;
  assign n19622 = n19620 | n19621 ;
  assign n19623 = ( n19610 & ~n19616 ) | ( n19610 & n19622 ) | ( ~n19616 & n19622 ) ;
  assign n19624 = ( n19610 & ~n19622 ) | ( n19610 & n19616 ) | ( ~n19622 & n19616 ) ;
  assign n19625 = ( n19623 & ~n19610 ) | ( n19623 & n19624 ) | ( ~n19610 & n19624 ) ;
  assign n19600 = ( n19562 & n19591 ) | ( n19562 & n19592 ) | ( n19591 & n19592 ) ;
  assign n19626 = ( n19599 & ~n19625 ) | ( n19599 & n19600 ) | ( ~n19625 & n19600 ) ;
  assign n19627 = ( n19599 & ~n19600 ) | ( n19599 & n19625 ) | ( ~n19600 & n19625 ) ;
  assign n19628 = ( n19626 & ~n19599 ) | ( n19626 & n19627 ) | ( ~n19599 & n19627 ) ;
  assign n19629 = ( n19610 & n19616 ) | ( n19610 & n19622 ) | ( n19616 & n19622 ) ;
  assign n19630 = ( n19600 & ~n19599 ) | ( n19600 & n19625 ) | ( ~n19599 & n19625 ) ;
  assign n19631 = ( n19567 & ~n19613 ) | ( n19567 & n19578 ) | ( ~n19613 & n19578 ) ;
  assign n19641 = x125 &  n9457 ;
  assign n19638 = ( x127 & ~n9150 ) | ( x127 & 1'b0 ) | ( ~n9150 & 1'b0 ) ;
  assign n19639 = x126 &  n9145 ;
  assign n19640 = n19638 | n19639 ;
  assign n19642 = ( x125 & ~n19641 ) | ( x125 & n19640 ) | ( ~n19641 & n19640 ) ;
  assign n19643 = n9153 | n9941 ;
  assign n19644 = ~n19642 & n19643 ;
  assign n19632 = x123 &  n10104 ;
  assign n19633 = ( x124 & ~n9760 ) | ( x124 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n19634 = n19632 | n19633 ;
  assign n19635 = ( x59 & n19613 ) | ( x59 & n19634 ) | ( n19613 & n19634 ) ;
  assign n19636 = ( x59 & ~n19613 ) | ( x59 & n19634 ) | ( ~n19613 & n19634 ) ;
  assign n19637 = ( n19613 & ~n19635 ) | ( n19613 & n19636 ) | ( ~n19635 & n19636 ) ;
  assign n19645 = ( x62 & ~n19644 ) | ( x62 & n19637 ) | ( ~n19644 & n19637 ) ;
  assign n19646 = ( n19637 & ~x62 ) | ( n19637 & n19644 ) | ( ~x62 & n19644 ) ;
  assign n19647 = ( n19645 & ~n19637 ) | ( n19645 & n19646 ) | ( ~n19637 & n19646 ) ;
  assign n19648 = n19631 &  n19647 ;
  assign n19649 = n19631 | n19647 ;
  assign n19650 = ~n19648 & n19649 ;
  assign n19651 = ( n19629 & ~n19630 ) | ( n19629 & n19650 ) | ( ~n19630 & n19650 ) ;
  assign n19652 = ( n19629 & ~n19650 ) | ( n19629 & n19630 ) | ( ~n19650 & n19630 ) ;
  assign n19653 = ( n19651 & ~n19629 ) | ( n19651 & n19652 ) | ( ~n19629 & n19652 ) ;
  assign n19654 = ~x62 & n19644 ;
  assign n19655 = ( n19645 & ~n19648 ) | ( n19645 & n19654 ) | ( ~n19648 & n19654 ) ;
  assign n19656 = ( n19613 & ~x59 ) | ( n19613 & n19634 ) | ( ~x59 & n19634 ) ;
  assign n19657 = x124 &  n10104 ;
  assign n19658 = ( x125 & ~n9760 ) | ( x125 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n19659 = n19657 | n19658 ;
  assign n19660 = ( x126 & ~n9457 ) | ( x126 & 1'b0 ) | ( ~n9457 & 1'b0 ) ;
  assign n19661 = x127 &  n9145 ;
  assign n19662 = n19660 | n19661 ;
  assign n19663 = n9153 | n9960 ;
  assign n19664 = ( n19662 & ~n9153 ) | ( n19662 & n19663 ) | ( ~n9153 & n19663 ) ;
  assign n19665 = x62 | n19664 ;
  assign n19666 = ( x62 & ~n19664 ) | ( x62 & 1'b0 ) | ( ~n19664 & 1'b0 ) ;
  assign n19667 = ( n19665 & ~x62 ) | ( n19665 & n19666 ) | ( ~x62 & n19666 ) ;
  assign n19668 = ( n19656 & ~n19659 ) | ( n19656 & n19667 ) | ( ~n19659 & n19667 ) ;
  assign n19669 = ( n19656 & ~n19667 ) | ( n19656 & n19659 ) | ( ~n19667 & n19659 ) ;
  assign n19670 = ( n19668 & ~n19656 ) | ( n19668 & n19669 ) | ( ~n19656 & n19669 ) ;
  assign n19672 = ( n19652 & n19655 ) | ( n19652 & n19670 ) | ( n19655 & n19670 ) ;
  assign n19671 = ( n19652 & ~n19655 ) | ( n19652 & n19670 ) | ( ~n19655 & n19670 ) ;
  assign n19673 = ( n19655 & ~n19672 ) | ( n19655 & n19671 ) | ( ~n19672 & n19671 ) ;
  assign n19674 = x125 &  n10104 ;
  assign n19675 = ( x126 & ~n9760 ) | ( x126 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n19676 = n19674 | n19675 ;
  assign n19677 = ( x127 & ~n9457 ) | ( x127 & 1'b0 ) | ( ~n9457 & 1'b0 ) ;
  assign n19678 = ( n9153 & ~n10258 ) | ( n9153 & n19677 ) | ( ~n10258 & n19677 ) ;
  assign n19679 = n10258 | n19678 ;
  assign n19680 = ( x62 & ~n19677 ) | ( x62 & n19679 ) | ( ~n19677 & n19679 ) ;
  assign n19681 = ( n19677 & ~x62 ) | ( n19677 & n19679 ) | ( ~x62 & n19679 ) ;
  assign n19682 = ( n19680 & ~n19679 ) | ( n19680 & n19681 ) | ( ~n19679 & n19681 ) ;
  assign n19684 = ( n19659 & n19676 ) | ( n19659 & n19682 ) | ( n19676 & n19682 ) ;
  assign n19683 = ( n19659 & ~n19676 ) | ( n19659 & n19682 ) | ( ~n19676 & n19682 ) ;
  assign n19685 = ( n19676 & ~n19684 ) | ( n19676 & n19683 ) | ( ~n19684 & n19683 ) ;
  assign n19686 = ( n19668 & ~n19685 ) | ( n19668 & n19672 ) | ( ~n19685 & n19672 ) ;
  assign n19687 = ( n19668 & ~n19672 ) | ( n19668 & n19685 ) | ( ~n19672 & n19685 ) ;
  assign n19688 = ( n19686 & ~n19668 ) | ( n19686 & n19687 ) | ( ~n19668 & n19687 ) ;
  assign n19689 = x126 &  n10104 ;
  assign n19690 = ( x127 & ~n9760 ) | ( x127 & 1'b0 ) | ( ~n9760 & 1'b0 ) ;
  assign n19691 = n19689 | n19690 ;
  assign n19692 = ( x62 & n19659 ) | ( x62 & n19691 ) | ( n19659 & n19691 ) ;
  assign n19693 = ( x62 & ~n19659 ) | ( x62 & n19691 ) | ( ~n19659 & n19691 ) ;
  assign n19694 = ( n19659 & ~n19692 ) | ( n19659 & n19693 ) | ( ~n19692 & n19693 ) ;
  assign n19695 = ( n19683 & ~n19694 ) | ( n19683 & n19687 ) | ( ~n19694 & n19687 ) ;
  assign n19696 = ( n19683 & ~n19687 ) | ( n19683 & n19694 ) | ( ~n19687 & n19694 ) ;
  assign n19697 = ( n19695 & ~n19683 ) | ( n19695 & n19696 ) | ( ~n19683 & n19696 ) ;
  assign n19698 = ( n19659 & ~x62 ) | ( n19659 & n19691 ) | ( ~x62 & n19691 ) ;
  assign n19699 = x127 &  n10104 ;
  assign n19701 = ( n19696 & n19698 ) | ( n19696 & n19699 ) | ( n19698 & n19699 ) ;
  assign n19700 = ( n19696 & ~n19698 ) | ( n19696 & n19699 ) | ( ~n19698 & n19699 ) ;
  assign n19702 = ( n19698 & ~n19701 ) | ( n19698 & n19700 ) | ( ~n19701 & n19700 ) ;
  assign y0 = n129 ;
  assign y1 = n147 ;
  assign y2 = n163 ;
  assign y3 = ~n188 ;
  assign y4 = n222 ;
  assign y5 = n254 ;
  assign y6 = ~n290 ;
  assign y7 = n337 ;
  assign y8 = n381 ;
  assign y9 = ~n431 ;
  assign y10 = n490 ;
  assign y11 = n548 ;
  assign y12 = ~n611 ;
  assign y13 = n685 ;
  assign y14 = n758 ;
  assign y15 = ~n834 ;
  assign y16 = n919 ;
  assign y17 = n1002 ;
  assign y18 = ~n1092 ;
  assign y19 = n1191 ;
  assign y20 = n1287 ;
  assign y21 = ~n1391 ;
  assign y22 = n1504 ;
  assign y23 = n1616 ;
  assign y24 = ~n1733 ;
  assign y25 = n1861 ;
  assign y26 = n1984 ;
  assign y27 = ~n2116 ;
  assign y28 = n2256 ;
  assign y29 = ~n2393 ;
  assign y30 = ~n2539 ;
  assign y31 = n2694 ;
  assign y32 = ~n2844 ;
  assign y33 = ~n3007 ;
  assign y34 = n3178 ;
  assign y35 = ~n3346 ;
  assign y36 = n3521 ;
  assign y37 = n3702 ;
  assign y38 = ~n3880 ;
  assign y39 = n4064 ;
  assign y40 = n4257 ;
  assign y41 = n4450 ;
  assign y42 = ~n4646 ;
  assign y43 = n4856 ;
  assign y44 = ~n5063 ;
  assign y45 = ~n5275 ;
  assign y46 = ~n5500 ;
  assign y47 = n5719 ;
  assign y48 = n5943 ;
  assign y49 = ~n6177 ;
  assign y50 = n6412 ;
  assign y51 = ~n6648 ;
  assign y52 = n6893 ;
  assign y53 = n7144 ;
  assign y54 = ~n7397 ;
  assign y55 = ~n7656 ;
  assign y56 = n7916 ;
  assign y57 = ~n8184 ;
  assign y58 = ~n8460 ;
  assign y59 = n8735 ;
  assign y60 = ~n9034 ;
  assign y61 = ~n9332 ;
  assign y62 = ~n9643 ;
  assign y63 = n9949 ;
  assign y64 = n10249 ;
  assign y65 = ~n10544 ;
  assign y66 = n10840 ;
  assign y67 = n11126 ;
  assign y68 = ~n11409 ;
  assign y69 = n11682 ;
  assign y70 = n11947 ;
  assign y71 = ~n12221 ;
  assign y72 = n12481 ;
  assign y73 = n12737 ;
  assign y74 = ~n12989 ;
  assign y75 = n13236 ;
  assign y76 = n13484 ;
  assign y77 = ~n13718 ;
  assign y78 = n13950 ;
  assign y79 = n14184 ;
  assign y80 = ~n14417 ;
  assign y81 = n14638 ;
  assign y82 = n14848 ;
  assign y83 = ~n15062 ;
  assign y84 = n15263 ;
  assign y85 = n15462 ;
  assign y86 = ~n15665 ;
  assign y87 = n15856 ;
  assign y88 = n16043 ;
  assign y89 = ~n16225 ;
  assign y90 = n16400 ;
  assign y91 = n16573 ;
  assign y92 = n16746 ;
  assign y93 = n16907 ;
  assign y94 = n17068 ;
  assign y95 = n17219 ;
  assign y96 = n17367 ;
  assign y97 = n17516 ;
  assign y98 = n17658 ;
  assign y99 = ~n17793 ;
  assign y100 = n17922 ;
  assign y101 = n18056 ;
  assign y102 = ~n18176 ;
  assign y103 = n18293 ;
  assign y104 = ~n18410 ;
  assign y105 = n18515 ;
  assign y106 = n18614 ;
  assign y107 = n18713 ;
  assign y108 = n18803 ;
  assign y109 = ~n18890 ;
  assign y110 = n18973 ;
  assign y111 = ~n19052 ;
  assign y112 = ~n19124 ;
  assign y113 = n19196 ;
  assign y114 = n19261 ;
  assign y115 = n19318 ;
  assign y116 = ~n19377 ;
  assign y117 = n19430 ;
  assign y118 = ~n19477 ;
  assign y119 = n19519 ;
  assign y120 = n19557 ;
  assign y121 = ~n19595 ;
  assign y122 = n19628 ;
  assign y123 = n19653 ;
  assign y124 = ~n19673 ;
  assign y125 = ~n19688 ;
  assign y126 = n19697 ;
  assign y127 = n19702 ;
endmodule
