module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 ;
  wire n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 ;
  assign n514 = ( x376 & ~x504 ) | ( x376 & 1'b0 ) | ( ~x504 & 1'b0 ) ;
  assign n515 = ( x377 & ~x505 ) | ( x377 & n514 ) | ( ~x505 & n514 ) ;
  assign n516 = ( x378 & ~x506 ) | ( x378 & n515 ) | ( ~x506 & n515 ) ;
  assign n517 = ( x379 & ~x507 ) | ( x379 & n516 ) | ( ~x507 & n516 ) ;
  assign n873 = ~x380 & x508 ;
  assign n877 = x383 &  x511 ;
  assign n874 = ~x382 & x510 ;
  assign n875 = ~x381 & x509 ;
  assign n876 = n874 | n875 ;
  assign n878 = ( x383 & ~n877 ) | ( x383 & n876 ) | ( ~n877 & n876 ) ;
  assign n879 = n873 | n878 ;
  assign n518 = ( x375 & ~x503 ) | ( x375 & 1'b0 ) | ( ~x503 & 1'b0 ) ;
  assign n513 = ~x379 & x507 ;
  assign n864 = ~x377 & x505 ;
  assign n865 = ~x378 & x506 ;
  assign n866 = ~x376 & x504 ;
  assign n867 = ( n865 & ~n864 ) | ( n865 & n866 ) | ( ~n864 & n866 ) ;
  assign n868 = ( n864 & ~n513 ) | ( n864 & n867 ) | ( ~n513 & n867 ) ;
  assign n869 = n513 | n868 ;
  assign n870 = n517 | n869 ;
  assign n526 = ~x367 & x495 ;
  assign n835 = ( x364 & ~x492 ) | ( x364 & 1'b0 ) | ( ~x492 & 1'b0 ) ;
  assign n836 = ( x365 & ~x493 ) | ( x365 & n835 ) | ( ~x493 & n835 ) ;
  assign n837 = ( x366 & ~x494 ) | ( x366 & n836 ) | ( ~x494 & n836 ) ;
  assign n838 = ~n526 & n837 ;
  assign n527 = ~x366 & x494 ;
  assign n528 = n526 | n527 ;
  assign n529 = ~x365 & x493 ;
  assign n530 = ~x364 & x492 ;
  assign n531 = ( n529 & ~n528 ) | ( n529 & n530 ) | ( ~n528 & n530 ) ;
  assign n532 = n528 | n531 ;
  assign n533 = ( x359 & ~x487 ) | ( x359 & 1'b0 ) | ( ~x487 & 1'b0 ) ;
  assign n821 = ~x363 & x491 ;
  assign n822 = ~x361 & x489 ;
  assign n823 = ~x362 & x490 ;
  assign n824 = ~x360 & x488 ;
  assign n825 = ( n823 & ~n822 ) | ( n823 & n824 ) | ( ~n822 & n824 ) ;
  assign n826 = ( n822 & ~n821 ) | ( n822 & n825 ) | ( ~n821 & n825 ) ;
  assign n827 = n821 | n826 ;
  assign n541 = ~x351 & x479 ;
  assign n792 = ( x348 & ~x476 ) | ( x348 & 1'b0 ) | ( ~x476 & 1'b0 ) ;
  assign n793 = ( x349 & ~x477 ) | ( x349 & n792 ) | ( ~x477 & n792 ) ;
  assign n794 = ( x350 & ~x478 ) | ( x350 & n793 ) | ( ~x478 & n793 ) ;
  assign n795 = ~n541 & n794 ;
  assign n542 = ~x350 & x478 ;
  assign n543 = n541 | n542 ;
  assign n544 = ~x349 & x477 ;
  assign n545 = ~x348 & x476 ;
  assign n546 = ( n544 & ~n543 ) | ( n544 & n545 ) | ( ~n543 & n545 ) ;
  assign n547 = n543 | n546 ;
  assign n548 = ( x343 & ~x471 ) | ( x343 & 1'b0 ) | ( ~x471 & 1'b0 ) ;
  assign n778 = ~x347 & x475 ;
  assign n779 = ~x345 & x473 ;
  assign n780 = ~x346 & x474 ;
  assign n781 = ~x344 & x472 ;
  assign n782 = ( n780 & ~n779 ) | ( n780 & n781 ) | ( ~n779 & n781 ) ;
  assign n783 = ( n779 & ~n778 ) | ( n779 & n782 ) | ( ~n778 & n782 ) ;
  assign n784 = n778 | n783 ;
  assign n556 = ~x335 & x463 ;
  assign n749 = ( x332 & ~x460 ) | ( x332 & 1'b0 ) | ( ~x460 & 1'b0 ) ;
  assign n750 = ( x333 & ~x461 ) | ( x333 & n749 ) | ( ~x461 & n749 ) ;
  assign n751 = ( x334 & ~x462 ) | ( x334 & n750 ) | ( ~x462 & n750 ) ;
  assign n752 = ~n556 & n751 ;
  assign n557 = ~x334 & x462 ;
  assign n558 = n556 | n557 ;
  assign n559 = ~x333 & x461 ;
  assign n560 = ~x332 & x460 ;
  assign n561 = ( n559 & ~n558 ) | ( n559 & n560 ) | ( ~n558 & n560 ) ;
  assign n562 = n558 | n561 ;
  assign n563 = ( x327 & ~x455 ) | ( x327 & 1'b0 ) | ( ~x455 & 1'b0 ) ;
  assign n735 = ~x331 & x459 ;
  assign n736 = ~x329 & x457 ;
  assign n737 = ~x330 & x458 ;
  assign n738 = ~x328 & x456 ;
  assign n739 = ( n737 & ~n736 ) | ( n737 & n738 ) | ( ~n736 & n738 ) ;
  assign n740 = ( n736 & ~n735 ) | ( n736 & n739 ) | ( ~n735 & n739 ) ;
  assign n741 = n735 | n740 ;
  assign n571 = ( x319 & ~x447 ) | ( x319 & 1'b0 ) | ( ~x447 & 1'b0 ) ;
  assign n714 = ~x321 & x449 ;
  assign n715 = ~x320 & x448 ;
  assign n716 = n714 | n715 ;
  assign n678 = x303 &  x431 ;
  assign n658 = x288 | x416 ;
  assign n612 = ( x256 & ~x384 ) | ( x256 & 1'b0 ) | ( ~x384 & 1'b0 ) ;
  assign n613 = ( x257 & ~x385 ) | ( x257 & n612 ) | ( ~x385 & n612 ) ;
  assign n614 = ( x258 & ~x386 ) | ( x258 & n613 ) | ( ~x386 & n613 ) ;
  assign n615 = ( x259 & ~x387 ) | ( x259 & n614 ) | ( ~x387 & n614 ) ;
  assign n616 = ( x260 & ~x388 ) | ( x260 & n615 ) | ( ~x388 & n615 ) ;
  assign n617 = ( x261 & ~x389 ) | ( x261 & n616 ) | ( ~x389 & n616 ) ;
  assign n618 = ( x262 & ~x390 ) | ( x262 & n617 ) | ( ~x390 & n617 ) ;
  assign n619 = ( x263 & ~x391 ) | ( x263 & n618 ) | ( ~x391 & n618 ) ;
  assign n620 = ( x264 & ~x392 ) | ( x264 & n619 ) | ( ~x392 & n619 ) ;
  assign n621 = ( x265 & ~x393 ) | ( x265 & n620 ) | ( ~x393 & n620 ) ;
  assign n622 = ( x266 & ~x394 ) | ( x266 & n621 ) | ( ~x394 & n621 ) ;
  assign n623 = ( x267 & ~x395 ) | ( x267 & n622 ) | ( ~x395 & n622 ) ;
  assign n624 = ( x268 & ~x396 ) | ( x268 & n623 ) | ( ~x396 & n623 ) ;
  assign n625 = ( x269 & ~x397 ) | ( x269 & n624 ) | ( ~x397 & n624 ) ;
  assign n626 = ( x270 & ~x398 ) | ( x270 & n625 ) | ( ~x398 & n625 ) ;
  assign n627 = ( x271 & ~x399 ) | ( x271 & n626 ) | ( ~x399 & n626 ) ;
  assign n628 = ( x272 & ~x400 ) | ( x272 & n627 ) | ( ~x400 & n627 ) ;
  assign n629 = ( x273 & ~x401 ) | ( x273 & n628 ) | ( ~x401 & n628 ) ;
  assign n630 = ( x274 & ~x402 ) | ( x274 & n629 ) | ( ~x402 & n629 ) ;
  assign n631 = ( x275 & ~x403 ) | ( x275 & n630 ) | ( ~x403 & n630 ) ;
  assign n632 = ( x276 & ~x404 ) | ( x276 & n631 ) | ( ~x404 & n631 ) ;
  assign n633 = ( x277 & ~x405 ) | ( x277 & n632 ) | ( ~x405 & n632 ) ;
  assign n634 = ( x278 & ~x406 ) | ( x278 & n633 ) | ( ~x406 & n633 ) ;
  assign n635 = ( x279 & ~x407 ) | ( x279 & n634 ) | ( ~x407 & n634 ) ;
  assign n636 = ( x280 & ~x408 ) | ( x280 & n635 ) | ( ~x408 & n635 ) ;
  assign n637 = ( x281 & ~x409 ) | ( x281 & n636 ) | ( ~x409 & n636 ) ;
  assign n638 = ( x282 & ~x410 ) | ( x282 & n637 ) | ( ~x410 & n637 ) ;
  assign n639 = ( x283 & ~x411 ) | ( x283 & n638 ) | ( ~x411 & n638 ) ;
  assign n640 = ( x284 & ~x412 ) | ( x284 & n639 ) | ( ~x412 & n639 ) ;
  assign n641 = ( x285 & ~x413 ) | ( x285 & n640 ) | ( ~x413 & n640 ) ;
  assign n642 = ( x286 & ~x414 ) | ( x286 & n641 ) | ( ~x414 & n641 ) ;
  assign n643 = ( x287 & ~x415 ) | ( x287 & n642 ) | ( ~x415 & n642 ) ;
  assign n644 = ~x295 & x423 ;
  assign n645 = ~x294 & x422 ;
  assign n646 = n644 | n645 ;
  assign n647 = ~x292 & x420 ;
  assign n648 = ~x293 & x421 ;
  assign n649 = ( n647 & ~n646 ) | ( n647 & n648 ) | ( ~n646 & n648 ) ;
  assign n650 = n646 | n649 ;
  assign n651 = x289 &  x417 ;
  assign n652 = ~x291 & x419 ;
  assign n653 = ~x290 & x418 ;
  assign n654 = n652 | n653 ;
  assign n655 = ( x417 & ~n651 ) | ( x417 & n654 ) | ( ~n651 & n654 ) ;
  assign n656 = n650 | n655 ;
  assign n657 = ( n643 & ~n656 ) | ( n643 & 1'b0 ) | ( ~n656 & 1'b0 ) ;
  assign n659 = ( x288 & ~n658 ) | ( x288 & n657 ) | ( ~n658 & n657 ) ;
  assign n660 = ( x288 & ~x416 ) | ( x288 & 1'b0 ) | ( ~x416 & 1'b0 ) ;
  assign n661 = ( x289 & ~x417 ) | ( x289 & n660 ) | ( ~x417 & n660 ) ;
  assign n662 = ( x290 & ~x418 ) | ( x290 & n661 ) | ( ~x418 & n661 ) ;
  assign n663 = ( x291 & ~x419 ) | ( x291 & n662 ) | ( ~x419 & n662 ) ;
  assign n668 = n663 | n650 ;
  assign n664 = ( x292 & ~x420 ) | ( x292 & 1'b0 ) | ( ~x420 & 1'b0 ) ;
  assign n665 = ( x293 & ~x421 ) | ( x293 & n664 ) | ( ~x421 & n664 ) ;
  assign n666 = ( x294 & ~x422 ) | ( x294 & n665 ) | ( ~x422 & n665 ) ;
  assign n667 = ( x295 & ~x423 ) | ( x295 & n666 ) | ( ~x423 & n666 ) ;
  assign n669 = ( n668 & ~n650 ) | ( n668 & n667 ) | ( ~n650 & n667 ) ;
  assign n670 = n659 | n669 ;
  assign n592 = ~x303 & x431 ;
  assign n593 = ~x302 & x430 ;
  assign n594 = n592 | n593 ;
  assign n595 = ~x300 & x428 ;
  assign n596 = ~x301 & x429 ;
  assign n597 = ( n595 & ~n594 ) | ( n595 & n596 ) | ( ~n594 & n596 ) ;
  assign n598 = n594 | n597 ;
  assign n599 = ~x299 & x427 ;
  assign n605 = ~x297 & x425 ;
  assign n606 = ~x298 & x426 ;
  assign n607 = ~x296 & x424 ;
  assign n608 = ( n606 & ~n605 ) | ( n606 & n607 ) | ( ~n605 & n607 ) ;
  assign n609 = ( n605 & ~n599 ) | ( n605 & n608 ) | ( ~n599 & n608 ) ;
  assign n610 = n599 | n609 ;
  assign n611 = n598 | n610 ;
  assign n676 = n670 | n611 ;
  assign n600 = ( x296 & ~x424 ) | ( x296 & 1'b0 ) | ( ~x424 & 1'b0 ) ;
  assign n601 = ( x297 & ~x425 ) | ( x297 & n600 ) | ( ~x425 & n600 ) ;
  assign n602 = ( x298 & ~x426 ) | ( x298 & n601 ) | ( ~x426 & n601 ) ;
  assign n603 = ( x299 & ~x427 ) | ( x299 & n602 ) | ( ~x427 & n602 ) ;
  assign n604 = ~n598 & n603 ;
  assign n671 = ( x300 & ~x428 ) | ( x300 & 1'b0 ) | ( ~x428 & 1'b0 ) ;
  assign n672 = ( x301 & ~x429 ) | ( x301 & n671 ) | ( ~x429 & n671 ) ;
  assign n673 = ( x302 & ~x430 ) | ( x302 & n672 ) | ( ~x430 & n672 ) ;
  assign n674 = ~n592 & n673 ;
  assign n675 = n604 | n674 ;
  assign n677 = ( n676 & ~n611 ) | ( n676 & n675 ) | ( ~n611 & n675 ) ;
  assign n679 = ( x303 & ~n678 ) | ( x303 & n677 ) | ( ~n678 & n677 ) ;
  assign n680 = ~x311 & x439 ;
  assign n681 = ~x309 & x437 ;
  assign n682 = ~x310 & x438 ;
  assign n683 = ~x308 & x436 ;
  assign n684 = ( n682 & ~n681 ) | ( n682 & n683 ) | ( ~n681 & n683 ) ;
  assign n685 = ( n681 & ~n680 ) | ( n681 & n684 ) | ( ~n680 & n684 ) ;
  assign n686 = n680 | n685 ;
  assign n687 = x305 &  x433 ;
  assign n688 = ~x307 & x435 ;
  assign n689 = ~x306 & x434 ;
  assign n690 = n688 | n689 ;
  assign n691 = ( x433 & ~n687 ) | ( x433 & n690 ) | ( ~n687 & n690 ) ;
  assign n692 = n686 | n691 ;
  assign n693 = x304 | x432 ;
  assign n694 = ( n692 & ~x304 ) | ( n692 & n693 ) | ( ~x304 & n693 ) ;
  assign n710 = n679 &  n694 ;
  assign n579 = ~x315 & x443 ;
  assign n585 = ~x314 & x442 ;
  assign n572 = ~x319 & x447 ;
  assign n573 = ~x318 & x446 ;
  assign n574 = n572 | n573 ;
  assign n575 = ~x316 & x444 ;
  assign n576 = ~x317 & x445 ;
  assign n577 = ( n575 & ~n574 ) | ( n575 & n576 ) | ( ~n574 & n576 ) ;
  assign n578 = n574 | n577 ;
  assign n586 = ~x313 & x441 ;
  assign n587 = ~x312 & x440 ;
  assign n588 = ( n586 & ~n578 ) | ( n586 & n587 ) | ( ~n578 & n587 ) ;
  assign n589 = n578 | n588 ;
  assign n590 = ( n585 & ~n579 ) | ( n585 & n589 ) | ( ~n579 & n589 ) ;
  assign n591 = n579 | n590 ;
  assign n699 = ( x308 & ~x436 ) | ( x308 & 1'b0 ) | ( ~x436 & 1'b0 ) ;
  assign n700 = ( x309 & ~x437 ) | ( x309 & n699 ) | ( ~x437 & n699 ) ;
  assign n701 = ( x310 & ~x438 ) | ( x310 & n700 ) | ( ~x438 & n700 ) ;
  assign n702 = ( x311 & ~x439 ) | ( x311 & n701 ) | ( ~x439 & n701 ) ;
  assign n695 = ( x304 & ~x432 ) | ( x304 & 1'b0 ) | ( ~x432 & 1'b0 ) ;
  assign n696 = ( x305 & ~x433 ) | ( x305 & n695 ) | ( ~x433 & n695 ) ;
  assign n697 = ( x306 & ~x434 ) | ( x306 & n696 ) | ( ~x434 & n696 ) ;
  assign n698 = ( x307 & ~x435 ) | ( x307 & n697 ) | ( ~x435 & n697 ) ;
  assign n703 = n686 | n698 ;
  assign n704 = ( n702 & ~n686 ) | ( n702 & n703 ) | ( ~n686 & n703 ) ;
  assign n709 = n591 | n704 ;
  assign n711 = ( n679 & ~n710 ) | ( n679 & n709 ) | ( ~n710 & n709 ) ;
  assign n580 = ( x312 & ~x440 ) | ( x312 & 1'b0 ) | ( ~x440 & 1'b0 ) ;
  assign n581 = ( x313 & ~x441 ) | ( x313 & n580 ) | ( ~x441 & n580 ) ;
  assign n582 = ( x314 & ~x442 ) | ( x314 & n581 ) | ( ~x442 & n581 ) ;
  assign n583 = ( x315 & ~x443 ) | ( x315 & n582 ) | ( ~x443 & n582 ) ;
  assign n584 = ~n578 & n583 ;
  assign n705 = ( x316 & ~x444 ) | ( x316 & 1'b0 ) | ( ~x444 & 1'b0 ) ;
  assign n706 = ( x317 & ~x445 ) | ( x317 & n705 ) | ( ~x445 & n705 ) ;
  assign n707 = ( x318 & ~x446 ) | ( x318 & n706 ) | ( ~x446 & n706 ) ;
  assign n708 = ~n572 & n707 ;
  assign n712 = n584 | n708 ;
  assign n713 = ( n711 & ~n591 ) | ( n711 & n712 ) | ( ~n591 & n712 ) ;
  assign n717 = ~n571 & n713 ;
  assign n718 = ( n571 & ~n716 ) | ( n571 & n717 ) | ( ~n716 & n717 ) ;
  assign n719 = ~x323 & x451 ;
  assign n720 = ~x322 & x450 ;
  assign n721 = n719 | n720 ;
  assign n726 = ~n716 & n721 ;
  assign n727 = ( n571 & n717 ) | ( n571 & n726 ) | ( n717 & n726 ) ;
  assign n564 = ~x327 & x455 ;
  assign n565 = ~x326 & x454 ;
  assign n566 = n564 | n565 ;
  assign n567 = ~x325 & x453 ;
  assign n568 = ~x324 & x452 ;
  assign n569 = ( n567 & ~n566 ) | ( n567 & n568 ) | ( ~n566 & n568 ) ;
  assign n570 = n566 | n569 ;
  assign n722 = ( x320 & ~x448 ) | ( x320 & 1'b0 ) | ( ~x448 & 1'b0 ) ;
  assign n723 = ( x321 & ~x449 ) | ( x321 & n722 ) | ( ~x449 & n722 ) ;
  assign n724 = ( x322 & ~x450 ) | ( x322 & n723 ) | ( ~x450 & n723 ) ;
  assign n725 = ( x323 & ~x451 ) | ( x323 & n724 ) | ( ~x451 & n724 ) ;
  assign n728 = n570 | n725 ;
  assign n729 = ( n718 & ~n727 ) | ( n718 & n728 ) | ( ~n727 & n728 ) ;
  assign n730 = ( x324 & ~x452 ) | ( x324 & 1'b0 ) | ( ~x452 & 1'b0 ) ;
  assign n731 = ( x325 & ~x453 ) | ( x325 & n730 ) | ( ~x453 & n730 ) ;
  assign n732 = ( x326 & ~x454 ) | ( x326 & n731 ) | ( ~x454 & n731 ) ;
  assign n733 = ~n564 & n732 ;
  assign n734 = ( n729 & ~n570 ) | ( n729 & n733 ) | ( ~n570 & n733 ) ;
  assign n742 = ~n563 & n734 ;
  assign n743 = ( n563 & ~n741 ) | ( n563 & n742 ) | ( ~n741 & n742 ) ;
  assign n744 = ( x328 & ~x456 ) | ( x328 & 1'b0 ) | ( ~x456 & 1'b0 ) ;
  assign n745 = ( x329 & ~x457 ) | ( x329 & n744 ) | ( ~x457 & n744 ) ;
  assign n746 = ( x330 & ~x458 ) | ( x330 & n745 ) | ( ~x458 & n745 ) ;
  assign n747 = ( x331 & ~x459 ) | ( x331 & n746 ) | ( ~x459 & n746 ) ;
  assign n748 = n743 | n747 ;
  assign n753 = n562 | n748 ;
  assign n754 = ( n752 & ~n562 ) | ( n752 & n753 ) | ( ~n562 & n753 ) ;
  assign n759 = ~x339 & x467 ;
  assign n760 = ~x338 & x466 ;
  assign n761 = n759 | n760 ;
  assign n762 = ~x337 & x465 ;
  assign n763 = n761 | n762 ;
  assign n757 = n748 | n562 ;
  assign n755 = ( x335 & ~x463 ) | ( x335 & 1'b0 ) | ( ~x463 & 1'b0 ) ;
  assign n756 = ~n752 & n755 ;
  assign n758 = ( n562 & ~n757 ) | ( n562 & n756 ) | ( ~n757 & n756 ) ;
  assign n764 = ( n754 & ~n763 ) | ( n754 & n758 ) | ( ~n763 & n758 ) ;
  assign n765 = ~x336 & x464 ;
  assign n771 = n765 &  n764 ;
  assign n549 = ~x343 & x471 ;
  assign n550 = ~x342 & x470 ;
  assign n551 = n549 | n550 ;
  assign n552 = ~x341 & x469 ;
  assign n553 = ~x340 & x468 ;
  assign n554 = ( n552 & ~n551 ) | ( n552 & n553 ) | ( ~n551 & n553 ) ;
  assign n555 = n551 | n554 ;
  assign n766 = ( x336 & ~x464 ) | ( x336 & 1'b0 ) | ( ~x464 & 1'b0 ) ;
  assign n767 = ( x337 & ~x465 ) | ( x337 & n766 ) | ( ~x465 & n766 ) ;
  assign n768 = ( x338 & ~x466 ) | ( x338 & n767 ) | ( ~x466 & n767 ) ;
  assign n769 = ( x339 & ~x467 ) | ( x339 & n768 ) | ( ~x467 & n768 ) ;
  assign n770 = n555 | n769 ;
  assign n772 = ( n764 & ~n771 ) | ( n764 & n770 ) | ( ~n771 & n770 ) ;
  assign n773 = ( x340 & ~x468 ) | ( x340 & 1'b0 ) | ( ~x468 & 1'b0 ) ;
  assign n774 = ( x341 & ~x469 ) | ( x341 & n773 ) | ( ~x469 & n773 ) ;
  assign n775 = ( x342 & ~x470 ) | ( x342 & n774 ) | ( ~x470 & n774 ) ;
  assign n776 = ~n549 & n775 ;
  assign n777 = ( n772 & ~n555 ) | ( n772 & n776 ) | ( ~n555 & n776 ) ;
  assign n785 = ~n548 & n777 ;
  assign n786 = ( n548 & ~n784 ) | ( n548 & n785 ) | ( ~n784 & n785 ) ;
  assign n787 = ( x344 & ~x472 ) | ( x344 & 1'b0 ) | ( ~x472 & 1'b0 ) ;
  assign n788 = ( x345 & ~x473 ) | ( x345 & n787 ) | ( ~x473 & n787 ) ;
  assign n789 = ( x346 & ~x474 ) | ( x346 & n788 ) | ( ~x474 & n788 ) ;
  assign n790 = ( x347 & ~x475 ) | ( x347 & n789 ) | ( ~x475 & n789 ) ;
  assign n791 = n786 | n790 ;
  assign n796 = n547 | n791 ;
  assign n797 = ( n795 & ~n547 ) | ( n795 & n796 ) | ( ~n547 & n796 ) ;
  assign n802 = ~x355 & x483 ;
  assign n803 = ~x354 & x482 ;
  assign n804 = n802 | n803 ;
  assign n805 = ~x353 & x481 ;
  assign n806 = n804 | n805 ;
  assign n800 = n791 | n547 ;
  assign n798 = ( x351 & ~x479 ) | ( x351 & 1'b0 ) | ( ~x479 & 1'b0 ) ;
  assign n799 = ~n795 & n798 ;
  assign n801 = ( n547 & ~n800 ) | ( n547 & n799 ) | ( ~n800 & n799 ) ;
  assign n807 = ( n797 & ~n806 ) | ( n797 & n801 ) | ( ~n806 & n801 ) ;
  assign n808 = ~x352 & x480 ;
  assign n814 = n808 &  n807 ;
  assign n534 = ~x359 & x487 ;
  assign n535 = ~x358 & x486 ;
  assign n536 = n534 | n535 ;
  assign n537 = ~x357 & x485 ;
  assign n538 = ~x356 & x484 ;
  assign n539 = ( n537 & ~n536 ) | ( n537 & n538 ) | ( ~n536 & n538 ) ;
  assign n540 = n536 | n539 ;
  assign n809 = ( x352 & ~x480 ) | ( x352 & 1'b0 ) | ( ~x480 & 1'b0 ) ;
  assign n810 = ( x353 & ~x481 ) | ( x353 & n809 ) | ( ~x481 & n809 ) ;
  assign n811 = ( x354 & ~x482 ) | ( x354 & n810 ) | ( ~x482 & n810 ) ;
  assign n812 = ( x355 & ~x483 ) | ( x355 & n811 ) | ( ~x483 & n811 ) ;
  assign n813 = n540 | n812 ;
  assign n815 = ( n807 & ~n814 ) | ( n807 & n813 ) | ( ~n814 & n813 ) ;
  assign n816 = ( x356 & ~x484 ) | ( x356 & 1'b0 ) | ( ~x484 & 1'b0 ) ;
  assign n817 = ( x357 & ~x485 ) | ( x357 & n816 ) | ( ~x485 & n816 ) ;
  assign n818 = ( x358 & ~x486 ) | ( x358 & n817 ) | ( ~x486 & n817 ) ;
  assign n819 = ~n534 & n818 ;
  assign n820 = ( n815 & ~n540 ) | ( n815 & n819 ) | ( ~n540 & n819 ) ;
  assign n828 = ~n533 & n820 ;
  assign n829 = ( n533 & ~n827 ) | ( n533 & n828 ) | ( ~n827 & n828 ) ;
  assign n830 = ( x360 & ~x488 ) | ( x360 & 1'b0 ) | ( ~x488 & 1'b0 ) ;
  assign n831 = ( x361 & ~x489 ) | ( x361 & n830 ) | ( ~x489 & n830 ) ;
  assign n832 = ( x362 & ~x490 ) | ( x362 & n831 ) | ( ~x490 & n831 ) ;
  assign n833 = ( x363 & ~x491 ) | ( x363 & n832 ) | ( ~x491 & n832 ) ;
  assign n834 = n829 | n833 ;
  assign n839 = n532 | n834 ;
  assign n840 = ( n838 & ~n532 ) | ( n838 & n839 ) | ( ~n532 & n839 ) ;
  assign n845 = ~x371 & x499 ;
  assign n846 = ~x370 & x498 ;
  assign n847 = n845 | n846 ;
  assign n848 = ~x369 & x497 ;
  assign n849 = n847 | n848 ;
  assign n843 = n834 | n532 ;
  assign n841 = ( x367 & ~x495 ) | ( x367 & 1'b0 ) | ( ~x495 & 1'b0 ) ;
  assign n842 = ~n838 & n841 ;
  assign n844 = ( n532 & ~n843 ) | ( n532 & n842 ) | ( ~n843 & n842 ) ;
  assign n850 = ( n840 & ~n849 ) | ( n840 & n844 ) | ( ~n849 & n844 ) ;
  assign n851 = ~x368 & x496 ;
  assign n857 = n851 &  n850 ;
  assign n519 = ~x375 & x503 ;
  assign n520 = ~x374 & x502 ;
  assign n521 = n519 | n520 ;
  assign n522 = ~x373 & x501 ;
  assign n523 = ~x372 & x500 ;
  assign n524 = ( n522 & ~n521 ) | ( n522 & n523 ) | ( ~n521 & n523 ) ;
  assign n525 = n521 | n524 ;
  assign n852 = ( x368 & ~x496 ) | ( x368 & 1'b0 ) | ( ~x496 & 1'b0 ) ;
  assign n853 = ( x369 & ~x497 ) | ( x369 & n852 ) | ( ~x497 & n852 ) ;
  assign n854 = ( x370 & ~x498 ) | ( x370 & n853 ) | ( ~x498 & n853 ) ;
  assign n855 = ( x371 & ~x499 ) | ( x371 & n854 ) | ( ~x499 & n854 ) ;
  assign n856 = n525 | n855 ;
  assign n858 = ( n850 & ~n857 ) | ( n850 & n856 ) | ( ~n857 & n856 ) ;
  assign n859 = ( x372 & ~x500 ) | ( x372 & 1'b0 ) | ( ~x500 & 1'b0 ) ;
  assign n860 = ( x373 & ~x501 ) | ( x373 & n859 ) | ( ~x501 & n859 ) ;
  assign n861 = ( x374 & ~x502 ) | ( x374 & n860 ) | ( ~x502 & n860 ) ;
  assign n862 = ~n519 & n861 ;
  assign n863 = ( n858 & ~n525 ) | ( n858 & n862 ) | ( ~n525 & n862 ) ;
  assign n871 = ~n518 & n863 ;
  assign n872 = ( n518 & ~n870 ) | ( n518 & n871 ) | ( ~n870 & n871 ) ;
  assign n880 = ( n517 & ~n879 ) | ( n517 & n872 ) | ( ~n879 & n872 ) ;
  assign n881 = ( x380 & ~x508 ) | ( x380 & 1'b0 ) | ( ~x508 & 1'b0 ) ;
  assign n882 = ( x381 & ~x509 ) | ( x381 & n881 ) | ( ~x509 & n881 ) ;
  assign n883 = ( x382 & ~x510 ) | ( x382 & n882 ) | ( ~x510 & n882 ) ;
  assign n884 = ( x511 & ~x383 ) | ( x511 & n883 ) | ( ~x383 & n883 ) ;
  assign n885 = n880 | n884 ;
  assign n886 = x384 | n885 ;
  assign n887 = ~x256 & n885 ;
  assign n888 = ( n886 & ~n887 ) | ( n886 & 1'b0 ) | ( ~n887 & 1'b0 ) ;
  assign n890 = ( x120 & ~x248 ) | ( x120 & 1'b0 ) | ( ~x248 & 1'b0 ) ;
  assign n891 = ( x121 & ~x249 ) | ( x121 & n890 ) | ( ~x249 & n890 ) ;
  assign n892 = ( x122 & ~x250 ) | ( x122 & n891 ) | ( ~x250 & n891 ) ;
  assign n893 = ( x123 & ~x251 ) | ( x123 & n892 ) | ( ~x251 & n892 ) ;
  assign n1249 = ~x124 & x252 ;
  assign n1253 = x127 &  x255 ;
  assign n1250 = ~x126 & x254 ;
  assign n1251 = ~x125 & x253 ;
  assign n1252 = n1250 | n1251 ;
  assign n1254 = ( x127 & ~n1253 ) | ( x127 & n1252 ) | ( ~n1253 & n1252 ) ;
  assign n1255 = n1249 | n1254 ;
  assign n894 = ( x119 & ~x247 ) | ( x119 & 1'b0 ) | ( ~x247 & 1'b0 ) ;
  assign n889 = ~x123 & x251 ;
  assign n1240 = ~x121 & x249 ;
  assign n1241 = ~x122 & x250 ;
  assign n1242 = ~x120 & x248 ;
  assign n1243 = ( n1241 & ~n1240 ) | ( n1241 & n1242 ) | ( ~n1240 & n1242 ) ;
  assign n1244 = ( n1240 & ~n889 ) | ( n1240 & n1243 ) | ( ~n889 & n1243 ) ;
  assign n1245 = n889 | n1244 ;
  assign n1246 = n893 | n1245 ;
  assign n902 = ~x111 & x239 ;
  assign n1211 = ( x108 & ~x236 ) | ( x108 & 1'b0 ) | ( ~x236 & 1'b0 ) ;
  assign n1212 = ( x109 & ~x237 ) | ( x109 & n1211 ) | ( ~x237 & n1211 ) ;
  assign n1213 = ( x110 & ~x238 ) | ( x110 & n1212 ) | ( ~x238 & n1212 ) ;
  assign n1214 = ~n902 & n1213 ;
  assign n903 = ~x110 & x238 ;
  assign n904 = n902 | n903 ;
  assign n905 = ~x109 & x237 ;
  assign n906 = ~x108 & x236 ;
  assign n907 = ( n905 & ~n904 ) | ( n905 & n906 ) | ( ~n904 & n906 ) ;
  assign n908 = n904 | n907 ;
  assign n909 = ( x103 & ~x231 ) | ( x103 & 1'b0 ) | ( ~x231 & 1'b0 ) ;
  assign n1197 = ~x107 & x235 ;
  assign n1198 = ~x105 & x233 ;
  assign n1199 = ~x106 & x234 ;
  assign n1200 = ~x104 & x232 ;
  assign n1201 = ( n1199 & ~n1198 ) | ( n1199 & n1200 ) | ( ~n1198 & n1200 ) ;
  assign n1202 = ( n1198 & ~n1197 ) | ( n1198 & n1201 ) | ( ~n1197 & n1201 ) ;
  assign n1203 = n1197 | n1202 ;
  assign n917 = ~x95 & x223 ;
  assign n1168 = ( x92 & ~x220 ) | ( x92 & 1'b0 ) | ( ~x220 & 1'b0 ) ;
  assign n1169 = ( x93 & ~x221 ) | ( x93 & n1168 ) | ( ~x221 & n1168 ) ;
  assign n1170 = ( x94 & ~x222 ) | ( x94 & n1169 ) | ( ~x222 & n1169 ) ;
  assign n1171 = ~n917 & n1170 ;
  assign n918 = ~x94 & x222 ;
  assign n919 = n917 | n918 ;
  assign n920 = ~x93 & x221 ;
  assign n921 = ~x92 & x220 ;
  assign n922 = ( n920 & ~n919 ) | ( n920 & n921 ) | ( ~n919 & n921 ) ;
  assign n923 = n919 | n922 ;
  assign n924 = ( x87 & ~x215 ) | ( x87 & 1'b0 ) | ( ~x215 & 1'b0 ) ;
  assign n1154 = ~x91 & x219 ;
  assign n1155 = ~x89 & x217 ;
  assign n1156 = ~x90 & x218 ;
  assign n1157 = ~x88 & x216 ;
  assign n1158 = ( n1156 & ~n1155 ) | ( n1156 & n1157 ) | ( ~n1155 & n1157 ) ;
  assign n1159 = ( n1155 & ~n1154 ) | ( n1155 & n1158 ) | ( ~n1154 & n1158 ) ;
  assign n1160 = n1154 | n1159 ;
  assign n932 = ~x79 & x207 ;
  assign n1125 = ( x76 & ~x204 ) | ( x76 & 1'b0 ) | ( ~x204 & 1'b0 ) ;
  assign n1126 = ( x77 & ~x205 ) | ( x77 & n1125 ) | ( ~x205 & n1125 ) ;
  assign n1127 = ( x78 & ~x206 ) | ( x78 & n1126 ) | ( ~x206 & n1126 ) ;
  assign n1128 = ~n932 & n1127 ;
  assign n933 = ~x78 & x206 ;
  assign n934 = n932 | n933 ;
  assign n935 = ~x77 & x205 ;
  assign n936 = ~x76 & x204 ;
  assign n937 = ( n935 & ~n934 ) | ( n935 & n936 ) | ( ~n934 & n936 ) ;
  assign n938 = n934 | n937 ;
  assign n939 = ( x71 & ~x199 ) | ( x71 & 1'b0 ) | ( ~x199 & 1'b0 ) ;
  assign n1111 = ~x75 & x203 ;
  assign n1112 = ~x73 & x201 ;
  assign n1113 = ~x74 & x202 ;
  assign n1114 = ~x72 & x200 ;
  assign n1115 = ( n1113 & ~n1112 ) | ( n1113 & n1114 ) | ( ~n1112 & n1114 ) ;
  assign n1116 = ( n1112 & ~n1111 ) | ( n1112 & n1115 ) | ( ~n1111 & n1115 ) ;
  assign n1117 = n1111 | n1116 ;
  assign n947 = ( x63 & ~x191 ) | ( x63 & 1'b0 ) | ( ~x191 & 1'b0 ) ;
  assign n1090 = ~x65 & x193 ;
  assign n1091 = ~x64 & x192 ;
  assign n1092 = n1090 | n1091 ;
  assign n1054 = x47 &  x175 ;
  assign n1034 = x32 | x160 ;
  assign n988 = ( x0 & ~x128 ) | ( x0 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n989 = ( x1 & ~x129 ) | ( x1 & n988 ) | ( ~x129 & n988 ) ;
  assign n990 = ( x2 & ~x130 ) | ( x2 & n989 ) | ( ~x130 & n989 ) ;
  assign n991 = ( x3 & ~x131 ) | ( x3 & n990 ) | ( ~x131 & n990 ) ;
  assign n992 = ( x4 & ~x132 ) | ( x4 & n991 ) | ( ~x132 & n991 ) ;
  assign n993 = ( x5 & ~x133 ) | ( x5 & n992 ) | ( ~x133 & n992 ) ;
  assign n994 = ( x6 & ~x134 ) | ( x6 & n993 ) | ( ~x134 & n993 ) ;
  assign n995 = ( x7 & ~x135 ) | ( x7 & n994 ) | ( ~x135 & n994 ) ;
  assign n996 = ( x8 & ~x136 ) | ( x8 & n995 ) | ( ~x136 & n995 ) ;
  assign n997 = ( x9 & ~x137 ) | ( x9 & n996 ) | ( ~x137 & n996 ) ;
  assign n998 = ( x10 & ~x138 ) | ( x10 & n997 ) | ( ~x138 & n997 ) ;
  assign n999 = ( x11 & ~x139 ) | ( x11 & n998 ) | ( ~x139 & n998 ) ;
  assign n1000 = ( x12 & ~x140 ) | ( x12 & n999 ) | ( ~x140 & n999 ) ;
  assign n1001 = ( x13 & ~x141 ) | ( x13 & n1000 ) | ( ~x141 & n1000 ) ;
  assign n1002 = ( x14 & ~x142 ) | ( x14 & n1001 ) | ( ~x142 & n1001 ) ;
  assign n1003 = ( x15 & ~x143 ) | ( x15 & n1002 ) | ( ~x143 & n1002 ) ;
  assign n1004 = ( x16 & ~x144 ) | ( x16 & n1003 ) | ( ~x144 & n1003 ) ;
  assign n1005 = ( x17 & ~x145 ) | ( x17 & n1004 ) | ( ~x145 & n1004 ) ;
  assign n1006 = ( x18 & ~x146 ) | ( x18 & n1005 ) | ( ~x146 & n1005 ) ;
  assign n1007 = ( x19 & ~x147 ) | ( x19 & n1006 ) | ( ~x147 & n1006 ) ;
  assign n1008 = ( x20 & ~x148 ) | ( x20 & n1007 ) | ( ~x148 & n1007 ) ;
  assign n1009 = ( x21 & ~x149 ) | ( x21 & n1008 ) | ( ~x149 & n1008 ) ;
  assign n1010 = ( x22 & ~x150 ) | ( x22 & n1009 ) | ( ~x150 & n1009 ) ;
  assign n1011 = ( x23 & ~x151 ) | ( x23 & n1010 ) | ( ~x151 & n1010 ) ;
  assign n1012 = ( x24 & ~x152 ) | ( x24 & n1011 ) | ( ~x152 & n1011 ) ;
  assign n1013 = ( x25 & ~x153 ) | ( x25 & n1012 ) | ( ~x153 & n1012 ) ;
  assign n1014 = ( x26 & ~x154 ) | ( x26 & n1013 ) | ( ~x154 & n1013 ) ;
  assign n1015 = ( x27 & ~x155 ) | ( x27 & n1014 ) | ( ~x155 & n1014 ) ;
  assign n1016 = ( x28 & ~x156 ) | ( x28 & n1015 ) | ( ~x156 & n1015 ) ;
  assign n1017 = ( x29 & ~x157 ) | ( x29 & n1016 ) | ( ~x157 & n1016 ) ;
  assign n1018 = ( x30 & ~x158 ) | ( x30 & n1017 ) | ( ~x158 & n1017 ) ;
  assign n1019 = ( x31 & ~x159 ) | ( x31 & n1018 ) | ( ~x159 & n1018 ) ;
  assign n1020 = ~x39 & x167 ;
  assign n1021 = ~x38 & x166 ;
  assign n1022 = n1020 | n1021 ;
  assign n1023 = ~x36 & x164 ;
  assign n1024 = ~x37 & x165 ;
  assign n1025 = ( n1023 & ~n1022 ) | ( n1023 & n1024 ) | ( ~n1022 & n1024 ) ;
  assign n1026 = n1022 | n1025 ;
  assign n1027 = x33 &  x161 ;
  assign n1028 = ~x35 & x163 ;
  assign n1029 = ~x34 & x162 ;
  assign n1030 = n1028 | n1029 ;
  assign n1031 = ( x161 & ~n1027 ) | ( x161 & n1030 ) | ( ~n1027 & n1030 ) ;
  assign n1032 = n1026 | n1031 ;
  assign n1033 = ( n1019 & ~n1032 ) | ( n1019 & 1'b0 ) | ( ~n1032 & 1'b0 ) ;
  assign n1035 = ( x32 & ~n1034 ) | ( x32 & n1033 ) | ( ~n1034 & n1033 ) ;
  assign n1036 = ( x32 & ~x160 ) | ( x32 & 1'b0 ) | ( ~x160 & 1'b0 ) ;
  assign n1037 = ( x33 & ~x161 ) | ( x33 & n1036 ) | ( ~x161 & n1036 ) ;
  assign n1038 = ( x34 & ~x162 ) | ( x34 & n1037 ) | ( ~x162 & n1037 ) ;
  assign n1039 = ( x35 & ~x163 ) | ( x35 & n1038 ) | ( ~x163 & n1038 ) ;
  assign n1044 = n1039 | n1026 ;
  assign n1040 = ( x36 & ~x164 ) | ( x36 & 1'b0 ) | ( ~x164 & 1'b0 ) ;
  assign n1041 = ( x37 & ~x165 ) | ( x37 & n1040 ) | ( ~x165 & n1040 ) ;
  assign n1042 = ( x38 & ~x166 ) | ( x38 & n1041 ) | ( ~x166 & n1041 ) ;
  assign n1043 = ( x39 & ~x167 ) | ( x39 & n1042 ) | ( ~x167 & n1042 ) ;
  assign n1045 = ( n1044 & ~n1026 ) | ( n1044 & n1043 ) | ( ~n1026 & n1043 ) ;
  assign n1046 = n1035 | n1045 ;
  assign n968 = ~x47 & x175 ;
  assign n969 = ~x46 & x174 ;
  assign n970 = n968 | n969 ;
  assign n971 = ~x44 & x172 ;
  assign n972 = ~x45 & x173 ;
  assign n973 = ( n971 & ~n970 ) | ( n971 & n972 ) | ( ~n970 & n972 ) ;
  assign n974 = n970 | n973 ;
  assign n975 = ~x43 & x171 ;
  assign n981 = ~x41 & x169 ;
  assign n982 = ~x42 & x170 ;
  assign n983 = ~x40 & x168 ;
  assign n984 = ( n982 & ~n981 ) | ( n982 & n983 ) | ( ~n981 & n983 ) ;
  assign n985 = ( n981 & ~n975 ) | ( n981 & n984 ) | ( ~n975 & n984 ) ;
  assign n986 = n975 | n985 ;
  assign n987 = n974 | n986 ;
  assign n1052 = n1046 | n987 ;
  assign n976 = ( x40 & ~x168 ) | ( x40 & 1'b0 ) | ( ~x168 & 1'b0 ) ;
  assign n977 = ( x41 & ~x169 ) | ( x41 & n976 ) | ( ~x169 & n976 ) ;
  assign n978 = ( x42 & ~x170 ) | ( x42 & n977 ) | ( ~x170 & n977 ) ;
  assign n979 = ( x43 & ~x171 ) | ( x43 & n978 ) | ( ~x171 & n978 ) ;
  assign n980 = ~n974 & n979 ;
  assign n1047 = ( x44 & ~x172 ) | ( x44 & 1'b0 ) | ( ~x172 & 1'b0 ) ;
  assign n1048 = ( x45 & ~x173 ) | ( x45 & n1047 ) | ( ~x173 & n1047 ) ;
  assign n1049 = ( x46 & ~x174 ) | ( x46 & n1048 ) | ( ~x174 & n1048 ) ;
  assign n1050 = ~n968 & n1049 ;
  assign n1051 = n980 | n1050 ;
  assign n1053 = ( n1052 & ~n987 ) | ( n1052 & n1051 ) | ( ~n987 & n1051 ) ;
  assign n1055 = ( x47 & ~n1054 ) | ( x47 & n1053 ) | ( ~n1054 & n1053 ) ;
  assign n1056 = ~x55 & x183 ;
  assign n1057 = ~x53 & x181 ;
  assign n1058 = ~x54 & x182 ;
  assign n1059 = ~x52 & x180 ;
  assign n1060 = ( n1058 & ~n1057 ) | ( n1058 & n1059 ) | ( ~n1057 & n1059 ) ;
  assign n1061 = ( n1057 & ~n1056 ) | ( n1057 & n1060 ) | ( ~n1056 & n1060 ) ;
  assign n1062 = n1056 | n1061 ;
  assign n1063 = x49 &  x177 ;
  assign n1064 = ~x51 & x179 ;
  assign n1065 = ~x50 & x178 ;
  assign n1066 = n1064 | n1065 ;
  assign n1067 = ( x177 & ~n1063 ) | ( x177 & n1066 ) | ( ~n1063 & n1066 ) ;
  assign n1068 = n1062 | n1067 ;
  assign n1069 = x48 | x176 ;
  assign n1070 = ( n1068 & ~x48 ) | ( n1068 & n1069 ) | ( ~x48 & n1069 ) ;
  assign n1086 = n1055 &  n1070 ;
  assign n955 = ~x59 & x187 ;
  assign n961 = ~x58 & x186 ;
  assign n948 = ~x63 & x191 ;
  assign n949 = ~x62 & x190 ;
  assign n950 = n948 | n949 ;
  assign n951 = ~x60 & x188 ;
  assign n952 = ~x61 & x189 ;
  assign n953 = ( n951 & ~n950 ) | ( n951 & n952 ) | ( ~n950 & n952 ) ;
  assign n954 = n950 | n953 ;
  assign n962 = ~x57 & x185 ;
  assign n963 = ~x56 & x184 ;
  assign n964 = ( n962 & ~n954 ) | ( n962 & n963 ) | ( ~n954 & n963 ) ;
  assign n965 = n954 | n964 ;
  assign n966 = ( n961 & ~n955 ) | ( n961 & n965 ) | ( ~n955 & n965 ) ;
  assign n967 = n955 | n966 ;
  assign n1075 = ( x52 & ~x180 ) | ( x52 & 1'b0 ) | ( ~x180 & 1'b0 ) ;
  assign n1076 = ( x53 & ~x181 ) | ( x53 & n1075 ) | ( ~x181 & n1075 ) ;
  assign n1077 = ( x54 & ~x182 ) | ( x54 & n1076 ) | ( ~x182 & n1076 ) ;
  assign n1078 = ( x55 & ~x183 ) | ( x55 & n1077 ) | ( ~x183 & n1077 ) ;
  assign n1071 = ( x48 & ~x176 ) | ( x48 & 1'b0 ) | ( ~x176 & 1'b0 ) ;
  assign n1072 = ( x49 & ~x177 ) | ( x49 & n1071 ) | ( ~x177 & n1071 ) ;
  assign n1073 = ( x50 & ~x178 ) | ( x50 & n1072 ) | ( ~x178 & n1072 ) ;
  assign n1074 = ( x51 & ~x179 ) | ( x51 & n1073 ) | ( ~x179 & n1073 ) ;
  assign n1079 = n1062 | n1074 ;
  assign n1080 = ( n1078 & ~n1062 ) | ( n1078 & n1079 ) | ( ~n1062 & n1079 ) ;
  assign n1085 = n967 | n1080 ;
  assign n1087 = ( n1055 & ~n1086 ) | ( n1055 & n1085 ) | ( ~n1086 & n1085 ) ;
  assign n956 = ( x56 & ~x184 ) | ( x56 & 1'b0 ) | ( ~x184 & 1'b0 ) ;
  assign n957 = ( x57 & ~x185 ) | ( x57 & n956 ) | ( ~x185 & n956 ) ;
  assign n958 = ( x58 & ~x186 ) | ( x58 & n957 ) | ( ~x186 & n957 ) ;
  assign n959 = ( x59 & ~x187 ) | ( x59 & n958 ) | ( ~x187 & n958 ) ;
  assign n960 = ~n954 & n959 ;
  assign n1081 = ( x60 & ~x188 ) | ( x60 & 1'b0 ) | ( ~x188 & 1'b0 ) ;
  assign n1082 = ( x61 & ~x189 ) | ( x61 & n1081 ) | ( ~x189 & n1081 ) ;
  assign n1083 = ( x62 & ~x190 ) | ( x62 & n1082 ) | ( ~x190 & n1082 ) ;
  assign n1084 = ~n948 & n1083 ;
  assign n1088 = n960 | n1084 ;
  assign n1089 = ( n1087 & ~n967 ) | ( n1087 & n1088 ) | ( ~n967 & n1088 ) ;
  assign n1093 = ~n947 & n1089 ;
  assign n1094 = ( n947 & ~n1092 ) | ( n947 & n1093 ) | ( ~n1092 & n1093 ) ;
  assign n1095 = ~x67 & x195 ;
  assign n1096 = ~x66 & x194 ;
  assign n1097 = n1095 | n1096 ;
  assign n1102 = ~n1092 & n1097 ;
  assign n1103 = ( n947 & n1093 ) | ( n947 & n1102 ) | ( n1093 & n1102 ) ;
  assign n940 = ~x71 & x199 ;
  assign n941 = ~x70 & x198 ;
  assign n942 = n940 | n941 ;
  assign n943 = ~x69 & x197 ;
  assign n944 = ~x68 & x196 ;
  assign n945 = ( n943 & ~n942 ) | ( n943 & n944 ) | ( ~n942 & n944 ) ;
  assign n946 = n942 | n945 ;
  assign n1098 = ( x64 & ~x192 ) | ( x64 & 1'b0 ) | ( ~x192 & 1'b0 ) ;
  assign n1099 = ( x65 & ~x193 ) | ( x65 & n1098 ) | ( ~x193 & n1098 ) ;
  assign n1100 = ( x66 & ~x194 ) | ( x66 & n1099 ) | ( ~x194 & n1099 ) ;
  assign n1101 = ( x67 & ~x195 ) | ( x67 & n1100 ) | ( ~x195 & n1100 ) ;
  assign n1104 = n946 | n1101 ;
  assign n1105 = ( n1094 & ~n1103 ) | ( n1094 & n1104 ) | ( ~n1103 & n1104 ) ;
  assign n1106 = ( x68 & ~x196 ) | ( x68 & 1'b0 ) | ( ~x196 & 1'b0 ) ;
  assign n1107 = ( x69 & ~x197 ) | ( x69 & n1106 ) | ( ~x197 & n1106 ) ;
  assign n1108 = ( x70 & ~x198 ) | ( x70 & n1107 ) | ( ~x198 & n1107 ) ;
  assign n1109 = ~n940 & n1108 ;
  assign n1110 = ( n1105 & ~n946 ) | ( n1105 & n1109 ) | ( ~n946 & n1109 ) ;
  assign n1118 = ~n939 & n1110 ;
  assign n1119 = ( n939 & ~n1117 ) | ( n939 & n1118 ) | ( ~n1117 & n1118 ) ;
  assign n1120 = ( x72 & ~x200 ) | ( x72 & 1'b0 ) | ( ~x200 & 1'b0 ) ;
  assign n1121 = ( x73 & ~x201 ) | ( x73 & n1120 ) | ( ~x201 & n1120 ) ;
  assign n1122 = ( x74 & ~x202 ) | ( x74 & n1121 ) | ( ~x202 & n1121 ) ;
  assign n1123 = ( x75 & ~x203 ) | ( x75 & n1122 ) | ( ~x203 & n1122 ) ;
  assign n1124 = n1119 | n1123 ;
  assign n1129 = n938 | n1124 ;
  assign n1130 = ( n1128 & ~n938 ) | ( n1128 & n1129 ) | ( ~n938 & n1129 ) ;
  assign n1135 = ~x83 & x211 ;
  assign n1136 = ~x82 & x210 ;
  assign n1137 = n1135 | n1136 ;
  assign n1138 = ~x81 & x209 ;
  assign n1139 = n1137 | n1138 ;
  assign n1133 = n1124 | n938 ;
  assign n1131 = ( x79 & ~x207 ) | ( x79 & 1'b0 ) | ( ~x207 & 1'b0 ) ;
  assign n1132 = ~n1128 & n1131 ;
  assign n1134 = ( n938 & ~n1133 ) | ( n938 & n1132 ) | ( ~n1133 & n1132 ) ;
  assign n1140 = ( n1130 & ~n1139 ) | ( n1130 & n1134 ) | ( ~n1139 & n1134 ) ;
  assign n1141 = ~x80 & x208 ;
  assign n1147 = n1141 &  n1140 ;
  assign n925 = ~x87 & x215 ;
  assign n926 = ~x86 & x214 ;
  assign n927 = n925 | n926 ;
  assign n928 = ~x85 & x213 ;
  assign n929 = ~x84 & x212 ;
  assign n930 = ( n928 & ~n927 ) | ( n928 & n929 ) | ( ~n927 & n929 ) ;
  assign n931 = n927 | n930 ;
  assign n1142 = ( x80 & ~x208 ) | ( x80 & 1'b0 ) | ( ~x208 & 1'b0 ) ;
  assign n1143 = ( x81 & ~x209 ) | ( x81 & n1142 ) | ( ~x209 & n1142 ) ;
  assign n1144 = ( x82 & ~x210 ) | ( x82 & n1143 ) | ( ~x210 & n1143 ) ;
  assign n1145 = ( x83 & ~x211 ) | ( x83 & n1144 ) | ( ~x211 & n1144 ) ;
  assign n1146 = n931 | n1145 ;
  assign n1148 = ( n1140 & ~n1147 ) | ( n1140 & n1146 ) | ( ~n1147 & n1146 ) ;
  assign n1149 = ( x84 & ~x212 ) | ( x84 & 1'b0 ) | ( ~x212 & 1'b0 ) ;
  assign n1150 = ( x85 & ~x213 ) | ( x85 & n1149 ) | ( ~x213 & n1149 ) ;
  assign n1151 = ( x86 & ~x214 ) | ( x86 & n1150 ) | ( ~x214 & n1150 ) ;
  assign n1152 = ~n925 & n1151 ;
  assign n1153 = ( n1148 & ~n931 ) | ( n1148 & n1152 ) | ( ~n931 & n1152 ) ;
  assign n1161 = ~n924 & n1153 ;
  assign n1162 = ( n924 & ~n1160 ) | ( n924 & n1161 ) | ( ~n1160 & n1161 ) ;
  assign n1163 = ( x88 & ~x216 ) | ( x88 & 1'b0 ) | ( ~x216 & 1'b0 ) ;
  assign n1164 = ( x89 & ~x217 ) | ( x89 & n1163 ) | ( ~x217 & n1163 ) ;
  assign n1165 = ( x90 & ~x218 ) | ( x90 & n1164 ) | ( ~x218 & n1164 ) ;
  assign n1166 = ( x91 & ~x219 ) | ( x91 & n1165 ) | ( ~x219 & n1165 ) ;
  assign n1167 = n1162 | n1166 ;
  assign n1172 = n923 | n1167 ;
  assign n1173 = ( n1171 & ~n923 ) | ( n1171 & n1172 ) | ( ~n923 & n1172 ) ;
  assign n1178 = ~x99 & x227 ;
  assign n1179 = ~x98 & x226 ;
  assign n1180 = n1178 | n1179 ;
  assign n1181 = ~x97 & x225 ;
  assign n1182 = n1180 | n1181 ;
  assign n1176 = n1167 | n923 ;
  assign n1174 = ( x95 & ~x223 ) | ( x95 & 1'b0 ) | ( ~x223 & 1'b0 ) ;
  assign n1175 = ~n1171 & n1174 ;
  assign n1177 = ( n923 & ~n1176 ) | ( n923 & n1175 ) | ( ~n1176 & n1175 ) ;
  assign n1183 = ( n1173 & ~n1182 ) | ( n1173 & n1177 ) | ( ~n1182 & n1177 ) ;
  assign n1184 = ~x96 & x224 ;
  assign n1190 = n1184 &  n1183 ;
  assign n910 = ~x103 & x231 ;
  assign n911 = ~x102 & x230 ;
  assign n912 = n910 | n911 ;
  assign n913 = ~x101 & x229 ;
  assign n914 = ~x100 & x228 ;
  assign n915 = ( n913 & ~n912 ) | ( n913 & n914 ) | ( ~n912 & n914 ) ;
  assign n916 = n912 | n915 ;
  assign n1185 = ( x96 & ~x224 ) | ( x96 & 1'b0 ) | ( ~x224 & 1'b0 ) ;
  assign n1186 = ( x97 & ~x225 ) | ( x97 & n1185 ) | ( ~x225 & n1185 ) ;
  assign n1187 = ( x98 & ~x226 ) | ( x98 & n1186 ) | ( ~x226 & n1186 ) ;
  assign n1188 = ( x99 & ~x227 ) | ( x99 & n1187 ) | ( ~x227 & n1187 ) ;
  assign n1189 = n916 | n1188 ;
  assign n1191 = ( n1183 & ~n1190 ) | ( n1183 & n1189 ) | ( ~n1190 & n1189 ) ;
  assign n1192 = ( x100 & ~x228 ) | ( x100 & 1'b0 ) | ( ~x228 & 1'b0 ) ;
  assign n1193 = ( x101 & ~x229 ) | ( x101 & n1192 ) | ( ~x229 & n1192 ) ;
  assign n1194 = ( x102 & ~x230 ) | ( x102 & n1193 ) | ( ~x230 & n1193 ) ;
  assign n1195 = ~n910 & n1194 ;
  assign n1196 = ( n1191 & ~n916 ) | ( n1191 & n1195 ) | ( ~n916 & n1195 ) ;
  assign n1204 = ~n909 & n1196 ;
  assign n1205 = ( n909 & ~n1203 ) | ( n909 & n1204 ) | ( ~n1203 & n1204 ) ;
  assign n1206 = ( x104 & ~x232 ) | ( x104 & 1'b0 ) | ( ~x232 & 1'b0 ) ;
  assign n1207 = ( x105 & ~x233 ) | ( x105 & n1206 ) | ( ~x233 & n1206 ) ;
  assign n1208 = ( x106 & ~x234 ) | ( x106 & n1207 ) | ( ~x234 & n1207 ) ;
  assign n1209 = ( x107 & ~x235 ) | ( x107 & n1208 ) | ( ~x235 & n1208 ) ;
  assign n1210 = n1205 | n1209 ;
  assign n1215 = n908 | n1210 ;
  assign n1216 = ( n1214 & ~n908 ) | ( n1214 & n1215 ) | ( ~n908 & n1215 ) ;
  assign n1221 = ~x115 & x243 ;
  assign n1222 = ~x114 & x242 ;
  assign n1223 = n1221 | n1222 ;
  assign n1224 = ~x113 & x241 ;
  assign n1225 = n1223 | n1224 ;
  assign n1219 = n1210 | n908 ;
  assign n1217 = ( x111 & ~x239 ) | ( x111 & 1'b0 ) | ( ~x239 & 1'b0 ) ;
  assign n1218 = ~n1214 & n1217 ;
  assign n1220 = ( n908 & ~n1219 ) | ( n908 & n1218 ) | ( ~n1219 & n1218 ) ;
  assign n1226 = ( n1216 & ~n1225 ) | ( n1216 & n1220 ) | ( ~n1225 & n1220 ) ;
  assign n1227 = ~x112 & x240 ;
  assign n1233 = n1227 &  n1226 ;
  assign n895 = ~x119 & x247 ;
  assign n896 = ~x118 & x246 ;
  assign n897 = n895 | n896 ;
  assign n898 = ~x117 & x245 ;
  assign n899 = ~x116 & x244 ;
  assign n900 = ( n898 & ~n897 ) | ( n898 & n899 ) | ( ~n897 & n899 ) ;
  assign n901 = n897 | n900 ;
  assign n1228 = ( x112 & ~x240 ) | ( x112 & 1'b0 ) | ( ~x240 & 1'b0 ) ;
  assign n1229 = ( x113 & ~x241 ) | ( x113 & n1228 ) | ( ~x241 & n1228 ) ;
  assign n1230 = ( x114 & ~x242 ) | ( x114 & n1229 ) | ( ~x242 & n1229 ) ;
  assign n1231 = ( x115 & ~x243 ) | ( x115 & n1230 ) | ( ~x243 & n1230 ) ;
  assign n1232 = n901 | n1231 ;
  assign n1234 = ( n1226 & ~n1233 ) | ( n1226 & n1232 ) | ( ~n1233 & n1232 ) ;
  assign n1235 = ( x116 & ~x244 ) | ( x116 & 1'b0 ) | ( ~x244 & 1'b0 ) ;
  assign n1236 = ( x117 & ~x245 ) | ( x117 & n1235 ) | ( ~x245 & n1235 ) ;
  assign n1237 = ( x118 & ~x246 ) | ( x118 & n1236 ) | ( ~x246 & n1236 ) ;
  assign n1238 = ~n895 & n1237 ;
  assign n1239 = ( n1234 & ~n901 ) | ( n1234 & n1238 ) | ( ~n901 & n1238 ) ;
  assign n1247 = ~n894 & n1239 ;
  assign n1248 = ( n894 & ~n1246 ) | ( n894 & n1247 ) | ( ~n1246 & n1247 ) ;
  assign n1256 = ( n893 & ~n1255 ) | ( n893 & n1248 ) | ( ~n1255 & n1248 ) ;
  assign n1257 = ( x124 & ~x252 ) | ( x124 & 1'b0 ) | ( ~x252 & 1'b0 ) ;
  assign n1258 = ( x125 & ~x253 ) | ( x125 & n1257 ) | ( ~x253 & n1257 ) ;
  assign n1259 = ( x126 & ~x254 ) | ( x126 & n1258 ) | ( ~x254 & n1258 ) ;
  assign n1260 = ( x255 & ~x127 ) | ( x255 & n1259 ) | ( ~x127 & n1259 ) ;
  assign n1261 = n1256 | n1260 ;
  assign n1293 = x247 | n1261 ;
  assign n1294 = ~x119 & n1261 ;
  assign n1295 = ( n1293 & ~n1294 ) | ( n1293 & 1'b0 ) | ( ~n1294 & 1'b0 ) ;
  assign n1296 = ( x503 & ~n885 ) | ( x503 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1297 = x375 &  n885 ;
  assign n1298 = n1296 | n1297 ;
  assign n2349 = n1295 &  n1298 ;
  assign n1299 = ~n1295 & n1298 ;
  assign n1303 = ( x246 & ~n1261 ) | ( x246 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1304 = x118 &  n1261 ;
  assign n1305 = n1303 | n1304 ;
  assign n1300 = ( x502 & ~n885 ) | ( x502 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1301 = x374 &  n885 ;
  assign n1302 = n1300 | n1301 ;
  assign n1308 = ( x245 & ~n1261 ) | ( x245 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1309 = x117 &  n1261 ;
  assign n1310 = n1308 | n1309 ;
  assign n1311 = ( x501 & ~n885 ) | ( x501 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1312 = x373 &  n885 ;
  assign n1313 = n1311 | n1312 ;
  assign n1315 = ( x244 & ~n1261 ) | ( x244 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1316 = x116 &  n1261 ;
  assign n1317 = n1315 | n1316 ;
  assign n1318 = ( x500 & ~n885 ) | ( x500 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1319 = x372 &  n885 ;
  assign n1320 = n1318 | n1319 ;
  assign n2343 = ( n1317 & ~n1320 ) | ( n1317 & 1'b0 ) | ( ~n1320 & 1'b0 ) ;
  assign n2344 = ( n1310 & ~n1313 ) | ( n1310 & n2343 ) | ( ~n1313 & n2343 ) ;
  assign n2345 = ( n1305 & ~n1302 ) | ( n1305 & n2344 ) | ( ~n1302 & n2344 ) ;
  assign n2346 = ~n1299 & n2345 ;
  assign n1306 = n1302 | n1305 ;
  assign n1307 = ( n1299 & ~n1305 ) | ( n1299 & n1306 ) | ( ~n1305 & n1306 ) ;
  assign n1314 = ~n1310 & n1313 ;
  assign n1321 = ~n1317 & n1320 ;
  assign n1322 = n1314 | n1321 ;
  assign n1323 = n1307 | n1322 ;
  assign n1327 = ( x240 & ~n1261 ) | ( x240 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1328 = x112 &  n1261 ;
  assign n1329 = n1327 | n1328 ;
  assign n1324 = ( x496 & ~n885 ) | ( x496 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1325 = x368 &  n885 ;
  assign n1326 = n1324 | n1325 ;
  assign n2336 = n1329 &  n1326 ;
  assign n1392 = ( x231 & ~n1261 ) | ( x231 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1393 = x103 &  n1261 ;
  assign n1394 = n1392 | n1393 ;
  assign n1395 = ( x487 & ~n885 ) | ( x487 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1396 = x359 &  n885 ;
  assign n1397 = n1395 | n1396 ;
  assign n2296 = n1394 &  n1397 ;
  assign n1398 = ~n1394 & n1397 ;
  assign n1402 = ( x230 & ~n1261 ) | ( x230 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1403 = x102 &  n1261 ;
  assign n1404 = n1402 | n1403 ;
  assign n1399 = ( x486 & ~n885 ) | ( x486 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1400 = x358 &  n885 ;
  assign n1401 = n1399 | n1400 ;
  assign n1407 = ( x229 & ~n1261 ) | ( x229 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1408 = x101 &  n1261 ;
  assign n1409 = n1407 | n1408 ;
  assign n1410 = ( x485 & ~n885 ) | ( x485 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1411 = x357 &  n885 ;
  assign n1412 = n1410 | n1411 ;
  assign n1414 = ( x228 & ~n1261 ) | ( x228 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1415 = x100 &  n1261 ;
  assign n1416 = n1414 | n1415 ;
  assign n1417 = ( x484 & ~n885 ) | ( x484 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1418 = x356 &  n885 ;
  assign n1419 = n1417 | n1418 ;
  assign n2290 = ( n1416 & ~n1419 ) | ( n1416 & 1'b0 ) | ( ~n1419 & 1'b0 ) ;
  assign n2291 = ( n1409 & ~n1412 ) | ( n1409 & n2290 ) | ( ~n1412 & n2290 ) ;
  assign n2292 = ( n1404 & ~n1401 ) | ( n1404 & n2291 ) | ( ~n1401 & n2291 ) ;
  assign n2293 = ~n1398 & n2292 ;
  assign n1405 = n1401 | n1404 ;
  assign n1406 = ( n1398 & ~n1404 ) | ( n1398 & n1405 ) | ( ~n1404 & n1405 ) ;
  assign n1413 = ~n1409 & n1412 ;
  assign n1420 = ~n1416 & n1419 ;
  assign n1421 = n1413 | n1420 ;
  assign n1422 = n1406 | n1421 ;
  assign n1426 = ( x224 & ~n1261 ) | ( x224 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1427 = x96 &  n1261 ;
  assign n1428 = n1426 | n1427 ;
  assign n1423 = ( x480 & ~n885 ) | ( x480 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1424 = x352 &  n885 ;
  assign n1425 = n1423 | n1424 ;
  assign n2283 = n1428 &  n1425 ;
  assign n1491 = ( x215 & ~n1261 ) | ( x215 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1492 = x87 &  n1261 ;
  assign n1493 = n1491 | n1492 ;
  assign n1494 = ( x471 & ~n885 ) | ( x471 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1495 = x343 &  n885 ;
  assign n1496 = n1494 | n1495 ;
  assign n2243 = n1493 &  n1496 ;
  assign n1497 = ~n1493 & n1496 ;
  assign n1501 = ( x214 & ~n1261 ) | ( x214 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1502 = x86 &  n1261 ;
  assign n1503 = n1501 | n1502 ;
  assign n1498 = ( x470 & ~n885 ) | ( x470 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1499 = x342 &  n885 ;
  assign n1500 = n1498 | n1499 ;
  assign n1506 = ( x213 & ~n1261 ) | ( x213 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1507 = x85 &  n1261 ;
  assign n1508 = n1506 | n1507 ;
  assign n1509 = ( x469 & ~n885 ) | ( x469 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1510 = x341 &  n885 ;
  assign n1511 = n1509 | n1510 ;
  assign n1513 = ( x212 & ~n1261 ) | ( x212 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1514 = x84 &  n1261 ;
  assign n1515 = n1513 | n1514 ;
  assign n1516 = ( x468 & ~n885 ) | ( x468 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1517 = x340 &  n885 ;
  assign n1518 = n1516 | n1517 ;
  assign n2237 = ( n1515 & ~n1518 ) | ( n1515 & 1'b0 ) | ( ~n1518 & 1'b0 ) ;
  assign n2238 = ( n1508 & ~n1511 ) | ( n1508 & n2237 ) | ( ~n1511 & n2237 ) ;
  assign n2239 = ( n1503 & ~n1500 ) | ( n1503 & n2238 ) | ( ~n1500 & n2238 ) ;
  assign n2240 = ~n1497 & n2239 ;
  assign n1504 = n1500 | n1503 ;
  assign n1505 = ( n1497 & ~n1503 ) | ( n1497 & n1504 ) | ( ~n1503 & n1504 ) ;
  assign n1512 = ~n1508 & n1511 ;
  assign n1519 = ~n1515 & n1518 ;
  assign n1520 = n1512 | n1519 ;
  assign n1521 = n1505 | n1520 ;
  assign n1525 = ( x208 & ~n1261 ) | ( x208 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1526 = x80 &  n1261 ;
  assign n1527 = n1525 | n1526 ;
  assign n1522 = ( x464 & ~n885 ) | ( x464 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1523 = x336 &  n885 ;
  assign n1524 = n1522 | n1523 ;
  assign n2230 = n1527 &  n1524 ;
  assign n1590 = ( x199 & ~n1261 ) | ( x199 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1591 = x71 &  n1261 ;
  assign n1592 = n1590 | n1591 ;
  assign n1593 = ( x455 & ~n885 ) | ( x455 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1594 = x327 &  n885 ;
  assign n1595 = n1593 | n1594 ;
  assign n2190 = n1592 &  n1595 ;
  assign n1688 = ( x175 & ~n1261 ) | ( x175 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1689 = x47 &  n1261 ;
  assign n1690 = n1688 | n1689 ;
  assign n1691 = ( x431 & ~n885 ) | ( x431 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1692 = x303 &  n885 ;
  assign n1693 = n1691 | n1692 ;
  assign n2059 = n1690 &  n1693 ;
  assign n1755 = ( x416 & ~n885 ) | ( x416 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1756 = x288 &  n885 ;
  assign n1757 = n1755 | n1756 ;
  assign n1758 = ( x160 & ~n1261 ) | ( x160 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1759 = x32 &  n1261 ;
  assign n1760 = n1758 | n1759 ;
  assign n1761 = n1757 &  n1760 ;
  assign n1762 = ( x159 & ~n1261 ) | ( x159 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1763 = x31 &  n1261 ;
  assign n1764 = n1762 | n1763 ;
  assign n1765 = ( x415 & ~n885 ) | ( x415 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1766 = x287 &  n885 ;
  assign n1767 = n1765 | n1766 ;
  assign n1768 = ( x158 & ~n1261 ) | ( x158 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1769 = x30 &  n1261 ;
  assign n1770 = n1768 | n1769 ;
  assign n1771 = ( x414 & ~n885 ) | ( x414 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1772 = x286 &  n885 ;
  assign n1773 = n1771 | n1772 ;
  assign n1774 = ( x157 & ~n1261 ) | ( x157 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1775 = x29 &  n1261 ;
  assign n1776 = n1774 | n1775 ;
  assign n1777 = ( x413 & ~n885 ) | ( x413 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1778 = x285 &  n885 ;
  assign n1779 = n1777 | n1778 ;
  assign n1780 = ( x156 & ~n1261 ) | ( x156 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1781 = x28 &  n1261 ;
  assign n1782 = n1780 | n1781 ;
  assign n1783 = ( x412 & ~n885 ) | ( x412 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1784 = x284 &  n885 ;
  assign n1785 = n1783 | n1784 ;
  assign n1786 = ( x155 & ~n1261 ) | ( x155 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1787 = x27 &  n1261 ;
  assign n1788 = n1786 | n1787 ;
  assign n1789 = ( x411 & ~n885 ) | ( x411 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1790 = x283 &  n885 ;
  assign n1791 = n1789 | n1790 ;
  assign n1792 = ( x154 & ~n1261 ) | ( x154 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1793 = x26 &  n1261 ;
  assign n1794 = n1792 | n1793 ;
  assign n1795 = ( x410 & ~n885 ) | ( x410 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1796 = x282 &  n885 ;
  assign n1797 = n1795 | n1796 ;
  assign n1804 = ( x151 & ~n1261 ) | ( x151 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1805 = x23 &  n1261 ;
  assign n1806 = n1804 | n1805 ;
  assign n1807 = ( x407 & ~n885 ) | ( x407 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1808 = x279 &  n885 ;
  assign n1809 = n1807 | n1808 ;
  assign n1810 = ( x150 & ~n1261 ) | ( x150 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1811 = x22 &  n1261 ;
  assign n1812 = n1810 | n1811 ;
  assign n1813 = ( x406 & ~n885 ) | ( x406 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1814 = x278 &  n885 ;
  assign n1815 = n1813 | n1814 ;
  assign n1816 = ( x149 & ~n1261 ) | ( x149 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1817 = x21 &  n1261 ;
  assign n1818 = n1816 | n1817 ;
  assign n1819 = ( x405 & ~n885 ) | ( x405 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1820 = x277 &  n885 ;
  assign n1821 = n1819 | n1820 ;
  assign n1822 = ( x148 & ~n1261 ) | ( x148 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1823 = x20 &  n1261 ;
  assign n1824 = n1822 | n1823 ;
  assign n1825 = ( x404 & ~n885 ) | ( x404 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1826 = x276 &  n885 ;
  assign n1827 = n1825 | n1826 ;
  assign n1828 = ( x147 & ~n1261 ) | ( x147 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1829 = x19 &  n1261 ;
  assign n1830 = n1828 | n1829 ;
  assign n1831 = ( x403 & ~n885 ) | ( x403 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1832 = x275 &  n885 ;
  assign n1833 = n1831 | n1832 ;
  assign n1834 = ( x146 & ~n1261 ) | ( x146 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1835 = x18 &  n1261 ;
  assign n1836 = n1834 | n1835 ;
  assign n1837 = ( x402 & ~n885 ) | ( x402 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1838 = x274 &  n885 ;
  assign n1839 = n1837 | n1838 ;
  assign n1846 = ( x143 & ~n1261 ) | ( x143 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1847 = x15 &  n1261 ;
  assign n1848 = n1846 | n1847 ;
  assign n1849 = ( x399 & ~n885 ) | ( x399 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1850 = x271 &  n885 ;
  assign n1851 = n1849 | n1850 ;
  assign n1852 = ( x142 & ~n1261 ) | ( x142 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1853 = x14 &  n1261 ;
  assign n1854 = n1852 | n1853 ;
  assign n1855 = ( x398 & ~n885 ) | ( x398 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1856 = x270 &  n885 ;
  assign n1857 = n1855 | n1856 ;
  assign n1858 = ( x141 & ~n1261 ) | ( x141 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1859 = x13 &  n1261 ;
  assign n1860 = n1858 | n1859 ;
  assign n1861 = ( x397 & ~n885 ) | ( x397 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1862 = x269 &  n885 ;
  assign n1863 = n1861 | n1862 ;
  assign n1864 = ( x140 & ~n1261 ) | ( x140 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1865 = x12 &  n1261 ;
  assign n1866 = n1864 | n1865 ;
  assign n1867 = ( x396 & ~n885 ) | ( x396 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1868 = x268 &  n885 ;
  assign n1869 = n1867 | n1868 ;
  assign n1870 = ( x139 & ~n1261 ) | ( x139 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1871 = x11 &  n1261 ;
  assign n1872 = n1870 | n1871 ;
  assign n1873 = ( x395 & ~n885 ) | ( x395 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1874 = x267 &  n885 ;
  assign n1875 = n1873 | n1874 ;
  assign n1876 = ( x138 & ~n1261 ) | ( x138 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1877 = x10 &  n1261 ;
  assign n1878 = n1876 | n1877 ;
  assign n1879 = ( x394 & ~n885 ) | ( x394 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1880 = x266 &  n885 ;
  assign n1881 = n1879 | n1880 ;
  assign n1888 = ( x135 & ~n1261 ) | ( x135 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1889 = x7 &  n1261 ;
  assign n1890 = n1888 | n1889 ;
  assign n1891 = ( x391 & ~n885 ) | ( x391 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1892 = x263 &  n885 ;
  assign n1893 = n1891 | n1892 ;
  assign n1897 = ( x134 & ~n1261 ) | ( x134 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1898 = x6 &  n1261 ;
  assign n1899 = n1897 | n1898 ;
  assign n1894 = ( x390 & ~n885 ) | ( x390 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1895 = x262 &  n885 ;
  assign n1896 = n1894 | n1895 ;
  assign n1903 = ( x133 & ~n1261 ) | ( x133 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1904 = x5 &  n1261 ;
  assign n1905 = n1903 | n1904 ;
  assign n1900 = ( x389 & ~n885 ) | ( x389 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1901 = x261 &  n885 ;
  assign n1902 = n1900 | n1901 ;
  assign n1909 = ( x132 & ~n1261 ) | ( x132 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1910 = x4 &  n1261 ;
  assign n1911 = n1909 | n1910 ;
  assign n1906 = ( x388 & ~n885 ) | ( x388 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1907 = x260 &  n885 ;
  assign n1908 = n1906 | n1907 ;
  assign n1912 = ( x131 & ~n1261 ) | ( x131 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1913 = x3 &  n1261 ;
  assign n1914 = n1912 | n1913 ;
  assign n1915 = ( x387 & ~n885 ) | ( x387 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1916 = x259 &  n885 ;
  assign n1917 = n1915 | n1916 ;
  assign n1918 = ( x130 & ~n1261 ) | ( x130 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1919 = x2 &  n1261 ;
  assign n1920 = n1918 | n1919 ;
  assign n1921 = ( x386 & ~n885 ) | ( x386 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1922 = x258 &  n885 ;
  assign n1923 = n1921 | n1922 ;
  assign n1927 = ( x128 & ~n1261 ) | ( x128 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1928 = x0 &  n1261 ;
  assign n1929 = n1927 | n1928 ;
  assign n1930 = ~n888 & n1929 ;
  assign n1924 = ( x385 & ~n885 ) | ( x385 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1925 = x257 &  n885 ;
  assign n1926 = n1924 | n1925 ;
  assign n1931 = ( x129 & ~n1261 ) | ( x129 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1932 = x1 &  n1261 ;
  assign n1933 = n1931 | n1932 ;
  assign n1934 = ( n1930 & ~n1926 ) | ( n1930 & n1933 ) | ( ~n1926 & n1933 ) ;
  assign n1935 = ( n1920 & ~n1923 ) | ( n1920 & n1934 ) | ( ~n1923 & n1934 ) ;
  assign n1936 = ( n1914 & ~n1917 ) | ( n1914 & n1935 ) | ( ~n1917 & n1935 ) ;
  assign n1937 = ( n1911 & ~n1908 ) | ( n1911 & n1936 ) | ( ~n1908 & n1936 ) ;
  assign n1938 = ( n1905 & ~n1902 ) | ( n1905 & n1937 ) | ( ~n1902 & n1937 ) ;
  assign n1939 = ( n1899 & ~n1896 ) | ( n1899 & n1938 ) | ( ~n1896 & n1938 ) ;
  assign n1940 = ( n1890 & ~n1893 ) | ( n1890 & n1939 ) | ( ~n1893 & n1939 ) ;
  assign n1885 = ( x392 & ~n885 ) | ( x392 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1886 = x264 &  n885 ;
  assign n1887 = n1885 | n1886 ;
  assign n1941 = ( x136 & ~n1261 ) | ( x136 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1942 = x8 &  n1261 ;
  assign n1943 = n1941 | n1942 ;
  assign n1944 = ( n1940 & ~n1887 ) | ( n1940 & n1943 ) | ( ~n1887 & n1943 ) ;
  assign n1882 = ( x393 & ~n885 ) | ( x393 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1883 = x265 &  n885 ;
  assign n1884 = n1882 | n1883 ;
  assign n1945 = ( x137 & ~n1261 ) | ( x137 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1946 = x9 &  n1261 ;
  assign n1947 = n1945 | n1946 ;
  assign n1948 = ( n1944 & ~n1884 ) | ( n1944 & n1947 ) | ( ~n1884 & n1947 ) ;
  assign n1949 = ( n1878 & ~n1881 ) | ( n1878 & n1948 ) | ( ~n1881 & n1948 ) ;
  assign n1950 = ( n1872 & ~n1875 ) | ( n1872 & n1949 ) | ( ~n1875 & n1949 ) ;
  assign n1951 = ( n1866 & ~n1869 ) | ( n1866 & n1950 ) | ( ~n1869 & n1950 ) ;
  assign n1952 = ( n1860 & ~n1863 ) | ( n1860 & n1951 ) | ( ~n1863 & n1951 ) ;
  assign n1953 = ( n1854 & ~n1857 ) | ( n1854 & n1952 ) | ( ~n1857 & n1952 ) ;
  assign n1954 = ( n1848 & ~n1851 ) | ( n1848 & n1953 ) | ( ~n1851 & n1953 ) ;
  assign n1843 = ( x400 & ~n885 ) | ( x400 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1844 = x272 &  n885 ;
  assign n1845 = n1843 | n1844 ;
  assign n1955 = ( x144 & ~n1261 ) | ( x144 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1956 = x16 &  n1261 ;
  assign n1957 = n1955 | n1956 ;
  assign n1958 = ( n1954 & ~n1845 ) | ( n1954 & n1957 ) | ( ~n1845 & n1957 ) ;
  assign n1840 = ( x401 & ~n885 ) | ( x401 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1841 = x273 &  n885 ;
  assign n1842 = n1840 | n1841 ;
  assign n1959 = ( x145 & ~n1261 ) | ( x145 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1960 = x17 &  n1261 ;
  assign n1961 = n1959 | n1960 ;
  assign n1962 = ( n1958 & ~n1842 ) | ( n1958 & n1961 ) | ( ~n1842 & n1961 ) ;
  assign n1963 = ( n1836 & ~n1839 ) | ( n1836 & n1962 ) | ( ~n1839 & n1962 ) ;
  assign n1964 = ( n1830 & ~n1833 ) | ( n1830 & n1963 ) | ( ~n1833 & n1963 ) ;
  assign n1965 = ( n1824 & ~n1827 ) | ( n1824 & n1964 ) | ( ~n1827 & n1964 ) ;
  assign n1966 = ( n1818 & ~n1821 ) | ( n1818 & n1965 ) | ( ~n1821 & n1965 ) ;
  assign n1967 = ( n1812 & ~n1815 ) | ( n1812 & n1966 ) | ( ~n1815 & n1966 ) ;
  assign n1968 = ( n1806 & ~n1809 ) | ( n1806 & n1967 ) | ( ~n1809 & n1967 ) ;
  assign n1801 = ( x408 & ~n885 ) | ( x408 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1802 = x280 &  n885 ;
  assign n1803 = n1801 | n1802 ;
  assign n1969 = ( x152 & ~n1261 ) | ( x152 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1970 = x24 &  n1261 ;
  assign n1971 = n1969 | n1970 ;
  assign n1972 = ( n1968 & ~n1803 ) | ( n1968 & n1971 ) | ( ~n1803 & n1971 ) ;
  assign n1798 = ( x409 & ~n885 ) | ( x409 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1799 = x281 &  n885 ;
  assign n1800 = n1798 | n1799 ;
  assign n1973 = ( x153 & ~n1261 ) | ( x153 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1974 = x25 &  n1261 ;
  assign n1975 = n1973 | n1974 ;
  assign n1976 = ( n1972 & ~n1800 ) | ( n1972 & n1975 ) | ( ~n1800 & n1975 ) ;
  assign n1977 = ( n1794 & ~n1797 ) | ( n1794 & n1976 ) | ( ~n1797 & n1976 ) ;
  assign n1978 = ( n1788 & ~n1791 ) | ( n1788 & n1977 ) | ( ~n1791 & n1977 ) ;
  assign n1979 = ( n1782 & ~n1785 ) | ( n1782 & n1978 ) | ( ~n1785 & n1978 ) ;
  assign n1980 = ( n1776 & ~n1779 ) | ( n1776 & n1979 ) | ( ~n1779 & n1979 ) ;
  assign n1981 = ( n1770 & ~n1773 ) | ( n1770 & n1980 ) | ( ~n1773 & n1980 ) ;
  assign n1982 = ( n1764 & ~n1767 ) | ( n1764 & n1981 ) | ( ~n1767 & n1981 ) ;
  assign n1986 = ( x417 & ~n885 ) | ( x417 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1987 = x289 &  n885 ;
  assign n1988 = n1986 | n1987 ;
  assign n1983 = ( x161 & ~n1261 ) | ( x161 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1984 = x33 &  n1261 ;
  assign n1985 = n1983 | n1984 ;
  assign n2036 = n1988 | n1985 ;
  assign n1989 = ( x167 & ~n1261 ) | ( x167 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1990 = x39 &  n1261 ;
  assign n1991 = n1989 | n1990 ;
  assign n1992 = ( x423 & ~n885 ) | ( x423 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1993 = x295 &  n885 ;
  assign n1994 = n1992 | n1993 ;
  assign n1995 = ~n1991 & n1994 ;
  assign n1999 = ( x166 & ~n1261 ) | ( x166 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2000 = x38 &  n1261 ;
  assign n2001 = n1999 | n2000 ;
  assign n1996 = ( x422 & ~n885 ) | ( x422 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1997 = x294 &  n885 ;
  assign n1998 = n1996 | n1997 ;
  assign n2002 = n1998 | n2001 ;
  assign n2003 = ( n1995 & ~n2001 ) | ( n1995 & n2002 ) | ( ~n2001 & n2002 ) ;
  assign n2004 = ( x164 & ~n1261 ) | ( x164 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2005 = x36 &  n1261 ;
  assign n2006 = n2004 | n2005 ;
  assign n2007 = ( x420 & ~n885 ) | ( x420 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2008 = x292 &  n885 ;
  assign n2009 = n2007 | n2008 ;
  assign n2010 = ~n2006 & n2009 ;
  assign n2011 = ( x165 & ~n1261 ) | ( x165 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2012 = x37 &  n1261 ;
  assign n2013 = n2011 | n2012 ;
  assign n2014 = ( x421 & ~n885 ) | ( x421 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2015 = x293 &  n885 ;
  assign n2016 = n2014 | n2015 ;
  assign n2017 = ~n2013 & n2016 ;
  assign n2018 = n2010 | n2017 ;
  assign n2019 = n2003 | n2018 ;
  assign n2020 = ( x163 & ~n1261 ) | ( x163 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2021 = x35 &  n1261 ;
  assign n2022 = n2020 | n2021 ;
  assign n2023 = ( x419 & ~n885 ) | ( x419 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2024 = x291 &  n885 ;
  assign n2025 = n2023 | n2024 ;
  assign n2026 = ~n2022 & n2025 ;
  assign n2030 = ( x162 & ~n1261 ) | ( x162 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2031 = x34 &  n1261 ;
  assign n2032 = n2030 | n2031 ;
  assign n2027 = ( x418 & ~n885 ) | ( x418 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2028 = x290 &  n885 ;
  assign n2029 = n2027 | n2028 ;
  assign n2033 = n2029 | n2032 ;
  assign n2034 = ( n2026 & ~n2032 ) | ( n2026 & n2033 ) | ( ~n2032 & n2033 ) ;
  assign n2035 = n2019 | n2034 ;
  assign n2037 = ( n2036 & ~n1985 ) | ( n2036 & n2035 ) | ( ~n1985 & n2035 ) ;
  assign n2038 = ( n1982 & ~n2037 ) | ( n1982 & 1'b0 ) | ( ~n2037 & 1'b0 ) ;
  assign n2039 = ( n1761 & ~n1757 ) | ( n1761 & n2038 ) | ( ~n1757 & n2038 ) ;
  assign n2044 = ( n2006 & ~n2009 ) | ( n2006 & 1'b0 ) | ( ~n2009 & 1'b0 ) ;
  assign n2045 = ( n2013 & ~n2016 ) | ( n2013 & n2044 ) | ( ~n2016 & n2044 ) ;
  assign n2046 = ( n2001 & ~n1998 ) | ( n2001 & n2045 ) | ( ~n1998 & n2045 ) ;
  assign n2047 = ( n1991 & ~n1994 ) | ( n1991 & n2046 ) | ( ~n1994 & n2046 ) ;
  assign n2040 = ~n1757 & n1760 ;
  assign n2041 = ( n1985 & ~n1988 ) | ( n1985 & n2040 ) | ( ~n1988 & n2040 ) ;
  assign n2042 = ( n2032 & ~n2029 ) | ( n2032 & n2041 ) | ( ~n2029 & n2041 ) ;
  assign n2043 = ( n2022 & ~n2025 ) | ( n2022 & n2042 ) | ( ~n2025 & n2042 ) ;
  assign n2048 = n2019 | n2043 ;
  assign n2049 = ( n2047 & ~n2019 ) | ( n2047 & n2048 ) | ( ~n2019 & n2048 ) ;
  assign n2050 = n2039 | n2049 ;
  assign n1694 = ~n1690 & n1693 ;
  assign n1698 = ( x174 & ~n1261 ) | ( x174 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1699 = x46 &  n1261 ;
  assign n1700 = n1698 | n1699 ;
  assign n1695 = ( x430 & ~n885 ) | ( x430 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1696 = x302 &  n885 ;
  assign n1697 = n1695 | n1696 ;
  assign n1701 = n1697 | n1700 ;
  assign n1702 = ( n1694 & ~n1700 ) | ( n1694 & n1701 ) | ( ~n1700 & n1701 ) ;
  assign n1703 = ( x172 & ~n1261 ) | ( x172 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1704 = x44 &  n1261 ;
  assign n1705 = n1703 | n1704 ;
  assign n1706 = ( x428 & ~n885 ) | ( x428 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1707 = x300 &  n885 ;
  assign n1708 = n1706 | n1707 ;
  assign n1709 = ~n1705 & n1708 ;
  assign n1710 = ( x173 & ~n1261 ) | ( x173 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1711 = x45 &  n1261 ;
  assign n1712 = n1710 | n1711 ;
  assign n1713 = ( x429 & ~n885 ) | ( x429 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1714 = x301 &  n885 ;
  assign n1715 = n1713 | n1714 ;
  assign n1716 = ~n1712 & n1715 ;
  assign n1717 = n1709 | n1716 ;
  assign n1718 = n1702 | n1717 ;
  assign n1719 = ( x171 & ~n1261 ) | ( x171 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1720 = x43 &  n1261 ;
  assign n1721 = n1719 | n1720 ;
  assign n1722 = ( x427 & ~n885 ) | ( x427 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1723 = x299 &  n885 ;
  assign n1724 = n1722 | n1723 ;
  assign n1725 = ~n1721 & n1724 ;
  assign n1726 = ( x170 & ~n1261 ) | ( x170 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1727 = x42 &  n1261 ;
  assign n1728 = n1726 | n1727 ;
  assign n1729 = ( x426 & ~n885 ) | ( x426 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1730 = x298 &  n885 ;
  assign n1731 = n1729 | n1730 ;
  assign n1748 = n1728 &  n1731 ;
  assign n1749 = ( n1725 & ~n1748 ) | ( n1725 & n1731 ) | ( ~n1748 & n1731 ) ;
  assign n1732 = ( x169 & ~n1261 ) | ( x169 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1733 = x41 &  n1261 ;
  assign n1734 = n1732 | n1733 ;
  assign n1735 = ( x425 & ~n885 ) | ( x425 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1736 = x297 &  n885 ;
  assign n1737 = n1735 | n1736 ;
  assign n1750 = ~n1734 & n1737 ;
  assign n1738 = ( x168 & ~n1261 ) | ( x168 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1739 = x40 &  n1261 ;
  assign n1740 = n1738 | n1739 ;
  assign n1741 = ( x424 & ~n885 ) | ( x424 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1742 = x296 &  n885 ;
  assign n1743 = n1741 | n1742 ;
  assign n1751 = ~n1740 & n1743 ;
  assign n1752 = n1750 | n1751 ;
  assign n1753 = ( n1749 & ~n1718 ) | ( n1749 & n1752 ) | ( ~n1718 & n1752 ) ;
  assign n1754 = n1718 | n1753 ;
  assign n2055 = n2050 | n1754 ;
  assign n2051 = ( n1705 & ~n1708 ) | ( n1705 & 1'b0 ) | ( ~n1708 & 1'b0 ) ;
  assign n2052 = ( n1712 & ~n1715 ) | ( n1712 & n2051 ) | ( ~n1715 & n2051 ) ;
  assign n2053 = ( n1700 & ~n1697 ) | ( n1700 & n2052 ) | ( ~n1697 & n2052 ) ;
  assign n2054 = ~n1694 & n2053 ;
  assign n2056 = ( n2055 & ~n1754 ) | ( n2055 & n2054 ) | ( ~n1754 & n2054 ) ;
  assign n1744 = ( n1740 & ~n1743 ) | ( n1740 & 1'b0 ) | ( ~n1743 & 1'b0 ) ;
  assign n1745 = ( n1734 & ~n1737 ) | ( n1734 & n1744 ) | ( ~n1737 & n1744 ) ;
  assign n1746 = ( n1728 & ~n1731 ) | ( n1728 & n1745 ) | ( ~n1731 & n1745 ) ;
  assign n1747 = ( n1721 & ~n1724 ) | ( n1721 & n1746 ) | ( ~n1724 & n1746 ) ;
  assign n2057 = n1718 | n1747 ;
  assign n2058 = ( n2056 & ~n1718 ) | ( n2056 & n2057 ) | ( ~n1718 & n2057 ) ;
  assign n2060 = ( n1690 & ~n2059 ) | ( n1690 & n2058 ) | ( ~n2059 & n2058 ) ;
  assign n2061 = ( x432 & ~n885 ) | ( x432 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2062 = x304 &  n885 ;
  assign n2063 = n2061 | n2062 ;
  assign n2064 = ( x176 & ~n1261 ) | ( x176 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2065 = x48 &  n1261 ;
  assign n2066 = n2064 | n2065 ;
  assign n2067 = n2063 &  n2066 ;
  assign n2071 = ( x433 & ~n885 ) | ( x433 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2072 = x305 &  n885 ;
  assign n2073 = n2071 | n2072 ;
  assign n2068 = ( x177 & ~n1261 ) | ( x177 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2069 = x49 &  n1261 ;
  assign n2070 = n2068 | n2069 ;
  assign n2121 = n2073 | n2070 ;
  assign n2074 = ( x183 & ~n1261 ) | ( x183 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2075 = x55 &  n1261 ;
  assign n2076 = n2074 | n2075 ;
  assign n2077 = ( x439 & ~n885 ) | ( x439 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2078 = x311 &  n885 ;
  assign n2079 = n2077 | n2078 ;
  assign n2080 = ~n2076 & n2079 ;
  assign n2084 = ( x182 & ~n1261 ) | ( x182 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2085 = x54 &  n1261 ;
  assign n2086 = n2084 | n2085 ;
  assign n2081 = ( x438 & ~n885 ) | ( x438 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2082 = x310 &  n885 ;
  assign n2083 = n2081 | n2082 ;
  assign n2087 = n2083 | n2086 ;
  assign n2088 = ( n2080 & ~n2086 ) | ( n2080 & n2087 ) | ( ~n2086 & n2087 ) ;
  assign n2089 = ( x181 & ~n1261 ) | ( x181 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2090 = x53 &  n1261 ;
  assign n2091 = n2089 | n2090 ;
  assign n2092 = ( x437 & ~n885 ) | ( x437 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2093 = x309 &  n885 ;
  assign n2094 = n2092 | n2093 ;
  assign n2095 = ~n2091 & n2094 ;
  assign n2096 = ( x436 & ~n885 ) | ( x436 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2097 = x308 &  n885 ;
  assign n2098 = n2096 | n2097 ;
  assign n2099 = ( x180 & ~n1261 ) | ( x180 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2100 = x52 &  n1261 ;
  assign n2101 = n2099 | n2100 ;
  assign n2102 = ( n2098 & ~n2101 ) | ( n2098 & 1'b0 ) | ( ~n2101 & 1'b0 ) ;
  assign n2103 = n2095 | n2102 ;
  assign n2104 = n2088 | n2103 ;
  assign n2105 = ( x179 & ~n1261 ) | ( x179 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2106 = x51 &  n1261 ;
  assign n2107 = n2105 | n2106 ;
  assign n2108 = ( x435 & ~n885 ) | ( x435 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2109 = x307 &  n885 ;
  assign n2110 = n2108 | n2109 ;
  assign n2111 = ~n2107 & n2110 ;
  assign n2115 = ( x178 & ~n1261 ) | ( x178 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2116 = x50 &  n1261 ;
  assign n2117 = n2115 | n2116 ;
  assign n2112 = ( x434 & ~n885 ) | ( x434 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2113 = x306 &  n885 ;
  assign n2114 = n2112 | n2113 ;
  assign n2118 = n2114 | n2117 ;
  assign n2119 = ( n2111 & ~n2117 ) | ( n2111 & n2118 ) | ( ~n2117 & n2118 ) ;
  assign n2120 = n2104 | n2119 ;
  assign n2122 = ( n2121 & ~n2070 ) | ( n2121 & n2120 ) | ( ~n2070 & n2120 ) ;
  assign n2123 = ( n2063 & ~n2067 ) | ( n2063 & n2122 ) | ( ~n2067 & n2122 ) ;
  assign n2135 = n2060 &  n2123 ;
  assign n1652 = ( x187 & ~n1261 ) | ( x187 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1653 = x59 &  n1261 ;
  assign n1654 = n1652 | n1653 ;
  assign n1655 = ( x443 & ~n885 ) | ( x443 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1656 = x315 &  n885 ;
  assign n1657 = n1655 | n1656 ;
  assign n1658 = ~n1654 & n1657 ;
  assign n1659 = ( x186 & ~n1261 ) | ( x186 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1660 = x58 &  n1261 ;
  assign n1661 = n1659 | n1660 ;
  assign n1662 = ( x442 & ~n885 ) | ( x442 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1663 = x314 &  n885 ;
  assign n1664 = n1662 | n1663 ;
  assign n1681 = n1661 &  n1664 ;
  assign n1682 = ( n1658 & ~n1681 ) | ( n1658 & n1664 ) | ( ~n1681 & n1664 ) ;
  assign n1621 = ( x191 & ~n1261 ) | ( x191 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1622 = x63 &  n1261 ;
  assign n1623 = n1621 | n1622 ;
  assign n1624 = ( x447 & ~n885 ) | ( x447 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1625 = x319 &  n885 ;
  assign n1626 = n1624 | n1625 ;
  assign n1627 = ~n1623 & n1626 ;
  assign n1631 = ( x190 & ~n1261 ) | ( x190 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1632 = x62 &  n1261 ;
  assign n1633 = n1631 | n1632 ;
  assign n1628 = ( x446 & ~n885 ) | ( x446 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1629 = x318 &  n885 ;
  assign n1630 = n1628 | n1629 ;
  assign n1634 = n1630 | n1633 ;
  assign n1635 = ( n1627 & ~n1633 ) | ( n1627 & n1634 ) | ( ~n1633 & n1634 ) ;
  assign n1636 = ( x188 & ~n1261 ) | ( x188 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1637 = x60 &  n1261 ;
  assign n1638 = n1636 | n1637 ;
  assign n1639 = ( x444 & ~n885 ) | ( x444 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1640 = x316 &  n885 ;
  assign n1641 = n1639 | n1640 ;
  assign n1642 = ~n1638 & n1641 ;
  assign n1643 = ( x189 & ~n1261 ) | ( x189 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1644 = x61 &  n1261 ;
  assign n1645 = n1643 | n1644 ;
  assign n1646 = ( x445 & ~n885 ) | ( x445 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1647 = x317 &  n885 ;
  assign n1648 = n1646 | n1647 ;
  assign n1649 = ~n1645 & n1648 ;
  assign n1650 = n1642 | n1649 ;
  assign n1651 = n1635 | n1650 ;
  assign n1665 = ( x185 & ~n1261 ) | ( x185 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1666 = x57 &  n1261 ;
  assign n1667 = n1665 | n1666 ;
  assign n1668 = ( x441 & ~n885 ) | ( x441 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1669 = x313 &  n885 ;
  assign n1670 = n1668 | n1669 ;
  assign n1683 = ~n1667 & n1670 ;
  assign n1671 = ( x184 & ~n1261 ) | ( x184 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1672 = x56 &  n1261 ;
  assign n1673 = n1671 | n1672 ;
  assign n1674 = ( x440 & ~n885 ) | ( x440 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1675 = x312 &  n885 ;
  assign n1676 = n1674 | n1675 ;
  assign n1684 = ~n1673 & n1676 ;
  assign n1685 = n1683 | n1684 ;
  assign n1686 = n1651 | n1685 ;
  assign n1687 = n1682 | n1686 ;
  assign n2124 = ~n2063 & n2066 ;
  assign n2125 = ( n2070 & ~n2073 ) | ( n2070 & n2124 ) | ( ~n2073 & n2124 ) ;
  assign n2126 = ( n2117 & ~n2114 ) | ( n2117 & n2125 ) | ( ~n2114 & n2125 ) ;
  assign n2127 = ( n2107 & ~n2110 ) | ( n2107 & n2126 ) | ( ~n2110 & n2126 ) ;
  assign n2132 = n2127 | n2104 ;
  assign n2128 = ~n2098 & n2101 ;
  assign n2129 = ( n2091 & ~n2094 ) | ( n2091 & n2128 ) | ( ~n2094 & n2128 ) ;
  assign n2130 = ( n2086 & ~n2083 ) | ( n2086 & n2129 ) | ( ~n2083 & n2129 ) ;
  assign n2131 = ( n2076 & ~n2079 ) | ( n2076 & n2130 ) | ( ~n2079 & n2130 ) ;
  assign n2133 = ( n2132 & ~n2104 ) | ( n2132 & n2131 ) | ( ~n2104 & n2131 ) ;
  assign n2134 = n1687 | n2133 ;
  assign n2136 = ( n2060 & ~n2135 ) | ( n2060 & n2134 ) | ( ~n2135 & n2134 ) ;
  assign n2137 = ( n1638 & ~n1641 ) | ( n1638 & 1'b0 ) | ( ~n1641 & 1'b0 ) ;
  assign n2138 = ( n1645 & ~n1648 ) | ( n1645 & n2137 ) | ( ~n1648 & n2137 ) ;
  assign n2139 = ( n1633 & ~n1630 ) | ( n1633 & n2138 ) | ( ~n1630 & n2138 ) ;
  assign n2140 = ~n1627 & n2139 ;
  assign n2141 = ( n2136 & ~n1687 ) | ( n2136 & n2140 ) | ( ~n1687 & n2140 ) ;
  assign n1677 = ( n1673 & ~n1676 ) | ( n1673 & 1'b0 ) | ( ~n1676 & 1'b0 ) ;
  assign n1678 = ( n1667 & ~n1670 ) | ( n1667 & n1677 ) | ( ~n1670 & n1677 ) ;
  assign n1679 = ( n1661 & ~n1664 ) | ( n1661 & n1678 ) | ( ~n1664 & n1678 ) ;
  assign n1680 = ( n1654 & ~n1657 ) | ( n1654 & n1679 ) | ( ~n1657 & n1679 ) ;
  assign n2142 = n1651 | n1680 ;
  assign n2143 = ( n2141 & ~n1651 ) | ( n2141 & n2142 ) | ( ~n1651 & n2142 ) ;
  assign n2145 = ( x448 & ~n885 ) | ( x448 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2146 = x320 &  n885 ;
  assign n2147 = n2145 | n2146 ;
  assign n2148 = ( x192 & ~n1261 ) | ( x192 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2149 = x64 &  n1261 ;
  assign n2150 = n2148 | n2149 ;
  assign n2151 = ( n2147 & ~n2150 ) | ( n2147 & 1'b0 ) | ( ~n2150 & 1'b0 ) ;
  assign n2152 = ( x193 & ~n1261 ) | ( x193 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2153 = x65 &  n1261 ;
  assign n2154 = n2152 | n2153 ;
  assign n2155 = ( x449 & ~n885 ) | ( x449 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2156 = x321 &  n885 ;
  assign n2157 = n2155 | n2156 ;
  assign n2158 = ~n2154 & n2157 ;
  assign n2159 = n2151 | n2158 ;
  assign n2144 = ( n1623 & ~n1626 ) | ( n1623 & 1'b0 ) | ( ~n1626 & 1'b0 ) ;
  assign n2160 = ~n2143 & n2144 ;
  assign n2161 = ( n2143 & ~n2159 ) | ( n2143 & n2160 ) | ( ~n2159 & n2160 ) ;
  assign n2162 = ( x195 & ~n1261 ) | ( x195 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2163 = x67 &  n1261 ;
  assign n2164 = n2162 | n2163 ;
  assign n2165 = ( x451 & ~n885 ) | ( x451 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2166 = x323 &  n885 ;
  assign n2167 = n2165 | n2166 ;
  assign n2168 = ~n2164 & n2167 ;
  assign n2172 = ( x194 & ~n1261 ) | ( x194 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2173 = x66 &  n1261 ;
  assign n2174 = n2172 | n2173 ;
  assign n2169 = ( x450 & ~n885 ) | ( x450 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2170 = x322 &  n885 ;
  assign n2171 = n2169 | n2170 ;
  assign n2175 = n2171 | n2174 ;
  assign n2176 = ( n2168 & ~n2174 ) | ( n2168 & n2175 ) | ( ~n2174 & n2175 ) ;
  assign n2181 = ~n2159 & n2176 ;
  assign n2182 = ( n2143 & n2160 ) | ( n2143 & n2181 ) | ( n2160 & n2181 ) ;
  assign n1596 = ~n1592 & n1595 ;
  assign n1600 = ( x198 & ~n1261 ) | ( x198 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1601 = x70 &  n1261 ;
  assign n1602 = n1600 | n1601 ;
  assign n1597 = ( x454 & ~n885 ) | ( x454 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1598 = x326 &  n885 ;
  assign n1599 = n1597 | n1598 ;
  assign n1603 = n1599 | n1602 ;
  assign n1604 = ( n1596 & ~n1602 ) | ( n1596 & n1603 ) | ( ~n1602 & n1603 ) ;
  assign n1605 = ( x197 & ~n1261 ) | ( x197 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1606 = x69 &  n1261 ;
  assign n1607 = n1605 | n1606 ;
  assign n1608 = ( x453 & ~n885 ) | ( x453 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1609 = x325 &  n885 ;
  assign n1610 = n1608 | n1609 ;
  assign n1611 = ~n1607 & n1610 ;
  assign n1612 = ( x196 & ~n1261 ) | ( x196 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1613 = x68 &  n1261 ;
  assign n1614 = n1612 | n1613 ;
  assign n1615 = ( x452 & ~n885 ) | ( x452 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1616 = x324 &  n885 ;
  assign n1617 = n1615 | n1616 ;
  assign n1618 = ~n1614 & n1617 ;
  assign n1619 = n1611 | n1618 ;
  assign n1620 = n1604 | n1619 ;
  assign n2177 = ~n2147 & n2150 ;
  assign n2178 = ( n2154 & ~n2157 ) | ( n2154 & n2177 ) | ( ~n2157 & n2177 ) ;
  assign n2179 = ( n2174 & ~n2171 ) | ( n2174 & n2178 ) | ( ~n2171 & n2178 ) ;
  assign n2180 = ( n2164 & ~n2167 ) | ( n2164 & n2179 ) | ( ~n2167 & n2179 ) ;
  assign n2183 = n1620 | n2180 ;
  assign n2184 = ( n2161 & ~n2182 ) | ( n2161 & n2183 ) | ( ~n2182 & n2183 ) ;
  assign n2185 = ( n1614 & ~n1617 ) | ( n1614 & 1'b0 ) | ( ~n1617 & 1'b0 ) ;
  assign n2186 = ( n1607 & ~n1610 ) | ( n1607 & n2185 ) | ( ~n1610 & n2185 ) ;
  assign n2187 = ( n1602 & ~n1599 ) | ( n1602 & n2186 ) | ( ~n1599 & n2186 ) ;
  assign n2188 = ~n1596 & n2187 ;
  assign n2189 = ( n2184 & ~n1620 ) | ( n2184 & n2188 ) | ( ~n1620 & n2188 ) ;
  assign n2191 = ( n1592 & ~n2190 ) | ( n1592 & n2189 ) | ( ~n2190 & n2189 ) ;
  assign n1559 = ( x203 & ~n1261 ) | ( x203 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1560 = x75 &  n1261 ;
  assign n1561 = n1559 | n1560 ;
  assign n1562 = ( x459 & ~n885 ) | ( x459 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1563 = x331 &  n885 ;
  assign n1564 = n1562 | n1563 ;
  assign n1565 = ~n1561 & n1564 ;
  assign n1569 = ( x202 & ~n1261 ) | ( x202 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1570 = x74 &  n1261 ;
  assign n1571 = n1569 | n1570 ;
  assign n1566 = ( x458 & ~n885 ) | ( x458 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1567 = x330 &  n885 ;
  assign n1568 = n1566 | n1567 ;
  assign n1572 = n1568 | n1571 ;
  assign n1573 = ( n1565 & ~n1571 ) | ( n1565 & n1572 ) | ( ~n1571 & n1572 ) ;
  assign n1574 = ( x201 & ~n1261 ) | ( x201 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1575 = x73 &  n1261 ;
  assign n1576 = n1574 | n1575 ;
  assign n1577 = ( x457 & ~n885 ) | ( x457 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1578 = x329 &  n885 ;
  assign n1579 = n1577 | n1578 ;
  assign n1580 = ~n1576 & n1579 ;
  assign n1581 = ( x456 & ~n885 ) | ( x456 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1582 = x328 &  n885 ;
  assign n1583 = n1581 | n1582 ;
  assign n1584 = ( x200 & ~n1261 ) | ( x200 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1585 = x72 &  n1261 ;
  assign n1586 = n1584 | n1585 ;
  assign n1587 = ( n1583 & ~n1586 ) | ( n1583 & 1'b0 ) | ( ~n1586 & 1'b0 ) ;
  assign n1588 = n1580 | n1587 ;
  assign n1589 = n1573 | n1588 ;
  assign n2197 = n2191 | n1589 ;
  assign n1528 = ( x207 & ~n1261 ) | ( x207 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1529 = x79 &  n1261 ;
  assign n1530 = n1528 | n1529 ;
  assign n1531 = ( x463 & ~n885 ) | ( x463 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1532 = x335 &  n885 ;
  assign n1533 = n1531 | n1532 ;
  assign n1534 = ~n1530 & n1533 ;
  assign n1538 = ( x206 & ~n1261 ) | ( x206 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1539 = x78 &  n1261 ;
  assign n1540 = n1538 | n1539 ;
  assign n1535 = ( x462 & ~n885 ) | ( x462 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1536 = x334 &  n885 ;
  assign n1537 = n1535 | n1536 ;
  assign n1541 = n1537 | n1540 ;
  assign n1542 = ( n1534 & ~n1540 ) | ( n1534 & n1541 ) | ( ~n1540 & n1541 ) ;
  assign n1543 = ( x205 & ~n1261 ) | ( x205 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1544 = x77 &  n1261 ;
  assign n1545 = n1543 | n1544 ;
  assign n1546 = ( x461 & ~n885 ) | ( x461 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1547 = x333 &  n885 ;
  assign n1548 = n1546 | n1547 ;
  assign n1549 = ~n1545 & n1548 ;
  assign n1550 = ( x204 & ~n1261 ) | ( x204 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1551 = x76 &  n1261 ;
  assign n1552 = n1550 | n1551 ;
  assign n1553 = ( x460 & ~n885 ) | ( x460 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1554 = x332 &  n885 ;
  assign n1555 = n1553 | n1554 ;
  assign n1556 = ~n1552 & n1555 ;
  assign n1557 = n1549 | n1556 ;
  assign n1558 = n1542 | n1557 ;
  assign n2192 = ~n1583 & n1586 ;
  assign n2193 = ( n1576 & ~n1579 ) | ( n1576 & n2192 ) | ( ~n1579 & n2192 ) ;
  assign n2194 = ( n1571 & ~n1568 ) | ( n1571 & n2193 ) | ( ~n1568 & n2193 ) ;
  assign n2195 = ( n1561 & ~n1564 ) | ( n1561 & n2194 ) | ( ~n1564 & n2194 ) ;
  assign n2196 = n1558 | n2195 ;
  assign n2198 = ( n2197 & ~n1589 ) | ( n2197 & n2196 ) | ( ~n1589 & n2196 ) ;
  assign n2199 = ( n1552 & ~n1555 ) | ( n1552 & 1'b0 ) | ( ~n1555 & 1'b0 ) ;
  assign n2200 = ( n1545 & ~n1548 ) | ( n1545 & n2199 ) | ( ~n1548 & n2199 ) ;
  assign n2201 = ( n1540 & ~n1537 ) | ( n1540 & n2200 ) | ( ~n1537 & n2200 ) ;
  assign n2202 = ~n1534 & n2201 ;
  assign n2203 = ( n2198 & ~n1558 ) | ( n2198 & n2202 ) | ( ~n1558 & n2202 ) ;
  assign n2205 = ( x211 & ~n1261 ) | ( x211 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2206 = x83 &  n1261 ;
  assign n2207 = n2205 | n2206 ;
  assign n2208 = ( x467 & ~n885 ) | ( x467 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2209 = x339 &  n885 ;
  assign n2210 = n2208 | n2209 ;
  assign n2211 = ~n2207 & n2210 ;
  assign n2215 = ( x210 & ~n1261 ) | ( x210 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2216 = x82 &  n1261 ;
  assign n2217 = n2215 | n2216 ;
  assign n2212 = ( x466 & ~n885 ) | ( x466 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2213 = x338 &  n885 ;
  assign n2214 = n2212 | n2213 ;
  assign n2218 = n2214 | n2217 ;
  assign n2219 = ( n2211 & ~n2217 ) | ( n2211 & n2218 ) | ( ~n2217 & n2218 ) ;
  assign n2220 = ( x209 & ~n1261 ) | ( x209 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2221 = x81 &  n1261 ;
  assign n2222 = n2220 | n2221 ;
  assign n2223 = ( x465 & ~n885 ) | ( x465 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2224 = x337 &  n885 ;
  assign n2225 = n2223 | n2224 ;
  assign n2226 = ~n2222 & n2225 ;
  assign n2227 = n2219 | n2226 ;
  assign n2204 = ( n1530 & ~n1533 ) | ( n1530 & 1'b0 ) | ( ~n1533 & 1'b0 ) ;
  assign n2228 = ~n2203 & n2204 ;
  assign n2229 = ( n2203 & ~n2227 ) | ( n2203 & n2228 ) | ( ~n2227 & n2228 ) ;
  assign n2231 = ( n2230 & ~n1524 ) | ( n2230 & n2229 ) | ( ~n1524 & n2229 ) ;
  assign n2232 = ~n1524 & n1527 ;
  assign n2233 = ( n2222 & ~n2225 ) | ( n2222 & n2232 ) | ( ~n2225 & n2232 ) ;
  assign n2234 = ( n2217 & ~n2214 ) | ( n2217 & n2233 ) | ( ~n2214 & n2233 ) ;
  assign n2235 = ( n2207 & ~n2210 ) | ( n2207 & n2234 ) | ( ~n2210 & n2234 ) ;
  assign n2236 = n2231 | n2235 ;
  assign n2241 = n1521 | n2236 ;
  assign n2242 = ( n2240 & ~n1521 ) | ( n2240 & n2241 ) | ( ~n1521 & n2241 ) ;
  assign n2244 = ( n1493 & ~n2243 ) | ( n1493 & n2242 ) | ( ~n2243 & n2242 ) ;
  assign n1460 = ( x219 & ~n1261 ) | ( x219 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1461 = x91 &  n1261 ;
  assign n1462 = n1460 | n1461 ;
  assign n1463 = ( x475 & ~n885 ) | ( x475 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1464 = x347 &  n885 ;
  assign n1465 = n1463 | n1464 ;
  assign n1466 = ~n1462 & n1465 ;
  assign n1470 = ( x218 & ~n1261 ) | ( x218 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1471 = x90 &  n1261 ;
  assign n1472 = n1470 | n1471 ;
  assign n1467 = ( x474 & ~n885 ) | ( x474 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1468 = x346 &  n885 ;
  assign n1469 = n1467 | n1468 ;
  assign n1473 = n1469 | n1472 ;
  assign n1474 = ( n1466 & ~n1472 ) | ( n1466 & n1473 ) | ( ~n1472 & n1473 ) ;
  assign n1475 = ( x217 & ~n1261 ) | ( x217 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1476 = x89 &  n1261 ;
  assign n1477 = n1475 | n1476 ;
  assign n1478 = ( x473 & ~n885 ) | ( x473 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1479 = x345 &  n885 ;
  assign n1480 = n1478 | n1479 ;
  assign n1481 = ~n1477 & n1480 ;
  assign n1482 = ( x472 & ~n885 ) | ( x472 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1483 = x344 &  n885 ;
  assign n1484 = n1482 | n1483 ;
  assign n1485 = ( x216 & ~n1261 ) | ( x216 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1486 = x88 &  n1261 ;
  assign n1487 = n1485 | n1486 ;
  assign n1488 = ( n1484 & ~n1487 ) | ( n1484 & 1'b0 ) | ( ~n1487 & 1'b0 ) ;
  assign n1489 = n1481 | n1488 ;
  assign n1490 = n1474 | n1489 ;
  assign n2250 = n2244 | n1490 ;
  assign n1429 = ( x223 & ~n1261 ) | ( x223 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1430 = x95 &  n1261 ;
  assign n1431 = n1429 | n1430 ;
  assign n1432 = ( x479 & ~n885 ) | ( x479 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1433 = x351 &  n885 ;
  assign n1434 = n1432 | n1433 ;
  assign n1435 = ~n1431 & n1434 ;
  assign n1439 = ( x222 & ~n1261 ) | ( x222 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1440 = x94 &  n1261 ;
  assign n1441 = n1439 | n1440 ;
  assign n1436 = ( x478 & ~n885 ) | ( x478 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1437 = x350 &  n885 ;
  assign n1438 = n1436 | n1437 ;
  assign n1442 = n1438 | n1441 ;
  assign n1443 = ( n1435 & ~n1441 ) | ( n1435 & n1442 ) | ( ~n1441 & n1442 ) ;
  assign n1444 = ( x221 & ~n1261 ) | ( x221 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1445 = x93 &  n1261 ;
  assign n1446 = n1444 | n1445 ;
  assign n1447 = ( x477 & ~n885 ) | ( x477 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1448 = x349 &  n885 ;
  assign n1449 = n1447 | n1448 ;
  assign n1450 = ~n1446 & n1449 ;
  assign n1451 = ( x220 & ~n1261 ) | ( x220 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1452 = x92 &  n1261 ;
  assign n1453 = n1451 | n1452 ;
  assign n1454 = ( x476 & ~n885 ) | ( x476 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1455 = x348 &  n885 ;
  assign n1456 = n1454 | n1455 ;
  assign n1457 = ~n1453 & n1456 ;
  assign n1458 = n1450 | n1457 ;
  assign n1459 = n1443 | n1458 ;
  assign n2245 = ~n1484 & n1487 ;
  assign n2246 = ( n1477 & ~n1480 ) | ( n1477 & n2245 ) | ( ~n1480 & n2245 ) ;
  assign n2247 = ( n1472 & ~n1469 ) | ( n1472 & n2246 ) | ( ~n1469 & n2246 ) ;
  assign n2248 = ( n1462 & ~n1465 ) | ( n1462 & n2247 ) | ( ~n1465 & n2247 ) ;
  assign n2249 = n1459 | n2248 ;
  assign n2251 = ( n2250 & ~n1490 ) | ( n2250 & n2249 ) | ( ~n1490 & n2249 ) ;
  assign n2252 = ( n1453 & ~n1456 ) | ( n1453 & 1'b0 ) | ( ~n1456 & 1'b0 ) ;
  assign n2253 = ( n1446 & ~n1449 ) | ( n1446 & n2252 ) | ( ~n1449 & n2252 ) ;
  assign n2254 = ( n1441 & ~n1438 ) | ( n1441 & n2253 ) | ( ~n1438 & n2253 ) ;
  assign n2255 = ~n1435 & n2254 ;
  assign n2256 = ( n2251 & ~n1459 ) | ( n2251 & n2255 ) | ( ~n1459 & n2255 ) ;
  assign n2258 = ( x227 & ~n1261 ) | ( x227 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2259 = x99 &  n1261 ;
  assign n2260 = n2258 | n2259 ;
  assign n2261 = ( x483 & ~n885 ) | ( x483 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2262 = x355 &  n885 ;
  assign n2263 = n2261 | n2262 ;
  assign n2264 = ~n2260 & n2263 ;
  assign n2268 = ( x226 & ~n1261 ) | ( x226 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2269 = x98 &  n1261 ;
  assign n2270 = n2268 | n2269 ;
  assign n2265 = ( x482 & ~n885 ) | ( x482 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2266 = x354 &  n885 ;
  assign n2267 = n2265 | n2266 ;
  assign n2271 = n2267 | n2270 ;
  assign n2272 = ( n2264 & ~n2270 ) | ( n2264 & n2271 ) | ( ~n2270 & n2271 ) ;
  assign n2273 = ( x225 & ~n1261 ) | ( x225 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2274 = x97 &  n1261 ;
  assign n2275 = n2273 | n2274 ;
  assign n2276 = ( x481 & ~n885 ) | ( x481 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2277 = x353 &  n885 ;
  assign n2278 = n2276 | n2277 ;
  assign n2279 = ~n2275 & n2278 ;
  assign n2280 = n2272 | n2279 ;
  assign n2257 = ( n1431 & ~n1434 ) | ( n1431 & 1'b0 ) | ( ~n1434 & 1'b0 ) ;
  assign n2281 = ~n2256 & n2257 ;
  assign n2282 = ( n2256 & ~n2280 ) | ( n2256 & n2281 ) | ( ~n2280 & n2281 ) ;
  assign n2284 = ( n2283 & ~n1425 ) | ( n2283 & n2282 ) | ( ~n1425 & n2282 ) ;
  assign n2285 = ~n1425 & n1428 ;
  assign n2286 = ( n2275 & ~n2278 ) | ( n2275 & n2285 ) | ( ~n2278 & n2285 ) ;
  assign n2287 = ( n2270 & ~n2267 ) | ( n2270 & n2286 ) | ( ~n2267 & n2286 ) ;
  assign n2288 = ( n2260 & ~n2263 ) | ( n2260 & n2287 ) | ( ~n2263 & n2287 ) ;
  assign n2289 = n2284 | n2288 ;
  assign n2294 = n1422 | n2289 ;
  assign n2295 = ( n2293 & ~n1422 ) | ( n2293 & n2294 ) | ( ~n1422 & n2294 ) ;
  assign n2297 = ( n1394 & ~n2296 ) | ( n1394 & n2295 ) | ( ~n2296 & n2295 ) ;
  assign n1361 = ( x235 & ~n1261 ) | ( x235 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1362 = x107 &  n1261 ;
  assign n1363 = n1361 | n1362 ;
  assign n1364 = ( x491 & ~n885 ) | ( x491 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1365 = x363 &  n885 ;
  assign n1366 = n1364 | n1365 ;
  assign n1367 = ~n1363 & n1366 ;
  assign n1371 = ( x234 & ~n1261 ) | ( x234 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1372 = x106 &  n1261 ;
  assign n1373 = n1371 | n1372 ;
  assign n1368 = ( x490 & ~n885 ) | ( x490 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1369 = x362 &  n885 ;
  assign n1370 = n1368 | n1369 ;
  assign n1374 = n1370 | n1373 ;
  assign n1375 = ( n1367 & ~n1373 ) | ( n1367 & n1374 ) | ( ~n1373 & n1374 ) ;
  assign n1376 = ( x233 & ~n1261 ) | ( x233 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1377 = x105 &  n1261 ;
  assign n1378 = n1376 | n1377 ;
  assign n1379 = ( x489 & ~n885 ) | ( x489 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1380 = x361 &  n885 ;
  assign n1381 = n1379 | n1380 ;
  assign n1382 = ~n1378 & n1381 ;
  assign n1383 = ( x488 & ~n885 ) | ( x488 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1384 = x360 &  n885 ;
  assign n1385 = n1383 | n1384 ;
  assign n1386 = ( x232 & ~n1261 ) | ( x232 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1387 = x104 &  n1261 ;
  assign n1388 = n1386 | n1387 ;
  assign n1389 = ( n1385 & ~n1388 ) | ( n1385 & 1'b0 ) | ( ~n1388 & 1'b0 ) ;
  assign n1390 = n1382 | n1389 ;
  assign n1391 = n1375 | n1390 ;
  assign n2303 = n2297 | n1391 ;
  assign n1330 = ( x239 & ~n1261 ) | ( x239 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1331 = x111 &  n1261 ;
  assign n1332 = n1330 | n1331 ;
  assign n1333 = ( x495 & ~n885 ) | ( x495 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1334 = x367 &  n885 ;
  assign n1335 = n1333 | n1334 ;
  assign n1336 = ~n1332 & n1335 ;
  assign n1340 = ( x238 & ~n1261 ) | ( x238 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1341 = x110 &  n1261 ;
  assign n1342 = n1340 | n1341 ;
  assign n1337 = ( x494 & ~n885 ) | ( x494 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1338 = x366 &  n885 ;
  assign n1339 = n1337 | n1338 ;
  assign n1343 = n1339 | n1342 ;
  assign n1344 = ( n1336 & ~n1342 ) | ( n1336 & n1343 ) | ( ~n1342 & n1343 ) ;
  assign n1345 = ( x237 & ~n1261 ) | ( x237 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1346 = x109 &  n1261 ;
  assign n1347 = n1345 | n1346 ;
  assign n1348 = ( x493 & ~n885 ) | ( x493 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1349 = x365 &  n885 ;
  assign n1350 = n1348 | n1349 ;
  assign n1351 = ~n1347 & n1350 ;
  assign n1352 = ( x236 & ~n1261 ) | ( x236 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1353 = x108 &  n1261 ;
  assign n1354 = n1352 | n1353 ;
  assign n1355 = ( x492 & ~n885 ) | ( x492 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1356 = x364 &  n885 ;
  assign n1357 = n1355 | n1356 ;
  assign n1358 = ~n1354 & n1357 ;
  assign n1359 = n1351 | n1358 ;
  assign n1360 = n1344 | n1359 ;
  assign n2298 = ~n1385 & n1388 ;
  assign n2299 = ( n1378 & ~n1381 ) | ( n1378 & n2298 ) | ( ~n1381 & n2298 ) ;
  assign n2300 = ( n1373 & ~n1370 ) | ( n1373 & n2299 ) | ( ~n1370 & n2299 ) ;
  assign n2301 = ( n1363 & ~n1366 ) | ( n1363 & n2300 ) | ( ~n1366 & n2300 ) ;
  assign n2302 = n1360 | n2301 ;
  assign n2304 = ( n2303 & ~n1391 ) | ( n2303 & n2302 ) | ( ~n1391 & n2302 ) ;
  assign n2305 = ( n1354 & ~n1357 ) | ( n1354 & 1'b0 ) | ( ~n1357 & 1'b0 ) ;
  assign n2306 = ( n1347 & ~n1350 ) | ( n1347 & n2305 ) | ( ~n1350 & n2305 ) ;
  assign n2307 = ( n1342 & ~n1339 ) | ( n1342 & n2306 ) | ( ~n1339 & n2306 ) ;
  assign n2308 = ~n1336 & n2307 ;
  assign n2309 = ( n2304 & ~n1360 ) | ( n2304 & n2308 ) | ( ~n1360 & n2308 ) ;
  assign n2311 = ( x243 & ~n1261 ) | ( x243 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2312 = x115 &  n1261 ;
  assign n2313 = n2311 | n2312 ;
  assign n2314 = ( x499 & ~n885 ) | ( x499 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2315 = x371 &  n885 ;
  assign n2316 = n2314 | n2315 ;
  assign n2317 = ~n2313 & n2316 ;
  assign n2321 = ( x242 & ~n1261 ) | ( x242 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2322 = x114 &  n1261 ;
  assign n2323 = n2321 | n2322 ;
  assign n2318 = ( x498 & ~n885 ) | ( x498 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2319 = x370 &  n885 ;
  assign n2320 = n2318 | n2319 ;
  assign n2324 = n2320 | n2323 ;
  assign n2325 = ( n2317 & ~n2323 ) | ( n2317 & n2324 ) | ( ~n2323 & n2324 ) ;
  assign n2326 = ( x241 & ~n1261 ) | ( x241 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2327 = x113 &  n1261 ;
  assign n2328 = n2326 | n2327 ;
  assign n2329 = ( x497 & ~n885 ) | ( x497 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2330 = x369 &  n885 ;
  assign n2331 = n2329 | n2330 ;
  assign n2332 = ~n2328 & n2331 ;
  assign n2333 = n2325 | n2332 ;
  assign n2310 = ( n1332 & ~n1335 ) | ( n1332 & 1'b0 ) | ( ~n1335 & 1'b0 ) ;
  assign n2334 = ~n2309 & n2310 ;
  assign n2335 = ( n2309 & ~n2333 ) | ( n2309 & n2334 ) | ( ~n2333 & n2334 ) ;
  assign n2337 = ( n2336 & ~n1326 ) | ( n2336 & n2335 ) | ( ~n1326 & n2335 ) ;
  assign n2338 = ~n1326 & n1329 ;
  assign n2339 = ( n2328 & ~n2331 ) | ( n2328 & n2338 ) | ( ~n2331 & n2338 ) ;
  assign n2340 = ( n2323 & ~n2320 ) | ( n2323 & n2339 ) | ( ~n2320 & n2339 ) ;
  assign n2341 = ( n2313 & ~n2316 ) | ( n2313 & n2340 ) | ( ~n2316 & n2340 ) ;
  assign n2342 = n2337 | n2341 ;
  assign n2347 = n1323 | n2342 ;
  assign n2348 = ( n2346 & ~n1323 ) | ( n2346 & n2347 ) | ( ~n1323 & n2347 ) ;
  assign n2350 = ( n1295 & ~n2349 ) | ( n1295 & n2348 ) | ( ~n2349 & n2348 ) ;
  assign n1262 = ( x251 & ~n1261 ) | ( x251 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1263 = x123 &  n1261 ;
  assign n1264 = n1262 | n1263 ;
  assign n1265 = ( x507 & ~n885 ) | ( x507 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1266 = x379 &  n885 ;
  assign n1267 = n1265 | n1266 ;
  assign n1268 = ~n1264 & n1267 ;
  assign n1272 = ( x250 & ~n1261 ) | ( x250 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1273 = x122 &  n1261 ;
  assign n1274 = n1272 | n1273 ;
  assign n1269 = ( x506 & ~n885 ) | ( x506 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1270 = x378 &  n885 ;
  assign n1271 = n1269 | n1270 ;
  assign n1275 = n1271 | n1274 ;
  assign n1276 = ( n1268 & ~n1274 ) | ( n1268 & n1275 ) | ( ~n1274 & n1275 ) ;
  assign n1277 = ( x249 & ~n1261 ) | ( x249 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1278 = x121 &  n1261 ;
  assign n1279 = n1277 | n1278 ;
  assign n1280 = ( x505 & ~n885 ) | ( x505 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1281 = x377 &  n885 ;
  assign n1282 = n1280 | n1281 ;
  assign n1283 = ~n1279 & n1282 ;
  assign n1284 = ( x504 & ~n885 ) | ( x504 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n1285 = x376 &  n885 ;
  assign n1286 = n1284 | n1285 ;
  assign n1287 = ( x248 & ~n1261 ) | ( x248 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n1288 = x120 &  n1261 ;
  assign n1289 = n1287 | n1288 ;
  assign n1290 = ( n1286 & ~n1289 ) | ( n1286 & 1'b0 ) | ( ~n1289 & 1'b0 ) ;
  assign n1291 = n1283 | n1290 ;
  assign n1292 = n1276 | n1291 ;
  assign n2355 = n2350 | n1292 ;
  assign n2351 = ~n1286 & n1289 ;
  assign n2352 = ( n1279 & ~n1282 ) | ( n1279 & n2351 ) | ( ~n1282 & n2351 ) ;
  assign n2353 = ( n1274 & ~n1271 ) | ( n1274 & n2352 ) | ( ~n1271 & n2352 ) ;
  assign n2354 = ( n1264 & ~n1267 ) | ( n1264 & n2353 ) | ( ~n1267 & n2353 ) ;
  assign n2356 = ( n2355 & ~n1292 ) | ( n2355 & n2354 ) | ( ~n1292 & n2354 ) ;
  assign n2360 = ( x508 & ~n885 ) | ( x508 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2361 = x380 &  n885 ;
  assign n2362 = n2360 | n2361 ;
  assign n2357 = ( x252 & ~n1261 ) | ( x252 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2358 = x124 &  n1261 ;
  assign n2359 = n2357 | n2358 ;
  assign n2384 = n2362 | n2359 ;
  assign n2365 = ~n1256 & x255 ;
  assign n2366 = ( x127 & n2365 ) | ( x127 & n1256 ) | ( n2365 & n1256 ) ;
  assign n2363 = ~n880 & x511 ;
  assign n2364 = ( x383 & n2363 ) | ( x383 & n880 ) | ( n2363 & n880 ) ;
  assign n2382 = n2366 | n2364 ;
  assign n2367 = ( x254 & ~n1261 ) | ( x254 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2368 = x126 &  n1261 ;
  assign n2369 = n2367 | n2368 ;
  assign n2370 = ( x510 & ~n885 ) | ( x510 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2371 = x382 &  n885 ;
  assign n2372 = n2370 | n2371 ;
  assign n2373 = ~n2369 & n2372 ;
  assign n2374 = ( x253 & ~n1261 ) | ( x253 & 1'b0 ) | ( ~n1261 & 1'b0 ) ;
  assign n2375 = x125 &  n1261 ;
  assign n2376 = n2374 | n2375 ;
  assign n2377 = ( x509 & ~n885 ) | ( x509 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n2378 = x381 &  n885 ;
  assign n2379 = n2377 | n2378 ;
  assign n2380 = n2376 &  n2379 ;
  assign n2381 = ( n2373 & ~n2380 ) | ( n2373 & n2379 ) | ( ~n2380 & n2379 ) ;
  assign n2383 = ( n2382 & ~n2364 ) | ( n2382 & n2381 ) | ( ~n2364 & n2381 ) ;
  assign n2385 = ( n2384 & ~n2359 ) | ( n2384 & n2383 ) | ( ~n2359 & n2383 ) ;
  assign n2386 = ( n2356 & ~n2385 ) | ( n2356 & 1'b0 ) | ( ~n2385 & 1'b0 ) ;
  assign n2387 = ( n2359 & ~n2362 ) | ( n2359 & 1'b0 ) | ( ~n2362 & 1'b0 ) ;
  assign n2388 = ( n2376 & ~n2379 ) | ( n2376 & n2387 ) | ( ~n2379 & n2387 ) ;
  assign n2389 = ( n2369 & ~n2372 ) | ( n2369 & n2388 ) | ( ~n2372 & n2388 ) ;
  assign n2390 = ( n2364 & ~n2366 ) | ( n2364 & n2389 ) | ( ~n2366 & n2389 ) ;
  assign n2391 = n2386 | n2390 ;
  assign n2392 = ( n888 & ~n2391 ) | ( n888 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2393 = n1929 &  n2391 ;
  assign n2394 = n2392 | n2393 ;
  assign n2395 = ( n1926 & ~n2391 ) | ( n1926 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2396 = n1933 &  n2391 ;
  assign n2397 = n2395 | n2396 ;
  assign n2398 = ( n1923 & ~n2391 ) | ( n1923 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2399 = n1920 &  n2391 ;
  assign n2400 = n2398 | n2399 ;
  assign n2401 = ( n1917 & ~n2391 ) | ( n1917 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2402 = n1914 &  n2391 ;
  assign n2403 = n2401 | n2402 ;
  assign n2404 = ( n1908 & ~n2391 ) | ( n1908 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2405 = n1911 &  n2391 ;
  assign n2406 = n2404 | n2405 ;
  assign n2407 = ( n1902 & ~n2391 ) | ( n1902 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2408 = n1905 &  n2391 ;
  assign n2409 = n2407 | n2408 ;
  assign n2410 = ( n1896 & ~n2391 ) | ( n1896 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2411 = n1899 &  n2391 ;
  assign n2412 = n2410 | n2411 ;
  assign n2413 = ( n1893 & ~n2391 ) | ( n1893 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2414 = n1890 &  n2391 ;
  assign n2415 = n2413 | n2414 ;
  assign n2416 = ( n1887 & ~n2391 ) | ( n1887 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2417 = n1943 &  n2391 ;
  assign n2418 = n2416 | n2417 ;
  assign n2419 = ( n1884 & ~n2391 ) | ( n1884 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2420 = n1947 &  n2391 ;
  assign n2421 = n2419 | n2420 ;
  assign n2422 = ( n1881 & ~n2391 ) | ( n1881 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2423 = n1878 &  n2391 ;
  assign n2424 = n2422 | n2423 ;
  assign n2425 = ( n1875 & ~n2391 ) | ( n1875 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2426 = n1872 &  n2391 ;
  assign n2427 = n2425 | n2426 ;
  assign n2428 = ( n1869 & ~n2391 ) | ( n1869 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2429 = n1866 &  n2391 ;
  assign n2430 = n2428 | n2429 ;
  assign n2431 = ( n1863 & ~n2391 ) | ( n1863 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2432 = n1860 &  n2391 ;
  assign n2433 = n2431 | n2432 ;
  assign n2434 = ( n1857 & ~n2391 ) | ( n1857 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2435 = n1854 &  n2391 ;
  assign n2436 = n2434 | n2435 ;
  assign n2437 = ( n1851 & ~n2391 ) | ( n1851 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2438 = n1848 &  n2391 ;
  assign n2439 = n2437 | n2438 ;
  assign n2440 = ( n1845 & ~n2391 ) | ( n1845 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2441 = n1957 &  n2391 ;
  assign n2442 = n2440 | n2441 ;
  assign n2443 = ( n1842 & ~n2391 ) | ( n1842 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2444 = n1961 &  n2391 ;
  assign n2445 = n2443 | n2444 ;
  assign n2446 = ( n1839 & ~n2391 ) | ( n1839 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2447 = n1836 &  n2391 ;
  assign n2448 = n2446 | n2447 ;
  assign n2449 = ( n1833 & ~n2391 ) | ( n1833 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2450 = n1830 &  n2391 ;
  assign n2451 = n2449 | n2450 ;
  assign n2452 = ( n1827 & ~n2391 ) | ( n1827 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2453 = n1824 &  n2391 ;
  assign n2454 = n2452 | n2453 ;
  assign n2455 = ( n1821 & ~n2391 ) | ( n1821 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2456 = n1818 &  n2391 ;
  assign n2457 = n2455 | n2456 ;
  assign n2458 = ( n1815 & ~n2391 ) | ( n1815 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2459 = n1812 &  n2391 ;
  assign n2460 = n2458 | n2459 ;
  assign n2461 = ( n1809 & ~n2391 ) | ( n1809 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2462 = n1806 &  n2391 ;
  assign n2463 = n2461 | n2462 ;
  assign n2464 = ( n1803 & ~n2391 ) | ( n1803 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2465 = n1971 &  n2391 ;
  assign n2466 = n2464 | n2465 ;
  assign n2467 = ( n1800 & ~n2391 ) | ( n1800 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2468 = n1975 &  n2391 ;
  assign n2469 = n2467 | n2468 ;
  assign n2470 = ( n1797 & ~n2391 ) | ( n1797 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2471 = n1794 &  n2391 ;
  assign n2472 = n2470 | n2471 ;
  assign n2473 = ( n1791 & ~n2391 ) | ( n1791 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2474 = n1788 &  n2391 ;
  assign n2475 = n2473 | n2474 ;
  assign n2476 = ( n1785 & ~n2391 ) | ( n1785 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2477 = n1782 &  n2391 ;
  assign n2478 = n2476 | n2477 ;
  assign n2479 = ( n1779 & ~n2391 ) | ( n1779 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2480 = n1776 &  n2391 ;
  assign n2481 = n2479 | n2480 ;
  assign n2482 = ( n1773 & ~n2391 ) | ( n1773 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2483 = n1770 &  n2391 ;
  assign n2484 = n2482 | n2483 ;
  assign n2485 = ( n1767 & ~n2391 ) | ( n1767 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2486 = n1764 &  n2391 ;
  assign n2487 = n2485 | n2486 ;
  assign n2488 = ( n1757 & ~n2391 ) | ( n1757 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2489 = n1760 &  n2391 ;
  assign n2490 = n2488 | n2489 ;
  assign n2491 = ( n1988 & ~n2391 ) | ( n1988 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2492 = n1985 &  n2391 ;
  assign n2493 = n2491 | n2492 ;
  assign n2494 = ( n2029 & ~n2391 ) | ( n2029 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2495 = n2032 &  n2391 ;
  assign n2496 = n2494 | n2495 ;
  assign n2497 = ( n2025 & ~n2391 ) | ( n2025 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2498 = n2022 &  n2391 ;
  assign n2499 = n2497 | n2498 ;
  assign n2500 = ( n2009 & ~n2391 ) | ( n2009 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2501 = n2006 &  n2391 ;
  assign n2502 = n2500 | n2501 ;
  assign n2503 = ( n2016 & ~n2391 ) | ( n2016 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2504 = n2013 &  n2391 ;
  assign n2505 = n2503 | n2504 ;
  assign n2506 = ( n1998 & ~n2391 ) | ( n1998 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2507 = n2001 &  n2391 ;
  assign n2508 = n2506 | n2507 ;
  assign n2509 = ( n1994 & ~n2391 ) | ( n1994 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2510 = n1991 &  n2391 ;
  assign n2511 = n2509 | n2510 ;
  assign n2512 = ( n1743 & ~n2391 ) | ( n1743 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2513 = n1740 &  n2391 ;
  assign n2514 = n2512 | n2513 ;
  assign n2515 = ( n1737 & ~n2391 ) | ( n1737 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2516 = n1734 &  n2391 ;
  assign n2517 = n2515 | n2516 ;
  assign n2518 = ( n1731 & ~n2391 ) | ( n1731 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2519 = n1728 &  n2391 ;
  assign n2520 = n2518 | n2519 ;
  assign n2521 = ( n1724 & ~n2391 ) | ( n1724 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2522 = n1721 &  n2391 ;
  assign n2523 = n2521 | n2522 ;
  assign n2524 = ( n1708 & ~n2391 ) | ( n1708 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2525 = n1705 &  n2391 ;
  assign n2526 = n2524 | n2525 ;
  assign n2527 = ( n1715 & ~n2391 ) | ( n1715 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2528 = n1712 &  n2391 ;
  assign n2529 = n2527 | n2528 ;
  assign n2530 = ( n1697 & ~n2391 ) | ( n1697 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2531 = n1700 &  n2391 ;
  assign n2532 = n2530 | n2531 ;
  assign n2533 = ( n1693 & ~n2391 ) | ( n1693 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2534 = n1690 &  n2391 ;
  assign n2535 = n2533 | n2534 ;
  assign n2536 = ( n2063 & ~n2391 ) | ( n2063 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2537 = n2066 &  n2391 ;
  assign n2538 = n2536 | n2537 ;
  assign n2539 = ( n2073 & ~n2391 ) | ( n2073 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2540 = n2070 &  n2391 ;
  assign n2541 = n2539 | n2540 ;
  assign n2542 = ( n2114 & ~n2391 ) | ( n2114 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2543 = n2117 &  n2391 ;
  assign n2544 = n2542 | n2543 ;
  assign n2545 = ( n2110 & ~n2391 ) | ( n2110 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2546 = n2107 &  n2391 ;
  assign n2547 = n2545 | n2546 ;
  assign n2548 = ( n2098 & ~n2391 ) | ( n2098 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2549 = n2101 &  n2391 ;
  assign n2550 = n2548 | n2549 ;
  assign n2551 = ( n2094 & ~n2391 ) | ( n2094 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2552 = n2091 &  n2391 ;
  assign n2553 = n2551 | n2552 ;
  assign n2554 = ( n2083 & ~n2391 ) | ( n2083 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2555 = n2086 &  n2391 ;
  assign n2556 = n2554 | n2555 ;
  assign n2557 = ( n2079 & ~n2391 ) | ( n2079 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2558 = n2076 &  n2391 ;
  assign n2559 = n2557 | n2558 ;
  assign n2560 = ( n1676 & ~n2391 ) | ( n1676 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2561 = n1673 &  n2391 ;
  assign n2562 = n2560 | n2561 ;
  assign n2563 = ( n1670 & ~n2391 ) | ( n1670 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2564 = n1667 &  n2391 ;
  assign n2565 = n2563 | n2564 ;
  assign n2566 = ( n1664 & ~n2391 ) | ( n1664 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2567 = n1661 &  n2391 ;
  assign n2568 = n2566 | n2567 ;
  assign n2569 = ( n1657 & ~n2391 ) | ( n1657 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2570 = n1654 &  n2391 ;
  assign n2571 = n2569 | n2570 ;
  assign n2572 = ( n1641 & ~n2391 ) | ( n1641 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2573 = n1638 &  n2391 ;
  assign n2574 = n2572 | n2573 ;
  assign n2575 = ( n1648 & ~n2391 ) | ( n1648 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2576 = n1645 &  n2391 ;
  assign n2577 = n2575 | n2576 ;
  assign n2578 = ( n1630 & ~n2391 ) | ( n1630 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2579 = n1633 &  n2391 ;
  assign n2580 = n2578 | n2579 ;
  assign n2581 = ( n1626 & ~n2391 ) | ( n1626 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2582 = n1623 &  n2391 ;
  assign n2583 = n2581 | n2582 ;
  assign n2584 = ( n2147 & ~n2391 ) | ( n2147 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2585 = n2150 &  n2391 ;
  assign n2586 = n2584 | n2585 ;
  assign n2587 = ( n2157 & ~n2391 ) | ( n2157 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2588 = n2154 &  n2391 ;
  assign n2589 = n2587 | n2588 ;
  assign n2590 = ( n2171 & ~n2391 ) | ( n2171 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2591 = n2174 &  n2391 ;
  assign n2592 = n2590 | n2591 ;
  assign n2593 = ( n2167 & ~n2391 ) | ( n2167 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2594 = n2164 &  n2391 ;
  assign n2595 = n2593 | n2594 ;
  assign n2596 = ( n1617 & ~n2391 ) | ( n1617 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2597 = n1614 &  n2391 ;
  assign n2598 = n2596 | n2597 ;
  assign n2599 = ( n1610 & ~n2391 ) | ( n1610 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2600 = n1607 &  n2391 ;
  assign n2601 = n2599 | n2600 ;
  assign n2602 = ( n1599 & ~n2391 ) | ( n1599 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2603 = n1602 &  n2391 ;
  assign n2604 = n2602 | n2603 ;
  assign n2605 = ( n1595 & ~n2391 ) | ( n1595 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2606 = n1592 &  n2391 ;
  assign n2607 = n2605 | n2606 ;
  assign n2608 = ( n1583 & ~n2391 ) | ( n1583 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2609 = n1586 &  n2391 ;
  assign n2610 = n2608 | n2609 ;
  assign n2611 = ( n1579 & ~n2391 ) | ( n1579 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2612 = n1576 &  n2391 ;
  assign n2613 = n2611 | n2612 ;
  assign n2614 = ( n1568 & ~n2391 ) | ( n1568 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2615 = n1571 &  n2391 ;
  assign n2616 = n2614 | n2615 ;
  assign n2617 = ( n1564 & ~n2391 ) | ( n1564 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2618 = n1561 &  n2391 ;
  assign n2619 = n2617 | n2618 ;
  assign n2620 = ( n1555 & ~n2391 ) | ( n1555 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2621 = n1552 &  n2391 ;
  assign n2622 = n2620 | n2621 ;
  assign n2623 = ( n1548 & ~n2391 ) | ( n1548 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2624 = n1545 &  n2391 ;
  assign n2625 = n2623 | n2624 ;
  assign n2626 = ( n1537 & ~n2391 ) | ( n1537 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2627 = n1540 &  n2391 ;
  assign n2628 = n2626 | n2627 ;
  assign n2629 = ( n1533 & ~n2391 ) | ( n1533 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2630 = n1530 &  n2391 ;
  assign n2631 = n2629 | n2630 ;
  assign n2632 = ( n1524 & ~n2391 ) | ( n1524 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2633 = n1527 &  n2391 ;
  assign n2634 = n2632 | n2633 ;
  assign n2635 = ( n2225 & ~n2391 ) | ( n2225 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2636 = n2222 &  n2391 ;
  assign n2637 = n2635 | n2636 ;
  assign n2638 = ( n2214 & ~n2391 ) | ( n2214 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2639 = n2217 &  n2391 ;
  assign n2640 = n2638 | n2639 ;
  assign n2641 = ( n2210 & ~n2391 ) | ( n2210 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2642 = n2207 &  n2391 ;
  assign n2643 = n2641 | n2642 ;
  assign n2644 = ( n1518 & ~n2391 ) | ( n1518 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2645 = n1515 &  n2391 ;
  assign n2646 = n2644 | n2645 ;
  assign n2647 = ( n1511 & ~n2391 ) | ( n1511 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2648 = n1508 &  n2391 ;
  assign n2649 = n2647 | n2648 ;
  assign n2650 = ( n1500 & ~n2391 ) | ( n1500 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2651 = n1503 &  n2391 ;
  assign n2652 = n2650 | n2651 ;
  assign n2653 = ( n1496 & ~n2391 ) | ( n1496 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2654 = n1493 &  n2391 ;
  assign n2655 = n2653 | n2654 ;
  assign n2656 = ( n1484 & ~n2391 ) | ( n1484 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2657 = n1487 &  n2391 ;
  assign n2658 = n2656 | n2657 ;
  assign n2659 = ( n1480 & ~n2391 ) | ( n1480 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2660 = n1477 &  n2391 ;
  assign n2661 = n2659 | n2660 ;
  assign n2662 = ( n1469 & ~n2391 ) | ( n1469 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2663 = n1472 &  n2391 ;
  assign n2664 = n2662 | n2663 ;
  assign n2665 = ( n1465 & ~n2391 ) | ( n1465 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2666 = n1462 &  n2391 ;
  assign n2667 = n2665 | n2666 ;
  assign n2668 = ( n1456 & ~n2391 ) | ( n1456 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2669 = n1453 &  n2391 ;
  assign n2670 = n2668 | n2669 ;
  assign n2671 = ( n1449 & ~n2391 ) | ( n1449 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2672 = n1446 &  n2391 ;
  assign n2673 = n2671 | n2672 ;
  assign n2674 = ( n1438 & ~n2391 ) | ( n1438 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2675 = n1441 &  n2391 ;
  assign n2676 = n2674 | n2675 ;
  assign n2677 = ( n1434 & ~n2391 ) | ( n1434 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2678 = n1431 &  n2391 ;
  assign n2679 = n2677 | n2678 ;
  assign n2680 = ( n1425 & ~n2391 ) | ( n1425 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2681 = n1428 &  n2391 ;
  assign n2682 = n2680 | n2681 ;
  assign n2683 = ( n2278 & ~n2391 ) | ( n2278 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2684 = n2275 &  n2391 ;
  assign n2685 = n2683 | n2684 ;
  assign n2686 = ( n2267 & ~n2391 ) | ( n2267 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2687 = n2270 &  n2391 ;
  assign n2688 = n2686 | n2687 ;
  assign n2689 = ( n2263 & ~n2391 ) | ( n2263 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2690 = n2260 &  n2391 ;
  assign n2691 = n2689 | n2690 ;
  assign n2692 = ( n1419 & ~n2391 ) | ( n1419 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2693 = n1416 &  n2391 ;
  assign n2694 = n2692 | n2693 ;
  assign n2695 = ( n1412 & ~n2391 ) | ( n1412 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2696 = n1409 &  n2391 ;
  assign n2697 = n2695 | n2696 ;
  assign n2698 = ( n1401 & ~n2391 ) | ( n1401 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2699 = n1404 &  n2391 ;
  assign n2700 = n2698 | n2699 ;
  assign n2701 = ( n1397 & ~n2391 ) | ( n1397 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2702 = n1394 &  n2391 ;
  assign n2703 = n2701 | n2702 ;
  assign n2704 = ( n1385 & ~n2391 ) | ( n1385 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2705 = n1388 &  n2391 ;
  assign n2706 = n2704 | n2705 ;
  assign n2707 = ( n1381 & ~n2391 ) | ( n1381 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2708 = n1378 &  n2391 ;
  assign n2709 = n2707 | n2708 ;
  assign n2710 = ( n1370 & ~n2391 ) | ( n1370 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2711 = n1373 &  n2391 ;
  assign n2712 = n2710 | n2711 ;
  assign n2713 = ( n1366 & ~n2391 ) | ( n1366 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2714 = n1363 &  n2391 ;
  assign n2715 = n2713 | n2714 ;
  assign n2716 = ( n1357 & ~n2391 ) | ( n1357 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2717 = n1354 &  n2391 ;
  assign n2718 = n2716 | n2717 ;
  assign n2719 = ( n1350 & ~n2391 ) | ( n1350 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2720 = n1347 &  n2391 ;
  assign n2721 = n2719 | n2720 ;
  assign n2722 = ( n1339 & ~n2391 ) | ( n1339 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2723 = n1342 &  n2391 ;
  assign n2724 = n2722 | n2723 ;
  assign n2725 = ( n1335 & ~n2391 ) | ( n1335 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2726 = n1332 &  n2391 ;
  assign n2727 = n2725 | n2726 ;
  assign n2728 = ( n1326 & ~n2391 ) | ( n1326 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2729 = n1329 &  n2391 ;
  assign n2730 = n2728 | n2729 ;
  assign n2731 = ( n2331 & ~n2391 ) | ( n2331 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2732 = n2328 &  n2391 ;
  assign n2733 = n2731 | n2732 ;
  assign n2734 = ( n2320 & ~n2391 ) | ( n2320 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2735 = n2323 &  n2391 ;
  assign n2736 = n2734 | n2735 ;
  assign n2737 = ( n2316 & ~n2391 ) | ( n2316 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2738 = n2313 &  n2391 ;
  assign n2739 = n2737 | n2738 ;
  assign n2740 = ( n1320 & ~n2391 ) | ( n1320 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2741 = n1317 &  n2391 ;
  assign n2742 = n2740 | n2741 ;
  assign n2743 = ( n1313 & ~n2391 ) | ( n1313 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2744 = n1310 &  n2391 ;
  assign n2745 = n2743 | n2744 ;
  assign n2746 = ( n1302 & ~n2391 ) | ( n1302 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2747 = n1305 &  n2391 ;
  assign n2748 = n2746 | n2747 ;
  assign n2749 = ( n1298 & ~n2391 ) | ( n1298 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2750 = n1295 &  n2391 ;
  assign n2751 = n2749 | n2750 ;
  assign n2752 = ( n1286 & ~n2391 ) | ( n1286 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2753 = n1289 &  n2391 ;
  assign n2754 = n2752 | n2753 ;
  assign n2755 = ( n1282 & ~n2391 ) | ( n1282 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2756 = n1279 &  n2391 ;
  assign n2757 = n2755 | n2756 ;
  assign n2758 = ( n1271 & ~n2391 ) | ( n1271 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2759 = n1274 &  n2391 ;
  assign n2760 = n2758 | n2759 ;
  assign n2761 = ( n1267 & ~n2391 ) | ( n1267 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2762 = n1264 &  n2391 ;
  assign n2763 = n2761 | n2762 ;
  assign n2764 = ( n2362 & ~n2391 ) | ( n2362 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2765 = n2359 &  n2391 ;
  assign n2766 = n2764 | n2765 ;
  assign n2767 = ( n2379 & ~n2391 ) | ( n2379 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2768 = n2376 &  n2391 ;
  assign n2769 = n2767 | n2768 ;
  assign n2770 = ( n2372 & ~n2391 ) | ( n2372 & 1'b0 ) | ( ~n2391 & 1'b0 ) ;
  assign n2771 = n2369 &  n2391 ;
  assign n2772 = n2770 | n2771 ;
  assign n2773 = ~n2364 & n2386 ;
  assign n2774 = ( n2364 & n2773 ) | ( n2364 & n2366 ) | ( n2773 & n2366 ) ;
  assign n2775 = n885 | n2391 ;
  assign n2776 = ~n1261 & n2391 ;
  assign n2777 = ( n2775 & ~n2776 ) | ( n2775 & 1'b0 ) | ( ~n2776 & 1'b0 ) ;
  assign y0 = n2394 ;
  assign y1 = n2397 ;
  assign y2 = n2400 ;
  assign y3 = n2403 ;
  assign y4 = n2406 ;
  assign y5 = n2409 ;
  assign y6 = n2412 ;
  assign y7 = n2415 ;
  assign y8 = n2418 ;
  assign y9 = n2421 ;
  assign y10 = n2424 ;
  assign y11 = n2427 ;
  assign y12 = n2430 ;
  assign y13 = n2433 ;
  assign y14 = n2436 ;
  assign y15 = n2439 ;
  assign y16 = n2442 ;
  assign y17 = n2445 ;
  assign y18 = n2448 ;
  assign y19 = n2451 ;
  assign y20 = n2454 ;
  assign y21 = n2457 ;
  assign y22 = n2460 ;
  assign y23 = n2463 ;
  assign y24 = n2466 ;
  assign y25 = n2469 ;
  assign y26 = n2472 ;
  assign y27 = n2475 ;
  assign y28 = n2478 ;
  assign y29 = n2481 ;
  assign y30 = n2484 ;
  assign y31 = n2487 ;
  assign y32 = n2490 ;
  assign y33 = n2493 ;
  assign y34 = n2496 ;
  assign y35 = n2499 ;
  assign y36 = n2502 ;
  assign y37 = n2505 ;
  assign y38 = n2508 ;
  assign y39 = n2511 ;
  assign y40 = n2514 ;
  assign y41 = n2517 ;
  assign y42 = n2520 ;
  assign y43 = n2523 ;
  assign y44 = n2526 ;
  assign y45 = n2529 ;
  assign y46 = n2532 ;
  assign y47 = n2535 ;
  assign y48 = n2538 ;
  assign y49 = n2541 ;
  assign y50 = n2544 ;
  assign y51 = n2547 ;
  assign y52 = n2550 ;
  assign y53 = n2553 ;
  assign y54 = n2556 ;
  assign y55 = n2559 ;
  assign y56 = n2562 ;
  assign y57 = n2565 ;
  assign y58 = n2568 ;
  assign y59 = n2571 ;
  assign y60 = n2574 ;
  assign y61 = n2577 ;
  assign y62 = n2580 ;
  assign y63 = n2583 ;
  assign y64 = n2586 ;
  assign y65 = n2589 ;
  assign y66 = n2592 ;
  assign y67 = n2595 ;
  assign y68 = n2598 ;
  assign y69 = n2601 ;
  assign y70 = n2604 ;
  assign y71 = n2607 ;
  assign y72 = n2610 ;
  assign y73 = n2613 ;
  assign y74 = n2616 ;
  assign y75 = n2619 ;
  assign y76 = n2622 ;
  assign y77 = n2625 ;
  assign y78 = n2628 ;
  assign y79 = n2631 ;
  assign y80 = n2634 ;
  assign y81 = n2637 ;
  assign y82 = n2640 ;
  assign y83 = n2643 ;
  assign y84 = n2646 ;
  assign y85 = n2649 ;
  assign y86 = n2652 ;
  assign y87 = n2655 ;
  assign y88 = n2658 ;
  assign y89 = n2661 ;
  assign y90 = n2664 ;
  assign y91 = n2667 ;
  assign y92 = n2670 ;
  assign y93 = n2673 ;
  assign y94 = n2676 ;
  assign y95 = n2679 ;
  assign y96 = n2682 ;
  assign y97 = n2685 ;
  assign y98 = n2688 ;
  assign y99 = n2691 ;
  assign y100 = n2694 ;
  assign y101 = n2697 ;
  assign y102 = n2700 ;
  assign y103 = n2703 ;
  assign y104 = n2706 ;
  assign y105 = n2709 ;
  assign y106 = n2712 ;
  assign y107 = n2715 ;
  assign y108 = n2718 ;
  assign y109 = n2721 ;
  assign y110 = n2724 ;
  assign y111 = n2727 ;
  assign y112 = n2730 ;
  assign y113 = n2733 ;
  assign y114 = n2736 ;
  assign y115 = n2739 ;
  assign y116 = n2742 ;
  assign y117 = n2745 ;
  assign y118 = n2748 ;
  assign y119 = n2751 ;
  assign y120 = n2754 ;
  assign y121 = n2757 ;
  assign y122 = n2760 ;
  assign y123 = n2763 ;
  assign y124 = n2766 ;
  assign y125 = n2769 ;
  assign y126 = n2772 ;
  assign y127 = n2774 ;
  assign y128 = ~n2777 ;
  assign y129 = ~n2391 ;
endmodule
