module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 ;
  assign n33 = x23 | x26 ;
  assign n34 = x24 &  x25 ;
  assign n35 = ~n33 & n34 ;
  assign n36 = x27 &  x28 ;
  assign n37 = ( x29 & ~x30 ) | ( x29 & 1'b0 ) | ( ~x30 & 1'b0 ) ;
  assign n38 = n36 &  n37 ;
  assign n39 = n35 &  n38 ;
  assign n40 = ~x27 & x28 ;
  assign n41 = x29 | x30 ;
  assign n42 = ( n40 & ~n41 ) | ( n40 & 1'b0 ) | ( ~n41 & 1'b0 ) ;
  assign n43 = n35 &  n42 ;
  assign n44 = x27 | x28 ;
  assign n45 = n41 | n44 ;
  assign n46 = ~x23 & x26 ;
  assign n47 = ( x24 & ~x25 ) | ( x24 & 1'b0 ) | ( ~x25 & 1'b0 ) ;
  assign n48 = n46 &  n47 ;
  assign n49 = ~n45 & n48 ;
  assign n50 = x29 &  x30 ;
  assign n51 = n40 &  n50 ;
  assign n52 = n48 &  n51 ;
  assign n53 = ( x27 & ~x28 ) | ( x27 & 1'b0 ) | ( ~x28 & 1'b0 ) ;
  assign n54 = ~x29 & x30 ;
  assign n55 = n53 &  n54 ;
  assign n56 = ( x23 & ~x26 ) | ( x23 & 1'b0 ) | ( ~x26 & 1'b0 ) ;
  assign n57 = n47 &  n56 ;
  assign n58 = n55 &  n57 ;
  assign n59 = n34 &  n56 ;
  assign n60 = n40 &  n54 ;
  assign n61 = n59 &  n60 ;
  assign n62 = n58 | n61 ;
  assign n63 = n34 &  n46 ;
  assign n64 = ~n44 & n54 ;
  assign n65 = n63 &  n64 ;
  assign n66 = ~x24 & x25 ;
  assign n67 = x23 &  x26 ;
  assign n68 = n66 &  n67 ;
  assign n69 = n60 &  n68 ;
  assign n70 = n65 | n69 ;
  assign n71 = n36 &  n54 ;
  assign n72 = n35 &  n71 ;
  assign n73 = ( n36 & ~n41 ) | ( n36 & 1'b0 ) | ( ~n41 & 1'b0 ) ;
  assign n74 = n35 &  n73 ;
  assign n75 = n72 | n74 ;
  assign n76 = n37 &  n40 ;
  assign n77 = n35 &  n76 ;
  assign n78 = x24 | x25 ;
  assign n79 = n33 | n78 ;
  assign n80 = ( n42 & ~n79 ) | ( n42 & 1'b0 ) | ( ~n79 & 1'b0 ) ;
  assign n81 = n77 | n80 ;
  assign n82 = n56 &  n66 ;
  assign n83 = n38 &  n82 ;
  assign n84 = ( n56 & ~n78 ) | ( n56 & 1'b0 ) | ( ~n78 & 1'b0 ) ;
  assign n85 = ( n37 & ~n44 ) | ( n37 & 1'b0 ) | ( ~n44 & 1'b0 ) ;
  assign n86 = n84 &  n85 ;
  assign n87 = ~n33 & n47 ;
  assign n88 = n76 &  n87 ;
  assign n89 = n59 &  n73 ;
  assign n90 = ~n41 & n53 ;
  assign n91 = n59 &  n90 ;
  assign n92 = n47 &  n67 ;
  assign n93 = n85 &  n92 ;
  assign n94 = n46 &  n66 ;
  assign n95 = n85 &  n94 ;
  assign n96 = n93 | n95 ;
  assign n97 = n37 &  n53 ;
  assign n98 = ( n67 & ~n78 ) | ( n67 & 1'b0 ) | ( ~n78 & 1'b0 ) ;
  assign n99 = n97 &  n98 ;
  assign n100 = n50 &  n53 ;
  assign n101 = n98 &  n100 ;
  assign n102 = n99 | n101 ;
  assign n103 = ~n33 & n66 ;
  assign n104 = n97 &  n103 ;
  assign n105 = n35 &  n51 ;
  assign n106 = n48 &  n71 ;
  assign n107 = n105 | n106 ;
  assign n108 = n104 | n107 ;
  assign n109 = ( n102 & ~n96 ) | ( n102 & n108 ) | ( ~n96 & n108 ) ;
  assign n110 = n96 | n109 ;
  assign n111 = ( n91 & ~n89 ) | ( n91 & n110 ) | ( ~n89 & n110 ) ;
  assign n112 = n89 | n111 ;
  assign n113 = ( n88 & ~n86 ) | ( n88 & n112 ) | ( ~n86 & n112 ) ;
  assign n114 = n86 | n113 ;
  assign n115 = n83 | n114 ;
  assign n116 = ( n46 & ~n78 ) | ( n46 & 1'b0 ) | ( ~n78 & 1'b0 ) ;
  assign n117 = n76 &  n116 ;
  assign n118 = n42 &  n92 ;
  assign n119 = n34 &  n67 ;
  assign n120 = n73 &  n119 ;
  assign n121 = ~n44 & n50 ;
  assign n122 = n48 &  n121 ;
  assign n123 = n87 &  n100 ;
  assign n124 = n60 &  n87 ;
  assign n125 = ( n60 & ~n79 ) | ( n60 & 1'b0 ) | ( ~n79 & 1'b0 ) ;
  assign n126 = n71 &  n116 ;
  assign n127 = n71 &  n98 ;
  assign n128 = n126 | n127 ;
  assign n129 = n63 &  n97 ;
  assign n130 = n51 &  n103 ;
  assign n131 = n36 &  n50 ;
  assign n132 = n59 &  n131 ;
  assign n133 = n130 | n132 ;
  assign n134 = n129 | n133 ;
  assign n135 = n76 &  n84 ;
  assign n136 = ~n45 & n116 ;
  assign n137 = n97 &  n116 ;
  assign n138 = n35 &  n55 ;
  assign n139 = n90 &  n116 ;
  assign n140 = n68 &  n85 ;
  assign n141 = ~n79 & n85 ;
  assign n142 = n140 | n141 ;
  assign n143 = ( n139 & ~n138 ) | ( n139 & n142 ) | ( ~n138 & n142 ) ;
  assign n144 = n138 | n143 ;
  assign n145 = ( n137 & ~n136 ) | ( n137 & n144 ) | ( ~n136 & n144 ) ;
  assign n146 = n136 | n145 ;
  assign n147 = n135 | n146 ;
  assign n148 = n42 &  n82 ;
  assign n149 = n82 &  n97 ;
  assign n150 = n71 &  n82 ;
  assign n151 = ~n45 & n59 ;
  assign n152 = n150 | n151 ;
  assign n153 = ( n149 & ~n148 ) | ( n149 & n152 ) | ( ~n148 & n152 ) ;
  assign n154 = n148 | n153 ;
  assign n155 = n38 &  n59 ;
  assign n156 = n76 &  n92 ;
  assign n157 = n60 &  n63 ;
  assign n158 = n156 | n157 ;
  assign n159 = n155 | n158 ;
  assign n160 = n42 &  n119 ;
  assign n161 = n90 &  n94 ;
  assign n162 = n90 &  n92 ;
  assign n163 = n161 | n162 ;
  assign n164 = n160 | n163 ;
  assign n165 = n48 &  n131 ;
  assign n166 = n85 &  n98 ;
  assign n167 = n68 &  n97 ;
  assign n168 = n35 &  n121 ;
  assign n169 = n92 &  n97 ;
  assign n170 = n168 | n169 ;
  assign n171 = n167 | n170 ;
  assign n172 = ( n166 & ~n165 ) | ( n166 & n171 ) | ( ~n165 & n171 ) ;
  assign n173 = n165 | n172 ;
  assign n174 = n164 | n173 ;
  assign n175 = ( n159 & ~n154 ) | ( n159 & n174 ) | ( ~n154 & n174 ) ;
  assign n176 = ( n154 & ~n147 ) | ( n154 & n175 ) | ( ~n147 & n175 ) ;
  assign n177 = n147 | n176 ;
  assign n178 = ( n134 & ~n128 ) | ( n134 & n177 ) | ( ~n128 & n177 ) ;
  assign n179 = n128 | n178 ;
  assign n180 = ( n125 & ~n124 ) | ( n125 & n179 ) | ( ~n124 & n179 ) ;
  assign n181 = n124 | n180 ;
  assign n182 = ( n123 & ~n122 ) | ( n123 & n181 ) | ( ~n122 & n181 ) ;
  assign n183 = n122 | n182 ;
  assign n184 = ( n120 & ~n118 ) | ( n120 & n183 ) | ( ~n118 & n183 ) ;
  assign n185 = n118 | n184 ;
  assign n186 = n117 | n185 ;
  assign n187 = n48 &  n100 ;
  assign n188 = n94 &  n100 ;
  assign n189 = n187 | n188 ;
  assign n205 = ~n45 & n94 ;
  assign n206 = n68 &  n121 ;
  assign n207 = n51 &  n57 ;
  assign n208 = n64 &  n119 ;
  assign n209 = n207 | n208 ;
  assign n210 = ( n206 & ~n205 ) | ( n206 & n209 ) | ( ~n205 & n209 ) ;
  assign n211 = n205 | n210 ;
  assign n212 = n38 &  n87 ;
  assign n213 = n76 &  n98 ;
  assign n214 = n90 &  n119 ;
  assign n215 = n213 | n214 ;
  assign n216 = n63 &  n100 ;
  assign n217 = n51 &  n92 ;
  assign n218 = n216 | n217 ;
  assign n219 = n215 | n218 ;
  assign n220 = n212 | n219 ;
  assign n221 = n42 &  n87 ;
  assign n222 = ~n79 & n100 ;
  assign n223 = n221 | n222 ;
  assign n224 = n55 &  n92 ;
  assign n225 = n38 &  n63 ;
  assign n226 = n82 &  n131 ;
  assign n227 = n225 | n226 ;
  assign n228 = n84 &  n97 ;
  assign n229 = n57 &  n85 ;
  assign n230 = ~n79 & n131 ;
  assign n231 = n100 &  n119 ;
  assign n232 = n98 &  n121 ;
  assign n233 = n51 &  n63 ;
  assign n234 = n64 &  n92 ;
  assign n235 = n71 &  n119 ;
  assign n236 = ~n79 & n97 ;
  assign n237 = n68 &  n73 ;
  assign n238 = n236 | n237 ;
  assign n239 = n42 &  n94 ;
  assign n240 = n42 &  n103 ;
  assign n241 = n51 &  n87 ;
  assign n242 = n64 &  n84 ;
  assign n243 = n64 &  n82 ;
  assign n244 = n71 &  n87 ;
  assign n245 = n64 &  n103 ;
  assign n246 = n244 | n245 ;
  assign n247 = n243 | n246 ;
  assign n248 = ( n242 & ~n241 ) | ( n242 & n247 ) | ( ~n241 & n247 ) ;
  assign n249 = n241 | n248 ;
  assign n250 = ( n240 & ~n239 ) | ( n240 & n249 ) | ( ~n239 & n249 ) ;
  assign n251 = n239 | n250 ;
  assign n252 = n85 &  n103 ;
  assign n253 = n55 &  n59 ;
  assign n254 = n252 | n253 ;
  assign n255 = n84 &  n90 ;
  assign n256 = n48 &  n76 ;
  assign n257 = n55 &  n119 ;
  assign n258 = n71 &  n94 ;
  assign n259 = n60 &  n98 ;
  assign n260 = n60 &  n116 ;
  assign n261 = n259 | n260 ;
  assign n262 = ( n258 & ~n257 ) | ( n258 & n261 ) | ( ~n257 & n261 ) ;
  assign n263 = n257 | n262 ;
  assign n264 = ( n256 & ~n255 ) | ( n256 & n263 ) | ( ~n255 & n263 ) ;
  assign n265 = n255 | n264 ;
  assign n299 = n73 &  n87 ;
  assign n300 = n42 &  n57 ;
  assign n301 = n299 | n300 ;
  assign n266 = ~n45 & n68 ;
  assign n267 = ( n35 & ~n45 ) | ( n35 & 1'b0 ) | ( ~n45 & 1'b0 ) ;
  assign n268 = n90 &  n98 ;
  assign n269 = n119 &  n131 ;
  assign n270 = n63 &  n131 ;
  assign n271 = n100 &  n116 ;
  assign n272 = n92 &  n121 ;
  assign n273 = ~n79 & n121 ;
  assign n274 = n51 &  n94 ;
  assign n275 = n71 &  n92 ;
  assign n276 = n76 &  n82 ;
  assign n277 = n64 &  n94 ;
  assign n278 = n276 | n277 ;
  assign n279 = ~n45 & n84 ;
  assign n280 = n57 &  n64 ;
  assign n281 = ~n45 & n63 ;
  assign n282 = n280 | n281 ;
  assign n283 = n279 | n282 ;
  assign n284 = n116 &  n121 ;
  assign n285 = n76 &  n94 ;
  assign n286 = n284 | n285 ;
  assign n287 = n283 | n286 ;
  assign n288 = ( n278 & ~n275 ) | ( n278 & n287 ) | ( ~n275 & n287 ) ;
  assign n289 = n275 | n288 ;
  assign n290 = ( n274 & ~n273 ) | ( n274 & n289 ) | ( ~n273 & n289 ) ;
  assign n291 = n273 | n290 ;
  assign n292 = ( n272 & ~n271 ) | ( n272 & n291 ) | ( ~n271 & n291 ) ;
  assign n293 = n271 | n292 ;
  assign n294 = ( n270 & ~n269 ) | ( n270 & n293 ) | ( ~n269 & n293 ) ;
  assign n295 = n269 | n294 ;
  assign n296 = ( n268 & ~n267 ) | ( n268 & n295 ) | ( ~n267 & n295 ) ;
  assign n297 = n267 | n296 ;
  assign n298 = n266 | n297 ;
  assign n302 = ( n301 & ~n265 ) | ( n301 & n298 ) | ( ~n265 & n298 ) ;
  assign n303 = ( n265 & ~n254 ) | ( n265 & n302 ) | ( ~n254 & n302 ) ;
  assign n304 = n254 | n303 ;
  assign n305 = ( n251 & ~n238 ) | ( n251 & n304 ) | ( ~n238 & n304 ) ;
  assign n306 = n238 | n305 ;
  assign n307 = ( n235 & ~n234 ) | ( n235 & n306 ) | ( ~n234 & n306 ) ;
  assign n308 = n234 | n307 ;
  assign n309 = ( n233 & ~n232 ) | ( n233 & n308 ) | ( ~n232 & n308 ) ;
  assign n310 = n232 | n309 ;
  assign n311 = ( n231 & ~n230 ) | ( n231 & n310 ) | ( ~n230 & n310 ) ;
  assign n312 = n230 | n311 ;
  assign n313 = ( n229 & ~n228 ) | ( n229 & n312 ) | ( ~n228 & n312 ) ;
  assign n314 = n228 | n313 ;
  assign n315 = ( n227 & ~n224 ) | ( n227 & n314 ) | ( ~n224 & n314 ) ;
  assign n316 = n224 | n315 ;
  assign n317 = n223 | n316 ;
  assign n318 = ( n220 & ~n211 ) | ( n220 & n317 ) | ( ~n211 & n317 ) ;
  assign n319 = n211 | n318 ;
  assign n190 = n73 &  n82 ;
  assign n191 = n87 &  n121 ;
  assign n192 = n87 &  n90 ;
  assign n193 = ( n64 & ~n79 ) | ( n64 & 1'b0 ) | ( ~n79 & 1'b0 ) ;
  assign n194 = ( n71 & ~n79 ) | ( n71 & 1'b0 ) | ( ~n79 & 1'b0 ) ;
  assign n195 = n60 &  n94 ;
  assign n196 = n85 &  n119 ;
  assign n197 = n45 | n79 ;
  assign n198 = ~n196 & n197 ;
  assign n199 = ~n195 & n198 ;
  assign n200 = ( n193 & ~n194 ) | ( n193 & n199 ) | ( ~n194 & n199 ) ;
  assign n201 = ~n193 & n200 ;
  assign n202 = ( n191 & ~n192 ) | ( n191 & n201 ) | ( ~n192 & n201 ) ;
  assign n203 = ~n191 & n202 ;
  assign n204 = ~n190 & n203 ;
  assign n320 = ( n189 & ~n319 ) | ( n189 & n204 ) | ( ~n319 & n204 ) ;
  assign n321 = ~n189 & n320 ;
  assign n322 = ( n115 & ~n186 ) | ( n115 & n321 ) | ( ~n186 & n321 ) ;
  assign n323 = ~n115 & n322 ;
  assign n324 = ( n75 & ~n81 ) | ( n75 & n323 ) | ( ~n81 & n323 ) ;
  assign n325 = ~n75 & n324 ;
  assign n326 = ( n62 & ~n70 ) | ( n62 & n325 ) | ( ~n70 & n325 ) ;
  assign n327 = ~n62 & n326 ;
  assign n328 = ( n49 & ~n52 ) | ( n49 & n327 ) | ( ~n52 & n327 ) ;
  assign n329 = ~n49 & n328 ;
  assign n330 = ( n39 & ~n43 ) | ( n39 & n329 ) | ( ~n43 & n329 ) ;
  assign n331 = ~n39 & n330 ;
  assign n332 = n59 &  n97 ;
  assign n333 = n55 &  n68 ;
  assign n334 = n57 &  n76 ;
  assign n335 = n130 | n334 ;
  assign n336 = n85 &  n116 ;
  assign n337 = n156 | n336 ;
  assign n338 = n48 &  n90 ;
  assign n339 = n207 | n338 ;
  assign n340 = n57 &  n97 ;
  assign n341 = n280 | n340 ;
  assign n342 = n42 &  n68 ;
  assign n343 = ~n119 |  n45 ;
  assign n344 = ~n342 & n343 ;
  assign n347 = n38 &  n84 ;
  assign n348 = n84 &  n131 ;
  assign n349 = n63 &  n121 ;
  assign n350 = n119 &  n121 ;
  assign n351 = n38 &  n119 ;
  assign n352 = n350 | n351 ;
  assign n372 = n100 &  n103 ;
  assign n373 = n35 &  n100 ;
  assign n374 = n35 &  n60 ;
  assign n375 = n188 | n374 ;
  assign n376 = n57 &  n60 ;
  assign n377 = n229 | n376 ;
  assign n378 = n375 | n377 ;
  assign n379 = ( n373 & ~n372 ) | ( n373 & n378 ) | ( ~n372 & n378 ) ;
  assign n380 = n372 | n379 ;
  assign n381 = n267 | n380 ;
  assign n382 = n57 &  n131 ;
  assign n383 = n272 | n382 ;
  assign n384 = n57 &  n73 ;
  assign n385 = n244 | n384 ;
  assign n386 = ( n218 & ~n88 ) | ( n218 & n242 ) | ( ~n88 & n242 ) ;
  assign n387 = n88 | n386 ;
  assign n388 = n91 | n132 ;
  assign n389 = n221 | n388 ;
  assign n390 = ( n387 & ~n385 ) | ( n387 & n389 ) | ( ~n385 & n389 ) ;
  assign n391 = n385 | n390 ;
  assign n392 = ( n383 & ~n381 ) | ( n383 & n391 ) | ( ~n381 & n391 ) ;
  assign n393 = n381 | n392 ;
  assign n353 = n68 &  n76 ;
  assign n354 = ~n82 | ~n85 ;
  assign n355 = ~n151 & n354 ;
  assign n356 = n59 &  n76 ;
  assign n357 = n208 | n356 ;
  assign n358 = ( n38 & ~n79 ) | ( n38 & 1'b0 ) | ( ~n79 & 1'b0 ) ;
  assign n359 = n55 &  n82 ;
  assign n360 = n72 | n359 ;
  assign n361 = n358 | n360 ;
  assign n362 = n60 &  n84 ;
  assign n363 = n148 | n362 ;
  assign n364 = n361 | n363 ;
  assign n365 = ( n355 & n357 ) | ( n355 & n364 ) | ( n357 & n364 ) ;
  assign n366 = ( n355 & ~n365 ) | ( n355 & 1'b0 ) | ( ~n365 & 1'b0 ) ;
  assign n367 = ( n243 & ~n253 ) | ( n243 & n366 ) | ( ~n253 & n366 ) ;
  assign n368 = ~n243 & n367 ;
  assign n369 = ( n162 & ~n89 ) | ( n162 & n368 ) | ( ~n89 & n368 ) ;
  assign n370 = ~n162 & n369 ;
  assign n371 = ~n353 & n370 ;
  assign n394 = ( n352 & ~n393 ) | ( n352 & n371 ) | ( ~n393 & n371 ) ;
  assign n395 = ~n352 & n394 ;
  assign n396 = ( n349 & ~n257 ) | ( n349 & n395 ) | ( ~n257 & n395 ) ;
  assign n397 = ~n349 & n396 ;
  assign n398 = ( n161 & ~n348 ) | ( n161 & n397 ) | ( ~n348 & n397 ) ;
  assign n399 = ~n161 & n398 ;
  assign n400 = ( n285 & ~n129 ) | ( n285 & n399 ) | ( ~n129 & n399 ) ;
  assign n401 = ~n285 & n400 ;
  assign n402 = ~n347 & n401 ;
  assign n403 = n42 &  n59 ;
  assign n404 = n68 &  n131 ;
  assign n405 = ~n45 & n87 ;
  assign n406 = ~n45 & n57 ;
  assign n407 = n405 | n406 ;
  assign n408 = n60 &  n119 ;
  assign n409 = n191 | n408 ;
  assign n410 = n38 &  n92 ;
  assign n411 = n73 &  n103 ;
  assign n412 = n410 | n411 ;
  assign n413 = n139 | n237 ;
  assign n414 = n224 | n268 ;
  assign n415 = n55 &  n98 ;
  assign n416 = n269 | n415 ;
  assign n417 = ~n45 & n92 ;
  assign n418 = n51 &  n59 ;
  assign n419 = n417 | n418 ;
  assign n420 = ( n240 & ~n49 ) | ( n240 & n419 ) | ( ~n49 & n419 ) ;
  assign n421 = n49 | n420 ;
  assign n422 = ( n213 & ~n300 ) | ( n213 & n421 ) | ( ~n300 & n421 ) ;
  assign n423 = n300 | n422 ;
  assign n424 = n57 &  n100 ;
  assign n425 = n57 &  n71 ;
  assign n426 = n277 | n425 ;
  assign n427 = ( n424 & ~n168 ) | ( n424 & n426 ) | ( ~n168 & n426 ) ;
  assign n428 = n168 | n427 ;
  assign n429 = n64 &  n116 ;
  assign n430 = n65 | n429 ;
  assign n431 = n38 &  n68 ;
  assign n432 = n38 &  n48 ;
  assign n433 = n38 &  n94 ;
  assign n434 = n225 | n433 ;
  assign n435 = n432 | n434 ;
  assign n436 = n431 | n435 ;
  assign n437 = n430 | n436 ;
  assign n438 = ( n198 & n428 ) | ( n198 & n437 ) | ( n428 & n437 ) ;
  assign n439 = ( n198 & ~n438 ) | ( n198 & 1'b0 ) | ( ~n438 & 1'b0 ) ;
  assign n440 = ( n416 & ~n423 ) | ( n416 & n439 ) | ( ~n423 & n439 ) ;
  assign n441 = ~n416 & n440 ;
  assign n442 = ( n413 & ~n414 ) | ( n413 & n441 ) | ( ~n414 & n441 ) ;
  assign n443 = ~n413 & n442 ;
  assign n444 = ( n409 & ~n412 ) | ( n409 & n443 ) | ( ~n412 & n443 ) ;
  assign n445 = ~n409 & n444 ;
  assign n446 = ( n404 & ~n407 ) | ( n404 & n445 ) | ( ~n407 & n445 ) ;
  assign n447 = ~n404 & n446 ;
  assign n448 = ( n160 & ~n403 ) | ( n160 & n447 ) | ( ~n403 & n447 ) ;
  assign n449 = ~n160 & n448 ;
  assign n450 = ~n99 & n449 ;
  assign n451 = n116 &  n131 ;
  assign n452 = n68 &  n90 ;
  assign n453 = n87 &  n131 ;
  assign n456 = n103 &  n131 ;
  assign n457 = n68 &  n100 ;
  assign n458 = n456 | n457 ;
  assign n459 = n63 &  n85 ;
  assign n460 = n82 &  n90 ;
  assign n461 = n459 | n460 ;
  assign n462 = n77 | n232 ;
  assign n463 = n83 | n125 ;
  assign n464 = n462 | n463 ;
  assign n465 = ( n461 & ~n458 ) | ( n461 & n464 ) | ( ~n458 & n464 ) ;
  assign n466 = n458 | n465 ;
  assign n454 = n42 &  n48 ;
  assign n455 = n118 | n454 ;
  assign n467 = ( n466 & ~n106 ) | ( n466 & n455 ) | ( ~n106 & n455 ) ;
  assign n468 = n106 | n467 ;
  assign n469 = ( n453 & ~n122 ) | ( n453 & n468 ) | ( ~n122 & n468 ) ;
  assign n470 = n122 | n469 ;
  assign n471 = ( n452 & ~n451 ) | ( n452 & n470 ) | ( ~n451 & n470 ) ;
  assign n472 = n451 | n471 ;
  assign n473 = ( n266 & ~n137 ) | ( n266 & n472 ) | ( ~n137 & n472 ) ;
  assign n474 = n137 | n473 ;
  assign n475 = n55 &  n84 ;
  assign n476 = n85 &  n87 ;
  assign n477 = n192 | n476 ;
  assign n478 = ( n76 & ~n79 ) | ( n76 & 1'b0 ) | ( ~n79 & 1'b0 ) ;
  assign n479 = n193 | n478 ;
  assign n480 = ( n194 & ~n477 ) | ( n194 & n479 ) | ( ~n477 & n479 ) ;
  assign n481 = n477 | n480 ;
  assign n482 = ( n475 & ~n245 ) | ( n475 & n481 ) | ( ~n245 & n481 ) ;
  assign n483 = n245 | n482 ;
  assign n490 = n51 &  n82 ;
  assign n491 = n136 | n490 ;
  assign n492 = n87 &  n97 ;
  assign n493 = n63 &  n71 ;
  assign n494 = n103 &  n121 ;
  assign n495 = n493 | n494 ;
  assign n496 = ( n492 & ~n231 ) | ( n492 & n495 ) | ( ~n231 & n495 ) ;
  assign n497 = n231 | n496 ;
  assign n498 = n491 | n497 ;
  assign n484 = ~n73 |  n79 ;
  assign n485 = n35 &  n131 ;
  assign n486 = n150 | n241 ;
  assign n487 = n273 | n486 ;
  assign n488 = ( n484 & n485 ) | ( n484 & n487 ) | ( n485 & n487 ) ;
  assign n489 = ( n484 & ~n488 ) | ( n484 & 1'b0 ) | ( ~n488 & 1'b0 ) ;
  assign n499 = ( n483 & ~n498 ) | ( n483 & n489 ) | ( ~n498 & n489 ) ;
  assign n500 = ~n483 & n499 ;
  assign n501 = ( n474 & ~n500 ) | ( n474 & n450 ) | ( ~n500 & n450 ) ;
  assign n502 = ( n402 & ~n450 ) | ( n402 & n501 ) | ( ~n450 & n501 ) ;
  assign n503 = ( n402 & ~n502 ) | ( n402 & 1'b0 ) | ( ~n502 & 1'b0 ) ;
  assign n345 = n48 &  n60 ;
  assign n346 = n212 | n345 ;
  assign n504 = ( n344 & ~n503 ) | ( n344 & n346 ) | ( ~n503 & n346 ) ;
  assign n505 = ( n344 & ~n504 ) | ( n344 & 1'b0 ) | ( ~n504 & 1'b0 ) ;
  assign n506 = ( n339 & ~n341 ) | ( n339 & n505 ) | ( ~n341 & n505 ) ;
  assign n507 = ~n339 & n506 ;
  assign n508 = ( n335 & ~n337 ) | ( n335 & n507 ) | ( ~n337 & n507 ) ;
  assign n509 = ~n335 & n508 ;
  assign n510 = ( n333 & ~n69 ) | ( n333 & n509 ) | ( ~n69 & n509 ) ;
  assign n511 = ~n333 & n510 ;
  assign n512 = ( n299 & ~n214 ) | ( n299 & n511 ) | ( ~n214 & n511 ) ;
  assign n513 = ~n299 & n512 ;
  assign n514 = ~n332 & n513 ;
  assign n3643 = n37 | n54 ;
  assign n3644 = ~x31 | ~n3643 ;
  assign n516 = ( x28 & ~x29 ) | ( x28 & 1'b0 ) | ( ~x29 & 1'b0 ) ;
  assign n517 = ~x28 & x29 ;
  assign n518 = n516 | n517 ;
  assign n519 = ( x26 & ~x27 ) | ( x26 & 1'b0 ) | ( ~x27 & 1'b0 ) ;
  assign n520 = ~x26 & x27 ;
  assign n521 = n519 | n520 ;
  assign n522 = ( n518 & ~n521 ) | ( n518 & 1'b0 ) | ( ~n521 & 1'b0 ) ;
  assign n515 = ~n36 & n44 ;
  assign n523 = ~n522 |  n515 ;
  assign n526 = ~n45 & n103 ;
  assign n527 = n281 | n526 ;
  assign n528 = n136 | n407 ;
  assign n529 = ~n45 & n98 ;
  assign n530 = n279 | n529 ;
  assign n540 = ~n45 & n82 ;
  assign n541 = n267 | n540 ;
  assign n531 = n57 &  n90 ;
  assign n532 = n192 | n531 ;
  assign n533 = n417 | n532 ;
  assign n534 = ~n79 & n90 ;
  assign n535 = n255 | n534 ;
  assign n536 = ( n533 & ~n205 ) | ( n533 & n535 ) | ( ~n205 & n535 ) ;
  assign n537 = n205 | n536 ;
  assign n538 = ( n537 & ~n49 ) | ( n537 & n266 ) | ( ~n49 & n266 ) ;
  assign n539 = n49 | n538 ;
  assign n542 = ( n541 & ~n530 ) | ( n541 & n539 ) | ( ~n530 & n539 ) ;
  assign n543 = n530 | n542 ;
  assign n544 = ( n528 & ~n527 ) | ( n528 & n543 ) | ( ~n527 & n543 ) ;
  assign n545 = n527 | n544 ;
  assign n524 = ~n90 | ~n103 ;
  assign n525 = n343 &  n524 ;
  assign n546 = ( n151 & ~n545 ) | ( n151 & n525 ) | ( ~n545 & n525 ) ;
  assign n547 = ~n151 & n546 ;
  assign n548 = n197 &  n547 ;
  assign n549 = n35 &  n90 ;
  assign n550 = n139 | n549 ;
  assign n551 = ( n91 & ~n338 ) | ( n91 & n550 ) | ( ~n338 & n550 ) ;
  assign n552 = n338 | n551 ;
  assign n553 = n268 | n552 ;
  assign n554 = n73 &  n84 ;
  assign n555 = n384 | n411 ;
  assign n556 = n42 &  n84 ;
  assign n557 = n300 | n556 ;
  assign n558 = n73 &  n116 ;
  assign n559 = n73 &  n92 ;
  assign n560 = n48 &  n73 ;
  assign n561 = n73 &  n94 ;
  assign n562 = n560 | n561 ;
  assign n563 = n559 | n562 ;
  assign n564 = ( n74 & ~n558 ) | ( n74 & n563 ) | ( ~n558 & n563 ) ;
  assign n565 = n558 | n564 ;
  assign n566 = ( n89 & ~n190 ) | ( n89 & n565 ) | ( ~n190 & n565 ) ;
  assign n567 = n190 | n566 ;
  assign n568 = n73 &  n98 ;
  assign n569 = n63 &  n90 ;
  assign n570 = n568 | n569 ;
  assign n571 = n42 &  n116 ;
  assign n572 = n42 &  n98 ;
  assign n573 = n43 | n240 ;
  assign n574 = n42 &  n63 ;
  assign n575 = n452 | n574 ;
  assign n576 = n80 | n214 ;
  assign n577 = n160 | n221 ;
  assign n578 = n576 | n577 ;
  assign n579 = ( n575 & ~n573 ) | ( n575 & n578 ) | ( ~n573 & n578 ) ;
  assign n580 = n573 | n579 ;
  assign n581 = ( n299 & ~n580 ) | ( n299 & n484 ) | ( ~n580 & n484 ) ;
  assign n582 = ~n299 & n581 ;
  assign n583 = ( n572 & ~n239 ) | ( n572 & n582 ) | ( ~n239 & n582 ) ;
  assign n584 = ~n572 & n583 ;
  assign n585 = ( n148 & ~n571 ) | ( n148 & n584 ) | ( ~n571 & n584 ) ;
  assign n586 = ~n148 & n585 ;
  assign n587 = ( n567 & ~n570 ) | ( n567 & n586 ) | ( ~n570 & n586 ) ;
  assign n588 = ( n557 & ~n567 ) | ( n557 & n587 ) | ( ~n567 & n587 ) ;
  assign n589 = ~n557 & n588 ;
  assign n590 = ( n163 & ~n555 ) | ( n163 & n589 ) | ( ~n555 & n589 ) ;
  assign n591 = ~n163 & n590 ;
  assign n592 = ( n554 & ~n455 ) | ( n554 & n591 ) | ( ~n455 & n591 ) ;
  assign n593 = ~n554 & n592 ;
  assign n594 = ( n342 & ~n403 ) | ( n342 & n593 ) | ( ~n403 & n593 ) ;
  assign n595 = ~n342 & n594 ;
  assign n596 = ( n460 & ~n553 ) | ( n460 & n595 ) | ( ~n553 & n595 ) ;
  assign n597 = ~n460 & n596 ;
  assign n598 = ~n237 & n597 ;
  assign n599 = n548 &  n598 ;
  assign n600 = n523 | n599 ;
  assign n601 = ~n518 | ~n521 ;
  assign n602 = ( n55 & ~n79 ) | ( n55 & 1'b0 ) | ( ~n79 & 1'b0 ) ;
  assign n603 = n94 &  n97 ;
  assign n604 = n149 | n332 ;
  assign n605 = n117 | n285 ;
  assign n606 = n99 | n358 ;
  assign n607 = n88 | n492 ;
  assign n608 = n606 | n607 ;
  assign n609 = ( n605 & ~n604 ) | ( n605 & n608 ) | ( ~n604 & n608 ) ;
  assign n610 = n604 | n609 ;
  assign n611 = ( n340 & ~n167 ) | ( n340 & n610 ) | ( ~n167 & n610 ) ;
  assign n612 = n167 | n611 ;
  assign n613 = ( n603 & ~n356 ) | ( n603 & n612 ) | ( ~n356 & n612 ) ;
  assign n614 = n356 | n613 ;
  assign n615 = ( n156 & ~n213 ) | ( n156 & n614 ) | ( ~n213 & n614 ) ;
  assign n616 = n213 | n615 ;
  assign n617 = n48 &  n85 ;
  assign n618 = n97 &  n119 ;
  assign n619 = n135 | n478 ;
  assign n620 = n256 | n334 ;
  assign n621 = ( n104 & ~n129 ) | ( n104 & n620 ) | ( ~n129 & n620 ) ;
  assign n622 = n129 | n621 ;
  assign n627 = n48 &  n97 ;
  assign n628 = n76 &  n119 ;
  assign n629 = n228 | n628 ;
  assign n630 = n63 &  n76 ;
  assign n631 = n76 &  n103 ;
  assign n632 = n630 | n631 ;
  assign n633 = n629 | n632 ;
  assign n634 = n627 | n633 ;
  assign n623 = ~n35 | ~n97 ;
  assign n624 = ~n169 & n623 ;
  assign n625 = ~n276 & n624 ;
  assign n626 = ~n353 & n625 ;
  assign n635 = ( n622 & ~n634 ) | ( n622 & n626 ) | ( ~n634 & n626 ) ;
  assign n636 = ~n622 & n635 ;
  assign n637 = ( n618 & ~n619 ) | ( n618 & n636 ) | ( ~n619 & n636 ) ;
  assign n638 = ~n618 & n637 ;
  assign n639 = ( n77 & ~n137 ) | ( n77 & n638 ) | ( ~n137 & n638 ) ;
  assign n640 = ~n77 & n639 ;
  assign n641 = ( n617 & ~n236 ) | ( n617 & n640 ) | ( ~n236 & n640 ) ;
  assign n642 = ~n617 & n641 ;
  assign n643 = n35 &  n85 ;
  assign n644 = ~n63 | ~n73 ;
  assign n645 = ~n86 & n644 ;
  assign n646 = n59 &  n85 ;
  assign n647 = n196 | n646 ;
  assign n648 = ( n645 & ~n647 ) | ( n645 & 1'b0 ) | ( ~n647 & 1'b0 ) ;
  assign n649 = ( n141 & ~n120 ) | ( n141 & n648 ) | ( ~n120 & n648 ) ;
  assign n650 = ~n141 & n649 ;
  assign n651 = ( n229 & ~n650 ) | ( n229 & n354 ) | ( ~n650 & n354 ) ;
  assign n652 = ( n354 & ~n651 ) | ( n354 & 1'b0 ) | ( ~n651 & 1'b0 ) ;
  assign n653 = ~n166 & n652 ;
  assign n654 = n252 | n336 ;
  assign n655 = ( n653 & ~n654 ) | ( n653 & 1'b0 ) | ( ~n654 & 1'b0 ) ;
  assign n656 = ( n96 & ~n643 ) | ( n96 & n655 ) | ( ~n643 & n655 ) ;
  assign n657 = ~n96 & n656 ;
  assign n658 = ~n140 & n657 ;
  assign n659 = ( n616 & n642 ) | ( n616 & n658 ) | ( n642 & n658 ) ;
  assign n660 = ( n459 & ~n616 ) | ( n459 & n659 ) | ( ~n616 & n659 ) ;
  assign n661 = ~n459 & n660 ;
  assign n662 = ~n476 & n661 ;
  assign n666 = n38 &  n57 ;
  assign n667 = n347 | n666 ;
  assign n668 = n83 | n155 ;
  assign n669 = n39 | n668 ;
  assign n670 = n38 &  n98 ;
  assign n671 = n48 &  n64 ;
  assign n672 = n64 &  n98 ;
  assign n673 = n277 | n672 ;
  assign n674 = n35 &  n64 ;
  assign n675 = n242 | n674 ;
  assign n676 = n64 &  n68 ;
  assign n677 = n351 | n676 ;
  assign n678 = n59 &  n64 ;
  assign n679 = n64 &  n87 ;
  assign n680 = n208 | n234 ;
  assign n681 = n679 | n680 ;
  assign n682 = n678 | n681 ;
  assign n683 = n245 | n280 ;
  assign n684 = n430 | n683 ;
  assign n685 = ( n682 & ~n677 ) | ( n682 & n684 ) | ( ~n677 & n684 ) ;
  assign n686 = n677 | n685 ;
  assign n687 = ( n675 & ~n673 ) | ( n675 & n686 ) | ( ~n673 & n686 ) ;
  assign n688 = n673 | n687 ;
  assign n689 = ( n243 & ~n671 ) | ( n243 & n688 ) | ( ~n671 & n688 ) ;
  assign n690 = n671 | n689 ;
  assign n691 = n193 | n690 ;
  assign n692 = ( n436 & ~n410 ) | ( n436 & n691 ) | ( ~n410 & n691 ) ;
  assign n693 = n410 | n692 ;
  assign n694 = n670 | n693 ;
  assign n695 = ( n669 & ~n667 ) | ( n669 & n694 ) | ( ~n667 & n694 ) ;
  assign n696 = n667 | n695 ;
  assign n663 = n38 &  n103 ;
  assign n664 = n38 &  n116 ;
  assign n665 = n663 | n664 ;
  assign n697 = ( n696 & ~n212 ) | ( n696 & n665 ) | ( ~n212 & n665 ) ;
  assign n698 = n212 | n697 ;
  assign n699 = ( n662 & ~n698 ) | ( n662 & 1'b0 ) | ( ~n698 & 1'b0 ) ;
  assign n700 = ( n548 & n602 ) | ( n548 & n699 ) | ( n602 & n699 ) ;
  assign n701 = ~n602 & n700 ;
  assign n702 = ~n460 & n701 ;
  assign n703 = ~n233 & n624 ;
  assign n704 = ~n167 & n703 ;
  assign n705 = ~n541 & n704 ;
  assign n706 = ( n627 & ~n274 ) | ( n627 & n705 ) | ( ~n274 & n705 ) ;
  assign n707 = ~n627 & n706 ;
  assign n708 = ( n99 & ~n137 ) | ( n99 & n707 ) | ( ~n137 & n707 ) ;
  assign n709 = ~n99 & n708 ;
  assign n710 = ~n603 & n709 ;
  assign n711 = n59 &  n121 ;
  assign n712 = n68 &  n71 ;
  assign n713 = n711 | n712 ;
  assign n714 = n84 &  n121 ;
  assign n715 = n275 | n714 ;
  assign n716 = n52 | n241 ;
  assign n717 = n105 | n490 ;
  assign n718 = n51 &  n84 ;
  assign n719 = n188 | n718 ;
  assign n720 = n51 &  n116 ;
  assign n721 = n51 &  n98 ;
  assign n722 = ( n51 & ~n79 ) | ( n51 & 1'b0 ) | ( ~n79 & 1'b0 ) ;
  assign n723 = n207 | n722 ;
  assign n724 = ( n721 & ~n130 ) | ( n721 & n723 ) | ( ~n130 & n723 ) ;
  assign n725 = n130 | n724 ;
  assign n726 = ( n231 & ~n720 ) | ( n231 & n725 ) | ( ~n720 & n725 ) ;
  assign n727 = n720 | n726 ;
  assign n728 = n719 | n727 ;
  assign n729 = ( n717 & ~n716 ) | ( n717 & n728 ) | ( ~n716 & n728 ) ;
  assign n730 = n716 | n729 ;
  assign n731 = ( n218 & ~n418 ) | ( n218 & n730 ) | ( ~n418 & n730 ) ;
  assign n732 = n418 | n731 ;
  assign n733 = n457 | n732 ;
  assign n761 = n82 &  n121 ;
  assign n762 = n235 | n495 ;
  assign n763 = ( n258 & ~n761 ) | ( n258 & n762 ) | ( ~n761 & n762 ) ;
  assign n764 = n761 | n763 ;
  assign n765 = n57 &  n121 ;
  assign n766 = n168 | n273 ;
  assign n767 = n765 | n766 ;
  assign n768 = n191 | n767 ;
  assign n769 = n764 | n768 ;
  assign n734 = n84 &  n100 ;
  assign n735 = n94 &  n121 ;
  assign n736 = n222 | n424 ;
  assign n737 = n59 &  n100 ;
  assign n738 = n206 | n737 ;
  assign n739 = n284 | n738 ;
  assign n740 = n187 | n739 ;
  assign n741 = ( n736 & ~n735 ) | ( n736 & n740 ) | ( ~n735 & n740 ) ;
  assign n742 = n735 | n741 ;
  assign n743 = n271 | n742 ;
  assign n744 = n82 &  n100 ;
  assign n745 = n92 &  n100 ;
  assign n746 = n373 | n745 ;
  assign n747 = n123 | n349 ;
  assign n748 = n746 | n747 ;
  assign n749 = ( n272 & ~n122 ) | ( n272 & n748 ) | ( ~n122 & n748 ) ;
  assign n750 = n122 | n749 ;
  assign n751 = ( n372 & ~n350 ) | ( n372 & n750 ) | ( ~n350 & n750 ) ;
  assign n752 = n350 | n751 ;
  assign n753 = ( n101 & ~n744 ) | ( n101 & n752 ) | ( ~n744 & n752 ) ;
  assign n754 = n744 | n753 ;
  assign n755 = ( n743 & ~n407 ) | ( n743 & n754 ) | ( ~n407 & n754 ) ;
  assign n756 = n407 | n755 ;
  assign n757 = ( n232 & ~n734 ) | ( n232 & n756 ) | ( ~n734 & n756 ) ;
  assign n758 = n734 | n757 ;
  assign n759 = ( n197 & ~n758 ) | ( n197 & n279 ) | ( ~n758 & n279 ) ;
  assign n760 = ~n279 & n759 ;
  assign n770 = ( n733 & ~n769 ) | ( n733 & n760 ) | ( ~n769 & n760 ) ;
  assign n771 = ( n715 & ~n733 ) | ( n715 & n770 ) | ( ~n733 & n770 ) ;
  assign n772 = ( n771 & ~n715 ) | ( n771 & 1'b0 ) | ( ~n715 & 1'b0 ) ;
  assign n773 = ( n713 & ~n526 ) | ( n713 & n772 ) | ( ~n526 & n772 ) ;
  assign n774 = ~n713 & n773 ;
  assign n786 = ~n55 | ~n87 ;
  assign n788 = n71 &  n103 ;
  assign n789 = n60 &  n103 ;
  assign n790 = n259 | n475 ;
  assign n791 = n194 | n790 ;
  assign n792 = n48 &  n55 ;
  assign n793 = n55 &  n63 ;
  assign n794 = n125 | n253 ;
  assign n795 = n138 | n359 ;
  assign n796 = n55 &  n94 ;
  assign n797 = n55 &  n116 ;
  assign n798 = n257 | n797 ;
  assign n799 = n796 | n798 ;
  assign n800 = n55 &  n103 ;
  assign n801 = n333 | n800 ;
  assign n802 = n58 | n801 ;
  assign n803 = n799 | n802 ;
  assign n804 = ( n795 & ~n794 ) | ( n795 & n803 ) | ( ~n794 & n803 ) ;
  assign n805 = n794 | n804 ;
  assign n806 = ( n362 & ~n224 ) | ( n362 & n805 ) | ( ~n224 & n805 ) ;
  assign n807 = n224 | n806 ;
  assign n808 = ( n793 & ~n792 ) | ( n793 & n807 ) | ( ~n792 & n807 ) ;
  assign n809 = n792 | n808 ;
  assign n810 = n415 | n809 ;
  assign n811 = n345 | n408 ;
  assign n812 = n71 &  n84 ;
  assign n813 = ~n60 | ~n92 ;
  assign n814 = n60 &  n82 ;
  assign n815 = n157 | n374 ;
  assign n816 = ( n813 & n814 ) | ( n813 & n815 ) | ( n814 & n815 ) ;
  assign n817 = ( n813 & ~n816 ) | ( n813 & 1'b0 ) | ( ~n816 & 1'b0 ) ;
  assign n818 = ( n69 & ~n260 ) | ( n69 & n817 ) | ( ~n260 & n817 ) ;
  assign n819 = ~n69 & n818 ;
  assign n820 = ~n812 & n819 ;
  assign n821 = ( n811 & ~n195 ) | ( n811 & n820 ) | ( ~n195 & n820 ) ;
  assign n822 = ~n811 & n821 ;
  assign n823 = n128 | n150 ;
  assign n824 = n72 | n823 ;
  assign n825 = ( n822 & ~n824 ) | ( n822 & 1'b0 ) | ( ~n824 & 1'b0 ) ;
  assign n826 = ( n791 & ~n810 ) | ( n791 & n825 ) | ( ~n810 & n825 ) ;
  assign n827 = ~n791 & n826 ;
  assign n828 = ( n124 & ~n376 ) | ( n124 & n827 ) | ( ~n376 & n827 ) ;
  assign n829 = ~n124 & n828 ;
  assign n830 = ( n61 & ~n789 ) | ( n61 & n829 ) | ( ~n789 & n829 ) ;
  assign n831 = ~n61 & n830 ;
  assign n832 = ( n106 & ~n788 ) | ( n106 & n831 ) | ( ~n788 & n831 ) ;
  assign n833 = ~n106 & n832 ;
  assign n834 = ( n244 & ~n425 ) | ( n244 & n833 ) | ( ~n425 & n833 ) ;
  assign n835 = ~n244 & n834 ;
  assign n787 = n59 &  n71 ;
  assign n836 = ( n786 & ~n835 ) | ( n786 & n787 ) | ( ~n835 & n787 ) ;
  assign n837 = ( n786 & ~n836 ) | ( n786 & 1'b0 ) | ( ~n836 & 1'b0 ) ;
  assign n775 = n51 &  n119 ;
  assign n776 = n382 | n451 ;
  assign n777 = n132 | n776 ;
  assign n778 = n51 &  n68 ;
  assign n779 = n453 | n778 ;
  assign n780 = n777 | n779 ;
  assign n781 = ( n775 & ~n230 ) | ( n775 & n780 ) | ( ~n230 & n780 ) ;
  assign n782 = n230 | n781 ;
  assign n783 = ( n348 & ~n456 ) | ( n348 & n782 ) | ( ~n456 & n782 ) ;
  assign n784 = n456 | n783 ;
  assign n785 = n226 | n784 ;
  assign n838 = ( n774 & ~n837 ) | ( n774 & n785 ) | ( ~n837 & n785 ) ;
  assign n839 = ( n485 & ~n838 ) | ( n485 & n774 ) | ( ~n838 & n774 ) ;
  assign n840 = ~n485 & n839 ;
  assign n841 = ~n151 & n840 ;
  assign n842 = n148 | n617 ;
  assign n843 = n221 | n228 ;
  assign n844 = n576 | n843 ;
  assign n845 = ( n844 & ~n556 ) | ( n844 & n569 ) | ( ~n556 & n569 ) ;
  assign n846 = n556 | n845 ;
  assign n847 = ( n104 & ~n236 ) | ( n104 & n846 ) | ( ~n236 & n846 ) ;
  assign n848 = n236 | n847 ;
  assign n849 = ( n492 & ~n340 ) | ( n492 & n848 ) | ( ~n340 & n848 ) ;
  assign n850 = n340 | n849 ;
  assign n851 = n459 | n850 ;
  assign n852 = n452 | n476 ;
  assign n853 = ( n658 & ~n852 ) | ( n658 & 1'b0 ) | ( ~n852 & 1'b0 ) ;
  assign n854 = ( n573 & ~n851 ) | ( n573 & n853 ) | ( ~n851 & n853 ) ;
  assign n855 = ~n573 & n854 ;
  assign n856 = ( n842 & ~n163 ) | ( n842 & n855 ) | ( ~n163 & n855 ) ;
  assign n857 = ~n842 & n856 ;
  assign n858 = ~n300 & n857 ;
  assign n859 = ( n841 & ~n710 ) | ( n841 & n858 ) | ( ~n710 & n858 ) ;
  assign n860 = n710 &  n859 ;
  assign n861 = ( n604 & ~n553 ) | ( n604 & n860 ) | ( ~n553 & n860 ) ;
  assign n862 = ~n604 & n861 ;
  assign n863 = ~n403 &  n862 ;
  assign n864 = n88 | n787 ;
  assign n865 = n618 | n788 ;
  assign n866 = n49 | n628 ;
  assign n867 = ( n824 & ~n120 ) | ( n824 & n866 ) | ( ~n120 & n866 ) ;
  assign n868 = n120 | n867 ;
  assign n869 = ( n205 & ~n417 ) | ( n205 & n868 ) | ( ~n417 & n868 ) ;
  assign n870 = n417 | n869 ;
  assign n871 = ( n266 & ~n529 ) | ( n266 & n870 ) | ( ~n529 & n870 ) ;
  assign n872 = n529 | n871 ;
  assign n873 = ( n358 & ~n141 ) | ( n358 & n872 ) | ( ~n141 & n872 ) ;
  assign n874 = n141 | n873 ;
  assign n875 = ( n354 & ~n646 ) | ( n354 & 1'b0 ) | ( ~n646 & 1'b0 ) ;
  assign n876 = ( n875 & ~n338 ) | ( n875 & n376 ) | ( ~n338 & n376 ) ;
  assign n877 = ( n876 & ~n376 ) | ( n876 & 1'b0 ) | ( ~n376 & 1'b0 ) ;
  assign n878 = ( n554 & ~n643 ) | ( n554 & n877 ) | ( ~n643 & n877 ) ;
  assign n879 = ~n554 & n878 ;
  assign n880 = n61 | n91 ;
  assign n881 = ( n239 & ~n571 ) | ( n239 & n880 ) | ( ~n571 & n880 ) ;
  assign n882 = n571 | n881 ;
  assign n883 = n336 | n882 ;
  assign n884 = n93 | n356 ;
  assign n885 = n95 | n617 ;
  assign n886 = n139 | n789 ;
  assign n887 = n124 | n574 ;
  assign n888 = ~n117 & n484 ;
  assign n889 = n156 | n252 ;
  assign n890 = ( n888 & ~n889 ) | ( n888 & 1'b0 ) | ( ~n889 & 1'b0 ) ;
  assign n891 = ( n886 & ~n887 ) | ( n886 & n890 ) | ( ~n887 & n890 ) ;
  assign n892 = ~n886 & n891 ;
  assign n893 = ( n884 & ~n885 ) | ( n884 & n892 ) | ( ~n885 & n892 ) ;
  assign n894 = ( n244 & ~n884 ) | ( n244 & n893 ) | ( ~n884 & n893 ) ;
  assign n895 = ~n244 & n894 ;
  assign n896 = ( n270 & ~n194 ) | ( n270 & n895 ) | ( ~n194 & n895 ) ;
  assign n897 = ~n270 & n896 ;
  assign n898 = ( n160 & ~n549 ) | ( n160 & n897 ) | ( ~n549 & n897 ) ;
  assign n899 = ~n160 & n898 ;
  assign n900 = ( n899 & ~n334 ) | ( n899 & n454 ) | ( ~n334 & n454 ) ;
  assign n901 = ( n900 & ~n454 ) | ( n900 & 1'b0 ) | ( ~n454 & 1'b0 ) ;
  assign n902 = ( n77 & ~n353 ) | ( n77 & n901 ) | ( ~n353 & n901 ) ;
  assign n903 = ~n77 & n902 ;
  assign n904 = ~n166 & n903 ;
  assign n905 = n98 &  n131 ;
  assign n906 = n572 | n905 ;
  assign n907 = ( n213 & ~n276 ) | ( n213 & n906 ) | ( ~n276 & n906 ) ;
  assign n908 = n276 | n907 ;
  assign n909 = n94 &  n131 ;
  assign n910 = n165 | n909 ;
  assign n911 = n92 &  n131 ;
  assign n912 = n269 | n911 ;
  assign n913 = n910 | n912 ;
  assign n914 = ( n822 & ~n632 ) | ( n822 & n913 ) | ( ~n632 & n913 ) ;
  assign n915 = ( n908 & ~n913 ) | ( n908 & n914 ) | ( ~n913 & n914 ) ;
  assign n916 = ~n908 & n915 ;
  assign n917 = ( n883 & n904 ) | ( n883 & n916 ) | ( n904 & n916 ) ;
  assign n918 = ( n879 & ~n917 ) | ( n879 & n883 ) | ( ~n917 & n883 ) ;
  assign n919 = ( n879 & ~n918 ) | ( n879 & 1'b0 ) | ( ~n918 & 1'b0 ) ;
  assign n920 = ( n404 & ~n259 ) | ( n404 & n919 ) | ( ~n259 & n919 ) ;
  assign n921 = ~n404 & n920 ;
  assign n922 = ( n268 & ~n342 ) | ( n268 & n921 ) | ( ~n342 & n921 ) ;
  assign n923 = ~n268 & n922 ;
  assign n924 = ( n118 & ~n285 ) | ( n118 & n923 ) | ( ~n285 & n923 ) ;
  assign n925 = ~n118 & n924 ;
  assign n926 = ( n256 & ~n229 ) | ( n256 & n925 ) | ( ~n229 & n925 ) ;
  assign n927 = ~n256 & n926 ;
  assign n928 = ~n476 & n927 ;
  assign n929 = ~n475 & n786 ;
  assign n930 = ( n197 & ~n667 ) | ( n197 & 1'b0 ) | ( ~n667 & 1'b0 ) ;
  assign n931 = ~n212 & n930 ;
  assign n932 = ( n929 & n810 ) | ( n929 & n931 ) | ( n810 & n931 ) ;
  assign n933 = ( n619 & ~n810 ) | ( n619 & n932 ) | ( ~n810 & n932 ) ;
  assign n934 = ~n619 & n933 ;
  assign n935 = ( n928 & n874 ) | ( n928 & n934 ) | ( n874 & n934 ) ;
  assign n936 = ( n163 & ~n874 ) | ( n163 & n935 ) | ( ~n874 & n935 ) ;
  assign n937 = ~n163 & n936 ;
  assign n938 = ( n864 & ~n865 ) | ( n864 & n937 ) | ( ~n865 & n937 ) ;
  assign n939 = ~n864 & n938 ;
  assign n940 = ( n425 & ~n939 ) | ( n425 & n645 ) | ( ~n939 & n645 ) ;
  assign n941 = ( n645 & ~n940 ) | ( n645 & 1'b0 ) | ( ~n940 & 1'b0 ) ;
  assign n942 = ( n281 & ~n452 ) | ( n281 & n941 ) | ( ~n452 & n941 ) ;
  assign n943 = ~n281 & n942 ;
  assign n944 = ( n279 & ~n136 ) | ( n279 & n943 ) | ( ~n136 & n943 ) ;
  assign n945 = ~n279 & n944 ;
  assign n946 = ~n129 &  n945 ;
  assign n947 = n140 | n534 ;
  assign n998 = n255 | n526 ;
  assign n999 = n138 | n735 ;
  assign n1000 = ( n270 & ~n478 ) | ( n270 & n999 ) | ( ~n478 & n999 ) ;
  assign n1001 = n478 | n1000 ;
  assign n1002 = n715 | n793 ;
  assign n1003 = n571 | n765 ;
  assign n1004 = n224 | n665 ;
  assign n1005 = n1003 | n1004 ;
  assign n1006 = ( n434 & ~n761 ) | ( n434 & n1005 ) | ( ~n761 & n1005 ) ;
  assign n1007 = n761 | n1006 ;
  assign n1008 = n123 | n1007 ;
  assign n1009 = n549 | n797 ;
  assign n1010 = n120 | n712 ;
  assign n1011 = ( n1009 & ~n232 ) | ( n1009 & n1010 ) | ( ~n232 & n1010 ) ;
  assign n1012 = n232 | n1011 ;
  assign n1013 = ( n88 & ~n734 ) | ( n88 & n1012 ) | ( ~n734 & n1012 ) ;
  assign n1014 = n734 | n1013 ;
  assign n1015 = n49 | n910 ;
  assign n1016 = ( n135 & ~n476 ) | ( n135 & n1015 ) | ( ~n476 & n1015 ) ;
  assign n1017 = n476 | n1016 ;
  assign n1018 = ( n1014 & ~n1008 ) | ( n1014 & n1017 ) | ( ~n1008 & n1017 ) ;
  assign n1019 = ( n1008 & ~n1002 ) | ( n1008 & n1018 ) | ( ~n1002 & n1018 ) ;
  assign n1020 = n1002 | n1019 ;
  assign n1021 = ( n1001 & ~n362 ) | ( n1001 & n1020 ) | ( ~n362 & n1020 ) ;
  assign n1022 = n362 | n1021 ;
  assign n1023 = ( n206 & ~n257 ) | ( n206 & n1022 ) | ( ~n257 & n1022 ) ;
  assign n1024 = n257 | n1023 ;
  assign n1025 = ( n239 & ~n252 ) | ( n239 & n1024 ) | ( ~n252 & n1024 ) ;
  assign n1026 = n252 | n1025 ;
  assign n1027 = ( n39 & ~n141 ) | ( n39 & n1026 ) | ( ~n141 & n1026 ) ;
  assign n1028 = n141 | n1027 ;
  assign n1029 = n89 | n299 ;
  assign n1030 = ( n343 & ~n1029 ) | ( n343 & 1'b0 ) | ( ~n1029 & 1'b0 ) ;
  assign n1031 = ( n851 & ~n1028 ) | ( n851 & n1030 ) | ( ~n1028 & n1030 ) ;
  assign n1032 = ( n998 & ~n851 ) | ( n998 & n1031 ) | ( ~n851 & n1031 ) ;
  assign n1033 = ~n998 & n1032 ;
  assign n990 = n74 | n424 ;
  assign n991 = n242 | n990 ;
  assign n992 = ( n190 & ~n276 ) | ( n190 & n991 ) | ( ~n276 & n991 ) ;
  assign n993 = n276 | n992 ;
  assign n994 = ( n631 & ~n334 ) | ( n631 & n993 ) | ( ~n334 & n993 ) ;
  assign n995 = n334 | n994 ;
  assign n996 = ( n117 & ~n77 ) | ( n117 & n995 ) | ( ~n77 & n995 ) ;
  assign n997 = n77 | n996 ;
  assign n1034 = ( n929 & ~n1033 ) | ( n929 & n997 ) | ( ~n1033 & n997 ) ;
  assign n1035 = ( n929 & ~n1034 ) | ( n929 & 1'b0 ) | ( ~n1034 & 1'b0 ) ;
  assign n949 = ( n493 & ~n122 ) | ( n493 & n802 ) | ( ~n122 & n802 ) ;
  assign n950 = n122 | n949 ;
  assign n951 = ( n529 & ~n404 ) | ( n529 & n950 ) | ( ~n404 & n950 ) ;
  assign n952 = n404 | n951 ;
  assign n953 = n136 | n273 ;
  assign n954 = n125 | n953 ;
  assign n955 = ( n258 & ~n235 ) | ( n258 & n954 ) | ( ~n235 & n954 ) ;
  assign n956 = n235 | n955 ;
  assign n957 = ( n193 & ~n350 ) | ( n193 & n956 ) | ( ~n350 & n956 ) ;
  assign n958 = n350 | n957 ;
  assign n959 = n618 | n958 ;
  assign n974 = n222 | n359 ;
  assign n975 = n349 | n410 ;
  assign n976 = n974 | n975 ;
  assign n960 = n91 | n911 ;
  assign n961 = n351 | n792 ;
  assign n962 = n269 | n494 ;
  assign n963 = n139 | n962 ;
  assign n964 = ( n961 & ~n272 ) | ( n961 & n963 ) | ( ~n272 & n963 ) ;
  assign n965 = n272 | n964 ;
  assign n966 = ( n711 & ~n191 ) | ( n711 & n965 ) | ( ~n191 & n965 ) ;
  assign n967 = n191 | n966 ;
  assign n968 = ( n229 & ~n432 ) | ( n229 & n967 ) | ( ~n432 & n967 ) ;
  assign n969 = n432 | n968 ;
  assign n970 = n960 | n969 ;
  assign n971 = ( n970 & ~n124 ) | ( n970 & n796 ) | ( ~n124 & n796 ) ;
  assign n972 = n124 | n971 ;
  assign n973 = n431 | n972 ;
  assign n977 = ( n976 & ~n959 ) | ( n976 & n973 ) | ( ~n959 & n973 ) ;
  assign n978 = n959 | n977 ;
  assign n979 = ( n952 & ~n668 ) | ( n952 & n978 ) | ( ~n668 & n978 ) ;
  assign n980 = n668 | n979 ;
  assign n948 = n129 | n670 ;
  assign n981 = ( n645 & n980 ) | ( n645 & n948 ) | ( n980 & n948 ) ;
  assign n982 = ( n645 & ~n981 ) | ( n645 & 1'b0 ) | ( ~n981 & 1'b0 ) ;
  assign n983 = ( n906 & ~n455 ) | ( n906 & n982 ) | ( ~n455 & n982 ) ;
  assign n984 = ~n906 & n983 ;
  assign n985 = ( n415 & ~n253 ) | ( n415 & n984 ) | ( ~n253 & n984 ) ;
  assign n986 = ~n415 & n985 ;
  assign n987 = ( n284 & ~n168 ) | ( n284 & n986 ) | ( ~n168 & n986 ) ;
  assign n988 = ~n284 & n987 ;
  assign n989 = ~n268 & n988 ;
  assign n1036 = ( n555 & ~n1035 ) | ( n555 & n989 ) | ( ~n1035 & n989 ) ;
  assign n1037 = ( n947 & ~n1036 ) | ( n947 & n989 ) | ( ~n1036 & n989 ) ;
  assign n1038 = ~n947 & n1037 ;
  assign n1039 = ( n106 & ~n407 ) | ( n106 & n1038 ) | ( ~n407 & n1038 ) ;
  assign n1040 = ~n106 & n1039 ;
  assign n1041 = ( n356 & ~n372 ) | ( n356 & n1040 ) | ( ~n372 & n1040 ) ;
  assign n1042 = ~n356 & n1041 ;
  assign n1043 = ~n196 & n1042 ;
  assign n1044 = n404 | n643 ;
  assign n1045 = n618 | n722 ;
  assign n1046 = n162 | n205 ;
  assign n1047 = n256 | n909 ;
  assign n1048 = n231 | n718 ;
  assign n1049 = n406 | n1048 ;
  assign n1050 = n490 | n814 ;
  assign n1051 = n135 | n1050 ;
  assign n1052 = ( n1049 & ~n1047 ) | ( n1049 & n1051 ) | ( ~n1047 & n1051 ) ;
  assign n1053 = n1047 | n1052 ;
  assign n1054 = ( n789 & ~n376 ) | ( n789 & n1053 ) | ( ~n376 & n1053 ) ;
  assign n1055 = n376 | n1054 ;
  assign n1056 = ( n130 & ~n558 ) | ( n130 & n1055 ) | ( ~n558 & n1055 ) ;
  assign n1057 = n558 | n1056 ;
  assign n1058 = ( n529 & ~n574 ) | ( n529 & n1057 ) | ( ~n574 & n1057 ) ;
  assign n1059 = n574 | n1058 ;
  assign n1060 = n299 | n679 ;
  assign n1061 = n429 | n664 ;
  assign n1062 = n271 | n674 ;
  assign n1071 = n253 | n411 ;
  assign n1072 = n678 | n800 ;
  assign n1073 = ( n813 & ~n1072 ) | ( n813 & 1'b0 ) | ( ~n1072 & 1'b0 ) ;
  assign n1074 = n141 | n604 ;
  assign n1075 = n83 | n1074 ;
  assign n1076 = n62 | n906 ;
  assign n1077 = ( n1073 & n1075 ) | ( n1073 & n1076 ) | ( n1075 & n1076 ) ;
  assign n1078 = ( n1073 & ~n1077 ) | ( n1073 & 1'b0 ) | ( ~n1077 & 1'b0 ) ;
  assign n1079 = ( n1071 & ~n576 ) | ( n1071 & n1078 ) | ( ~n576 & n1078 ) ;
  assign n1080 = ~n1071 & n1079 ;
  assign n1063 = n267 | n714 ;
  assign n1064 = n69 | n540 ;
  assign n1065 = n1063 | n1064 ;
  assign n1066 = ( n795 & ~n195 ) | ( n795 & n1065 ) | ( ~n195 & n1065 ) ;
  assign n1067 = n195 | n1066 ;
  assign n1068 = ( n188 & n1067 ) | ( n188 & n343 ) | ( n1067 & n343 ) ;
  assign n1069 = ( n343 & ~n1068 ) | ( n343 & 1'b0 ) | ( ~n1068 & 1'b0 ) ;
  assign n1070 = ~n137 & n1069 ;
  assign n1081 = ( n764 & ~n1080 ) | ( n764 & n1070 ) | ( ~n1080 & n1070 ) ;
  assign n1082 = ( n1062 & ~n1081 ) | ( n1062 & n1070 ) | ( ~n1081 & n1070 ) ;
  assign n1083 = ~n1062 & n1082 ;
  assign n1084 = ( n1060 & ~n1061 ) | ( n1060 & n1083 ) | ( ~n1061 & n1083 ) ;
  assign n1085 = ~n1060 & n1084 ;
  assign n1086 = ( n273 & n645 ) | ( n273 & n1085 ) | ( n645 & n1085 ) ;
  assign n1087 = ~n273 & n1086 ;
  assign n1088 = ( n744 & ~n101 ) | ( n744 & n1087 ) | ( ~n101 & n1087 ) ;
  assign n1089 = ~n744 & n1088 ;
  assign n1090 = ( n165 & ~n187 ) | ( n165 & n1089 ) | ( ~n187 & n1089 ) ;
  assign n1091 = ~n165 & n1090 ;
  assign n1092 = ~n549 & n1091 ;
  assign n1093 = n243 | n737 ;
  assign n1094 = n260 | n1010 ;
  assign n1095 = ( n191 & ~n275 ) | ( n191 & n1094 ) | ( ~n275 & n1094 ) ;
  assign n1096 = n275 | n1095 ;
  assign n1097 = n136 | n745 ;
  assign n1098 = n39 | n1097 ;
  assign n1099 = ( n415 & ~n374 ) | ( n415 & n1098 ) | ( ~n374 & n1098 ) ;
  assign n1100 = n374 | n1099 ;
  assign n1101 = ( n569 & ~n216 ) | ( n569 & n1100 ) | ( ~n216 & n1100 ) ;
  assign n1102 = n216 | n1101 ;
  assign n1103 = ( n384 & n1102 ) | ( n384 & n623 ) | ( n1102 & n623 ) ;
  assign n1104 = ( n623 & ~n1103 ) | ( n623 & 1'b0 ) | ( ~n1103 & 1'b0 ) ;
  assign n1105 = ( n197 & ~n345 ) | ( n197 & 1'b0 ) | ( ~n345 & 1'b0 ) ;
  assign n1106 = ~n213 & n1105 ;
  assign n1107 = n91 | n245 ;
  assign n1108 = n947 | n1107 ;
  assign n1109 = n797 | n1108 ;
  assign n1110 = n336 | n457 ;
  assign n1111 = n1003 | n1110 ;
  assign n1112 = ( n1106 & n1109 ) | ( n1106 & n1111 ) | ( n1109 & n1111 ) ;
  assign n1113 = ( n1106 & ~n1112 ) | ( n1106 & 1'b0 ) | ( ~n1112 & 1'b0 ) ;
  assign n1114 = ( n1096 & n1104 ) | ( n1096 & n1113 ) | ( n1104 & n1113 ) ;
  assign n1115 = ( n1093 & ~n1096 ) | ( n1093 & n1114 ) | ( ~n1096 & n1114 ) ;
  assign n1116 = ( n1115 & ~n1093 ) | ( n1115 & 1'b0 ) | ( ~n1093 & 1'b0 ) ;
  assign n1117 = ( n280 & ~n259 ) | ( n280 & n1116 ) | ( ~n259 & n1116 ) ;
  assign n1118 = ~n280 & n1117 ;
  assign n1119 = ( n99 & ~n373 ) | ( n99 & n1118 ) | ( ~n373 & n1118 ) ;
  assign n1120 = ~n99 & n1119 ;
  assign n1121 = ( n1120 & ~n155 ) | ( n1120 & n663 ) | ( ~n155 & n663 ) ;
  assign n1122 = ( n1121 & ~n663 ) | ( n1121 & 1'b0 ) | ( ~n663 & 1'b0 ) ;
  assign n1123 = n353 | n568 ;
  assign n1124 = n647 | n1123 ;
  assign n1125 = ( n342 & ~n300 ) | ( n342 & n1124 ) | ( ~n300 & n1124 ) ;
  assign n1126 = n300 | n1125 ;
  assign n1127 = ( n156 & n354 ) | ( n156 & n1126 ) | ( n354 & n1126 ) ;
  assign n1128 = ( n354 & ~n1127 ) | ( n354 & 1'b0 ) | ( ~n1127 & 1'b0 ) ;
  assign n1129 = ~n432 & n1128 ;
  assign n1130 = n459 | n560 ;
  assign n1131 = n241 | n948 ;
  assign n1132 = ( n240 & ~n405 ) | ( n240 & n1131 ) | ( ~n405 & n1131 ) ;
  assign n1133 = n405 | n1132 ;
  assign n1134 = ( n1130 & ~n533 ) | ( n1130 & n1133 ) | ( ~n533 & n1133 ) ;
  assign n1135 = ( n533 & n1129 ) | ( n533 & n1134 ) | ( n1129 & n1134 ) ;
  assign n1136 = ( n1129 & ~n1135 ) | ( n1129 & 1'b0 ) | ( ~n1135 & 1'b0 ) ;
  assign n1137 = ( n1122 & ~n1092 ) | ( n1122 & n1136 ) | ( ~n1092 & n1136 ) ;
  assign n1138 = ( n1092 & ~n929 ) | ( n1092 & n1137 ) | ( ~n929 & n1137 ) ;
  assign n1139 = n929 &  n1138 ;
  assign n1140 = ( n1046 & ~n1059 ) | ( n1046 & n1139 ) | ( ~n1059 & n1139 ) ;
  assign n1141 = ~n1046 & n1140 ;
  assign n1142 = ( n1044 & ~n1045 ) | ( n1044 & n1141 ) | ( ~n1045 & n1141 ) ;
  assign n1143 = ( n1142 & ~n1044 ) | ( n1142 & 1'b0 ) | ( ~n1044 & 1'b0 ) ;
  assign n1144 = ( n339 & ~n912 ) | ( n339 & n1143 ) | ( ~n912 & n1143 ) ;
  assign n1145 = ~n339 & n1144 ;
  assign n1146 = ( n106 & ~n270 ) | ( n106 & n1145 ) | ( ~n270 & n1145 ) ;
  assign n1147 = ~n106 & n1146 ;
  assign n1148 = ( n236 & ~n478 ) | ( n236 & n1147 ) | ( ~n478 & n1147 ) ;
  assign n1149 = ~n236 & n1148 ;
  assign n1150 = ( n285 & ~n88 ) | ( n285 & n1149 ) | ( ~n88 & n1149 ) ;
  assign n1151 = ~n285 &  n1150 ;
  assign n1152 = n275 | n735 ;
  assign n1153 = n454 | n475 ;
  assign n1154 = ( n168 & n484 ) | ( n168 & n778 ) | ( n484 & n778 ) ;
  assign n1155 = ( n484 & ~n1154 ) | ( n484 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n1156 = ( n493 & ~n1153 ) | ( n493 & n1155 ) | ( ~n1153 & n1155 ) ;
  assign n1157 = ~n493 & n1156 ;
  assign n1158 = ( n161 & ~n224 ) | ( n161 & n1157 ) | ( ~n224 & n1157 ) ;
  assign n1159 = ~n161 & n1158 ;
  assign n1160 = ( n561 & ~n1159 ) | ( n561 & n644 ) | ( ~n1159 & n644 ) ;
  assign n1161 = ( n644 & ~n1160 ) | ( n644 & 1'b0 ) | ( ~n1160 & 1'b0 ) ;
  assign n1162 = ( n276 & ~n160 ) | ( n276 & n1161 ) | ( ~n160 & n1161 ) ;
  assign n1163 = ~n276 & n1162 ;
  assign n1164 = ( n244 & ~n376 ) | ( n244 & n525 ) | ( ~n376 & n525 ) ;
  assign n1165 = ~n244 & n1164 ;
  assign n1166 = ~n333 & n1165 ;
  assign n1167 = ~n433 & n1166 ;
  assign n1168 = ~n217 & n624 ;
  assign n1169 = n165 | n190 ;
  assign n1170 = ( n1167 & ~n1168 ) | ( n1167 & n1169 ) | ( ~n1168 & n1169 ) ;
  assign n1171 = ( n1167 & ~n1170 ) | ( n1167 & 1'b0 ) | ( ~n1170 & 1'b0 ) ;
  assign n1172 = ( n842 & n1163 ) | ( n842 & n1171 ) | ( n1163 & n1171 ) ;
  assign n1173 = ~n842 & n1172 ;
  assign n1174 = ( n1152 & ~n245 ) | ( n1152 & n1173 ) | ( ~n245 & n1173 ) ;
  assign n1175 = ( n786 & ~n1174 ) | ( n786 & n1152 ) | ( ~n1174 & n1152 ) ;
  assign n1176 = ( n786 & ~n1175 ) | ( n786 & 1'b0 ) | ( ~n1175 & 1'b0 ) ;
  assign n1177 = ( n122 & ~n796 ) | ( n122 & n1176 ) | ( ~n796 & n1176 ) ;
  assign n1178 = ~n122 & n1177 ;
  assign n1179 = ( n1178 & ~n284 ) | ( n1178 & n745 ) | ( ~n284 & n745 ) ;
  assign n1180 = ( n1179 & ~n745 ) | ( n1179 & 1'b0 ) | ( ~n745 & 1'b0 ) ;
  assign n1181 = ( n299 & ~n558 ) | ( n299 & n1180 ) | ( ~n558 & n1180 ) ;
  assign n1182 = ~n299 & n1181 ;
  assign n1183 = ~n417 & n1182 ;
  assign n1184 = n206 | n720 ;
  assign n1185 = n256 | n671 ;
  assign n1186 = n814 | n911 ;
  assign n1187 = n140 | n1186 ;
  assign n1192 = n405 | n549 ;
  assign n1193 = ( n235 & ~n373 ) | ( n235 & n1192 ) | ( ~n373 & n1192 ) ;
  assign n1194 = n373 | n1193 ;
  assign n1195 = n300 | n1194 ;
  assign n1188 = n266 | n679 ;
  assign n1189 = ( n571 & ~n213 ) | ( n571 & n1188 ) | ( ~n213 & n1188 ) ;
  assign n1190 = n213 | n1189 ;
  assign n1191 = n476 | n1190 ;
  assign n1196 = n156 | n744 ;
  assign n1197 = ( n1195 & ~n1191 ) | ( n1195 & n1196 ) | ( ~n1191 & n1196 ) ;
  assign n1198 = ( n1197 & ~n1187 ) | ( n1197 & n1191 ) | ( ~n1187 & n1191 ) ;
  assign n1199 = n1187 | n1198 ;
  assign n1200 = ( n1185 & ~n1184 ) | ( n1185 & n1199 ) | ( ~n1184 & n1199 ) ;
  assign n1201 = ( n1184 & ~n886 ) | ( n1184 & n1200 ) | ( ~n886 & n1200 ) ;
  assign n1202 = n886 | n1201 ;
  assign n1203 = ( n713 & ~n277 ) | ( n713 & n1202 ) | ( ~n277 & n1202 ) ;
  assign n1204 = n277 | n1203 ;
  assign n1205 = ( n618 & ~n105 ) | ( n618 & n1204 ) | ( ~n105 & n1204 ) ;
  assign n1206 = n105 | n1205 ;
  assign n1207 = n374 | n909 ;
  assign n1208 = n492 | n559 ;
  assign n1209 = n410 | n1208 ;
  assign n1210 = ( n189 & ~n1207 ) | ( n189 & n1209 ) | ( ~n1207 & n1209 ) ;
  assign n1211 = n1207 | n1210 ;
  assign n1212 = ( n272 & ~n408 ) | ( n272 & n1211 ) | ( ~n408 & n1211 ) ;
  assign n1213 = n408 | n1212 ;
  assign n1214 = ( n232 & ~n737 ) | ( n232 & n1213 ) | ( ~n737 & n1213 ) ;
  assign n1215 = n737 | n1214 ;
  assign n1216 = ( n260 & ~n418 ) | ( n260 & n269 ) | ( ~n418 & n269 ) ;
  assign n1217 = ( n418 & ~n62 ) | ( n418 & n1216 ) | ( ~n62 & n1216 ) ;
  assign n1218 = n62 | n1217 ;
  assign n1219 = ( n192 & ~n338 ) | ( n192 & n1218 ) | ( ~n338 & n1218 ) ;
  assign n1220 = n338 | n1219 ;
  assign n1221 = n49 | n1220 ;
  assign n1222 = n234 | n258 ;
  assign n1223 = ( n793 & ~n568 ) | ( n793 & n1222 ) | ( ~n568 & n1222 ) ;
  assign n1224 = n568 | n1223 ;
  assign n1225 = n672 | n792 ;
  assign n1226 = ( n149 & ~n271 ) | ( n149 & n1225 ) | ( ~n271 & n1225 ) ;
  assign n1227 = n271 | n1226 ;
  assign n1228 = n233 | n274 ;
  assign n1229 = ( n270 & ~n905 ) | ( n270 & n1228 ) | ( ~n905 & n1228 ) ;
  assign n1230 = n905 | n1229 ;
  assign n1231 = n404 | n1230 ;
  assign n1232 = n342 | n540 ;
  assign n1233 = n334 | n425 ;
  assign n1234 = ( n634 & ~n1233 ) | ( n634 & n669 ) | ( ~n1233 & n669 ) ;
  assign n1235 = n1233 | n1234 ;
  assign n1236 = ( n1232 & ~n1231 ) | ( n1232 & n1235 ) | ( ~n1231 & n1235 ) ;
  assign n1237 = ( n1231 & ~n106 ) | ( n1231 & n1236 ) | ( ~n106 & n1236 ) ;
  assign n1238 = n106 | n1237 ;
  assign n1239 = ( n1238 & ~n136 ) | ( n1238 & n569 ) | ( ~n136 & n569 ) ;
  assign n1240 = n136 | n1239 ;
  assign n1241 = ( n129 & ~n556 ) | ( n129 & n1240 ) | ( ~n556 & n1240 ) ;
  assign n1242 = n556 | n1241 ;
  assign n1243 = n663 | n1242 ;
  assign n1244 = n194 | n229 ;
  assign n1245 = n120 | n431 ;
  assign n1246 = n1244 | n1245 ;
  assign n1247 = ( n354 & n812 ) | ( n354 & n1246 ) | ( n812 & n1246 ) ;
  assign n1248 = ( n354 & ~n1247 ) | ( n354 & 1'b0 ) | ( ~n1247 & 1'b0 ) ;
  assign n1249 = ~n166 & n1248 ;
  assign n1250 = ( n1227 & ~n1243 ) | ( n1227 & n1249 ) | ( ~n1243 & n1249 ) ;
  assign n1251 = ( n1224 & ~n1227 ) | ( n1224 & n1250 ) | ( ~n1227 & n1250 ) ;
  assign n1252 = ~n1224 & n1251 ;
  assign n1253 = ~n1221 & n1252 ;
  assign n1254 = ( n1206 & ~n1215 ) | ( n1206 & n1253 ) | ( ~n1215 & n1253 ) ;
  assign n1255 = ( n1206 & ~n1254 ) | ( n1206 & n1183 ) | ( ~n1254 & n1183 ) ;
  assign n1256 = ( n1183 & ~n1255 ) | ( n1183 & 1'b0 ) | ( ~n1255 & 1'b0 ) ;
  assign n1257 = ( n280 & ~n157 ) | ( n280 & n1256 ) | ( ~n157 & n1256 ) ;
  assign n1258 = ~n280 & n1257 ;
  assign n1259 = ( n1258 & ~n52 ) | ( n1258 & n800 ) | ( ~n52 & n800 ) ;
  assign n1260 = ( n1259 & ~n800 ) | ( n1259 & 1'b0 ) | ( ~n800 & 1'b0 ) ;
  assign n1261 = ( n101 & ~n721 ) | ( n101 & n1260 ) | ( ~n721 & n1260 ) ;
  assign n1262 = ~n101 & n1261 ;
  assign n1263 = ( n478 & ~n384 ) | ( n478 & n1262 ) | ( ~n384 & n1262 ) ;
  assign n1264 = ~n478 & n1263 ;
  assign n1265 = ( n459 & ~n643 ) | ( n459 & n1264 ) | ( ~n643 & n1264 ) ;
  assign n1266 = ~n459 & n1265 ;
  assign n1267 = ~n1266 |  n358 ;
  assign n1268 = n376 | n404 ;
  assign n1269 = n299 | n338 ;
  assign n1270 = n253 | n1269 ;
  assign n1271 = n224 | n266 ;
  assign n1272 = n463 | n1271 ;
  assign n1273 = ( n52 & ~n460 ) | ( n52 & n1272 ) | ( ~n460 & n1272 ) ;
  assign n1274 = n460 | n1273 ;
  assign n1275 = ( n452 & ~n618 ) | ( n452 & n1274 ) | ( ~n618 & n1274 ) ;
  assign n1276 = n618 | n1275 ;
  assign n1277 = n628 | n1276 ;
  assign n1278 = n417 | n559 ;
  assign n1279 = ~n775 & n786 ;
  assign n1283 = n157 | n168 ;
  assign n1280 = n679 | n721 ;
  assign n1281 = n214 | n1280 ;
  assign n1282 = n526 | n1281 ;
  assign n1284 = n453 | n603 ;
  assign n1285 = n409 | n814 ;
  assign n1286 = n631 | n1285 ;
  assign n1287 = ( n258 & ~n275 ) | ( n258 & n569 ) | ( ~n275 & n569 ) ;
  assign n1288 = n275 | n1287 ;
  assign n1289 = n382 | n720 ;
  assign n1290 = n1288 | n1289 ;
  assign n1291 = ( n1286 & ~n975 ) | ( n1286 & n1290 ) | ( ~n975 & n1290 ) ;
  assign n1292 = n975 | n1291 ;
  assign n1293 = ( n1284 & ~n462 ) | ( n1284 & n1292 ) | ( ~n462 & n1292 ) ;
  assign n1294 = n462 | n1293 ;
  assign n1295 = ( n1283 & ~n1282 ) | ( n1283 & n1294 ) | ( ~n1282 & n1294 ) ;
  assign n1296 = ( n1279 & n1295 ) | ( n1279 & n1282 ) | ( n1295 & n1282 ) ;
  assign n1297 = ( n1279 & ~n1296 ) | ( n1279 & 1'b0 ) | ( ~n1296 & 1'b0 ) ;
  assign n1298 = ( n1277 & ~n1278 ) | ( n1277 & n1297 ) | ( ~n1278 & n1297 ) ;
  assign n1299 = ( n163 & ~n1277 ) | ( n163 & n1298 ) | ( ~n1277 & n1298 ) ;
  assign n1300 = ~n163 & n1299 ;
  assign n1301 = ( n150 & ~n477 ) | ( n150 & n1300 ) | ( ~n477 & n1300 ) ;
  assign n1302 = ~n150 & n1301 ;
  assign n1303 = ( n644 & ~n1302 ) | ( n644 & n909 ) | ( ~n1302 & n909 ) ;
  assign n1304 = ( n644 & ~n1303 ) | ( n644 & 1'b0 ) | ( ~n1303 & 1'b0 ) ;
  assign n1305 = n148 | n722 ;
  assign n1306 = n166 | n905 ;
  assign n1307 = ( n257 & ~n1306 ) | ( n257 & n573 ) | ( ~n1306 & n573 ) ;
  assign n1308 = n1306 | n1307 ;
  assign n1309 = ( n1308 & ~n457 ) | ( n1308 & n714 ) | ( ~n457 & n714 ) ;
  assign n1310 = n457 | n1309 ;
  assign n1311 = ( n237 & ~n74 ) | ( n237 & n1310 ) | ( ~n74 & n1310 ) ;
  assign n1312 = n74 | n1311 ;
  assign n1313 = ( n149 & ~n574 ) | ( n149 & n1312 ) | ( ~n574 & n1312 ) ;
  assign n1314 = n574 | n1313 ;
  assign n1315 = ( n334 & ~n228 ) | ( n334 & n1314 ) | ( ~n228 & n1314 ) ;
  assign n1316 = n228 | n1315 ;
  assign n1317 = n744 | n788 ;
  assign n1318 = n974 | n1317 ;
  assign n1319 = ( n647 & ~n672 ) | ( n647 & n1318 ) | ( ~n672 & n1318 ) ;
  assign n1320 = n672 | n1319 ;
  assign n1321 = ( n270 & ~n671 ) | ( n270 & n1320 ) | ( ~n671 & n1320 ) ;
  assign n1322 = n671 | n1321 ;
  assign n1323 = ( n627 & ~n165 ) | ( n627 & n1322 ) | ( ~n165 & n1322 ) ;
  assign n1324 = n165 | n1323 ;
  assign n1325 = n160 | n531 ;
  assign n1326 = n118 | n418 ;
  assign n1327 = n151 | n347 ;
  assign n1328 = n286 | n1327 ;
  assign n1329 = ( n1326 & ~n1192 ) | ( n1326 & n1328 ) | ( ~n1192 & n1328 ) ;
  assign n1330 = n1192 | n1329 ;
  assign n1331 = ( n1325 & ~n1324 ) | ( n1325 & n1330 ) | ( ~n1324 & n1330 ) ;
  assign n1332 = ( n1324 & ~n1316 ) | ( n1324 & n1331 ) | ( ~n1316 & n1331 ) ;
  assign n1333 = n1316 | n1332 ;
  assign n1334 = ( n346 & ~n1093 ) | ( n346 & n1333 ) | ( ~n1093 & n1333 ) ;
  assign n1335 = n1093 | n1334 ;
  assign n1336 = ( n259 & ~n65 ) | ( n259 & n1335 ) | ( ~n65 & n1335 ) ;
  assign n1337 = n65 | n1336 ;
  assign n1338 = ( n711 & ~n1305 ) | ( n711 & n1337 ) | ( ~n1305 & n1337 ) ;
  assign n1339 = ( n1305 & ~n332 ) | ( n1305 & n1338 ) | ( ~n332 & n1338 ) ;
  assign n1340 = n332 | n1339 ;
  assign n1341 = n231 | n792 ;
  assign n1342 = n348 | n1341 ;
  assign n1344 = n665 | n718 ;
  assign n1345 = n268 | n1344 ;
  assign n1343 = ( n354 & ~n789 ) | ( n354 & 1'b0 ) | ( ~n789 & 1'b0 ) ;
  assign n1346 = ( n1342 & ~n1345 ) | ( n1342 & n1343 ) | ( ~n1345 & n1343 ) ;
  assign n1347 = ( n1153 & ~n1342 ) | ( n1153 & n1346 ) | ( ~n1342 & n1346 ) ;
  assign n1348 = ( n1347 & ~n1153 ) | ( n1347 & 1'b0 ) | ( ~n1153 & 1'b0 ) ;
  assign n1349 = ( n194 & ~n1340 ) | ( n194 & n1348 ) | ( ~n1340 & n1348 ) ;
  assign n1350 = ~n194 & n1349 ;
  assign n1351 = ( n205 & ~n540 ) | ( n205 & n1350 ) | ( ~n540 & n1350 ) ;
  assign n1352 = ~n205 & n1351 ;
  assign n1353 = ( n106 & ~n373 ) | ( n106 & n216 ) | ( ~n373 & n216 ) ;
  assign n1354 = n373 | n1353 ;
  assign n1355 = n279 | n1354 ;
  assign n1356 = n340 | n911 ;
  assign n1357 = n93 | n350 ;
  assign n1358 = n273 | n558 ;
  assign n1359 = n129 | n1358 ;
  assign n1360 = n91 | n230 ;
  assign n1361 = n190 | n1360 ;
  assign n1362 = n225 | n1361 ;
  assign n1363 = n213 | n255 ;
  assign n1364 = ( n1362 & ~n1359 ) | ( n1362 & n1363 ) | ( ~n1359 & n1363 ) ;
  assign n1365 = ( n1359 & ~n1357 ) | ( n1359 & n1364 ) | ( ~n1357 & n1364 ) ;
  assign n1366 = n1357 | n1365 ;
  assign n1367 = ( n1356 & ~n1355 ) | ( n1356 & n1366 ) | ( ~n1355 & n1366 ) ;
  assign n1368 = n1355 | n1367 ;
  assign n1369 = ( n1304 & ~n1352 ) | ( n1304 & n1368 ) | ( ~n1352 & n1368 ) ;
  assign n1370 = ( n1304 & ~n1369 ) | ( n1304 & 1'b0 ) | ( ~n1369 & 1'b0 ) ;
  assign n1371 = ( n1270 & ~n147 ) | ( n1270 & n1370 ) | ( ~n147 & n1370 ) ;
  assign n1372 = ~n1270 & n1371 ;
  assign n1373 = ( n677 & ~n1062 ) | ( n677 & n1372 ) | ( ~n1062 & n1372 ) ;
  assign n1374 = ~n677 & n1373 ;
  assign n1375 = ( n105 & ~n1268 ) | ( n105 & n1374 ) | ( ~n1268 & n1374 ) ;
  assign n1376 = ~n105 & n1375 ;
  assign n1377 = ( n524 & ~n1376 ) | ( n524 & n630 ) | ( ~n1376 & n630 ) ;
  assign n1378 = ( n524 & ~n1377 ) | ( n524 & 1'b0 ) | ( ~n1377 & 1'b0 ) ;
  assign n1381 = n300 | n332 ;
  assign n1382 = n122 | n1381 ;
  assign n1383 = ( n192 & ~n151 ) | ( n192 & n1382 ) | ( ~n151 & n1382 ) ;
  assign n1384 = n151 | n1383 ;
  assign n1379 = n274 | n376 ;
  assign n1380 = n485 | n1379 ;
  assign n1398 = n43 | n89 ;
  assign n1399 = n348 | n457 ;
  assign n1400 = n1398 | n1399 ;
  assign n1385 = n417 | n797 ;
  assign n1386 = n165 | n775 ;
  assign n1387 = ( n666 & ~n342 ) | ( n666 & n1386 ) | ( ~n342 & n1386 ) ;
  assign n1388 = n342 | n1387 ;
  assign n1389 = ( n1385 & ~n195 ) | ( n1385 & n1388 ) | ( ~n195 & n1388 ) ;
  assign n1390 = n195 | n1389 ;
  assign n1391 = ( n193 & ~n792 ) | ( n193 & n1390 ) | ( ~n792 & n1390 ) ;
  assign n1392 = n792 | n1391 ;
  assign n1393 = ( n494 & ~n572 ) | ( n494 & n1392 ) | ( ~n572 & n1392 ) ;
  assign n1394 = n572 | n1393 ;
  assign n1395 = ( n353 & ~n663 ) | ( n353 & n1394 ) | ( ~n663 & n1394 ) ;
  assign n1396 = n663 | n1395 ;
  assign n1397 = n358 | n1396 ;
  assign n1401 = ( n1400 & ~n1384 ) | ( n1400 & n1397 ) | ( ~n1384 & n1397 ) ;
  assign n1402 = ( n1384 & ~n1380 ) | ( n1384 & n1401 ) | ( ~n1380 & n1401 ) ;
  assign n1403 = n1402 | n1380 ;
  assign n1404 = ( n341 & ~n374 ) | ( n341 & n1403 ) | ( ~n374 & n1403 ) ;
  assign n1405 = n374 | n1404 ;
  assign n1406 = ( n672 & ~n362 ) | ( n672 & n1405 ) | ( ~n362 & n1405 ) ;
  assign n1407 = n362 | n1406 ;
  assign n1408 = ( n911 & ~n359 ) | ( n911 & n1407 ) | ( ~n359 & n1407 ) ;
  assign n1409 = n359 | n1408 ;
  assign n1410 = ( n559 & ~n554 ) | ( n559 & n1409 ) | ( ~n554 & n1409 ) ;
  assign n1411 = n554 | n1410 ;
  assign n1412 = ( n356 & ~n560 ) | ( n356 & n1411 ) | ( ~n560 & n1411 ) ;
  assign n1413 = n560 | n1412 ;
  assign n1414 = n252 | n1413 ;
  assign n1415 = n118 | n734 ;
  assign n1416 = ( n336 & ~n39 ) | ( n336 & n1415 ) | ( ~n39 & n1415 ) ;
  assign n1417 = n39 | n1416 ;
  assign n1418 = n475 | n1417 ;
  assign n1419 = ( n101 & ~n456 ) | ( n101 & n1418 ) | ( ~n456 & n1418 ) ;
  assign n1420 = n456 | n1419 ;
  assign n1421 = ( n214 & ~n279 ) | ( n214 & n1420 ) | ( ~n279 & n1420 ) ;
  assign n1422 = n279 | n1421 ;
  assign n1423 = ( n135 & n197 ) | ( n135 & n1422 ) | ( n197 & n1422 ) ;
  assign n1424 = ( n197 & ~n1423 ) | ( n197 & 1'b0 ) | ( ~n1423 & 1'b0 ) ;
  assign n1425 = ~n88 & n1424 ;
  assign n1426 = n259 | n676 ;
  assign n1427 = n187 | n257 ;
  assign n1428 = n226 | n255 ;
  assign n1429 = n207 | n789 ;
  assign n1430 = n77 | n529 ;
  assign n1431 = n1429 | n1430 ;
  assign n1432 = ( n452 & ~n106 ) | ( n452 & n1431 ) | ( ~n106 & n1431 ) ;
  assign n1433 = n106 | n1432 ;
  assign n1434 = n157 | n373 ;
  assign n1435 = n120 | n787 ;
  assign n1436 = n670 | n1435 ;
  assign n1437 = ~n230 & n644 ;
  assign n1438 = ~n1436 & n1437 ;
  assign n1439 = ~n1434 & n1438 ;
  assign n1440 = ( n682 & ~n1433 ) | ( n682 & n1439 ) | ( ~n1433 & n1439 ) ;
  assign n1441 = ( n747 & ~n682 ) | ( n747 & n1440 ) | ( ~n682 & n1440 ) ;
  assign n1442 = ~n747 & n1441 ;
  assign n1443 = ( n1428 & ~n1325 ) | ( n1428 & n1442 ) | ( ~n1325 & n1442 ) ;
  assign n1444 = ~n1428 & n1443 ;
  assign n1445 = ( n620 & ~n1427 ) | ( n620 & n1444 ) | ( ~n1427 & n1444 ) ;
  assign n1446 = ~n620 & n1445 ;
  assign n1447 = ( n272 & ~n1426 ) | ( n272 & n1446 ) | ( ~n1426 & n1446 ) ;
  assign n1448 = ~n272 & n1447 ;
  assign n1449 = ( n149 & ~n603 ) | ( n149 & n1448 ) | ( ~n603 & n1448 ) ;
  assign n1450 = ~n149 & n1449 ;
  assign n1451 = ( n643 & ~n646 ) | ( n643 & n1450 ) | ( ~n646 & n1450 ) ;
  assign n1452 = ( n1451 & ~n643 ) | ( n1451 & 1'b0 ) | ( ~n643 & 1'b0 ) ;
  assign n1453 = ~n347 & n1452 ;
  assign n1454 = n105 | n765 ;
  assign n1455 = n527 | n1454 ;
  assign n1456 = ( n492 & ~n569 ) | ( n492 & n1455 ) | ( ~n569 & n1455 ) ;
  assign n1457 = n569 | n1456 ;
  assign n1458 = ( n354 & ~n1457 ) | ( n354 & 1'b0 ) | ( ~n1457 & 1'b0 ) ;
  assign n1465 = ( n766 & ~n58 ) | ( n766 & n812 ) | ( ~n58 & n812 ) ;
  assign n1466 = n58 | n1465 ;
  assign n1467 = n1317 | n1466 ;
  assign n1459 = n241 | n713 ;
  assign n1460 = n129 | n1459 ;
  assign n1461 = n167 | n796 ;
  assign n1462 = n412 | n1461 ;
  assign n1463 = ( n104 & ~n243 ) | ( n104 & n1462 ) | ( ~n243 & n1462 ) ;
  assign n1464 = n243 | n1463 ;
  assign n1468 = ( n1467 & ~n1460 ) | ( n1467 & n1464 ) | ( ~n1460 & n1464 ) ;
  assign n1469 = ( n1458 & n1468 ) | ( n1458 & n1460 ) | ( n1468 & n1460 ) ;
  assign n1470 = ( n1458 & ~n1469 ) | ( n1458 & 1'b0 ) | ( ~n1469 & 1'b0 ) ;
  assign n1471 = ( n1453 & ~n1425 ) | ( n1453 & n1470 ) | ( ~n1425 & n1470 ) ;
  assign n1472 = ( n75 & n1425 ) | ( n75 & n1471 ) | ( n1425 & n1471 ) ;
  assign n1473 = ~n75 & n1472 ;
  assign n1474 = ( n434 & ~n1414 ) | ( n434 & n1473 ) | ( ~n1414 & n1473 ) ;
  assign n1475 = ~n434 & n1474 ;
  assign n1476 = ( n218 & ~n1475 ) | ( n218 & n813 ) | ( ~n1475 & n813 ) ;
  assign n1477 = ( n813 & ~n1476 ) | ( n813 & 1'b0 ) | ( ~n1476 & 1'b0 ) ;
  assign n1478 = ( n905 & ~n418 ) | ( n905 & n1477 ) | ( ~n418 & n1477 ) ;
  assign n1479 = ~n905 & n1478 ;
  assign n1480 = ( n269 & ~n221 ) | ( n269 & n1479 ) | ( ~n221 & n1479 ) ;
  assign n1481 = ~n269 & n1480 ;
  assign n1482 = ( n623 & ~n1481 ) | ( n623 & n630 ) | ( ~n1481 & n630 ) ;
  assign n1483 = ~n623 |  n1482 ;
  assign n1484 = n140 | n761 ;
  assign n1485 = ~n280 & n813 ;
  assign n1486 = ( n557 & ~n96 ) | ( n557 & n1485 ) | ( ~n96 & n1485 ) ;
  assign n1487 = ( n124 & ~n557 ) | ( n124 & n1486 ) | ( ~n557 & n1486 ) ;
  assign n1488 = ~n124 & n1487 ;
  assign n1489 = ~n273 & n1488 ;
  assign n1490 = n236 | n744 ;
  assign n1491 = n126 | n453 ;
  assign n1492 = ( n234 & ~n431 ) | ( n234 & n720 ) | ( ~n431 & n720 ) ;
  assign n1493 = n431 | n1492 ;
  assign n1494 = n157 | n627 ;
  assign n1495 = n349 | n560 ;
  assign n1496 = n231 | n347 ;
  assign n1497 = n86 | n167 ;
  assign n1498 = n138 | n676 ;
  assign n1499 = ( n1497 & ~n1496 ) | ( n1497 & n1498 ) | ( ~n1496 & n1498 ) ;
  assign n1500 = n1496 | n1499 ;
  assign n1501 = ( n1046 & ~n75 ) | ( n1046 & n1500 ) | ( ~n75 & n1500 ) ;
  assign n1502 = n75 | n1501 ;
  assign n1503 = ( n1495 & ~n1494 ) | ( n1495 & n1502 ) | ( ~n1494 & n1502 ) ;
  assign n1504 = n1494 | n1503 ;
  assign n1505 = ( n1493 & ~n1491 ) | ( n1493 & n1504 ) | ( ~n1491 & n1504 ) ;
  assign n1506 = n1491 | n1505 ;
  assign n1507 = ( n1490 & ~n65 ) | ( n1490 & n1506 ) | ( ~n65 & n1506 ) ;
  assign n1508 = n65 | n1507 ;
  assign n1509 = ( n350 & ~n225 ) | ( n350 & n1508 ) | ( ~n225 & n1508 ) ;
  assign n1510 = n225 | n1509 ;
  assign n1512 = n196 | n734 ;
  assign n1513 = n285 | n460 ;
  assign n1514 = ( n101 & ~n478 ) | ( n101 & n572 ) | ( ~n478 & n572 ) ;
  assign n1515 = n478 | n1514 ;
  assign n1516 = ( n1207 & ~n1063 ) | ( n1207 & n1515 ) | ( ~n1063 & n1515 ) ;
  assign n1517 = n1063 | n1516 ;
  assign n1518 = ( n1513 & ~n1512 ) | ( n1513 & n1517 ) | ( ~n1512 & n1517 ) ;
  assign n1519 = n1512 | n1518 ;
  assign n1520 = ( n1093 & ~n1428 ) | ( n1093 & n1519 ) | ( ~n1428 & n1519 ) ;
  assign n1521 = n1428 | n1520 ;
  assign n1511 = n279 | n671 ;
  assign n1522 = ( n1521 & ~n1072 ) | ( n1521 & n1511 ) | ( ~n1072 & n1511 ) ;
  assign n1523 = n1072 | n1522 ;
  assign n1524 = ( n357 & ~n362 ) | ( n357 & n1523 ) | ( ~n362 & n1523 ) ;
  assign n1525 = n362 | n1524 ;
  assign n1526 = ( n765 & ~n554 ) | ( n765 & n1525 ) | ( ~n554 & n1525 ) ;
  assign n1527 = n554 | n1526 ;
  assign n1528 = ( n118 & ~n228 ) | ( n118 & n1527 ) | ( ~n228 & n1527 ) ;
  assign n1529 = n228 | n1528 ;
  assign n1530 = ( n141 & ~n670 ) | ( n141 & n1529 ) | ( ~n670 & n1529 ) ;
  assign n1531 = n670 | n1530 ;
  assign n1532 = n105 | n359 ;
  assign n1533 = ( n129 & ~n663 ) | ( n129 & n335 ) | ( ~n663 & n335 ) ;
  assign n1534 = n663 | n1533 ;
  assign n1535 = ( n215 & ~n1532 ) | ( n215 & n1534 ) | ( ~n1532 & n1534 ) ;
  assign n1536 = ( n1532 & ~n150 ) | ( n1532 & n1535 ) | ( ~n150 & n1535 ) ;
  assign n1537 = n150 | n1536 ;
  assign n1538 = ( n602 & ~n429 ) | ( n602 & n1537 ) | ( ~n429 & n1537 ) ;
  assign n1539 = ( n429 & ~n775 ) | ( n429 & n1538 ) | ( ~n775 & n1538 ) ;
  assign n1540 = n775 | n1539 ;
  assign n1541 = n269 | n1540 ;
  assign n1542 = n252 | n1541 ;
  assign n1543 = ( n673 & ~n674 ) | ( n673 & n1306 ) | ( ~n674 & n1306 ) ;
  assign n1544 = n674 | n1543 ;
  assign n1545 = n241 | n1544 ;
  assign n1546 = n83 | n408 ;
  assign n1547 = ( n197 & ~n630 ) | ( n197 & 1'b0 ) | ( ~n630 & 1'b0 ) ;
  assign n1548 = ( n406 & ~n332 ) | ( n406 & n424 ) | ( ~n332 & n424 ) ;
  assign n1549 = n332 | n1548 ;
  assign n1550 = n132 | n571 ;
  assign n1551 = ( n1547 & n1549 ) | ( n1547 & n1550 ) | ( n1549 & n1550 ) ;
  assign n1552 = ( n1546 & ~n1551 ) | ( n1546 & n1547 ) | ( ~n1551 & n1547 ) ;
  assign n1553 = ~n1546 & n1552 ;
  assign n1554 = ( n1542 & ~n1545 ) | ( n1542 & n1553 ) | ( ~n1545 & n1553 ) ;
  assign n1555 = ( n1554 & ~n1542 ) | ( n1554 & 1'b0 ) | ( ~n1542 & 1'b0 ) ;
  assign n1556 = ( n1510 & ~n1531 ) | ( n1510 & n1555 ) | ( ~n1531 & n1555 ) ;
  assign n1557 = ~n1510 & n1556 ;
  assign n1558 = ( n1183 & ~n1489 ) | ( n1183 & n1557 ) | ( ~n1489 & n1557 ) ;
  assign n1559 = n1489 &  n1558 ;
  assign n1560 = ( n62 & ~n1484 ) | ( n62 & n1559 ) | ( ~n1484 & n1559 ) ;
  assign n1561 = ~n62 & n1560 ;
  assign n1562 = ( n355 & n458 ) | ( n355 & n1561 ) | ( n458 & n1561 ) ;
  assign n1563 = ( n230 & ~n458 ) | ( n230 & n1562 ) | ( ~n458 & n1562 ) ;
  assign n1564 = ~n230 & n1563 ;
  assign n1565 = ( n664 & ~n459 ) | ( n664 & n1564 ) | ( ~n459 & n1564 ) ;
  assign n1566 = ~n664 &  n1565 ;
  assign n1567 = n775 | n812 ;
  assign n1568 = n187 | n372 ;
  assign n1569 = n571 | n1568 ;
  assign n1570 = ( n1567 & ~n974 ) | ( n1567 & n1569 ) | ( ~n974 & n1569 ) ;
  assign n1571 = ( n974 & ~n61 ) | ( n974 & n1570 ) | ( ~n61 & n1570 ) ;
  assign n1572 = n61 | n1571 ;
  assign n1573 = ( n69 & ~n168 ) | ( n69 & n1572 ) | ( ~n168 & n1572 ) ;
  assign n1574 = n168 | n1573 ;
  assign n1575 = ( n271 & ~n714 ) | ( n271 & n1574 ) | ( ~n714 & n1574 ) ;
  assign n1576 = n714 | n1575 ;
  assign n1577 = ( n382 & ~n252 ) | ( n382 & n1576 ) | ( ~n252 & n1576 ) ;
  assign n1578 = n252 | n1577 ;
  assign n1579 = n196 | n1578 ;
  assign n1580 = n49 | n745 ;
  assign n1581 = n141 | n212 ;
  assign n1595 = ( n527 & ~n243 ) | ( n527 & n734 ) | ( ~n243 & n734 ) ;
  assign n1596 = n243 | n1595 ;
  assign n1597 = ( n255 & ~n236 ) | ( n255 & n1596 ) | ( ~n236 & n1596 ) ;
  assign n1598 = n236 | n1597 ;
  assign n1599 = n99 | n1598 ;
  assign n1600 = n89 | n720 ;
  assign n1601 = ( n604 & ~n342 ) | ( n604 & n814 ) | ( ~n342 & n814 ) ;
  assign n1602 = n342 | n1601 ;
  assign n1603 = n433 | n631 ;
  assign n1604 = ( n1602 & ~n1600 ) | ( n1602 & n1603 ) | ( ~n1600 & n1603 ) ;
  assign n1605 = n1600 | n1604 ;
  assign n1606 = ( n1355 & ~n1599 ) | ( n1355 & n1605 ) | ( ~n1599 & n1605 ) ;
  assign n1607 = n1599 | n1606 ;
  assign n1582 = ( n432 & ~n169 ) | ( n432 & n1269 ) | ( ~n169 & n1269 ) ;
  assign n1583 = n169 | n1582 ;
  assign n1584 = n39 | n1583 ;
  assign n1585 = n534 | n630 ;
  assign n1586 = ( n462 & ~n1584 ) | ( n462 & n1585 ) | ( ~n1584 & n1585 ) ;
  assign n1587 = n1584 | n1586 ;
  assign n1588 = ( n345 & ~n376 ) | ( n345 & n1587 ) | ( ~n376 & n1587 ) ;
  assign n1589 = n376 | n1588 ;
  assign n1590 = ( n792 & ~n800 ) | ( n792 & n1589 ) | ( ~n800 & n1589 ) ;
  assign n1591 = n800 | n1590 ;
  assign n1592 = ( n268 & ~n424 ) | ( n268 & n1591 ) | ( ~n424 & n1591 ) ;
  assign n1593 = n424 | n1592 ;
  assign n1594 = n411 | n1593 ;
  assign n1608 = ( n1607 & ~n1581 ) | ( n1607 & n1594 ) | ( ~n1581 & n1594 ) ;
  assign n1609 = ( n1581 & ~n842 ) | ( n1581 & n1608 ) | ( ~n842 & n1608 ) ;
  assign n1610 = n842 | n1609 ;
  assign n1611 = ( n1580 & ~n713 ) | ( n1580 & n1610 ) | ( ~n713 & n1610 ) ;
  assign n1612 = n713 | n1611 ;
  assign n1613 = ( n409 & ~n138 ) | ( n409 & n1612 ) | ( ~n138 & n1612 ) ;
  assign n1614 = n138 | n1613 ;
  assign n1615 = ( n451 & ~n663 ) | ( n451 & n1614 ) | ( ~n663 & n1614 ) ;
  assign n1616 = n663 | n1615 ;
  assign n1625 = n418 | n664 ;
  assign n1626 = n280 | n788 ;
  assign n1627 = n231 | n415 ;
  assign n1628 = ( n721 & ~n908 ) | ( n721 & n864 ) | ( ~n908 & n864 ) ;
  assign n1629 = ( n908 & ~n188 ) | ( n908 & n1628 ) | ( ~n188 & n1628 ) ;
  assign n1630 = n188 | n1629 ;
  assign n1631 = n554 | n1630 ;
  assign n1632 = n58 | n101 ;
  assign n1633 = n123 | n1632 ;
  assign n1634 = ( n166 & ~n267 ) | ( n166 & n528 ) | ( ~n267 & n528 ) ;
  assign n1635 = n267 | n1634 ;
  assign n1636 = ( n622 & ~n1357 ) | ( n622 & n1635 ) | ( ~n1357 & n1635 ) ;
  assign n1637 = n1357 | n1636 ;
  assign n1638 = ( n1633 & ~n629 ) | ( n1633 & n1637 ) | ( ~n629 & n1637 ) ;
  assign n1639 = n629 | n1638 ;
  assign n1640 = ( n1631 & ~n1627 ) | ( n1631 & n1639 ) | ( ~n1627 & n1639 ) ;
  assign n1641 = n1627 | n1640 ;
  assign n1642 = ( n1626 & ~n1454 ) | ( n1626 & n1641 ) | ( ~n1454 & n1641 ) ;
  assign n1643 = n1454 | n1642 ;
  assign n1644 = ( n1625 & ~n458 ) | ( n1625 & n1643 ) | ( ~n458 & n1643 ) ;
  assign n1645 = n458 | n1644 ;
  assign n1646 = ( n493 & ~n284 ) | ( n493 & n1645 ) | ( ~n284 & n1645 ) ;
  assign n1647 = n284 | n1646 ;
  assign n1648 = ( n91 & ~n120 ) | ( n91 & n1647 ) | ( ~n120 & n1647 ) ;
  assign n1649 = n120 | n1648 ;
  assign n1650 = n205 | n1649 ;
  assign n1617 = n43 | n161 ;
  assign n1618 = n139 | n233 ;
  assign n1619 = ( n1617 & ~n72 ) | ( n1617 & n1618 ) | ( ~n72 & n1618 ) ;
  assign n1620 = n72 | n1619 ;
  assign n1621 = ( n1620 & ~n333 ) | ( n1620 & n737 ) | ( ~n333 & n737 ) ;
  assign n1622 = n333 | n1621 ;
  assign n1623 = ( n549 & ~n431 ) | ( n549 & n1622 ) | ( ~n431 & n1622 ) ;
  assign n1624 = n431 | n1623 ;
  assign n1651 = ( n125 & ~n744 ) | ( n125 & n193 ) | ( ~n744 & n193 ) ;
  assign n1652 = n744 | n1651 ;
  assign n1653 = n356 | n1652 ;
  assign n1656 = n477 | n722 ;
  assign n1657 = n529 | n1656 ;
  assign n1654 = ( n117 & ~n351 ) | ( n117 & n569 ) | ( ~n351 & n569 ) ;
  assign n1655 = n351 | n1654 ;
  assign n1658 = ( n1657 & ~n1653 ) | ( n1657 & n1655 ) | ( ~n1653 & n1655 ) ;
  assign n1659 = n1653 | n1658 ;
  assign n1660 = ( n1650 & ~n1624 ) | ( n1650 & n1659 ) | ( ~n1624 & n1659 ) ;
  assign n1661 = n1660 | n1624 ;
  assign n1662 = ( n1044 & ~n1616 ) | ( n1044 & n1661 ) | ( ~n1616 & n1661 ) ;
  assign n1663 = n1616 | n1662 ;
  assign n1664 = ( n1579 & n1663 ) | ( n1579 & n525 ) | ( n1663 & n525 ) ;
  assign n1665 = ( n525 & ~n1664 ) | ( n525 & 1'b0 ) | ( ~n1664 & 1'b0 ) ;
  assign n1666 = ( n245 & ~n909 ) | ( n245 & n1665 ) | ( ~n909 & n1665 ) ;
  assign n1667 = ~n245 & n1666 ;
  assign n1668 = ( n74 & ~n239 ) | ( n74 & n1667 ) | ( ~n239 & n1667 ) ;
  assign n1669 = ~n74 & n1668 ;
  assign n1670 = ( n347 & ~n574 ) | ( n347 & n1669 ) | ( ~n574 & n1669 ) ;
  assign n1671 = ~n347 & n1670 ;
  assign n1672 = n190 | n272 ;
  assign n1673 = n1284 | n1672 ;
  assign n1674 = ( n168 & n813 ) | ( n168 & n1673 ) | ( n813 & n1673 ) ;
  assign n1675 = ( n813 & ~n1674 ) | ( n813 & 1'b0 ) | ( ~n1674 & 1'b0 ) ;
  assign n1676 = ( n140 & ~n239 ) | ( n140 & n1675 ) | ( ~n239 & n1675 ) ;
  assign n1677 = ~n140 & n1676 ;
  assign n1678 = n242 | n274 ;
  assign n1679 = n628 | n778 ;
  assign n1687 = n72 | n456 ;
  assign n1688 = ( n222 & ~n275 ) | ( n222 & n412 ) | ( ~n275 & n412 ) ;
  assign n1689 = n275 | n1688 ;
  assign n1690 = n494 | n722 ;
  assign n1691 = ( n960 & ~n1690 ) | ( n960 & n1009 ) | ( ~n1690 & n1009 ) ;
  assign n1692 = n1690 | n1691 ;
  assign n1693 = ( n1689 & ~n1687 ) | ( n1689 & n1692 ) | ( ~n1687 & n1692 ) ;
  assign n1694 = n1687 | n1693 ;
  assign n1680 = ( n359 & ~n796 ) | ( n359 & n683 ) | ( ~n796 & n683 ) ;
  assign n1681 = n796 | n1680 ;
  assign n1682 = ( n231 & n1681 ) | ( n231 & n644 ) | ( n1681 & n644 ) ;
  assign n1683 = ( n644 & ~n1682 ) | ( n644 & 1'b0 ) | ( ~n1682 & 1'b0 ) ;
  assign n1684 = ( n256 & ~n618 ) | ( n256 & n1683 ) | ( ~n618 & n1683 ) ;
  assign n1685 = ~n256 & n1684 ;
  assign n1686 = ~n459 & n1685 ;
  assign n1695 = ( n1679 & ~n1694 ) | ( n1679 & n1686 ) | ( ~n1694 & n1686 ) ;
  assign n1696 = ~n1679 & n1695 ;
  assign n1697 = ( n1678 & ~n790 ) | ( n1678 & n1696 ) | ( ~n790 & n1696 ) ;
  assign n1698 = ( n812 & ~n1678 ) | ( n812 & n1697 ) | ( ~n1678 & n1697 ) ;
  assign n1699 = ~n812 & n1698 ;
  assign n1700 = ( n122 & ~n350 ) | ( n122 & n1699 ) | ( ~n350 & n1699 ) ;
  assign n1701 = ~n122 & n1700 ;
  assign n1703 = n95 | n124 ;
  assign n1704 = n281 | n340 ;
  assign n1705 = ( n345 & ~n674 ) | ( n345 & n1704 ) | ( ~n674 & n1704 ) ;
  assign n1706 = n674 | n1705 ;
  assign n1707 = ( n792 & ~n490 ) | ( n792 & n1706 ) | ( ~n490 & n1706 ) ;
  assign n1708 = ( n490 & ~n734 ) | ( n490 & n1707 ) | ( ~n734 & n1707 ) ;
  assign n1709 = n734 | n1708 ;
  assign n1710 = n666 | n1709 ;
  assign n1711 = n235 | n678 ;
  assign n1712 = ( n88 & ~n338 ) | ( n88 & n1711 ) | ( ~n338 & n1711 ) ;
  assign n1713 = n338 | n1712 ;
  assign n1714 = n646 | n1713 ;
  assign n1715 = n192 | n299 ;
  assign n1716 = ( n1123 & ~n1714 ) | ( n1123 & n1715 ) | ( ~n1714 & n1715 ) ;
  assign n1717 = n1714 | n1716 ;
  assign n1718 = ( n530 & ~n1710 ) | ( n530 & n1717 ) | ( ~n1710 & n1717 ) ;
  assign n1719 = n1710 | n1718 ;
  assign n1720 = ( n1703 & ~n1581 ) | ( n1703 & n1719 ) | ( ~n1581 & n1719 ) ;
  assign n1721 = n1581 | n1720 ;
  assign n1722 = ( n711 & ~n150 ) | ( n711 & n1721 ) | ( ~n150 & n1721 ) ;
  assign n1723 = n150 | n1722 ;
  assign n1724 = ( n123 & ~n216 ) | ( n123 & n1723 ) | ( ~n216 & n1723 ) ;
  assign n1725 = n216 | n1724 ;
  assign n1726 = ( n49 & ~n454 ) | ( n49 & n1725 ) | ( ~n454 & n1725 ) ;
  assign n1727 = n454 | n1726 ;
  assign n1728 = n351 | n1727 ;
  assign n1729 = n130 | n429 ;
  assign n1730 = n136 | n712 ;
  assign n1731 = n342 | n1730 ;
  assign n1732 = n138 | n558 ;
  assign n1733 = ( n1731 & ~n1729 ) | ( n1731 & n1732 ) | ( ~n1729 & n1732 ) ;
  assign n1734 = n1729 | n1733 ;
  assign n1735 = ( n385 & ~n1728 ) | ( n385 & n1734 ) | ( ~n1728 & n1734 ) ;
  assign n1736 = n1728 | n1735 ;
  assign n1702 = n126 | n1550 ;
  assign n1737 = ( n1701 & n1736 ) | ( n1701 & n1702 ) | ( n1736 & n1702 ) ;
  assign n1738 = ( n215 & ~n1737 ) | ( n215 & n1701 ) | ( ~n1737 & n1701 ) ;
  assign n1739 = ~n215 & n1738 ;
  assign n1740 = ( n1279 & n1316 ) | ( n1279 & n1739 ) | ( n1316 & n1739 ) ;
  assign n1741 = ~n1316 & n1740 ;
  assign n1742 = ( n1268 & ~n1741 ) | ( n1268 & n1677 ) | ( ~n1741 & n1677 ) ;
  assign n1743 = ( n624 & ~n1677 ) | ( n624 & n1742 ) | ( ~n1677 & n1742 ) ;
  assign n1744 = ( n624 & ~n1743 ) | ( n624 & 1'b0 ) | ( ~n1743 & 1'b0 ) ;
  assign n1745 = ( n721 & ~n434 ) | ( n721 & n1744 ) | ( ~n434 & n1744 ) ;
  assign n1746 = ~n721 & n1745 ;
  assign n1747 = ( n269 & ~n403 ) | ( n269 & n1746 ) | ( ~n403 & n1746 ) ;
  assign n1748 = ~n269 & n1747 ;
  assign n1749 = ( n424 & ~n106 ) | ( n424 & n531 ) | ( ~n106 & n531 ) ;
  assign n1750 = ( n106 & n1485 ) | ( n106 & n1749 ) | ( n1485 & n1749 ) ;
  assign n1751 = ( n1485 & ~n1750 ) | ( n1485 & 1'b0 ) | ( ~n1750 & 1'b0 ) ;
  assign n1752 = n735 | n814 ;
  assign n1753 = n132 | n1752 ;
  assign n1754 = n284 | n373 ;
  assign n1755 = ( n1753 & ~n672 ) | ( n1753 & n1754 ) | ( ~n672 & n1754 ) ;
  assign n1756 = n672 | n1755 ;
  assign n1757 = ( n255 & ~n745 ) | ( n255 & n1756 ) | ( ~n745 & n1756 ) ;
  assign n1758 = n745 | n1757 ;
  assign n1759 = ( n529 & ~n574 ) | ( n529 & n1758 ) | ( ~n574 & n1758 ) ;
  assign n1760 = n574 | n1759 ;
  assign n1761 = n129 | n1760 ;
  assign n1762 = n558 | n722 ;
  assign n1763 = ~n88 & n484 ;
  assign n1764 = ~n617 & n1763 ;
  assign n1765 = ( n491 & n632 ) | ( n491 & n1764 ) | ( n632 & n1764 ) ;
  assign n1766 = ( n72 & ~n1765 ) | ( n72 & n1764 ) | ( ~n1765 & n1764 ) ;
  assign n1767 = ~n72 & n1766 ;
  assign n1768 = ( n243 & ~n101 ) | ( n243 & n1767 ) | ( ~n101 & n1767 ) ;
  assign n1769 = ~n243 & n1768 ;
  assign n1770 = ( n231 & ~n526 ) | ( n231 & n1769 ) | ( ~n526 & n1769 ) ;
  assign n1771 = ~n231 & n1770 ;
  assign n1772 = ( n239 & ~n1771 ) | ( n239 & n354 ) | ( ~n1771 & n354 ) ;
  assign n1773 = ( n354 & ~n1772 ) | ( n354 & 1'b0 ) | ( ~n1772 & 1'b0 ) ;
  assign n1774 = ~n83 & n1773 ;
  assign n1775 = ( n789 & ~n268 ) | ( n789 & n910 ) | ( ~n268 & n910 ) ;
  assign n1776 = n268 | n1775 ;
  assign n1777 = ( n603 & ~n151 ) | ( n603 & n1776 ) | ( ~n151 & n1776 ) ;
  assign n1778 = n151 | n1777 ;
  assign n1779 = ( n404 & ~n478 ) | ( n404 & n627 ) | ( ~n478 & n627 ) ;
  assign n1780 = ( n478 & n525 ) | ( n478 & n1779 ) | ( n525 & n1779 ) ;
  assign n1781 = ( n525 & ~n1780 ) | ( n525 & 1'b0 ) | ( ~n1780 & 1'b0 ) ;
  assign n1782 = ( n1778 & ~n1288 ) | ( n1778 & n1781 ) | ( ~n1288 & n1781 ) ;
  assign n1783 = ~n1778 & n1782 ;
  assign n1784 = ( n1762 & n1774 ) | ( n1762 & n1783 ) | ( n1774 & n1783 ) ;
  assign n1785 = ~n1762 & n1784 ;
  assign n1786 = ( n1761 & ~n1785 ) | ( n1761 & n645 ) | ( ~n1785 & n645 ) ;
  assign n1787 = ( n645 & ~n1786 ) | ( n645 & 1'b0 ) | ( ~n1786 & 1'b0 ) ;
  assign n1788 = ( n1490 & n1751 ) | ( n1490 & n1787 ) | ( n1751 & n1787 ) ;
  assign n1789 = ~n1490 & n1788 ;
  assign n1790 = ( n348 & ~n559 ) | ( n348 & n1789 ) | ( ~n559 & n1789 ) ;
  assign n1791 = ( n217 & ~n348 ) | ( n217 & n1790 ) | ( ~n348 & n1790 ) ;
  assign n1792 = ~n217 & n1791 ;
  assign n1793 = ( n561 & ~n432 ) | ( n561 & n1792 ) | ( ~n432 & n1792 ) ;
  assign n1794 = ~n561 & n1793 ;
  assign n1795 = n43 | n459 ;
  assign n1796 = n149 | n235 ;
  assign n1797 = n205 | n276 ;
  assign n1798 = ( n1797 & ~n189 ) | ( n1797 & n1271 ) | ( ~n189 & n1271 ) ;
  assign n1799 = n189 | n1798 ;
  assign n1800 = ( n1796 & ~n1679 ) | ( n1796 & n1799 ) | ( ~n1679 & n1799 ) ;
  assign n1801 = n1679 | n1800 ;
  assign n1802 = ( n271 & ~n168 ) | ( n271 & n1801 ) | ( ~n168 & n1801 ) ;
  assign n1803 = n168 | n1802 ;
  assign n1804 = ( n212 & ~n1795 ) | ( n212 & n1803 ) | ( ~n1795 & n1803 ) ;
  assign n1805 = ( n1795 & ~n356 ) | ( n1795 & n1804 ) | ( ~n356 & n1804 ) ;
  assign n1806 = n356 | n1805 ;
  assign n1808 = n244 | n560 ;
  assign n1807 = n166 | n372 ;
  assign n1809 = n208 | n602 ;
  assign n1810 = n270 | n663 ;
  assign n1811 = ( n1809 & ~n811 ) | ( n1809 & n1810 ) | ( ~n811 & n1810 ) ;
  assign n1812 = n811 | n1811 ;
  assign n1813 = ( n1808 & ~n1807 ) | ( n1808 & n1812 ) | ( ~n1807 & n1812 ) ;
  assign n1814 = ( n1813 & ~n737 ) | ( n1813 & n1807 ) | ( ~n737 & n1807 ) ;
  assign n1815 = n737 | n1814 ;
  assign n1816 = ( n451 & ~n905 ) | ( n451 & n1815 ) | ( ~n905 & n1815 ) ;
  assign n1817 = n905 | n1816 ;
  assign n1818 = ( n141 & ~n1817 ) | ( n141 & n197 ) | ( ~n1817 & n197 ) ;
  assign n1819 = ~n141 & n1818 ;
  assign n1820 = n233 | n721 ;
  assign n1821 = n460 | n549 ;
  assign n1822 = ( n49 & ~n571 ) | ( n49 & n1821 ) | ( ~n571 & n1821 ) ;
  assign n1823 = n571 | n1822 ;
  assign n1824 = n162 | n712 ;
  assign n1825 = ( n605 & ~n273 ) | ( n605 & n1824 ) | ( ~n273 & n1824 ) ;
  assign n1826 = n273 | n1825 ;
  assign n1827 = n485 | n1826 ;
  assign n1828 = n671 | n796 ;
  assign n1829 = n122 | n191 ;
  assign n1830 = n618 | n797 ;
  assign n1831 = n646 | n1830 ;
  assign n1832 = n242 | n493 ;
  assign n1833 = n353 | n1832 ;
  assign n1834 = ( n1831 & ~n1829 ) | ( n1831 & n1833 ) | ( ~n1829 & n1833 ) ;
  assign n1835 = n1829 | n1834 ;
  assign n1836 = ( n339 & ~n1828 ) | ( n339 & n1835 ) | ( ~n1828 & n1835 ) ;
  assign n1837 = ( n1836 & ~n453 ) | ( n1836 & n1828 ) | ( ~n453 & n1828 ) ;
  assign n1838 = n453 | n1837 ;
  assign n1839 = ( n332 & ~n74 ) | ( n332 & n1838 ) | ( ~n74 & n1838 ) ;
  assign n1840 = n74 | n1839 ;
  assign n1841 = n351 | n1840 ;
  assign n1842 = ( n1436 & ~n1827 ) | ( n1436 & n1841 ) | ( ~n1827 & n1841 ) ;
  assign n1843 = ( n1827 & ~n1600 ) | ( n1827 & n1842 ) | ( ~n1600 & n1842 ) ;
  assign n1844 = n1600 | n1843 ;
  assign n1845 = ( n1823 & ~n1820 ) | ( n1823 & n1844 ) | ( ~n1820 & n1844 ) ;
  assign n1846 = n1820 | n1845 ;
  assign n1847 = ( n416 & ~n788 ) | ( n416 & n1846 ) | ( ~n788 & n1846 ) ;
  assign n1848 = n788 | n1847 ;
  assign n1849 = ( n193 & ~n138 ) | ( n193 & n1848 ) | ( ~n138 & n1848 ) ;
  assign n1850 = n138 | n1849 ;
  assign n1851 = ( n253 & ~n800 ) | ( n253 & n1850 ) | ( ~n800 & n1850 ) ;
  assign n1852 = n800 | n1851 ;
  assign n1853 = n256 | n1852 ;
  assign n1854 = n1484 | n1703 ;
  assign n1855 = n333 | n1854 ;
  assign n1856 = n125 | n194 ;
  assign n1857 = n350 | n1856 ;
  assign n1858 = ( n259 & ~n674 ) | ( n259 & n1857 ) | ( ~n674 & n1857 ) ;
  assign n1859 = n674 | n1858 ;
  assign n1860 = ( n1855 & ~n1853 ) | ( n1855 & n1859 ) | ( ~n1853 & n1859 ) ;
  assign n1861 = n1853 | n1860 ;
  assign n1862 = ( n1819 & ~n1861 ) | ( n1819 & n1806 ) | ( ~n1861 & n1806 ) ;
  assign n1863 = ( n606 & ~n1806 ) | ( n606 & n1862 ) | ( ~n1806 & n1862 ) ;
  assign n1864 = ~n606 & n1863 ;
  assign n1865 = ( n679 & n1794 ) | ( n679 & n1864 ) | ( n1794 & n1864 ) ;
  assign n1866 = ~n679 & n1865 ;
  assign n1867 = ( n714 & ~n1866 ) | ( n714 & n786 ) | ( ~n1866 & n786 ) ;
  assign n1868 = ( n786 & ~n1867 ) | ( n786 & 1'b0 ) | ( ~n1867 & 1'b0 ) ;
  assign n1869 = ( n139 & ~n911 ) | ( n139 & n1868 ) | ( ~n911 & n1868 ) ;
  assign n1870 = ~n139 & n1869 ;
  assign n1871 = ( n417 & ~n342 ) | ( n417 & n1870 ) | ( ~n342 & n1870 ) ;
  assign n1872 = ~n417 & n1871 ;
  assign n1873 = ( n1872 & ~n137 ) | ( n1872 & n643 ) | ( ~n137 & n643 ) ;
  assign n1874 = ( n1873 & ~n643 ) | ( n1873 & 1'b0 ) | ( ~n643 & 1'b0 ) ;
  assign n1875 = ~n433 &  n1874 ;
  assign n1876 = n65 | n74 ;
  assign n1877 = n150 | n348 ;
  assign n1878 = ( n375 & ~n257 ) | ( n375 & n1877 ) | ( ~n257 & n1877 ) ;
  assign n1879 = n257 | n1878 ;
  assign n1880 = ( n252 & ~n190 ) | ( n252 & n1879 ) | ( ~n190 & n1879 ) ;
  assign n1881 = n190 | n1880 ;
  assign n1882 = n155 | n1881 ;
  assign n1883 = n157 | n228 ;
  assign n1884 = n268 | n643 ;
  assign n1885 = n129 | n345 ;
  assign n1886 = ~n277 & n1751 ;
  assign n1887 = ~n574 & n1886 ;
  assign n1888 = ( n1859 & ~n1885 ) | ( n1859 & n1887 ) | ( ~n1885 & n1887 ) ;
  assign n1889 = ~n1859 & n1888 ;
  assign n1890 = ( n96 & ~n528 ) | ( n96 & n1889 ) | ( ~n528 & n1889 ) ;
  assign n1891 = ~n96 & n1890 ;
  assign n1892 = ( n1567 & ~n1884 ) | ( n1567 & n1891 ) | ( ~n1884 & n1891 ) ;
  assign n1893 = ~n1567 & n1892 ;
  assign n1894 = ( n1625 & ~n969 ) | ( n1625 & n1893 ) | ( ~n969 & n1893 ) ;
  assign n1895 = ~n1625 & n1894 ;
  assign n1896 = ( n126 & ~n461 ) | ( n126 & n1895 ) | ( ~n461 & n1895 ) ;
  assign n1897 = ~n126 & n1896 ;
  assign n1898 = ( n1656 & ~n274 ) | ( n1656 & n1897 ) | ( ~n274 & n1897 ) ;
  assign n1899 = ~n1656 & n1898 ;
  assign n1900 = ( n485 & ~n206 ) | ( n485 & n1899 ) | ( ~n206 & n1899 ) ;
  assign n1901 = ~n485 & n1900 ;
  assign n1902 = ( n214 & ~n336 ) | ( n214 & n1901 ) | ( ~n336 & n1901 ) ;
  assign n1903 = ~n214 & n1902 ;
  assign n1904 = ~n39 & n1903 ;
  assign n1905 = n376 | n403 ;
  assign n1906 = ( n410 & ~n300 ) | ( n410 & n1905 ) | ( ~n300 & n1905 ) ;
  assign n1907 = n300 | n1906 ;
  assign n1908 = ( n676 & ~n361 ) | ( n676 & n1907 ) | ( ~n361 & n1907 ) ;
  assign n1909 = ( n361 & n1908 ) | ( n361 & n1155 ) | ( n1908 & n1155 ) ;
  assign n1910 = ( n1155 & ~n1909 ) | ( n1155 & 1'b0 ) | ( ~n1909 & 1'b0 ) ;
  assign n1911 = ( n333 & ~n602 ) | ( n333 & n1910 ) | ( ~n602 & n1910 ) ;
  assign n1912 = ~n333 & n1911 ;
  assign n1913 = ( n216 & ~n207 ) | ( n216 & n1912 ) | ( ~n207 & n1912 ) ;
  assign n1914 = ~n216 & n1913 ;
  assign n1915 = ( n558 & ~n382 ) | ( n558 & n1914 ) | ( ~n382 & n1914 ) ;
  assign n1916 = ~n558 & n1915 ;
  assign n1917 = ~n86 & n1916 ;
  assign n1918 = ( n241 & ~n678 ) | ( n241 & n947 ) | ( ~n678 & n947 ) ;
  assign n1919 = n678 | n1918 ;
  assign n1920 = n618 | n1919 ;
  assign n1921 = ( n81 & ~n1493 ) | ( n81 & n527 ) | ( ~n1493 & n527 ) ;
  assign n1922 = n1493 | n1921 ;
  assign n1923 = n417 | n1922 ;
  assign n1924 = ( n286 & ~n1920 ) | ( n286 & n1923 ) | ( ~n1920 & n1923 ) ;
  assign n1925 = ( n1920 & ~n1603 ) | ( n1920 & n1924 ) | ( ~n1603 & n1924 ) ;
  assign n1926 = n1603 | n1925 ;
  assign n1927 = ( n1904 & ~n1917 ) | ( n1904 & n1926 ) | ( ~n1917 & n1926 ) ;
  assign n1928 = ( n1904 & ~n1927 ) | ( n1904 & 1'b0 ) | ( ~n1927 & 1'b0 ) ;
  assign n1929 = ( n1882 & ~n1883 ) | ( n1882 & n1928 ) | ( ~n1883 & n1928 ) ;
  assign n1930 = ( n1060 & ~n1882 ) | ( n1060 & n1929 ) | ( ~n1882 & n1929 ) ;
  assign n1931 = ~n1060 & n1930 ;
  assign n1932 = ( n1931 & ~n1001 ) | ( n1931 & n1580 ) | ( ~n1001 & n1580 ) ;
  assign n1933 = ( n1932 & ~n1580 ) | ( n1932 & 1'b0 ) | ( ~n1580 & 1'b0 ) ;
  assign n1934 = ( n789 & ~n1876 ) | ( n789 & n1933 ) | ( ~n1876 & n1933 ) ;
  assign n1935 = ~n789 & n1934 ;
  assign n1936 = ( n672 & ~n222 ) | ( n672 & n1935 ) | ( ~n222 & n1935 ) ;
  assign n1937 = ~n672 & n1936 ;
  assign n1938 = ( n132 & ~n549 ) | ( n132 & n1937 ) | ( ~n549 & n1937 ) ;
  assign n1939 = ~n132 & n1938 ;
  assign n1940 = ~n617 & n1939 ;
  assign n1941 = ( n665 & ~n362 ) | ( n665 & n714 ) | ( ~n362 & n714 ) ;
  assign n1942 = n362 | n1941 ;
  assign n1943 = ( n188 & ~n561 ) | ( n188 & n1942 ) | ( ~n561 & n1942 ) ;
  assign n1944 = n561 | n1943 ;
  assign n1945 = ( n266 & ~n104 ) | ( n266 & n1944 ) | ( ~n104 & n1944 ) ;
  assign n1946 = n104 | n1945 ;
  assign n1947 = ( n336 & ~n643 ) | ( n336 & n1946 ) | ( ~n643 & n1946 ) ;
  assign n1948 = n643 | n1947 ;
  assign n1949 = n61 | n138 ;
  assign n1950 = ( n1064 & ~n241 ) | ( n1064 & n1949 ) | ( ~n241 & n1949 ) ;
  assign n1951 = n241 | n1950 ;
  assign n1952 = ( n206 & ~n456 ) | ( n206 & n1951 ) | ( ~n456 & n1951 ) ;
  assign n1953 = n456 | n1952 ;
  assign n1954 = n560 | n1953 ;
  assign n1955 = n239 | n432 ;
  assign n1956 = n65 | n244 ;
  assign n1957 = ( n404 & ~n720 ) | ( n404 & n1956 ) | ( ~n720 & n1956 ) ;
  assign n1958 = n720 | n1957 ;
  assign n1959 = n347 | n1958 ;
  assign n1960 = n118 | n275 ;
  assign n1961 = ( n1959 & ~n1569 ) | ( n1959 & n1960 ) | ( ~n1569 & n1960 ) ;
  assign n1962 = n1569 | n1961 ;
  assign n1963 = n222 | n353 ;
  assign n1964 = ( n425 & ~n345 ) | ( n425 & n1963 ) | ( ~n345 & n1963 ) ;
  assign n1965 = n345 | n1964 ;
  assign n1966 = ( n80 & ~n232 ) | ( n80 & n1965 ) | ( ~n232 & n1965 ) ;
  assign n1967 = n232 | n1966 ;
  assign n1968 = ( n618 & ~n300 ) | ( n618 & n1967 ) | ( ~n300 & n1967 ) ;
  assign n1969 = n300 | n1968 ;
  assign n1970 = ( n135 & ~n117 ) | ( n135 & n1969 ) | ( ~n117 & n1969 ) ;
  assign n1971 = n117 | n1970 ;
  assign n1972 = ( n1270 & ~n1962 ) | ( n1270 & n1971 ) | ( ~n1962 & n1971 ) ;
  assign n1973 = ( n1962 & ~n75 ) | ( n1962 & n1972 ) | ( ~n75 & n1972 ) ;
  assign n1974 = n75 | n1973 ;
  assign n1975 = ( n1974 & ~n910 ) | ( n1974 & n1461 ) | ( ~n910 & n1461 ) ;
  assign n1976 = n910 | n1975 ;
  assign n1977 = ( n792 & ~n124 ) | ( n792 & n1976 ) | ( ~n124 & n1976 ) ;
  assign n1978 = n124 | n1977 ;
  assign n1979 = ( n451 & ~n417 ) | ( n451 & n1978 ) | ( ~n417 & n1978 ) ;
  assign n1980 = n417 | n1979 ;
  assign n1981 = ( n49 & ~n86 ) | ( n49 & n1980 ) | ( ~n86 & n1980 ) ;
  assign n1982 = n86 | n1981 ;
  assign n1991 = n77 | n403 ;
  assign n1992 = n122 | n259 ;
  assign n1993 = n485 | n1992 ;
  assign n1994 = ( n1398 & ~n1991 ) | ( n1398 & n1993 ) | ( ~n1991 & n1993 ) ;
  assign n1995 = n1991 | n1994 ;
  assign n1983 = n217 | n255 ;
  assign n1984 = n332 | n1983 ;
  assign n1985 = ( n906 & ~n130 ) | ( n906 & n1984 ) | ( ~n130 & n1984 ) ;
  assign n1986 = n130 | n1985 ;
  assign n1987 = ( n452 & ~n761 ) | ( n452 & n1986 ) | ( ~n761 & n1986 ) ;
  assign n1988 = n761 | n1987 ;
  assign n1989 = ( n484 & ~n524 ) | ( n484 & n1988 ) | ( ~n524 & n1988 ) ;
  assign n1990 = ( n484 & ~n1989 ) | ( n484 & 1'b0 ) | ( ~n1989 & 1'b0 ) ;
  assign n1996 = ( n1626 & ~n1995 ) | ( n1626 & n1990 ) | ( ~n1995 & n1990 ) ;
  assign n1997 = ~n1626 & n1996 ;
  assign n1998 = ( n1494 & ~n1512 ) | ( n1494 & n1997 ) | ( ~n1512 & n1997 ) ;
  assign n1999 = ~n1494 & n1998 ;
  assign n2000 = ( n675 & ~n912 ) | ( n675 & n1999 ) | ( ~n912 & n1999 ) ;
  assign n2001 = ( n1490 & ~n675 ) | ( n1490 & n2000 ) | ( ~n675 & n2000 ) ;
  assign n2002 = ~n1490 & n2001 ;
  assign n2003 = ( n409 & ~n789 ) | ( n409 & n2002 ) | ( ~n789 & n2002 ) ;
  assign n2004 = ~n409 & n2003 ;
  assign n2005 = ( n168 & ~n384 ) | ( n168 & n2004 ) | ( ~n384 & n2004 ) ;
  assign n2006 = ~n168 & n2005 ;
  assign n2007 = ( n129 & ~n2006 ) | ( n129 & n644 ) | ( ~n2006 & n644 ) ;
  assign n2008 = ( n644 & ~n2007 ) | ( n644 & 1'b0 ) | ( ~n2007 & 1'b0 ) ;
  assign n2009 = ~n95 & n2008 ;
  assign n2010 = ( n483 & ~n164 ) | ( n483 & n1073 ) | ( ~n164 & n1073 ) ;
  assign n2011 = ~n483 & n2010 ;
  assign n2012 = ( n2009 & n1982 ) | ( n2009 & n2011 ) | ( n1982 & n2011 ) ;
  assign n2013 = ( n1955 & ~n1982 ) | ( n1955 & n2012 ) | ( ~n1982 & n2012 ) ;
  assign n2014 = ~n1955 & n2013 ;
  assign n2015 = ( n1948 & ~n1954 ) | ( n1948 & n2014 ) | ( ~n1954 & n2014 ) ;
  assign n2016 = ( n1679 & ~n1948 ) | ( n1679 & n2015 ) | ( ~n1948 & n2015 ) ;
  assign n2017 = ~n1679 & n2016 ;
  assign n2018 = ( n257 & ~n461 ) | ( n257 & n2017 ) | ( ~n461 & n2017 ) ;
  assign n2019 = ~n257 & n2018 ;
  assign n2020 = ( n268 & ~n418 ) | ( n268 & n2019 ) | ( ~n418 & n2019 ) ;
  assign n2021 = ~n268 & n2020 ;
  assign n2022 = ~n148 & n2021 ;
  assign n2023 = n425 | n711 ;
  assign n2024 = n663 | n2023 ;
  assign n2025 = ( n222 & ~n812 ) | ( n222 & n2024 ) | ( ~n812 & n2024 ) ;
  assign n2026 = n812 | n2025 ;
  assign n2027 = ( n155 & ~n161 ) | ( n155 & n2026 ) | ( ~n161 & n2026 ) ;
  assign n2028 = n161 | n2027 ;
  assign n2029 = n168 | n451 ;
  assign n2030 = n333 | n460 ;
  assign n2031 = ( n405 & ~n49 ) | ( n405 & n2030 ) | ( ~n49 & n2030 ) ;
  assign n2032 = n49 | n2031 ;
  assign n2033 = n99 | n2032 ;
  assign n2044 = n104 | n554 ;
  assign n2034 = n561 | n627 ;
  assign n2035 = n167 | n788 ;
  assign n2036 = n195 | n735 ;
  assign n2037 = ( n2035 & ~n2034 ) | ( n2035 & n2036 ) | ( ~n2034 & n2036 ) ;
  assign n2038 = ( n2034 & ~n374 ) | ( n2034 & n2037 ) | ( ~n374 & n2037 ) ;
  assign n2039 = n374 | n2038 ;
  assign n2040 = ( n797 & ~n122 ) | ( n797 & n2039 ) | ( ~n122 & n2039 ) ;
  assign n2041 = n122 | n2040 ;
  assign n2042 = ( n457 & ~n2041 ) | ( n457 & n484 ) | ( ~n2041 & n484 ) ;
  assign n2043 = ~n457 & n2042 ;
  assign n2045 = ( n2033 & ~n2044 ) | ( n2033 & n2043 ) | ( ~n2044 & n2043 ) ;
  assign n2046 = ( n1498 & ~n2033 ) | ( n1498 & n2045 ) | ( ~n2033 & n2045 ) ;
  assign n2047 = ~n1498 & n2046 ;
  assign n2048 = ( n2028 & ~n2029 ) | ( n2028 & n2047 ) | ( ~n2029 & n2047 ) ;
  assign n2049 = ( n842 & ~n2028 ) | ( n842 & n2048 ) | ( ~n2028 & n2048 ) ;
  assign n2050 = ~n842 & n2049 ;
  assign n2051 = ( n58 & ~n477 ) | ( n58 & n2050 ) | ( ~n477 & n2050 ) ;
  assign n2052 = ~n58 & n2051 ;
  assign n2053 = ( n267 & ~n718 ) | ( n267 & n2052 ) | ( ~n718 & n2052 ) ;
  assign n2054 = ~n267 & n2053 ;
  assign n2055 = ( n332 & ~n403 ) | ( n332 & n2054 ) | ( ~n403 & n2054 ) ;
  assign n2056 = ~n332 & n2055 ;
  assign n2057 = ( n334 & ~n630 ) | ( n334 & n2056 ) | ( ~n630 & n2056 ) ;
  assign n2058 = ~n334 & n2057 ;
  assign n2059 = ~n141 & n2058 ;
  assign n2060 = ( n358 & ~n240 ) | ( n358 & n607 ) | ( ~n240 & n607 ) ;
  assign n2061 = n240 | n2060 ;
  assign n2062 = n89 | n793 ;
  assign n2063 = n258 | n475 ;
  assign n2064 = n137 | n2063 ;
  assign n2065 = ( n2062 & ~n2061 ) | ( n2062 & n2064 ) | ( ~n2061 & n2064 ) ;
  assign n2066 = ( n813 & n2061 ) | ( n813 & n2065 ) | ( n2061 & n2065 ) ;
  assign n2067 = ( n813 & ~n2066 ) | ( n813 & 1'b0 ) | ( ~n2066 & 1'b0 ) ;
  assign n2068 = ( n69 & ~n106 ) | ( n69 & n2067 ) | ( ~n106 & n2067 ) ;
  assign n2069 = ~n69 & n2068 ;
  assign n2070 = ( n194 & ~n52 ) | ( n194 & n2069 ) | ( ~n52 & n2069 ) ;
  assign n2071 = ~n194 & n2070 ;
  assign n2072 = ( n382 & ~n232 ) | ( n382 & n2071 ) | ( ~n232 & n2071 ) ;
  assign n2073 = ~n382 & n2072 ;
  assign n2074 = ~n93 & n2073 ;
  assign n2075 = n162 | n349 ;
  assign n2076 = n118 | n2075 ;
  assign n2077 = ( n531 & ~n372 ) | ( n531 & n2076 ) | ( ~n372 & n2076 ) ;
  assign n2078 = n372 | n2077 ;
  assign n2079 = ( n169 & ~n299 ) | ( n169 & n2078 ) | ( ~n299 & n2078 ) ;
  assign n2080 = n299 | n2079 ;
  assign n2081 = n213 | n2080 ;
  assign n2082 = n39 | n814 ;
  assign n2085 = n273 | n362 ;
  assign n2086 = ( n646 & ~n404 ) | ( n646 & n2085 ) | ( ~n404 & n2085 ) ;
  assign n2087 = n404 | n2086 ;
  assign n2088 = n714 | n792 ;
  assign n2089 = ( n568 & ~n239 ) | ( n568 & n2088 ) | ( ~n239 & n2088 ) ;
  assign n2090 = n239 | n2089 ;
  assign n2091 = n190 | n734 ;
  assign n2092 = n117 | n2091 ;
  assign n2093 = ( n765 & ~n160 ) | ( n765 & n948 ) | ( ~n160 & n948 ) ;
  assign n2094 = n160 | n2093 ;
  assign n2095 = ( n2092 & ~n2090 ) | ( n2092 & n2094 ) | ( ~n2090 & n2094 ) ;
  assign n2096 = n2090 | n2095 ;
  assign n2097 = ( n1071 & ~n2087 ) | ( n1071 & n2096 ) | ( ~n2087 & n2096 ) ;
  assign n2098 = ( n2087 & ~n1923 ) | ( n2087 & n2097 ) | ( ~n1923 & n2097 ) ;
  assign n2099 = n1923 | n2098 ;
  assign n2083 = ( n193 & n418 ) | ( n193 & n786 ) | ( n418 & n786 ) ;
  assign n2084 = ( n786 & ~n2083 ) | ( n786 & 1'b0 ) | ( ~n2083 & 1'b0 ) ;
  assign n2100 = ( n2082 & ~n2099 ) | ( n2082 & n2084 ) | ( ~n2099 & n2084 ) ;
  assign n2101 = ~n2082 & n2100 ;
  assign n2102 = ( n337 & ~n1703 ) | ( n337 & n2101 ) | ( ~n1703 & n2101 ) ;
  assign n2103 = ( n494 & ~n337 ) | ( n494 & n2102 ) | ( ~n337 & n2102 ) ;
  assign n2104 = ~n494 & n2103 ;
  assign n2105 = ~n424 & n2104 ;
  assign n2106 = n675 | n1808 ;
  assign n2107 = ( n666 & ~n556 ) | ( n666 & n2106 ) | ( ~n556 & n2106 ) ;
  assign n2108 = n556 | n2107 ;
  assign n2109 = n101 | n151 ;
  assign n2110 = n196 | n2109 ;
  assign n2111 = ( n344 & ~n678 ) | ( n344 & 1'b0 ) | ( ~n678 & 1'b0 ) ;
  assign n2112 = ~n559 & n2111 ;
  assign n2113 = ( n1809 & ~n2110 ) | ( n1809 & n2112 ) | ( ~n2110 & n2112 ) ;
  assign n2114 = ~n1809 & n2113 ;
  assign n2115 = ( n619 & ~n2108 ) | ( n619 & n2114 ) | ( ~n2108 & n2114 ) ;
  assign n2116 = ~n619 & n2115 ;
  assign n2117 = ( n2081 & n2105 ) | ( n2081 & n2116 ) | ( n2105 & n2116 ) ;
  assign n2118 = ~n2081 & n2117 ;
  assign n2119 = ( n530 & n2074 ) | ( n530 & n2118 ) | ( n2074 & n2118 ) ;
  assign n2120 = ~n530 & n2119 ;
  assign n2121 = ( n2059 & n1884 ) | ( n2059 & n2120 ) | ( n1884 & n2120 ) ;
  assign n2122 = ~n1884 & n2121 ;
  assign n2123 = ( n259 & ~n947 ) | ( n259 & n2122 ) | ( ~n947 & n2122 ) ;
  assign n2124 = ~n259 & n2123 ;
  assign n2125 = ( n373 & ~n233 ) | ( n373 & n2124 ) | ( ~n233 & n2124 ) ;
  assign n2126 = ~n373 & n2125 ;
  assign n2127 = ~n351 &  n2126 ;
  assign n2128 = n232 | n711 ;
  assign n2129 = n947 | n1494 ;
  assign n2130 = n376 | n2129 ;
  assign n2131 = ( n1778 & ~n1715 ) | ( n1778 & n2130 ) | ( ~n1715 & n2130 ) ;
  assign n2132 = n1715 | n2131 ;
  assign n2133 = n619 | n2132 ;
  assign n2134 = ( n1061 & ~n2128 ) | ( n1061 & n2133 ) | ( ~n2128 & n2133 ) ;
  assign n2135 = ( n1819 & n2134 ) | ( n1819 & n2128 ) | ( n2134 & n2128 ) ;
  assign n2136 = ( n1819 & ~n2135 ) | ( n1819 & 1'b0 ) | ( ~n2135 & 1'b0 ) ;
  assign n2137 = ( n374 & ~n2136 ) | ( n374 & n813 ) | ( ~n2136 & n813 ) ;
  assign n2138 = ( n813 & ~n2137 ) | ( n813 & 1'b0 ) | ( ~n2137 & 1'b0 ) ;
  assign n2139 = ( n61 & ~n277 ) | ( n61 & n2138 ) | ( ~n277 & n2138 ) ;
  assign n2140 = ~n61 & n2139 ;
  assign n2141 = ( n65 & ~n206 ) | ( n65 & n2140 ) | ( ~n206 & n2140 ) ;
  assign n2142 = ~n65 & n2141 ;
  assign n2143 = ( n484 & ~n644 ) | ( n484 & n2142 ) | ( ~n644 & n2142 ) ;
  assign n2144 = n644 &  n2143 ;
  assign n2145 = ( n136 & ~n240 ) | ( n136 & n2144 ) | ( ~n240 & n2144 ) ;
  assign n2146 = ~n136 & n2145 ;
  assign n2147 = ~n666 & n2146 ;
  assign n2158 = ( n222 & ~n138 ) | ( n222 & n275 ) | ( ~n138 & n275 ) ;
  assign n2159 = ( n138 & ~n456 ) | ( n138 & n2158 ) | ( ~n456 & n2158 ) ;
  assign n2160 = n456 | n2159 ;
  assign n2161 = ( n403 & ~n214 ) | ( n403 & n2160 ) | ( ~n214 & n2160 ) ;
  assign n2162 = n214 | n2161 ;
  assign n2155 = n161 | n569 ;
  assign n2156 = ( n572 & ~n86 ) | ( n572 & n2155 ) | ( ~n86 & n2155 ) ;
  assign n2157 = n86 | n2156 ;
  assign n2163 = n49 | n490 ;
  assign n2164 = n225 | n2163 ;
  assign n2165 = ( n2162 & ~n2157 ) | ( n2162 & n2164 ) | ( ~n2157 & n2164 ) ;
  assign n2166 = ( n2165 & ~n1984 ) | ( n2165 & n2157 ) | ( ~n1984 & n2157 ) ;
  assign n2167 = n1984 | n2166 ;
  assign n2168 = ( n2105 & ~n2167 ) | ( n2105 & n1806 ) | ( ~n2167 & n1806 ) ;
  assign n2169 = ~n1806 & n2168 ;
  assign n2148 = n123 | n334 ;
  assign n2149 = n155 | n2148 ;
  assign n2150 = ( n852 & ~n775 ) | ( n852 & n2149 ) | ( ~n775 & n2149 ) ;
  assign n2151 = n775 | n2150 ;
  assign n2152 = ( n221 & ~n453 ) | ( n221 & n2151 ) | ( ~n453 & n2151 ) ;
  assign n2153 = n453 | n2152 ;
  assign n2154 = n252 | n2153 ;
  assign n2170 = ( n2147 & ~n2169 ) | ( n2147 & n2154 ) | ( ~n2169 & n2154 ) ;
  assign n2171 = ( n2147 & ~n2170 ) | ( n2147 & 1'b0 ) | ( ~n2170 & 1'b0 ) ;
  assign n2172 = ( n341 & ~n1107 ) | ( n341 & n2171 ) | ( ~n1107 & n2171 ) ;
  assign n2173 = ~n341 & n2172 ;
  assign n2174 = ( n132 & ~n787 ) | ( n132 & n2173 ) | ( ~n787 & n2173 ) ;
  assign n2175 = ~n132 & n2174 ;
  assign n2176 = ( n237 & ~n2175 ) | ( n237 & n623 ) | ( ~n2175 & n623 ) ;
  assign n2177 = ( n623 & ~n2176 ) | ( n623 & 1'b0 ) | ( ~n2176 & 1'b0 ) ;
  assign n2178 = ~n285 &  n2177 ;
  assign n2179 = n191 | n796 ;
  assign n2180 = ( n132 & ~n101 ) | ( n132 & n2179 ) | ( ~n101 & n2179 ) ;
  assign n2181 = n101 | n2180 ;
  assign n2182 = ( n434 & ~n372 ) | ( n434 & n2181 ) | ( ~n372 & n2181 ) ;
  assign n2183 = n372 | n2182 ;
  assign n2184 = ( n139 & ~n411 ) | ( n139 & n2183 ) | ( ~n411 & n2183 ) ;
  assign n2185 = n411 | n2184 ;
  assign n2186 = n356 | n2185 ;
  assign n2187 = n554 | n814 ;
  assign n2188 = ~n86 & n524 ;
  assign n2189 = ~n1207 & n2188 ;
  assign n2190 = ~n568 & n2189 ;
  assign n2191 = n120 | n630 ;
  assign n2192 = n358 | n406 ;
  assign n2193 = ( n1327 & n1764 ) | ( n1327 & n1831 ) | ( n1764 & n1831 ) ;
  assign n2194 = ( n1764 & ~n2193 ) | ( n1764 & 1'b0 ) | ( ~n2193 & 1'b0 ) ;
  assign n2195 = ( n677 & ~n2192 ) | ( n677 & n2194 ) | ( ~n2192 & n2194 ) ;
  assign n2196 = ( n2191 & ~n677 ) | ( n2191 & n2195 ) | ( ~n677 & n2195 ) ;
  assign n2197 = ~n2191 & n2196 ;
  assign n2198 = ( n460 & ~n233 ) | ( n460 & n2197 ) | ( ~n233 & n2197 ) ;
  assign n2199 = ~n460 & n2198 ;
  assign n2200 = ( n529 & ~n540 ) | ( n529 & n2199 ) | ( ~n540 & n2199 ) ;
  assign n2201 = ~n529 & n2200 ;
  assign n2202 = ( n405 & ~n452 ) | ( n405 & n454 ) | ( ~n452 & n454 ) ;
  assign n2203 = ( n452 & ~n75 ) | ( n452 & n2202 ) | ( ~n75 & n2202 ) ;
  assign n2204 = n75 | n2203 ;
  assign n2205 = n459 | n2204 ;
  assign n2206 = n275 | n721 ;
  assign n2207 = ( n206 & ~n429 ) | ( n206 & n346 ) | ( ~n429 & n346 ) ;
  assign n2208 = n429 | n2207 ;
  assign n2209 = n259 | n620 ;
  assign n2210 = n812 | n2209 ;
  assign n2211 = ( n2208 & ~n2206 ) | ( n2208 & n2210 ) | ( ~n2206 & n2210 ) ;
  assign n2212 = ( n2206 & ~n2062 ) | ( n2206 & n2211 ) | ( ~n2062 & n2211 ) ;
  assign n2213 = n2062 | n2212 ;
  assign n2214 = ( n2201 & n2205 ) | ( n2201 & n2213 ) | ( n2205 & n2213 ) ;
  assign n2215 = ( n2201 & ~n2214 ) | ( n2201 & 1'b0 ) | ( ~n2214 & 1'b0 ) ;
  assign n2216 = ( n1493 & n2190 ) | ( n1493 & n2215 ) | ( n2190 & n2215 ) ;
  assign n2217 = ~n1493 & n2216 ;
  assign n2218 = ( n716 & ~n2187 ) | ( n716 & n2217 ) | ( ~n2187 & n2217 ) ;
  assign n2219 = ( n1511 & ~n716 ) | ( n1511 & n2218 ) | ( ~n716 & n2218 ) ;
  assign n2220 = ~n1511 & n2219 ;
  assign n2221 = ( n792 & ~n127 ) | ( n792 & n2220 ) | ( ~n127 & n2220 ) ;
  assign n2222 = ~n792 & n2221 ;
  assign n2223 = ( n333 & ~n373 ) | ( n333 & n2222 ) | ( ~n373 & n2222 ) ;
  assign n2224 = ~n333 & n2223 ;
  assign n2225 = ( n226 & ~n80 ) | ( n226 & n2224 ) | ( ~n80 & n2224 ) ;
  assign n2226 = ~n226 & n2225 ;
  assign n2227 = ~n476 & n2226 ;
  assign n2228 = n571 | n911 ;
  assign n2229 = n118 | n2228 ;
  assign n2230 = ( n491 & ~n1306 ) | ( n491 & n2229 ) | ( ~n1306 & n2229 ) ;
  assign n2231 = n1306 | n2230 ;
  assign n2232 = ( n788 & ~n244 ) | ( n788 & n2231 ) | ( ~n244 & n2231 ) ;
  assign n2233 = n244 | n2232 ;
  assign n2234 = ( n237 & ~n216 ) | ( n237 & n2233 ) | ( ~n216 & n2233 ) ;
  assign n2235 = n216 | n2234 ;
  assign n2236 = ( n77 & n343 ) | ( n77 & n2235 ) | ( n343 & n2235 ) ;
  assign n2237 = ( n343 & ~n2236 ) | ( n343 & 1'b0 ) | ( ~n2236 & 1'b0 ) ;
  assign n2238 = ( n664 & ~n95 ) | ( n664 & n2237 ) | ( ~n95 & n2237 ) ;
  assign n2239 = ~n664 & n2238 ;
  assign n2240 = ~n410 & n2239 ;
  assign n2241 = n382 | n384 ;
  assign n2242 = n526 | n2241 ;
  assign n2243 = ( n260 & ~n274 ) | ( n260 & n2242 ) | ( ~n274 & n2242 ) ;
  assign n2244 = n274 | n2243 ;
  assign n2245 = ( n214 & ~n737 ) | ( n214 & n2244 ) | ( ~n737 & n2244 ) ;
  assign n2246 = n737 | n2245 ;
  assign n2247 = n670 | n2246 ;
  assign n2248 = n192 | n787 ;
  assign n2249 = ( n149 & ~n148 ) | ( n149 & n2248 ) | ( ~n148 & n2248 ) ;
  assign n2250 = n148 | n2249 ;
  assign n2251 = ( n340 & ~n39 ) | ( n340 & n2250 ) | ( ~n39 & n2250 ) ;
  assign n2252 = n39 | n2251 ;
  assign n2253 = n239 | n271 ;
  assign n2254 = n99 | n2253 ;
  assign n2255 = ( n2091 & ~n150 ) | ( n2091 & n2254 ) | ( ~n150 & n2254 ) ;
  assign n2256 = n150 | n2255 ;
  assign n2257 = ( n130 & ~n745 ) | ( n130 & n2256 ) | ( ~n745 & n2256 ) ;
  assign n2258 = n745 | n2257 ;
  assign n2259 = ( n559 & ~n549 ) | ( n559 & n2258 ) | ( ~n549 & n2258 ) ;
  assign n2260 = n549 | n2259 ;
  assign n2261 = ( n663 & ~n478 ) | ( n663 & n2260 ) | ( ~n478 & n2260 ) ;
  assign n2262 = n478 | n2261 ;
  assign n2263 = n122 | n257 ;
  assign n2264 = n627 | n1244 ;
  assign n2265 = ( n623 & ~n714 ) | ( n623 & 1'b0 ) | ( ~n714 & 1'b0 ) ;
  assign n2266 = ~n276 & n2265 ;
  assign n2267 = ( n2263 & ~n2264 ) | ( n2263 & n2266 ) | ( ~n2264 & n2266 ) ;
  assign n2268 = ~n2263 & n2267 ;
  assign n2269 = ( n2252 & ~n2262 ) | ( n2252 & n2268 ) | ( ~n2262 & n2268 ) ;
  assign n2270 = ( n1762 & ~n2252 ) | ( n1762 & n2269 ) | ( ~n2252 & n2269 ) ;
  assign n2271 = ~n1762 & n2270 ;
  assign n2272 = ( n789 & ~n2247 ) | ( n789 & n2271 ) | ( ~n2247 & n2271 ) ;
  assign n2273 = ~n789 & n2272 ;
  assign n2274 = ( n678 & ~n359 ) | ( n678 & n2273 ) | ( ~n359 & n2273 ) ;
  assign n2275 = ~n678 & n2274 ;
  assign n2276 = ( n58 & ~n349 ) | ( n58 & n2275 ) | ( ~n349 & n2275 ) ;
  assign n2277 = ~n58 & n2276 ;
  assign n2278 = ~n744 & n2277 ;
  assign n2279 = n277 | n761 ;
  assign n2280 = ( n736 & ~n1827 ) | ( n736 & n2279 ) | ( ~n1827 & n2279 ) ;
  assign n2281 = n1827 | n2280 ;
  assign n2282 = ( n2240 & ~n2278 ) | ( n2240 & n2281 ) | ( ~n2278 & n2281 ) ;
  assign n2283 = ( n2240 & ~n2282 ) | ( n2240 & 1'b0 ) | ( ~n2282 & 1'b0 ) ;
  assign n2284 = ( n794 & ~n2283 ) | ( n794 & n2227 ) | ( ~n2283 & n2227 ) ;
  assign n2285 = ( n2227 & ~n2284 ) | ( n2227 & 1'b0 ) | ( ~n2284 & 1'b0 ) ;
  assign n2286 = ( n947 & ~n2186 ) | ( n947 & n2285 ) | ( ~n2186 & n2285 ) ;
  assign n2287 = ~n947 & n2286 ;
  assign n2288 = ( n2287 & ~n70 ) | ( n2287 & n376 ) | ( ~n70 & n376 ) ;
  assign n2289 = ( n2288 & ~n376 ) | ( n2288 & 1'b0 ) | ( ~n376 & 1'b0 ) ;
  assign n2290 = ( n778 & ~n602 ) | ( n778 & n2289 ) | ( ~n602 & n2289 ) ;
  assign n2291 = ~n778 & n2290 ;
  assign n2292 = ( n49 & ~n494 ) | ( n49 & n2291 ) | ( ~n494 & n2291 ) ;
  assign n2293 = ~n49 & n2292 ;
  assign n2294 = ( n342 & ~n104 ) | ( n342 & n2293 ) | ( ~n104 & n2293 ) ;
  assign n2295 = ~n342 & n2294 ;
  assign n2296 = ~n332 &  n2295 ;
  assign n2297 = ~n241 & n343 ;
  assign n2298 = ~n228 & n2297 ;
  assign n2299 = n101 | n418 ;
  assign n2300 = ( n137 & ~n162 ) | ( n137 & n2299 ) | ( ~n162 & n2299 ) ;
  assign n2301 = n162 | n2300 ;
  assign n2302 = ( n2298 & n455 ) | ( n2298 & n2301 ) | ( n455 & n2301 ) ;
  assign n2303 = ( n61 & ~n2302 ) | ( n61 & n2298 ) | ( ~n2302 & n2298 ) ;
  assign n2304 = ~n61 & n2303 ;
  assign n2305 = ( n284 & ~n206 ) | ( n284 & n2304 ) | ( ~n206 & n2304 ) ;
  assign n2306 = ~n284 & n2305 ;
  assign n2307 = ~n909 & n2306 ;
  assign n2308 = n104 | n260 ;
  assign n2309 = n429 | n631 ;
  assign n2310 = ( n277 & ~n126 ) | ( n277 & n2309 ) | ( ~n126 & n2309 ) ;
  assign n2311 = n126 | n2310 ;
  assign n2312 = ( n403 & ~n460 ) | ( n403 & n2311 ) | ( ~n460 & n2311 ) ;
  assign n2313 = n460 | n2312 ;
  assign n2314 = n150 | n253 ;
  assign n2315 = ( n197 & n266 ) | ( n197 & n2314 ) | ( n266 & n2314 ) ;
  assign n2316 = ( n197 & ~n2315 ) | ( n197 & 1'b0 ) | ( ~n2315 & 1'b0 ) ;
  assign n2317 = n187 | n793 ;
  assign n2318 = ( n623 & ~n2317 ) | ( n623 & 1'b0 ) | ( ~n2317 & 1'b0 ) ;
  assign n2319 = ( n1855 & ~n1003 ) | ( n1855 & n2318 ) | ( ~n1003 & n2318 ) ;
  assign n2320 = ~n1855 & n2319 ;
  assign n2321 = ( n576 & ~n387 ) | ( n576 & n2320 ) | ( ~n387 & n2320 ) ;
  assign n2322 = ~n576 & n2321 ;
  assign n2323 = ( n2313 & n2316 ) | ( n2313 & n2322 ) | ( n2316 & n2322 ) ;
  assign n2324 = ~n2313 & n2323 ;
  assign n2325 = ( n341 & ~n2308 ) | ( n341 & n2324 ) | ( ~n2308 & n2324 ) ;
  assign n2326 = ~n341 & n2325 ;
  assign n2327 = ( n106 & ~n337 ) | ( n106 & n2326 ) | ( ~n337 & n2326 ) ;
  assign n2328 = ~n106 & n2327 ;
  assign n2329 = ( n350 & ~n234 ) | ( n350 & n2328 ) | ( ~n234 & n2328 ) ;
  assign n2330 = ~n350 & n2329 ;
  assign n2331 = ~n618 & n2330 ;
  assign n2332 = n410 | n540 ;
  assign n2333 = ( n1399 & ~n1796 ) | ( n1399 & n2332 ) | ( ~n1796 & n2332 ) ;
  assign n2334 = n1796 | n2333 ;
  assign n2335 = ( n258 & ~n208 ) | ( n258 & n2334 ) | ( ~n208 & n2334 ) ;
  assign n2336 = n208 | n2335 ;
  assign n2337 = ( n404 & ~n269 ) | ( n404 & n2336 ) | ( ~n269 & n2336 ) ;
  assign n2338 = n269 | n2337 ;
  assign n2339 = ( n558 & ~n151 ) | ( n558 & n2338 ) | ( ~n151 & n2338 ) ;
  assign n2340 = n151 | n2339 ;
  assign n2341 = ( n353 & ~n141 ) | ( n353 & n2340 ) | ( ~n141 & n2340 ) ;
  assign n2342 = n141 | n2341 ;
  assign n2343 = n139 | n424 ;
  assign n2344 = ( n568 & ~n459 ) | ( n568 & n2343 ) | ( ~n459 & n2343 ) ;
  assign n2345 = n459 | n2344 ;
  assign n2346 = n233 | n561 ;
  assign n2347 = n274 | n358 ;
  assign n2348 = n362 | n603 ;
  assign n2349 = ( n384 & ~n432 ) | ( n384 & n2348 ) | ( ~n432 & n2348 ) ;
  assign n2350 = n432 | n2349 ;
  assign n2351 = ( n2347 & ~n2157 ) | ( n2347 & n2350 ) | ( ~n2157 & n2350 ) ;
  assign n2352 = n2157 | n2351 ;
  assign n2353 = ( n2346 & ~n2029 ) | ( n2346 & n2352 ) | ( ~n2029 & n2352 ) ;
  assign n2354 = n2029 | n2353 ;
  assign n2355 = ( n123 & ~n456 ) | ( n123 & n2354 ) | ( ~n456 & n2354 ) ;
  assign n2356 = n456 | n2355 ;
  assign n2357 = n431 | n2356 ;
  assign n2358 = n243 | n718 ;
  assign n2359 = n382 | n722 ;
  assign n2360 = n485 | n2359 ;
  assign n2361 = ( n799 & ~n2358 ) | ( n799 & n2360 ) | ( ~n2358 & n2360 ) ;
  assign n2362 = ( n2361 & ~n2024 ) | ( n2361 & n2358 ) | ( ~n2024 & n2358 ) ;
  assign n2363 = n2024 | n2362 ;
  assign n2364 = ( n2091 & ~n2357 ) | ( n2091 & n2363 ) | ( ~n2357 & n2363 ) ;
  assign n2365 = ( n2364 & ~n573 ) | ( n2364 & n2357 ) | ( ~n573 & n2357 ) ;
  assign n2366 = n573 | n2365 ;
  assign n2367 = ( n1884 & ~n605 ) | ( n1884 & n2366 ) | ( ~n605 & n2366 ) ;
  assign n2368 = n605 | n2367 ;
  assign n2369 = ( n70 & ~n194 ) | ( n70 & n2368 ) | ( ~n194 & n2368 ) ;
  assign n2370 = n194 | n2369 ;
  assign n2371 = ( n191 & ~n453 ) | ( n191 & n2370 ) | ( ~n453 & n2370 ) ;
  assign n2372 = n453 | n2371 ;
  assign n2373 = ( n354 & ~n484 ) | ( n354 & n2372 ) | ( ~n484 & n2372 ) ;
  assign n2374 = ( n354 & ~n2373 ) | ( n354 & 1'b0 ) | ( ~n2373 & 1'b0 ) ;
  assign n2375 = ( n527 & ~n911 ) | ( n527 & n2374 ) | ( ~n911 & n2374 ) ;
  assign n2376 = ~n527 & n2375 ;
  assign n2377 = n245 | n529 ;
  assign n2378 = n276 | n2377 ;
  assign n2379 = ( n1437 & ~n2376 ) | ( n1437 & n2378 ) | ( ~n2376 & n2378 ) ;
  assign n2380 = ( n1437 & ~n2379 ) | ( n1437 & 1'b0 ) | ( ~n2379 & 1'b0 ) ;
  assign n2381 = ( n2342 & ~n2345 ) | ( n2342 & n2380 ) | ( ~n2345 & n2380 ) ;
  assign n2382 = ~n2342 & n2381 ;
  assign n2383 = ( n2331 & ~n2307 ) | ( n2331 & n2382 ) | ( ~n2307 & n2382 ) ;
  assign n2384 = n2307 &  n2383 ;
  assign n2385 = ( n346 & ~n238 ) | ( n346 & n2384 ) | ( ~n238 & n2384 ) ;
  assign n2386 = ~n346 & n2385 ;
  assign n2387 = ( n788 & ~n125 ) | ( n788 & n2386 ) | ( ~n125 & n2386 ) ;
  assign n2388 = ~n788 & n2387 ;
  assign n2389 = ( n122 & ~n372 ) | ( n122 & n2388 ) | ( ~n372 & n2388 ) ;
  assign n2390 = ~n122 & n2389 ;
  assign n2391 = ( n556 & ~n270 ) | ( n556 & n2390 ) | ( ~n270 & n2390 ) ;
  assign n2392 = ~n556 &  n2391 ;
  assign n2393 = n192 | n345 ;
  assign n2394 = n279 | n2393 ;
  assign n2395 = n213 | n234 ;
  assign n2396 = n1497 | n2313 ;
  assign n2397 = ( n348 & ~n671 ) | ( n348 & n2396 ) | ( ~n671 & n2396 ) ;
  assign n2398 = n671 | n2397 ;
  assign n2399 = ( n239 & ~n556 ) | ( n239 & n2398 ) | ( ~n556 & n2398 ) ;
  assign n2400 = n556 | n2399 ;
  assign n2401 = ( n135 & ~n149 ) | ( n135 & n2400 ) | ( ~n149 & n2400 ) ;
  assign n2402 = n149 | n2401 ;
  assign n2403 = n617 | n2402 ;
  assign n2404 = n425 | n457 ;
  assign n2405 = n454 | n2404 ;
  assign n2406 = ( n206 & ~n232 ) | ( n206 & n2405 ) | ( ~n232 & n2405 ) ;
  assign n2407 = n232 | n2406 ;
  assign n2408 = ( n214 & ~n148 ) | ( n214 & n2407 ) | ( ~n148 & n2407 ) ;
  assign n2409 = n148 | n2408 ;
  assign n2410 = ( n285 & ~n93 ) | ( n285 & n2409 ) | ( ~n93 & n2409 ) ;
  assign n2411 = n93 | n2410 ;
  assign n2412 = n207 | n735 ;
  assign n2413 = n188 | n258 ;
  assign n2414 = n268 | n2413 ;
  assign n2415 = ( n2412 & ~n2411 ) | ( n2412 & n2414 ) | ( ~n2411 & n2414 ) ;
  assign n2416 = n2411 | n2415 ;
  assign n2417 = ( n2403 & ~n667 ) | ( n2403 & n2416 ) | ( ~n667 & n2416 ) ;
  assign n2418 = n667 | n2417 ;
  assign n2419 = ( n777 & ~n886 ) | ( n777 & n2418 ) | ( ~n886 & n2418 ) ;
  assign n2420 = ( n886 & ~n257 ) | ( n886 & n2419 ) | ( ~n257 & n2419 ) ;
  assign n2421 = n257 | n2420 ;
  assign n2422 = ( n105 & n2421 ) | ( n105 & n484 ) | ( n2421 & n484 ) ;
  assign n2423 = ( n484 & ~n2422 ) | ( n484 & 1'b0 ) | ( ~n2422 & 1'b0 ) ;
  assign n2424 = ( n476 & ~n340 ) | ( n476 & n2423 ) | ( ~n340 & n2423 ) ;
  assign n2425 = ~n476 & n2424 ;
  assign n2426 = ~n670 & n2425 ;
  assign n2427 = n122 | n267 ;
  assign n2428 = n233 | n745 ;
  assign n2429 = ( n240 & ~n161 ) | ( n240 & n2428 ) | ( ~n161 & n2428 ) ;
  assign n2430 = n161 | n2429 ;
  assign n2431 = n643 | n2430 ;
  assign n2432 = ( n212 & ~n269 ) | ( n212 & n1062 ) | ( ~n269 & n1062 ) ;
  assign n2433 = n269 | n2432 ;
  assign n2434 = ( n647 & ~n531 ) | ( n647 & n2082 ) | ( ~n531 & n2082 ) ;
  assign n2435 = n531 | n2434 ;
  assign n2436 = ( n2264 & ~n2433 ) | ( n2264 & n2435 ) | ( ~n2433 & n2435 ) ;
  assign n2437 = ( n2433 & ~n1754 ) | ( n2433 & n2436 ) | ( ~n1754 & n2436 ) ;
  assign n2438 = n1754 | n2437 ;
  assign n2439 = ( n607 & ~n2431 ) | ( n607 & n2438 ) | ( ~n2431 & n2438 ) ;
  assign n2440 = ( n2439 & ~n1585 ) | ( n2439 & n2431 ) | ( ~n1585 & n2431 ) ;
  assign n2441 = n1585 | n2440 ;
  assign n2442 = ( n2348 & ~n2427 ) | ( n2348 & n2441 ) | ( ~n2427 & n2441 ) ;
  assign n2443 = ( n2240 & n2442 ) | ( n2240 & n2427 ) | ( n2442 & n2427 ) ;
  assign n2444 = ( n2240 & ~n2443 ) | ( n2240 & 1'b0 ) | ( ~n2443 & 1'b0 ) ;
  assign n2445 = ( n352 & ~n434 ) | ( n352 & n2444 ) | ( ~n434 & n2444 ) ;
  assign n2446 = ( n130 & ~n352 ) | ( n130 & n2445 ) | ( ~n352 & n2445 ) ;
  assign n2447 = ~n130 & n2446 ;
  assign n2448 = ( n572 & ~n91 ) | ( n572 & n2447 ) | ( ~n91 & n2447 ) ;
  assign n2449 = ~n572 & n2448 ;
  assign n2450 = ( n478 & ~n628 ) | ( n478 & n2449 ) | ( ~n628 & n2449 ) ;
  assign n2451 = ~n478 & n2450 ;
  assign n2462 = n125 | n554 ;
  assign n2463 = ( n624 & ~n1072 ) | ( n624 & 1'b0 ) | ( ~n1072 & 1'b0 ) ;
  assign n2464 = ( n452 & ~n2462 ) | ( n452 & n2463 ) | ( ~n2462 & n2463 ) ;
  assign n2465 = ~n452 & n2464 ;
  assign n2466 = ( n356 & ~n526 ) | ( n356 & n2465 ) | ( ~n526 & n2465 ) ;
  assign n2467 = ~n356 & n2466 ;
  assign n2468 = n106 | n141 ;
  assign n2469 = ( n1381 & n2467 ) | ( n1381 & n2468 ) | ( n2467 & n2468 ) ;
  assign n2470 = ( n2467 & ~n2469 ) | ( n2467 & 1'b0 ) | ( ~n2469 & 1'b0 ) ;
  assign n2452 = n408 | n1949 ;
  assign n2453 = ( n679 & ~n124 ) | ( n679 & n2452 ) | ( ~n124 & n2452 ) ;
  assign n2454 = n124 | n2453 ;
  assign n2455 = ( n775 & ~n168 ) | ( n775 & n2454 ) | ( ~n168 & n2454 ) ;
  assign n2456 = n168 | n2455 ;
  assign n2457 = ( n485 & ~n765 ) | ( n485 & n2456 ) | ( ~n765 & n2456 ) ;
  assign n2458 = n765 | n2457 ;
  assign n2459 = ( n228 & ~n560 ) | ( n228 & n2458 ) | ( ~n560 & n2458 ) ;
  assign n2460 = n560 | n2459 ;
  assign n2461 = n358 | n2460 ;
  assign n2471 = ( n2451 & ~n2470 ) | ( n2451 & n2461 ) | ( ~n2470 & n2461 ) ;
  assign n2472 = ( n1686 & ~n2451 ) | ( n1686 & n2471 ) | ( ~n2451 & n2471 ) ;
  assign n2473 = ( n1686 & ~n2472 ) | ( n1686 & 1'b0 ) | ( ~n2472 & 1'b0 ) ;
  assign n2474 = ( n2395 & n2426 ) | ( n2395 & n2473 ) | ( n2426 & n2473 ) ;
  assign n2475 = ~n2395 & n2474 ;
  assign n2476 = ( n1428 & ~n2394 ) | ( n1428 & n2475 ) | ( ~n2394 & n2475 ) ;
  assign n2477 = ~n1428 & n2476 ;
  assign n2478 = ( n411 & ~n2308 ) | ( n411 & n2477 ) | ( ~n2308 & n2477 ) ;
  assign n2479 = ~n411 & n2478 ;
  assign n2480 = ( n190 & ~n405 ) | ( n190 & n2479 ) | ( ~n405 & n2479 ) ;
  assign n2481 = ~n190 & n2480 ;
  assign n2482 = ( n276 & ~n432 ) | ( n276 & n2481 ) | ( ~n432 & n2481 ) ;
  assign n2483 = ~n276 & n2482 ;
  assign n2484 = n454 | n602 ;
  assign n2485 = n281 | n606 ;
  assign n2486 = ( n843 & ~n1107 ) | ( n843 & n2485 ) | ( ~n1107 & n2485 ) ;
  assign n2487 = n1107 | n2486 ;
  assign n2488 = ( n1060 & ~n1493 ) | ( n1060 & n2487 ) | ( ~n1493 & n2487 ) ;
  assign n2489 = n1493 | n2488 ;
  assign n2490 = ( n259 & ~n765 ) | ( n259 & n2489 ) | ( ~n765 & n2489 ) ;
  assign n2491 = n765 | n2490 ;
  assign n2492 = n459 | n2491 ;
  assign n2493 = n120 | n554 ;
  assign n2494 = n169 | n2493 ;
  assign n2495 = n2350 | n2494 ;
  assign n2496 = ( n2492 & ~n1356 ) | ( n2492 & n2495 ) | ( ~n1356 & n2495 ) ;
  assign n2497 = ( n1356 & ~n667 ) | ( n1356 & n2496 ) | ( ~n667 & n2496 ) ;
  assign n2498 = n667 | n2497 ;
  assign n2499 = ( n1762 & ~n1278 ) | ( n1762 & n2498 ) | ( ~n1278 & n2498 ) ;
  assign n2500 = ( n1278 & ~n1484 ) | ( n1278 & n2499 ) | ( ~n1484 & n2499 ) ;
  assign n2501 = n1484 | n2500 ;
  assign n2502 = ( n138 & ~n1152 ) | ( n138 & n2501 ) | ( ~n1152 & n2501 ) ;
  assign n2503 = n1152 | n2502 ;
  assign n2504 = ( n797 & ~n475 ) | ( n797 & n2503 ) | ( ~n475 & n2503 ) ;
  assign n2505 = n475 | n2504 ;
  assign n2506 = n226 | n2505 ;
  assign n2508 = n240 | n425 ;
  assign n2507 = n244 | n800 ;
  assign n2509 = ( n2508 & ~n1512 ) | ( n2508 & n2507 ) | ( ~n1512 & n2507 ) ;
  assign n2510 = n1512 | n2509 ;
  assign n2511 = ( n222 & ~n456 ) | ( n222 & n2510 ) | ( ~n456 & n2510 ) ;
  assign n2512 = n456 | n2511 ;
  assign n2513 = ( n139 & ~n162 ) | ( n139 & n2512 ) | ( ~n162 & n2512 ) ;
  assign n2514 = n162 | n2513 ;
  assign n2515 = n135 | n549 ;
  assign n2516 = n127 | n2515 ;
  assign n2517 = ( n494 & ~n775 ) | ( n494 & n2516 ) | ( ~n775 & n2516 ) ;
  assign n2518 = n775 | n2517 ;
  assign n2519 = n534 | n2518 ;
  assign n2520 = n61 | n237 ;
  assign n2521 = n353 | n2520 ;
  assign n2522 = n242 | n429 ;
  assign n2523 = ( n452 & ~n663 ) | ( n452 & n2522 ) | ( ~n663 & n2522 ) ;
  assign n2524 = n663 | n2523 ;
  assign n2525 = n212 | n2524 ;
  assign n2526 = ( n2521 & ~n2519 ) | ( n2521 & n2525 ) | ( ~n2519 & n2525 ) ;
  assign n2527 = n2519 | n2526 ;
  assign n2528 = ( n2514 & ~n278 ) | ( n2514 & n2527 ) | ( ~n278 & n2527 ) ;
  assign n2529 = n278 | n2528 ;
  assign n2530 = ( n125 & ~n374 ) | ( n125 & n2529 ) | ( ~n374 & n2529 ) ;
  assign n2531 = n374 | n2530 ;
  assign n2532 = ( n216 & ~n230 ) | ( n216 & n2531 ) | ( ~n230 & n2531 ) ;
  assign n2533 = n230 | n2532 ;
  assign n2534 = ( n451 & ~n406 ) | ( n451 & n2533 ) | ( ~n406 & n2533 ) ;
  assign n2535 = n406 | n2534 ;
  assign n2536 = ( n618 & ~n342 ) | ( n618 & n2535 ) | ( ~n342 & n2535 ) ;
  assign n2537 = n342 | n2536 ;
  assign n2538 = ( n643 & ~n356 ) | ( n643 & n2537 ) | ( ~n356 & n2537 ) ;
  assign n2539 = n356 | n2538 ;
  assign n2540 = n260 | n411 ;
  assign n2541 = ( n274 & ~n208 ) | ( n274 & n2540 ) | ( ~n208 & n2540 ) ;
  assign n2542 = n208 | n2541 ;
  assign n2543 = ( n132 & ~n86 ) | ( n132 & n2542 ) | ( ~n86 & n2542 ) ;
  assign n2544 = n86 | n2543 ;
  assign n2545 = n130 | n345 ;
  assign n2546 = ( n137 & ~n118 ) | ( n137 & n2545 ) | ( ~n118 & n2545 ) ;
  assign n2547 = n118 | n2546 ;
  assign n2548 = n270 | n453 ;
  assign n2549 = n350 | n677 ;
  assign n2550 = n214 | n2549 ;
  assign n2551 = ( n2548 & ~n2547 ) | ( n2548 & n2550 ) | ( ~n2547 & n2550 ) ;
  assign n2552 = n2547 | n2551 ;
  assign n2553 = ( n2544 & ~n2539 ) | ( n2544 & n2552 ) | ( ~n2539 & n2552 ) ;
  assign n2554 = n2539 | n2553 ;
  assign n2555 = ( n1283 & ~n2506 ) | ( n1283 & n2554 ) | ( ~n2506 & n2554 ) ;
  assign n2556 = n2506 | n2555 ;
  assign n2557 = ( n2484 & ~n1580 ) | ( n2484 & n2556 ) | ( ~n1580 & n2556 ) ;
  assign n2558 = n1580 | n2557 ;
  assign n2559 = ( n716 & n2558 ) | ( n716 & n1774 ) | ( n2558 & n1774 ) ;
  assign n2560 = ( n1774 & ~n2559 ) | ( n1774 & 1'b0 ) | ( ~n2559 & 1'b0 ) ;
  assign n2561 = ( n1306 & ~n1185 ) | ( n1306 & n2560 ) | ( ~n1185 & n2560 ) ;
  assign n2562 = ~n1306 & n2561 ;
  assign n2563 = ( n269 & ~n2562 ) | ( n269 & n786 ) | ( ~n2562 & n786 ) ;
  assign n2564 = ( n786 & ~n2563 ) | ( n786 & 1'b0 ) | ( ~n2563 & 1'b0 ) ;
  assign n2565 = ( n255 & ~n192 ) | ( n255 & n2564 ) | ( ~n192 & n2564 ) ;
  assign n2566 = ~n255 & n2565 ;
  assign n2567 = ( n529 & ~n492 ) | ( n529 & n2566 ) | ( ~n492 & n2566 ) ;
  assign n2568 = ~n529 & n2567 ;
  assign n2569 = ~n141 &  n2568 ;
  assign n2570 = ~n281 & n623 ;
  assign n2571 = ~n88 & n2570 ;
  assign n2572 = ( n124 & ~n2229 ) | ( n124 & n2571 ) | ( ~n2229 & n2571 ) ;
  assign n2573 = ~n124 & n2572 ;
  assign n2574 = ( n672 & ~n127 ) | ( n672 & n2573 ) | ( ~n127 & n2573 ) ;
  assign n2575 = ~n672 & n2574 ;
  assign n2576 = n347 | n556 ;
  assign n2577 = n106 | n230 ;
  assign n2578 = n39 | n1795 ;
  assign n2579 = ( n81 & ~n1857 ) | ( n81 & n2578 ) | ( ~n1857 & n2578 ) ;
  assign n2580 = n1857 | n2579 ;
  assign n2581 = ( n2394 & ~n2577 ) | ( n2394 & n2580 ) | ( ~n2577 & n2580 ) ;
  assign n2582 = ( n2577 & ~n61 ) | ( n2577 & n2581 ) | ( ~n61 & n2581 ) ;
  assign n2583 = n61 | n2582 ;
  assign n2584 = ( n531 & ~n268 ) | ( n531 & n2583 ) | ( ~n268 & n2583 ) ;
  assign n2585 = n268 | n2584 ;
  assign n2586 = ( n403 & ~n104 ) | ( n403 & n2585 ) | ( ~n104 & n2585 ) ;
  assign n2587 = n104 | n2586 ;
  assign n2588 = n431 | n2587 ;
  assign n2589 = n333 | n493 ;
  assign n2590 = ( n237 & ~n382 ) | ( n237 & n2589 ) | ( ~n382 & n2589 ) ;
  assign n2591 = n382 | n2590 ;
  assign n2592 = n574 | n2591 ;
  assign n2593 = n432 | n787 ;
  assign n2597 = n406 | n735 ;
  assign n2598 = n83 | n2597 ;
  assign n2594 = ~n714 & n813 ;
  assign n2595 = ( n231 & ~n631 ) | ( n231 & n2594 ) | ( ~n631 & n2594 ) ;
  assign n2596 = ~n231 & n2595 ;
  assign n2599 = ( n1810 & ~n2598 ) | ( n1810 & n2596 ) | ( ~n2598 & n2596 ) ;
  assign n2600 = ( n2599 & ~n1810 ) | ( n2599 & 1'b0 ) | ( ~n1810 & 1'b0 ) ;
  assign n2601 = ( n2592 & ~n2593 ) | ( n2592 & n2600 ) | ( ~n2593 & n2600 ) ;
  assign n2602 = ~n2592 & n2601 ;
  assign n2603 = ( n2588 & ~n1215 ) | ( n2588 & n2602 ) | ( ~n1215 & n2602 ) ;
  assign n2604 = ~n2588 & n2603 ;
  assign n2605 = ( n224 & ~n2576 ) | ( n224 & n2604 ) | ( ~n2576 & n2604 ) ;
  assign n2606 = ~n224 & n2605 ;
  assign n2607 = ( n197 & n226 ) | ( n197 & n2606 ) | ( n226 & n2606 ) ;
  assign n2608 = ~n226 & n2607 ;
  assign n2609 = ~n334 & n2608 ;
  assign n2610 = n89 | n136 ;
  assign n2611 = ( n2263 & n2609 ) | ( n2263 & n2610 ) | ( n2609 & n2610 ) ;
  assign n2612 = ( n344 & ~n2609 ) | ( n344 & n2611 ) | ( ~n2609 & n2611 ) ;
  assign n2613 = ( n344 & ~n2612 ) | ( n344 & 1'b0 ) | ( ~n2612 & 1'b0 ) ;
  assign n2614 = ( n245 & ~n243 ) | ( n245 & n2613 ) | ( ~n243 & n2613 ) ;
  assign n2615 = ~n245 & n2614 ;
  assign n2616 = ( n2615 & ~n348 ) | ( n2615 & n745 ) | ( ~n348 & n745 ) ;
  assign n2617 = ( n2616 & ~n745 ) | ( n2616 & 1'b0 ) | ( ~n745 & 1'b0 ) ;
  assign n2618 = ( n165 & ~n205 ) | ( n165 & n2617 ) | ( ~n205 & n2617 ) ;
  assign n2619 = ~n165 & n2618 ;
  assign n2620 = ~n617 & n2619 ;
  assign n2621 = n258 | n720 ;
  assign n2622 = ( n266 & ~n299 ) | ( n266 & n2621 ) | ( ~n299 & n2621 ) ;
  assign n2623 = n299 | n2622 ;
  assign n2624 = ( n353 & ~n666 ) | ( n353 & n2623 ) | ( ~n666 & n2623 ) ;
  assign n2625 = n666 | n2624 ;
  assign n2648 = ( n555 & ~n65 ) | ( n555 & n814 ) | ( ~n65 & n814 ) ;
  assign n2649 = n65 | n2648 ;
  assign n2650 = ( n680 & ~n1732 ) | ( n680 & n2649 ) | ( ~n1732 & n2649 ) ;
  assign n2651 = n1732 | n2650 ;
  assign n2632 = n74 | n494 ;
  assign n2633 = n140 | n233 ;
  assign n2634 = ( n1110 & ~n2632 ) | ( n1110 & n2633 ) | ( ~n2632 & n2633 ) ;
  assign n2635 = n2632 | n2634 ;
  assign n2630 = n404 | n2507 ;
  assign n2631 = n86 | n2630 ;
  assign n2636 = ( n2635 & ~n2301 ) | ( n2635 & n2631 ) | ( ~n2301 & n2631 ) ;
  assign n2637 = n2301 | n2636 ;
  assign n2626 = n195 | n674 ;
  assign n2627 = ( n69 & ~n160 ) | ( n69 & n2626 ) | ( ~n160 & n2626 ) ;
  assign n2628 = n160 | n2627 ;
  assign n2629 = n212 | n2628 ;
  assign n2638 = ( n879 & n2637 ) | ( n879 & n2629 ) | ( n2637 & n2629 ) ;
  assign n2639 = ( n879 & ~n2638 ) | ( n879 & 1'b0 ) | ( ~n2638 & 1'b0 ) ;
  assign n2640 = ( n1490 & ~n779 ) | ( n1490 & n2639 ) | ( ~n779 & n2639 ) ;
  assign n2641 = ~n1490 & n2640 ;
  assign n2642 = ( n150 & ~n792 ) | ( n150 & n2641 ) | ( ~n792 & n2641 ) ;
  assign n2643 = ~n150 & n2642 ;
  assign n2644 = ( n475 & ~n52 ) | ( n475 & n2643 ) | ( ~n52 & n2643 ) ;
  assign n2645 = ~n475 & n2644 ;
  assign n2646 = ( n168 & ~n529 ) | ( n168 & n2645 ) | ( ~n529 & n2645 ) ;
  assign n2647 = ~n168 & n2646 ;
  assign n2652 = ( n2625 & ~n2651 ) | ( n2625 & n2647 ) | ( ~n2651 & n2647 ) ;
  assign n2653 = ( n1807 & ~n2625 ) | ( n1807 & n2652 ) | ( ~n2625 & n2652 ) ;
  assign n2654 = ~n1807 & n2653 ;
  assign n2655 = ( n2620 & ~n2575 ) | ( n2620 & n2654 ) | ( ~n2575 & n2654 ) ;
  assign n2656 = ( n1061 & n2575 ) | ( n1061 & n2655 ) | ( n2575 & n2655 ) ;
  assign n2657 = ~n1061 & n2656 ;
  assign n2658 = ( n280 & ~n434 ) | ( n280 & n2657 ) | ( ~n434 & n2657 ) ;
  assign n2659 = ~n280 & n2658 ;
  assign n2660 = ( n222 & ~n569 ) | ( n222 & n2659 ) | ( ~n569 & n2659 ) ;
  assign n2661 = ~n222 & n2660 ;
  assign n2662 = ( n120 & ~n2661 ) | ( n120 & n644 ) | ( ~n2661 & n644 ) ;
  assign n2663 = ( n644 & ~n2662 ) | ( n644 & 1'b0 ) | ( ~n2662 & 1'b0 ) ;
  assign n2664 = ( n252 & ~n155 ) | ( n252 & n2663 ) | ( ~n155 & n2663 ) ;
  assign n2665 = ~n252 &  n2664 ;
  assign n2666 = n485 | n666 ;
  assign n2687 = n333 | n603 ;
  assign n2688 = ( n577 & ~n1884 ) | ( n577 & n1002 ) | ( ~n1884 & n1002 ) ;
  assign n2689 = n1884 | n2688 ;
  assign n2690 = ( n2687 & ~n418 ) | ( n2687 & n2689 ) | ( ~n418 & n2689 ) ;
  assign n2691 = n418 | n2690 ;
  assign n2692 = ( n2621 & ~n373 ) | ( n2621 & n2691 ) | ( ~n373 & n2691 ) ;
  assign n2693 = n373 | n2692 ;
  assign n2694 = ( n123 & ~n214 ) | ( n123 & n2693 ) | ( ~n214 & n2693 ) ;
  assign n2695 = n214 | n2694 ;
  assign n2696 = n384 | n2695 ;
  assign n2697 = n797 | n814 ;
  assign n2698 = ( n101 & ~n217 ) | ( n101 & n2697 ) | ( ~n217 & n2697 ) ;
  assign n2699 = n217 | n2698 ;
  assign n2700 = ( n155 & ~n141 ) | ( n155 & n2699 ) | ( ~n141 & n2699 ) ;
  assign n2701 = n141 | n2700 ;
  assign n2734 = n126 | n424 ;
  assign n2735 = n631 | n2734 ;
  assign n2702 = n89 | n270 ;
  assign n2703 = n52 | n744 ;
  assign n2704 = ( n2702 & ~n2576 ) | ( n2702 & n2703 ) | ( ~n2576 & n2703 ) ;
  assign n2705 = n2576 | n2704 ;
  assign n2706 = ( n718 & ~n1268 ) | ( n718 & n2705 ) | ( ~n1268 & n2705 ) ;
  assign n2707 = n1268 | n2706 ;
  assign n2708 = ( n91 & ~n737 ) | ( n91 & n2707 ) | ( ~n737 & n2707 ) ;
  assign n2709 = n737 | n2708 ;
  assign n2710 = ( n104 & ~n630 ) | ( n104 & n2709 ) | ( ~n630 & n2709 ) ;
  assign n2711 = n630 | n2710 ;
  assign n2712 = ( n476 & ~n663 ) | ( n476 & n2711 ) | ( ~n663 & n2711 ) ;
  assign n2713 = n663 | n2712 ;
  assign n2714 = n953 | n1064 ;
  assign n2715 = ( n672 & ~n796 ) | ( n672 & n2714 ) | ( ~n796 & n2714 ) ;
  assign n2716 = n796 | n2715 ;
  assign n2717 = ( n240 & ~n711 ) | ( n240 & n2716 ) | ( ~n711 & n2716 ) ;
  assign n2718 = n711 | n2717 ;
  assign n2719 = ( n2718 & ~n2713 ) | ( n2718 & n1245 ) | ( ~n2713 & n1245 ) ;
  assign n2720 = ( n2713 & ~n864 ) | ( n2713 & n2719 ) | ( ~n864 & n2719 ) ;
  assign n2721 = n864 | n2720 ;
  assign n2722 = ( n1278 & ~n1824 ) | ( n1278 & n2721 ) | ( ~n1824 & n2721 ) ;
  assign n2723 = n1824 | n2722 ;
  assign n2724 = ( n885 & ~n1427 ) | ( n885 & n2723 ) | ( ~n1427 & n2723 ) ;
  assign n2725 = ( n1427 & ~n194 ) | ( n1427 & n2724 ) | ( ~n194 & n2724 ) ;
  assign n2726 = n194 | n2725 ;
  assign n2727 = ( n253 & ~n429 ) | ( n253 & n2726 ) | ( ~n429 & n2726 ) ;
  assign n2728 = n429 | n2727 ;
  assign n2729 = ( n722 & ~n233 ) | ( n722 & n2728 ) | ( ~n233 & n2728 ) ;
  assign n2730 = n233 | n2729 ;
  assign n2731 = ( n623 & ~n2730 ) | ( n623 & 1'b0 ) | ( ~n2730 & 1'b0 ) ;
  assign n2732 = ( n549 & ~n911 ) | ( n549 & n2731 ) | ( ~n911 & n2731 ) ;
  assign n2733 = ~n549 & n2732 ;
  assign n2736 = ( n1809 & ~n2735 ) | ( n1809 & n2733 ) | ( ~n2735 & n2733 ) ;
  assign n2737 = ~n1809 & n2736 ;
  assign n2738 = ( n1458 & n2701 ) | ( n1458 & n2737 ) | ( n2701 & n2737 ) ;
  assign n2739 = ~n2701 & n2738 ;
  assign n2667 = n241 | n721 ;
  assign n2668 = ( n188 & ~n350 ) | ( n188 & n2667 ) | ( ~n350 & n2667 ) ;
  assign n2669 = n350 | n2668 ;
  assign n2670 = n83 | n2669 ;
  assign n2671 = ( n274 & ~n359 ) | ( n274 & n534 ) | ( ~n359 & n534 ) ;
  assign n2672 = n359 | n2671 ;
  assign n2673 = n1399 | n2672 ;
  assign n2674 = ( n1971 & ~n2670 ) | ( n1971 & n2673 ) | ( ~n2670 & n2673 ) ;
  assign n2675 = ( n2670 & ~n1617 ) | ( n2670 & n2674 ) | ( ~n1617 & n2674 ) ;
  assign n2676 = n1617 | n2675 ;
  assign n2677 = ( n525 & n906 ) | ( n525 & n2676 ) | ( n906 & n2676 ) ;
  assign n2678 = ( n525 & ~n2677 ) | ( n525 & 1'b0 ) | ( ~n2677 & 1'b0 ) ;
  assign n2679 = ( n475 & ~n2678 ) | ( n475 & n813 ) | ( ~n2678 & n813 ) ;
  assign n2680 = ( n813 & ~n2679 ) | ( n813 & 1'b0 ) | ( ~n2679 & 1'b0 ) ;
  assign n2681 = ( n460 & ~n191 ) | ( n460 & n2680 ) | ( ~n191 & n2680 ) ;
  assign n2682 = ~n460 & n2681 ;
  assign n2683 = ( n197 & n554 ) | ( n197 & n2682 ) | ( n554 & n2682 ) ;
  assign n2684 = ~n554 & n2683 ;
  assign n2685 = ( n433 & ~n229 ) | ( n433 & n2684 ) | ( ~n229 & n2684 ) ;
  assign n2686 = ~n433 & n2685 ;
  assign n2740 = ( n2696 & ~n2739 ) | ( n2696 & n2686 ) | ( ~n2739 & n2686 ) ;
  assign n2741 = ( n647 & ~n2740 ) | ( n647 & n2686 ) | ( ~n2740 & n2686 ) ;
  assign n2742 = ~n647 & n2741 ;
  assign n2743 = ( n620 & ~n2666 ) | ( n620 & n2742 ) | ( ~n2666 & n2742 ) ;
  assign n2744 = ~n620 & n2743 ;
  assign n2745 = ( n1072 & ~n1567 ) | ( n1072 & n2744 ) | ( ~n1567 & n2744 ) ;
  assign n2746 = ( n2745 & ~n1072 ) | ( n2745 & 1'b0 ) | ( ~n1072 & 1'b0 ) ;
  assign n2747 = ( n245 & ~n479 ) | ( n245 & n2746 ) | ( ~n479 & n2746 ) ;
  assign n2748 = ~n245 & n2747 ;
  assign n2749 = ( n349 & ~n226 ) | ( n349 & n2748 ) | ( ~n226 & n2748 ) ;
  assign n2750 = ~n349 & n2749 ;
  assign n2751 = ~n86 &  n2750 ;
  assign n2752 = n281 | n561 ;
  assign n2753 = ( n2358 & ~n2187 ) | ( n2358 & n2752 ) | ( ~n2187 & n2752 ) ;
  assign n2754 = n2187 | n2753 ;
  assign n2755 = ( n812 & ~n151 ) | ( n812 & n2754 ) | ( ~n151 & n2754 ) ;
  assign n2756 = n151 | n2755 ;
  assign n2757 = n137 | n2756 ;
  assign n2758 = ~n226 & n813 ;
  assign n2759 = ( n169 & ~n267 ) | ( n169 & n2758 ) | ( ~n267 & n2758 ) ;
  assign n2760 = ~n169 & n2759 ;
  assign n2767 = n415 | n617 ;
  assign n2768 = n196 | n2767 ;
  assign n2764 = n235 | n800 ;
  assign n2765 = ( n790 & ~n284 ) | ( n790 & n2764 ) | ( ~n284 & n2764 ) ;
  assign n2766 = n284 | n2765 ;
  assign n2769 = ( n2768 & ~n2598 ) | ( n2768 & n2766 ) | ( ~n2598 & n2766 ) ;
  assign n2770 = n2598 | n2769 ;
  assign n2771 = ( n2154 & ~n2770 ) | ( n2154 & n2278 ) | ( ~n2770 & n2278 ) ;
  assign n2772 = ~n2154 & n2771 ;
  assign n2773 = ( n2772 & ~n1283 ) | ( n2772 & n1982 ) | ( ~n1283 & n1982 ) ;
  assign n2774 = ( n2773 & ~n1982 ) | ( n2773 & 1'b0 ) | ( ~n1982 & 1'b0 ) ;
  assign n2761 = ( n211 & ~n279 ) | ( n211 & n270 ) | ( ~n279 & n270 ) ;
  assign n2762 = n279 | n2761 ;
  assign n2763 = n93 | n2762 ;
  assign n2775 = ( n2760 & ~n2774 ) | ( n2760 & n2763 ) | ( ~n2774 & n2763 ) ;
  assign n2776 = ( n2395 & ~n2775 ) | ( n2395 & n2760 ) | ( ~n2775 & n2760 ) ;
  assign n2777 = ~n2395 & n2776 ;
  assign n2778 = ( n793 & ~n2757 ) | ( n793 & n2777 ) | ( ~n2757 & n2777 ) ;
  assign n2779 = ~n793 & n2778 ;
  assign n2780 = ( n711 & ~n272 ) | ( n711 & n2779 ) | ( ~n272 & n2779 ) ;
  assign n2781 = ~n711 & n2780 ;
  assign n2782 = ( n603 & ~n348 ) | ( n603 & n2781 ) | ( ~n348 & n2781 ) ;
  assign n2783 = ~n603 &  n2782 ;
  assign n2784 = n793 | n909 ;
  assign n2785 = n69 | n224 ;
  assign n2786 = n403 | n2785 ;
  assign n2787 = ( n2768 & ~n1797 ) | ( n2768 & n2786 ) | ( ~n1797 & n2786 ) ;
  assign n2788 = n1797 | n2787 ;
  assign n2789 = ( n2784 & ~n1513 ) | ( n2784 & n2788 ) | ( ~n1513 & n2788 ) ;
  assign n2790 = n1513 | n2789 ;
  assign n2791 = ( n52 & ~n190 ) | ( n52 & n2790 ) | ( ~n190 & n2790 ) ;
  assign n2792 = n190 | n2791 ;
  assign n2793 = ( n156 & n343 ) | ( n156 & n2792 ) | ( n343 & n2792 ) ;
  assign n2794 = ( n343 & ~n2793 ) | ( n343 & 1'b0 ) | ( ~n2793 & 1'b0 ) ;
  assign n2795 = ( n2794 & ~n155 ) | ( n2794 & n643 ) | ( ~n155 & n643 ) ;
  assign n2796 = ( n2795 & ~n643 ) | ( n2795 & 1'b0 ) | ( ~n643 & 1'b0 ) ;
  assign n2797 = n675 | n1532 ;
  assign n2798 = ( n197 & ~n2797 ) | ( n197 & 1'b0 ) | ( ~n2797 & 1'b0 ) ;
  assign n2799 = n672 | n788 ;
  assign n2800 = ( n630 & ~n284 ) | ( n630 & n2799 ) | ( ~n284 & n2799 ) ;
  assign n2801 = n284 | n2800 ;
  assign n2802 = ( n562 & ~n607 ) | ( n562 & n1233 ) | ( ~n607 & n1233 ) ;
  assign n2803 = n607 | n2802 ;
  assign n2804 = n526 | n2803 ;
  assign n2805 = n165 | n408 ;
  assign n2806 = ( n49 & ~n332 ) | ( n49 & n2805 ) | ( ~n332 & n2805 ) ;
  assign n2807 = n332 | n2806 ;
  assign n2808 = n225 | n534 ;
  assign n2809 = ( n2263 & ~n1633 ) | ( n2263 & n2808 ) | ( ~n1633 & n2808 ) ;
  assign n2810 = n1633 | n2809 ;
  assign n2811 = ( n2807 & ~n2592 ) | ( n2807 & n2810 ) | ( ~n2592 & n2810 ) ;
  assign n2812 = n2592 | n2811 ;
  assign n2813 = ( n1325 & n1343 ) | ( n1325 & n2812 ) | ( n1343 & n2812 ) ;
  assign n2814 = ( n1244 & ~n2813 ) | ( n1244 & n1343 ) | ( ~n2813 & n1343 ) ;
  assign n2815 = ~n1244 & n2814 ;
  assign n2816 = ( n1461 & ~n2577 ) | ( n1461 & n2815 ) | ( ~n2577 & n2815 ) ;
  assign n2817 = ( n2816 & ~n1461 ) | ( n2816 & 1'b0 ) | ( ~n1461 & 1'b0 ) ;
  assign n2818 = ( n274 & ~n2817 ) | ( n274 & n524 ) | ( ~n2817 & n524 ) ;
  assign n2819 = ( n524 & ~n2818 ) | ( n524 & 1'b0 ) | ( ~n2818 & 1'b0 ) ;
  assign n2820 = ( n77 & ~n342 ) | ( n77 & n2819 ) | ( ~n342 & n2819 ) ;
  assign n2821 = ~n77 & n2820 ;
  assign n2822 = ~n476 & n2821 ;
  assign n2823 = ( n2801 & ~n2804 ) | ( n2801 & n2822 ) | ( ~n2804 & n2822 ) ;
  assign n2824 = ( n2506 & ~n2801 ) | ( n2506 & n2823 ) | ( ~n2801 & n2823 ) ;
  assign n2825 = ~n2506 & n2824 ;
  assign n2826 = ( n2128 & n2798 ) | ( n2128 & n2825 ) | ( n2798 & n2825 ) ;
  assign n2827 = ~n2128 & n2826 ;
  assign n2828 = ( n1195 & n2796 ) | ( n1195 & n2827 ) | ( n2796 & n2827 ) ;
  assign n2829 = ( n645 & ~n2828 ) | ( n645 & n1195 ) | ( ~n2828 & n1195 ) ;
  assign n2830 = ( n645 & ~n2829 ) | ( n645 & 1'b0 ) | ( ~n2829 & 1'b0 ) ;
  assign n2831 = ( n671 & ~n125 ) | ( n671 & n2830 ) | ( ~n125 & n2830 ) ;
  assign n2832 = ~n671 & n2831 ;
  assign n2833 = ( n217 & ~n2667 ) | ( n217 & n2832 ) | ( ~n2667 & n2832 ) ;
  assign n2834 = ~n217 & n2833 ;
  assign n2835 = ( n456 & ~n737 ) | ( n456 & n2834 ) | ( ~n737 & n2834 ) ;
  assign n2836 = ~n456 & n2835 ;
  assign n2837 = ( n411 & ~n149 ) | ( n411 & n2836 ) | ( ~n149 & n2836 ) ;
  assign n2838 = ~n411 & n2837 ;
  assign n2839 = ~n351 &  n2838 ;
  assign n2840 = n65 | n104 ;
  assign n2841 = n195 | n679 ;
  assign n2842 = ( n429 & ~n207 ) | ( n429 & n2841 ) | ( ~n207 & n2841 ) ;
  assign n2843 = ( n207 & ~n909 ) | ( n207 & n2842 ) | ( ~n909 & n2842 ) ;
  assign n2844 = n909 | n2843 ;
  assign n2845 = ( n531 & ~n556 ) | ( n531 & n2844 ) | ( ~n556 & n2844 ) ;
  assign n2846 = n556 | n2845 ;
  assign n2847 = ( n478 & ~n167 ) | ( n478 & n2846 ) | ( ~n167 & n2846 ) ;
  assign n2848 = n167 | n2847 ;
  assign n2849 = n206 | n374 ;
  assign n2850 = n132 | n2849 ;
  assign n2863 = n300 | n714 ;
  assign n2864 = n492 | n2863 ;
  assign n2851 = ( n197 & ~n216 ) | ( n197 & n792 ) | ( ~n216 & n792 ) ;
  assign n2852 = ( n75 & ~n792 ) | ( n75 & n2851 ) | ( ~n792 & n2851 ) ;
  assign n2853 = ~n75 & n2852 ;
  assign n2854 = ( n1883 & ~n2468 ) | ( n1883 & n2853 ) | ( ~n2468 & n2853 ) ;
  assign n2855 = ~n1883 & n2854 ;
  assign n2856 = ( n797 & ~n2348 ) | ( n797 & n2855 ) | ( ~n2348 & n2855 ) ;
  assign n2857 = ~n797 & n2856 ;
  assign n2858 = ( n130 & ~n721 ) | ( n130 & n2857 ) | ( ~n721 & n2857 ) ;
  assign n2859 = ~n130 & n2858 ;
  assign n2860 = ( n118 & ~n356 ) | ( n118 & n2859 ) | ( ~n356 & n2859 ) ;
  assign n2861 = ~n118 & n2860 ;
  assign n2862 = ~n252 & n2861 ;
  assign n2865 = ( n2850 & ~n2864 ) | ( n2850 & n2862 ) | ( ~n2864 & n2862 ) ;
  assign n2866 = ( n1991 & ~n2850 ) | ( n1991 & n2865 ) | ( ~n2850 & n2865 ) ;
  assign n2867 = ~n1991 & n2866 ;
  assign n2868 = ( n1955 & ~n1224 ) | ( n1955 & n2867 ) | ( ~n1224 & n2867 ) ;
  assign n2869 = ~n1955 & n2868 ;
  assign n2870 = ( n761 & ~n407 ) | ( n761 & n2869 ) | ( ~n407 & n2869 ) ;
  assign n2871 = ~n761 & n2870 ;
  assign n2872 = ( n560 & ~n279 ) | ( n560 & n2871 ) | ( ~n279 & n2871 ) ;
  assign n2873 = ~n560 & n2872 ;
  assign n2874 = ( n2873 & ~n221 ) | ( n2873 & n266 ) | ( ~n221 & n266 ) ;
  assign n2875 = ( n2874 & ~n266 ) | ( n2874 & 1'b0 ) | ( ~n266 & 1'b0 ) ;
  assign n2876 = ( n664 & ~n135 ) | ( n664 & n2875 ) | ( ~n135 & n2875 ) ;
  assign n2877 = ~n664 & n2876 ;
  assign n2878 = ~n225 & n2877 ;
  assign n2879 = ( n606 & ~n1627 ) | ( n606 & n1187 ) | ( ~n1627 & n1187 ) ;
  assign n2880 = n1627 | n2879 ;
  assign n2881 = ( n2128 & ~n1884 ) | ( n2128 & n2880 ) | ( ~n1884 & n2880 ) ;
  assign n2882 = n1884 | n2881 ;
  assign n2883 = ( n382 & ~n259 ) | ( n382 & n2882 ) | ( ~n259 & n2882 ) ;
  assign n2884 = ( n259 & ~n424 ) | ( n259 & n2883 ) | ( ~n424 & n2883 ) ;
  assign n2885 = n424 | n2884 ;
  assign n2886 = ( n628 & ~n166 ) | ( n628 & n2885 ) | ( ~n166 & n2885 ) ;
  assign n2887 = n166 | n2886 ;
  assign n2888 = ~n273 & n1183 ;
  assign n2889 = ~n43 & n2888 ;
  assign n2890 = n409 | n716 ;
  assign n2891 = ( n354 & ~n2890 ) | ( n354 & 1'b0 ) | ( ~n2890 & 1'b0 ) ;
  assign n2892 = ( n1704 & n2889 ) | ( n1704 & n2891 ) | ( n2889 & n2891 ) ;
  assign n2893 = ~n1704 & n2892 ;
  assign n2894 = ( n1877 & ~n2887 ) | ( n1877 & n2893 ) | ( ~n2887 & n2893 ) ;
  assign n2895 = ~n1877 & n2894 ;
  assign n2896 = ( n2848 & n2878 ) | ( n2848 & n2895 ) | ( n2878 & n2895 ) ;
  assign n2897 = ~n2848 & n2896 ;
  assign n2898 = ( n747 & ~n1045 ) | ( n747 & n2897 ) | ( ~n1045 & n2897 ) ;
  assign n2899 = ~n747 & n2898 ;
  assign n2900 = ( n906 & ~n2840 ) | ( n906 & n2899 ) | ( ~n2840 & n2899 ) ;
  assign n2901 = ~n906 & n2900 ;
  assign n2902 = ( n125 & ~n1185 ) | ( n125 & n2901 ) | ( ~n1185 & n2901 ) ;
  assign n2903 = ~n125 & n2902 ;
  assign n2904 = ( n2903 & ~n451 ) | ( n2903 & n800 ) | ( ~n451 & n800 ) ;
  assign n2905 = ( n2904 & ~n800 ) | ( n2904 & 1'b0 ) | ( ~n800 & 1'b0 ) ;
  assign n2906 = ( n460 & ~n91 ) | ( n460 & n2905 ) | ( ~n91 & n2905 ) ;
  assign n2907 = ~n460 & n2906 ;
  assign n2908 = ( n196 & ~n411 ) | ( n196 & n2907 ) | ( ~n411 & n2907 ) ;
  assign n2909 = ~n196 & n2908 ;
  assign n2910 = ~n2909 |  n670 ;
  assign n2911 = n716 | n2191 ;
  assign n2912 = ( n243 & ~n676 ) | ( n243 & n2911 ) | ( ~n676 & n2911 ) ;
  assign n2913 = n676 | n2912 ;
  assign n2914 = n643 | n2913 ;
  assign n2915 = ( n246 & ~n1268 ) | ( n246 & n491 ) | ( ~n1268 & n491 ) ;
  assign n2916 = n1268 | n2915 ;
  assign n2917 = ( n207 & ~n234 ) | ( n207 & n2916 ) | ( ~n234 & n2916 ) ;
  assign n2918 = n234 | n2917 ;
  assign n2919 = ( n139 & ~n299 ) | ( n139 & n2918 ) | ( ~n299 & n2918 ) ;
  assign n2920 = n299 | n2919 ;
  assign n2921 = ( n663 & ~n267 ) | ( n663 & n2920 ) | ( ~n267 & n2920 ) ;
  assign n2922 = n267 | n2921 ;
  assign n2923 = n410 | n2922 ;
  assign n2924 = ( n1002 & ~n1829 ) | ( n1002 & n497 ) | ( ~n1829 & n497 ) ;
  assign n2925 = n1829 | n2924 ;
  assign n2926 = ( n1071 & ~n1169 ) | ( n1071 & n2925 ) | ( ~n1169 & n2925 ) ;
  assign n2927 = n1169 | n2926 ;
  assign n2928 = ( n2044 & ~n361 ) | ( n2044 & n2927 ) | ( ~n361 & n2927 ) ;
  assign n2929 = n361 | n2928 ;
  assign n2930 = ( n2923 & ~n2914 ) | ( n2923 & n2929 ) | ( ~n2914 & n2929 ) ;
  assign n2931 = ( n2914 & ~n906 ) | ( n2914 & n2930 ) | ( ~n906 & n2930 ) ;
  assign n2932 = n906 | n2931 ;
  assign n2933 = ( n193 & ~n711 ) | ( n193 & n2932 ) | ( ~n711 & n2932 ) ;
  assign n2934 = n711 | n2933 ;
  assign n2935 = ( n237 & ~n271 ) | ( n237 & n2934 ) | ( ~n271 & n2934 ) ;
  assign n2936 = n271 | n2935 ;
  assign n2937 = n126 | n235 ;
  assign n2938 = ( n257 & ~n792 ) | ( n257 & n2937 ) | ( ~n792 & n2937 ) ;
  assign n2939 = n792 | n2938 ;
  assign n2940 = ( n105 & ~n58 ) | ( n105 & n2939 ) | ( ~n58 & n2939 ) ;
  assign n2941 = n58 | n2940 ;
  assign n2942 = ( n162 & ~n454 ) | ( n162 & n2941 ) | ( ~n454 & n2941 ) ;
  assign n2943 = n454 | n2942 ;
  assign n2944 = n195 | n337 ;
  assign n2945 = n745 | n2944 ;
  assign n2946 = ( n1317 & ~n2547 ) | ( n1317 & n2945 ) | ( ~n2547 & n2945 ) ;
  assign n2947 = n2547 | n2946 ;
  assign n2948 = ( n2752 & ~n1963 ) | ( n2752 & n2947 ) | ( ~n1963 & n2947 ) ;
  assign n2949 = n1963 | n2948 ;
  assign n2950 = ( n2943 & ~n1325 ) | ( n2943 & n2949 ) | ( ~n1325 & n2949 ) ;
  assign n2951 = n1325 | n2950 ;
  assign n2952 = ( n2029 & ~n458 ) | ( n2029 & n2951 ) | ( ~n458 & n2951 ) ;
  assign n2953 = n458 | n2952 ;
  assign n2954 = ( n272 & ~n1280 ) | ( n272 & n2953 ) | ( ~n1280 & n2953 ) ;
  assign n2955 = ( n1280 & ~n217 ) | ( n1280 & n2954 ) | ( ~n217 & n2954 ) ;
  assign n2956 = n217 | n2955 ;
  assign n2957 = n226 | n2956 ;
  assign n2972 = n69 | n123 ;
  assign n2973 = ( n529 & ~n205 ) | ( n529 & n2972 ) | ( ~n205 & n2972 ) ;
  assign n2974 = n205 | n2973 ;
  assign n2975 = ( n618 & ~n129 ) | ( n618 & n2974 ) | ( ~n129 & n2974 ) ;
  assign n2976 = n129 | n2975 ;
  assign n2977 = n1233 | n1603 ;
  assign n2978 = ( n719 & ~n2976 ) | ( n719 & n2977 ) | ( ~n2976 & n2977 ) ;
  assign n2979 = n2976 | n2978 ;
  assign n2958 = n408 | n2082 ;
  assign n2959 = n161 | n418 ;
  assign n2960 = n151 | n350 ;
  assign n2961 = ( n463 & ~n2959 ) | ( n463 & n2960 ) | ( ~n2959 & n2960 ) ;
  assign n2962 = ( n2959 & ~n1385 ) | ( n2959 & n2961 ) | ( ~n1385 & n2961 ) ;
  assign n2963 = n1385 | n2962 ;
  assign n2964 = ( n2958 & ~n429 ) | ( n2958 & n2963 ) | ( ~n429 & n2963 ) ;
  assign n2965 = n429 | n2964 ;
  assign n2966 = ( n206 & ~n796 ) | ( n206 & n2965 ) | ( ~n796 & n2965 ) ;
  assign n2967 = n796 | n2966 ;
  assign n2968 = ( n644 & ~n197 ) | ( n644 & n2967 ) | ( ~n197 & n2967 ) ;
  assign n2969 = ( n644 & ~n2968 ) | ( n644 & 1'b0 ) | ( ~n2968 & 1'b0 ) ;
  assign n2970 = ( n574 & ~n628 ) | ( n574 & n2969 ) | ( ~n628 & n2969 ) ;
  assign n2971 = ~n574 & n2970 ;
  assign n2980 = ( n2957 & ~n2979 ) | ( n2957 & n2971 ) | ( ~n2979 & n2971 ) ;
  assign n2981 = ( n2190 & ~n2980 ) | ( n2190 & n2957 ) | ( ~n2980 & n2957 ) ;
  assign n2982 = ( n2190 & ~n2981 ) | ( n2190 & 1'b0 ) | ( ~n2981 & 1'b0 ) ;
  assign n2983 = ( n2982 & ~n673 ) | ( n2982 & n2936 ) | ( ~n673 & n2936 ) ;
  assign n2984 = ( n1484 & ~n2936 ) | ( n1484 & n2983 ) | ( ~n2936 & n2983 ) ;
  assign n2985 = ~n1484 & n2984 ;
  assign n2986 = ( n786 & ~n2985 ) | ( n786 & n787 ) | ( ~n2985 & n787 ) ;
  assign n2987 = ( n786 & ~n2986 ) | ( n786 & 1'b0 ) | ( ~n2986 & 1'b0 ) ;
  assign n2988 = ( n735 & ~n232 ) | ( n735 & n2987 ) | ( ~n232 & n2987 ) ;
  assign n2989 = ~n735 & n2988 ;
  assign n2990 = ( n269 & ~n216 ) | ( n269 & n2989 ) | ( ~n216 & n2989 ) ;
  assign n2991 = ~n269 & n2990 ;
  assign n2992 = ( n300 & ~n406 ) | ( n300 & n2991 ) | ( ~n406 & n2991 ) ;
  assign n2993 = ~n300 & n2992 ;
  assign n2994 = ( n476 & ~n666 ) | ( n476 & n2993 ) | ( ~n666 & n2993 ) ;
  assign n2995 = ~n476 & n2994 ;
  assign n2996 = n195 | n761 ;
  assign n2997 = ( n2763 & ~n2252 ) | ( n2763 & n2996 ) | ( ~n2252 & n2996 ) ;
  assign n2998 = n2252 | n2997 ;
  assign n2999 = ( n2308 & ~n337 ) | ( n2308 & n2998 ) | ( ~n337 & n2998 ) ;
  assign n3000 = n337 | n2999 ;
  assign n3001 = ( n495 & ~n335 ) | ( n495 & n3000 ) | ( ~n335 & n3000 ) ;
  assign n3002 = n335 | n3001 ;
  assign n3003 = ( n127 & ~n376 ) | ( n127 & n3002 ) | ( ~n376 & n3002 ) ;
  assign n3004 = n376 | n3003 ;
  assign n3005 = ( n253 & ~n232 ) | ( n253 & n3004 ) | ( ~n232 & n3004 ) ;
  assign n3006 = n232 | n3005 ;
  assign n3007 = ( n905 & ~n417 ) | ( n905 & n3006 ) | ( ~n417 & n3006 ) ;
  assign n3008 = n417 | n3007 ;
  assign n3009 = n141 | n3008 ;
  assign n3010 = n549 | n721 ;
  assign n3011 = n628 | n3010 ;
  assign n3012 = ~n1152 & n2760 ;
  assign n3013 = ~n778 & n3012 ;
  assign n3016 = n910 | n1808 ;
  assign n3017 = n948 | n3016 ;
  assign n3018 = ( n2376 & ~n3017 ) | ( n2376 & 1'b0 ) | ( ~n3017 & 1'b0 ) ;
  assign n3014 = ( n373 & ~n673 ) | ( n373 & n575 ) | ( ~n673 & n575 ) ;
  assign n3015 = n673 | n3014 ;
  assign n3019 = ( n3013 & ~n3018 ) | ( n3013 & n3015 ) | ( ~n3018 & n3015 ) ;
  assign n3020 = ( n1781 & ~n3013 ) | ( n1781 & n3019 ) | ( ~n3013 & n3019 ) ;
  assign n3021 = ( n1781 & ~n3020 ) | ( n1781 & 1'b0 ) | ( ~n3020 & 1'b0 ) ;
  assign n3022 = ( n3011 & ~n2577 ) | ( n3011 & n3021 ) | ( ~n2577 & n3021 ) ;
  assign n3023 = ( n1714 & ~n3011 ) | ( n1714 & n3022 ) | ( ~n3011 & n3022 ) ;
  assign n3024 = ~n1714 & n3023 ;
  assign n3025 = ( n3024 & ~n2187 ) | ( n3024 & n3009 ) | ( ~n2187 & n3009 ) ;
  assign n3026 = ( n1580 & ~n3009 ) | ( n1580 & n3025 ) | ( ~n3009 & n3025 ) ;
  assign n3027 = ( n3026 & ~n1580 ) | ( n3026 & 1'b0 ) | ( ~n1580 & 1'b0 ) ;
  assign n3028 = ( n1454 & ~n679 ) | ( n1454 & n3027 ) | ( ~n679 & n3027 ) ;
  assign n3029 = ~n1454 & n3028 ;
  assign n3030 = ~n74 &  n3029 ;
  assign n3031 = n52 | n299 ;
  assign n3032 = ( n363 & ~n2996 ) | ( n363 & n3031 ) | ( ~n2996 & n3031 ) ;
  assign n3033 = n2996 | n3032 ;
  assign n3034 = ( n1427 & ~n2462 ) | ( n1427 & n3033 ) | ( ~n2462 & n3033 ) ;
  assign n3035 = n2462 | n3034 ;
  assign n3036 = ( n495 & ~n244 ) | ( n495 & n3035 ) | ( ~n244 & n3035 ) ;
  assign n3037 = n244 | n3036 ;
  assign n3038 = ( n208 & ~n273 ) | ( n208 & n3037 ) | ( ~n273 & n3037 ) ;
  assign n3039 = n273 | n3038 ;
  assign n3040 = ( n484 & n765 ) | ( n484 & n3039 ) | ( n765 & n3039 ) ;
  assign n3041 = ( n484 & ~n3040 ) | ( n484 & 1'b0 ) | ( ~n3040 & 1'b0 ) ;
  assign n3042 = n540 | n559 ;
  assign n3043 = ~n284 & n524 ;
  assign n3044 = ( n961 & ~n3042 ) | ( n961 & n3043 ) | ( ~n3042 & n3043 ) ;
  assign n3045 = ~n961 & n3044 ;
  assign n3046 = ( n678 & ~n193 ) | ( n678 & n3045 ) | ( ~n193 & n3045 ) ;
  assign n3047 = ~n678 & n3046 ;
  assign n3048 = ( n453 & ~n722 ) | ( n453 & n3047 ) | ( ~n722 & n3047 ) ;
  assign n3049 = ~n453 & n3048 ;
  assign n3050 = ~n531 & n3049 ;
  assign n3051 = ( n1326 & ~n1672 ) | ( n1326 & n2960 ) | ( ~n1672 & n2960 ) ;
  assign n3052 = n1672 | n3051 ;
  assign n3053 = ( n3052 & ~n277 ) | ( n3052 & n2028 ) | ( ~n277 & n2028 ) ;
  assign n3054 = n277 | n3053 ;
  assign n3055 = ( n253 & ~n424 ) | ( n253 & n3054 ) | ( ~n424 & n3054 ) ;
  assign n3056 = n424 | n3055 ;
  assign n3057 = ( n255 & ~n745 ) | ( n255 & n3056 ) | ( ~n745 & n3056 ) ;
  assign n3058 = n745 | n3057 ;
  assign n3059 = n205 | n3058 ;
  assign n3060 = n557 | n1434 ;
  assign n3061 = ( n2850 & ~n258 ) | ( n2850 & n3060 ) | ( ~n258 & n3060 ) ;
  assign n3062 = n258 | n3061 ;
  assign n3063 = ( n191 & ~n333 ) | ( n191 & n3062 ) | ( ~n333 & n3062 ) ;
  assign n3064 = n333 | n3063 ;
  assign n3065 = ( n526 & ~n239 ) | ( n526 & n3064 ) | ( ~n239 & n3064 ) ;
  assign n3066 = n239 | n3065 ;
  assign n3067 = ( n91 & ~n241 ) | ( n91 & n712 ) | ( ~n241 & n712 ) ;
  assign n3068 = n241 | n3067 ;
  assign n3069 = n160 | n3068 ;
  assign n3070 = n457 | n569 ;
  assign n3071 = ( n3069 & ~n2649 ) | ( n3069 & n3070 ) | ( ~n2649 & n3070 ) ;
  assign n3072 = n2649 | n3071 ;
  assign n3073 = ( n3066 & ~n1823 ) | ( n3066 & n3072 ) | ( ~n1823 & n3072 ) ;
  assign n3074 = n1823 | n3073 ;
  assign n3075 = ( n3059 & ~n2784 ) | ( n3059 & n3074 ) | ( ~n2784 & n3074 ) ;
  assign n3076 = n2784 | n3075 ;
  assign n3077 = ( n1380 & ~n62 ) | ( n1380 & n3076 ) | ( ~n62 & n3076 ) ;
  assign n3078 = n62 | n3077 ;
  assign n3079 = ( n218 & n3078 ) | ( n218 & n813 ) | ( n3078 & n813 ) ;
  assign n3080 = ( n813 & ~n3079 ) | ( n813 & 1'b0 ) | ( ~n3079 & 1'b0 ) ;
  assign n3081 = ( n797 & ~n679 ) | ( n797 & n3080 ) | ( ~n679 & n3080 ) ;
  assign n3082 = ~n797 & n3081 ;
  assign n3083 = ( n734 & ~n271 ) | ( n734 & n3082 ) | ( ~n271 & n3082 ) ;
  assign n3084 = ~n734 & n3083 ;
  assign n3085 = ( n231 & ~n737 ) | ( n231 & n3084 ) | ( ~n737 & n3084 ) ;
  assign n3086 = ~n231 & n3085 ;
  assign n3087 = ~n529 & n3086 ;
  assign n3088 = n790 | n2702 ;
  assign n3089 = ( n188 & ~n349 ) | ( n188 & n3088 ) | ( ~n349 & n3088 ) ;
  assign n3090 = n349 | n3089 ;
  assign n3091 = n432 | n3090 ;
  assign n3092 = ( n413 & ~n245 ) | ( n413 & n905 ) | ( ~n245 & n905 ) ;
  assign n3093 = n245 | n3092 ;
  assign n3094 = ( n642 & ~n3093 ) | ( n642 & n1546 ) | ( ~n3093 & n1546 ) ;
  assign n3095 = ~n1546 & n3094 ;
  assign n3096 = ( n1429 & ~n3091 ) | ( n1429 & n3095 ) | ( ~n3091 & n3095 ) ;
  assign n3097 = ( n3096 & ~n1429 ) | ( n3096 & n2205 ) | ( ~n1429 & n2205 ) ;
  assign n3098 = ( n3097 & ~n2205 ) | ( n3097 & 1'b0 ) | ( ~n2205 & 1'b0 ) ;
  assign n3099 = ( n3087 & ~n3050 ) | ( n3087 & n3098 ) | ( ~n3050 & n3098 ) ;
  assign n3100 = n3050 &  n3099 ;
  assign n3101 = ( n3041 & ~n653 ) | ( n3041 & n3100 ) | ( ~n653 & n3100 ) ;
  assign n3102 = ( n653 & n1626 ) | ( n653 & n3101 ) | ( n1626 & n3101 ) ;
  assign n3103 = ~n1626 & n3102 ;
  assign n3104 = ( n676 & ~n672 ) | ( n676 & n3103 ) | ( ~n672 & n3103 ) ;
  assign n3105 = ~n676 & n3104 ;
  assign n3106 = ~n242 &  n3105 ;
  assign n3107 = n605 | n746 ;
  assign n3108 = ( n194 & ~n796 ) | ( n194 & n3107 ) | ( ~n796 & n3107 ) ;
  assign n3109 = n796 | n3108 ;
  assign n3110 = n737 | n3109 ;
  assign n3111 = ( n405 & ~n453 ) | ( n405 & n990 ) | ( ~n453 & n990 ) ;
  assign n3112 = n453 | n3111 ;
  assign n3113 = n149 | n3112 ;
  assign n3114 = ( n2084 & ~n2395 ) | ( n2084 & 1'b0 ) | ( ~n2395 & 1'b0 ) ;
  assign n3115 = ~n789 & n3114 ;
  assign n3116 = ( n1960 & ~n2435 ) | ( n1960 & n3115 ) | ( ~n2435 & n3115 ) ;
  assign n3117 = ~n1960 & n3116 ;
  assign n3118 = ( n1169 & ~n1833 ) | ( n1169 & n3117 ) | ( ~n1833 & n3117 ) ;
  assign n3119 = ~n1169 & n3118 ;
  assign n3120 = ( n3110 & ~n3113 ) | ( n3110 & n3119 ) | ( ~n3113 & n3119 ) ;
  assign n3121 = ( n463 & ~n3110 ) | ( n463 & n3120 ) | ( ~n3110 & n3120 ) ;
  assign n3122 = ~n463 & n3121 ;
  assign n3123 = ( n1427 & ~n3011 ) | ( n1427 & n3122 ) | ( ~n3011 & n3122 ) ;
  assign n3124 = ~n1427 & n3123 ;
  assign n3125 = ( n126 & ~n270 ) | ( n126 & n3124 ) | ( ~n270 & n3124 ) ;
  assign n3126 = ~n126 & n3125 ;
  assign n3127 = ( n226 & ~n240 ) | ( n226 & n3126 ) | ( ~n240 & n3126 ) ;
  assign n3128 = ~n226 & n3127 ;
  assign n3129 = ~n492 & n3128 ;
  assign n3130 = n277 | n475 ;
  assign n3131 = ( n3130 & ~n765 ) | ( n3130 & n800 ) | ( ~n765 & n800 ) ;
  assign n3132 = n765 | n3131 ;
  assign n3133 = ( n451 & ~n734 ) | ( n451 & n3132 ) | ( ~n734 & n3132 ) ;
  assign n3134 = n734 | n3133 ;
  assign n3135 = ( n644 & ~n524 ) | ( n644 & n3134 ) | ( ~n524 & n3134 ) ;
  assign n3136 = ( n644 & ~n3135 ) | ( n644 & 1'b0 ) | ( ~n3135 & 1'b0 ) ;
  assign n3137 = ~n529 & n3136 ;
  assign n3138 = n374 | n462 ;
  assign n3139 = ( n905 & ~n130 ) | ( n905 & n3138 ) | ( ~n130 & n3138 ) ;
  assign n3140 = n130 | n3139 ;
  assign n3141 = ( n340 & ~n433 ) | ( n340 & n3140 ) | ( ~n433 & n3140 ) ;
  assign n3142 = n433 | n3141 ;
  assign n3143 = n235 | n237 ;
  assign n3144 = n663 | n3143 ;
  assign n3145 = n161 | n214 ;
  assign n3146 = n167 | n3145 ;
  assign n3147 = ( n961 & ~n3144 ) | ( n961 & n3146 ) | ( ~n3144 & n3146 ) ;
  assign n3148 = ( n3147 & ~n1687 ) | ( n3147 & n3144 ) | ( ~n1687 & n3144 ) ;
  assign n3149 = n1687 | n3148 ;
  assign n3150 = ( n3142 & ~n1494 ) | ( n3142 & n3149 ) | ( ~n1494 & n3149 ) ;
  assign n3151 = n1494 | n3150 ;
  assign n3152 = ( n3137 & ~n3151 ) | ( n3137 & n1884 ) | ( ~n3151 & n1884 ) ;
  assign n3153 = ~n1884 & n3152 ;
  assign n3154 = ( n674 & ~n712 ) | ( n674 & n3153 ) | ( ~n712 & n3153 ) ;
  assign n3155 = ~n674 & n3154 ;
  assign n3156 = ( n735 & ~n156 ) | ( n735 & n3155 ) | ( ~n156 & n3155 ) ;
  assign n3157 = ~n735 & n3156 ;
  assign n3158 = n570 | n778 ;
  assign n3159 = n127 | n403 ;
  assign n3160 = n1110 | n2540 ;
  assign n3161 = ( n1232 & ~n3159 ) | ( n1232 & n3160 ) | ( ~n3159 & n3160 ) ;
  assign n3162 = ( n3159 & ~n1495 ) | ( n3159 & n3161 ) | ( ~n1495 & n3161 ) ;
  assign n3163 = n1495 | n3162 ;
  assign n3164 = ( n793 & ~n3158 ) | ( n793 & n3163 ) | ( ~n3158 & n3163 ) ;
  assign n3165 = ( n3164 & ~n775 ) | ( n3164 & n3158 ) | ( ~n775 & n3158 ) ;
  assign n3166 = n775 | n3165 ;
  assign n3167 = ( n272 & ~n338 ) | ( n272 & n3166 ) | ( ~n338 & n3166 ) ;
  assign n3168 = n338 | n3167 ;
  assign n3169 = ( n221 & ~n631 ) | ( n221 & n3168 ) | ( ~n631 & n3168 ) ;
  assign n3170 = n631 | n3169 ;
  assign n3171 = n476 | n602 ;
  assign n3181 = n953 | n1797 ;
  assign n3172 = n230 | n787 ;
  assign n3173 = n417 | n3172 ;
  assign n3174 = ( n1047 & ~n678 ) | ( n1047 & n3173 ) | ( ~n678 & n3173 ) ;
  assign n3175 = n678 | n3174 ;
  assign n3176 = ( n266 & ~n284 ) | ( n266 & n3175 ) | ( ~n284 & n3175 ) ;
  assign n3177 = n284 | n3176 ;
  assign n3178 = ( n43 & ~n166 ) | ( n43 & n3177 ) | ( ~n166 & n3177 ) ;
  assign n3179 = n166 | n3178 ;
  assign n3180 = n155 | n3179 ;
  assign n3182 = ( n3181 & ~n3171 ) | ( n3181 & n3180 ) | ( ~n3171 & n3180 ) ;
  assign n3183 = ( n3171 & ~n1515 ) | ( n3171 & n3182 ) | ( ~n1515 & n3182 ) ;
  assign n3184 = n1515 | n3183 ;
  assign n3185 = ( n3170 & n3184 ) | ( n3170 & n3157 ) | ( n3184 & n3157 ) ;
  assign n3186 = ( n3157 & ~n3185 ) | ( n3157 & 1'b0 ) | ( ~n3185 & 1'b0 ) ;
  assign n3187 = ( n2576 & n3129 ) | ( n2576 & n3186 ) | ( n3129 & n3186 ) ;
  assign n3188 = ~n2576 & n3187 ;
  assign n3189 = ( n947 & ~n2191 ) | ( n947 & n3188 ) | ( ~n2191 & n3188 ) ;
  assign n3190 = ~n947 & n3189 ;
  assign n3191 = ( n106 & ~n1956 ) | ( n106 & n3190 ) | ( ~n1956 & n3190 ) ;
  assign n3192 = ~n106 & n3191 ;
  assign n3193 = ( n148 & ~n348 ) | ( n148 & n3192 ) | ( ~n348 & n3192 ) ;
  assign n3194 = ~n148 & n3193 ;
  assign n3195 = ( n252 & ~n229 ) | ( n252 & n3194 ) | ( ~n229 & n3194 ) ;
  assign n3196 = ~n252 & n3195 ;
  assign n3197 = ~n431 &  n3196 ;
  assign n3213 = n99 | n151 ;
  assign n3244 = n137 | n374 ;
  assign n3245 = n266 | n3244 ;
  assign n3246 = n268 | n3245 ;
  assign n3247 = n340 | n3246 ;
  assign n3214 = n141 | n284 ;
  assign n3215 = ( n2248 & ~n911 ) | ( n2248 & n3214 ) | ( ~n911 & n3214 ) ;
  assign n3216 = n911 | n3215 ;
  assign n3217 = ( n485 & ~n558 ) | ( n485 & n3216 ) | ( ~n558 & n3216 ) ;
  assign n3218 = n558 | n3217 ;
  assign n3219 = ( n197 & ~n3218 ) | ( n197 & n560 ) | ( ~n3218 & n560 ) ;
  assign n3220 = ~n560 & n3219 ;
  assign n3221 = ~n403 & n3220 ;
  assign n3222 = n140 | n417 ;
  assign n3223 = n494 | n793 ;
  assign n3224 = ( n221 & ~n190 ) | ( n221 & n3223 ) | ( ~n190 & n3223 ) ;
  assign n3225 = n190 | n3224 ;
  assign n3226 = ( n603 & ~n149 ) | ( n603 & n3225 ) | ( ~n149 & n3225 ) ;
  assign n3227 = n149 | n3226 ;
  assign n3228 = n350 | n711 ;
  assign n3229 = n80 | n1152 ;
  assign n3230 = ( n1049 & ~n3228 ) | ( n1049 & n3229 ) | ( ~n3228 & n3229 ) ;
  assign n3231 = n3228 | n3230 ;
  assign n3232 = ( n3227 & ~n3222 ) | ( n3227 & n3231 ) | ( ~n3222 & n3231 ) ;
  assign n3233 = ( n2084 & n3222 ) | ( n2084 & n3232 ) | ( n3222 & n3232 ) ;
  assign n3234 = ( n2084 & ~n3233 ) | ( n2084 & 1'b0 ) | ( ~n3233 & 1'b0 ) ;
  assign n3235 = ( n2187 & n3221 ) | ( n2187 & n3234 ) | ( n3221 & n3234 ) ;
  assign n3236 = ~n2187 & n3235 ;
  assign n3237 = ( n157 & ~n72 ) | ( n157 & n3236 ) | ( ~n72 & n3236 ) ;
  assign n3238 = ~n157 & n3237 ;
  assign n3239 = ( n300 & ~n671 ) | ( n300 & n3238 ) | ( ~n671 & n3238 ) ;
  assign n3240 = ~n300 & n3239 ;
  assign n3241 = ~n212 & n3240 ;
  assign n3242 = ( n1428 & ~n432 ) | ( n1428 & n3241 ) | ( ~n432 & n3241 ) ;
  assign n3243 = ~n1428 & n3242 ;
  assign n3248 = ( n1417 & n3247 ) | ( n1417 & n3243 ) | ( n3247 & n3243 ) ;
  assign n3249 = ( n189 & ~n3248 ) | ( n189 & n3243 ) | ( ~n3248 & n3243 ) ;
  assign n3250 = ~n189 & n3249 ;
  assign n3251 = ( n530 & n2822 ) | ( n530 & n3250 ) | ( n2822 & n3250 ) ;
  assign n3252 = ~n530 & n3251 ;
  assign n3253 = ( n573 & ~n3213 ) | ( n573 & n3252 ) | ( ~n3213 & n3252 ) ;
  assign n3254 = ~n573 & n3253 ;
  assign n3255 = ( n1567 & ~n2576 ) | ( n1567 & n3254 ) | ( ~n2576 & n3254 ) ;
  assign n3256 = ~n1567 & n3255 ;
  assign n3198 = ( n888 & ~n2309 ) | ( n888 & n2752 ) | ( ~n2309 & n2752 ) ;
  assign n3199 = ( n1545 & ~n2752 ) | ( n1545 & n3198 ) | ( ~n2752 & n3198 ) ;
  assign n3200 = ~n1545 & n3199 ;
  assign n3201 = ( n124 & ~n555 ) | ( n124 & n3200 ) | ( ~n555 & n3200 ) ;
  assign n3202 = ~n124 & n3201 ;
  assign n3203 = ( n415 & ~n2063 ) | ( n415 & n3202 ) | ( ~n2063 & n3202 ) ;
  assign n3204 = ~n415 & n3203 ;
  assign n3205 = ( n761 & ~n191 ) | ( n761 & n3204 ) | ( ~n191 & n3204 ) ;
  assign n3206 = ~n761 & n3205 ;
  assign n3207 = ( n3206 & ~n270 ) | ( n3206 & n737 ) | ( ~n270 & n737 ) ;
  assign n3208 = ( n3207 & ~n737 ) | ( n3207 & 1'b0 ) | ( ~n737 & 1'b0 ) ;
  assign n3209 = ( n405 & ~n3208 ) | ( n405 & n623 ) | ( ~n3208 & n623 ) ;
  assign n3210 = ( n623 & ~n3209 ) | ( n623 & 1'b0 ) | ( ~n3209 & 1'b0 ) ;
  assign n3211 = ( n228 & ~n156 ) | ( n228 & n3210 ) | ( ~n156 & n3210 ) ;
  assign n3212 = ~n228 & n3211 ;
  assign n3257 = ( n2923 & ~n3256 ) | ( n2923 & n3212 ) | ( ~n3256 & n3212 ) ;
  assign n3258 = ( n679 & ~n3257 ) | ( n679 & n3212 ) | ( ~n3257 & n3212 ) ;
  assign n3259 = ~n679 & n3258 ;
  assign n3260 = ( n720 & ~n216 ) | ( n720 & n3259 ) | ( ~n216 & n3259 ) ;
  assign n3261 = ~n720 & n3260 ;
  assign n3262 = ( n148 & ~n618 ) | ( n148 & n3261 ) | ( ~n618 & n3261 ) ;
  assign n3263 = ~n148 & n3262 ;
  assign n3264 = ( n129 & ~n256 ) | ( n129 & n3263 ) | ( ~n256 & n3263 ) ;
  assign n3265 = ~n129 & n3264 ;
  assign n3266 = ~n3265 |  n646 ;
  assign n3267 = n332 | n384 ;
  assign n3268 = ( n704 & ~n1398 ) | ( n704 & 1'b0 ) | ( ~n1398 & 1'b0 ) ;
  assign n3269 = ( n3267 & ~n1232 ) | ( n3267 & n3268 ) | ( ~n1232 & n3268 ) ;
  assign n3270 = ( n1887 & ~n3269 ) | ( n1887 & n3267 ) | ( ~n3269 & n3267 ) ;
  assign n3271 = ( n1887 & ~n3270 ) | ( n1887 & 1'b0 ) | ( ~n3270 & 1'b0 ) ;
  assign n3272 = ( n102 & ~n3271 ) | ( n102 & n525 ) | ( ~n3271 & n525 ) ;
  assign n3273 = ( n525 & ~n3272 ) | ( n525 & 1'b0 ) | ( ~n3272 & 1'b0 ) ;
  assign n3274 = ( n271 & ~n1426 ) | ( n271 & n3273 ) | ( ~n1426 & n3273 ) ;
  assign n3275 = ~n271 & n3274 ;
  assign n3276 = ( n279 & ~n737 ) | ( n279 & n3275 ) | ( ~n737 & n3275 ) ;
  assign n3277 = ~n279 & n3276 ;
  assign n3278 = ( n617 & ~n628 ) | ( n617 & n3277 ) | ( ~n628 & n3277 ) ;
  assign n3279 = ~n617 & n3278 ;
  assign n3280 = ~n666 & n3279 ;
  assign n3288 = n404 | n721 ;
  assign n3289 = ( n240 & ~n132 ) | ( n240 & n3288 ) | ( ~n132 & n3288 ) ;
  assign n3290 = n132 | n3289 ;
  assign n3291 = n852 | n1546 ;
  assign n3292 = ( n2840 & ~n3290 ) | ( n2840 & n3291 ) | ( ~n3290 & n3291 ) ;
  assign n3293 = ( n3290 & ~n1063 ) | ( n3290 & n3292 ) | ( ~n1063 & n3292 ) ;
  assign n3294 = n1063 | n3293 ;
  assign n3295 = ( n1884 & ~n1678 ) | ( n1884 & n3294 ) | ( ~n1678 & n3294 ) ;
  assign n3296 = n1678 | n3295 ;
  assign n3297 = ( n195 & ~n461 ) | ( n195 & n3296 ) | ( ~n461 & n3296 ) ;
  assign n3298 = n461 | n3297 ;
  assign n3299 = ( n207 & ~n61 ) | ( n207 & n3298 ) | ( ~n61 & n3298 ) ;
  assign n3300 = n61 | n3299 ;
  assign n3301 = ( n135 & ~n273 ) | ( n135 & n3300 ) | ( ~n273 & n3300 ) ;
  assign n3302 = n273 | n3301 ;
  assign n3303 = n358 | n3302 ;
  assign n3282 = n272 | n373 ;
  assign n3283 = ( n74 & ~n165 ) | ( n74 & n3282 ) | ( ~n165 & n3282 ) ;
  assign n3284 = n165 | n3283 ;
  assign n3285 = ( n340 & ~n276 ) | ( n340 & n3284 ) | ( ~n276 & n3284 ) ;
  assign n3286 = n276 | n3285 ;
  assign n3287 = n353 | n3286 ;
  assign n3304 = n127 | n160 ;
  assign n3305 = n234 | n1072 ;
  assign n3306 = ( n679 & ~n431 ) | ( n679 & n3305 ) | ( ~n431 & n3305 ) ;
  assign n3307 = n431 | n3306 ;
  assign n3308 = ( n3304 & ~n1014 ) | ( n3304 & n3307 ) | ( ~n1014 & n3307 ) ;
  assign n3309 = ( n3308 & ~n1542 ) | ( n3308 & n1014 ) | ( ~n1542 & n1014 ) ;
  assign n3310 = n3309 | n1542 ;
  assign n3311 = ( n3303 & ~n3287 ) | ( n3303 & n3310 ) | ( ~n3287 & n3310 ) ;
  assign n3312 = ( n3241 & n3311 ) | ( n3241 & n3287 ) | ( n3311 & n3287 ) ;
  assign n3313 = ( n3241 & ~n3312 ) | ( n3241 & 1'b0 ) | ( ~n3312 & 1'b0 ) ;
  assign n3281 = n161 | n338 ;
  assign n3314 = ( n645 & ~n3313 ) | ( n645 & n3281 ) | ( ~n3313 & n3281 ) ;
  assign n3315 = ( n645 & ~n3314 ) | ( n645 & 1'b0 ) | ( ~n3314 & 1'b0 ) ;
  assign n3316 = ( n333 & n3280 ) | ( n333 & n3315 ) | ( n3280 & n3315 ) ;
  assign n3317 = ~n333 & n3316 ;
  assign n3318 = ( n349 & ~n191 ) | ( n349 & n3317 ) | ( ~n191 & n3317 ) ;
  assign n3319 = ~n349 & n3318 ;
  assign n3320 = ( n744 & ~n534 ) | ( n744 & n3319 ) | ( ~n534 & n3319 ) ;
  assign n3321 = ~n744 & n3320 ;
  assign n3322 = ( n569 & ~n266 ) | ( n569 & n3321 ) | ( ~n266 & n3321 ) ;
  assign n3323 = ~n569 & n3322 ;
  assign n3324 = ( n196 & ~n285 ) | ( n196 & n3323 ) | ( ~n285 & n3323 ) ;
  assign n3325 = ~n196 & n3324 ;
  assign n3326 = n272 | n812 ;
  assign n3327 = n72 | n91 ;
  assign n3328 = n148 | n3327 ;
  assign n3329 = ( n3229 & ~n3326 ) | ( n3229 & n3328 ) | ( ~n3326 & n3328 ) ;
  assign n3330 = ( n3326 & ~n575 ) | ( n3326 & n3329 ) | ( ~n575 & n3329 ) ;
  assign n3331 = n575 | n3330 ;
  assign n3332 = ( n274 & ~n676 ) | ( n274 & n3331 ) | ( ~n676 & n3331 ) ;
  assign n3333 = n676 | n3332 ;
  assign n3334 = ( n572 & ~n226 ) | ( n572 & n3333 ) | ( ~n226 & n3333 ) ;
  assign n3335 = n226 | n3334 ;
  assign n3336 = ( n630 & ~n431 ) | ( n630 & n3335 ) | ( ~n431 & n3335 ) ;
  assign n3337 = n431 | n3336 ;
  assign n3338 = n231 | n775 ;
  assign n3339 = ( n118 & ~n230 ) | ( n118 & n3338 ) | ( ~n230 & n3338 ) ;
  assign n3340 = n230 | n3339 ;
  assign n3341 = ( n540 & ~n683 ) | ( n540 & n3340 ) | ( ~n683 & n3340 ) ;
  assign n3342 = n683 | n3341 ;
  assign n3343 = ( n236 & ~n300 ) | ( n236 & n3342 ) | ( ~n300 & n3342 ) ;
  assign n3344 = n300 | n3343 ;
  assign n3345 = ( n167 & n354 ) | ( n167 & n3344 ) | ( n354 & n3344 ) ;
  assign n3346 = ( n354 & ~n3345 ) | ( n354 & 1'b0 ) | ( ~n3345 & 1'b0 ) ;
  assign n3347 = ( n975 & ~n1690 ) | ( n975 & n1991 ) | ( ~n1690 & n1991 ) ;
  assign n3348 = n1690 | n3347 ;
  assign n3349 = n2752 | n3348 ;
  assign n3350 = n1853 | n3349 ;
  assign n3351 = ( n2147 & ~n3350 ) | ( n2147 & 1'b0 ) | ( ~n3350 & 1'b0 ) ;
  assign n3352 = ( n3337 & n3346 ) | ( n3337 & n3351 ) | ( n3346 & n3351 ) ;
  assign n3353 = ( n2308 & ~n3337 ) | ( n2308 & n3352 ) | ( ~n3337 & n3352 ) ;
  assign n3354 = ~n2308 & n3353 ;
  assign n3355 = ( n69 & ~n218 ) | ( n69 & n3354 ) | ( ~n218 & n3354 ) ;
  assign n3356 = ~n69 & n3355 ;
  assign n3357 = ( n105 & ~n258 ) | ( n105 & n3356 ) | ( ~n258 & n3356 ) ;
  assign n3358 = ~n105 & n3357 ;
  assign n3359 = ( n457 & ~n531 ) | ( n457 & n3358 ) | ( ~n531 & n3358 ) ;
  assign n3360 = ~n457 & n3359 ;
  assign n3361 = ~n476 & n3360 ;
  assign n3362 = ( x26 & ~n66 ) | ( x26 & 1'b0 ) | ( ~n66 & 1'b0 ) ;
  assign n3363 = ( n38 & ~x26 ) | ( n38 & n3362 ) | ( ~x26 & n3362 ) ;
  assign n3364 = ( n76 & ~n59 ) | ( n76 & n116 ) | ( ~n59 & n116 ) ;
  assign n3365 = ~n116 & n3364 ;
  assign n3366 = ( n60 & ~n94 ) | ( n60 & n82 ) | ( ~n94 & n82 ) ;
  assign n3367 = ~n82 & n3366 ;
  assign n3368 = ( n73 & ~n98 ) | ( n73 & n103 ) | ( ~n98 & n103 ) ;
  assign n3369 = ~n103 & n3368 ;
  assign n3370 = n342 | n812 ;
  assign n3371 = ( n1385 & ~n194 ) | ( n1385 & n3370 ) | ( ~n194 & n3370 ) ;
  assign n3372 = n194 | n3371 ;
  assign n3373 = ( n350 & ~n778 ) | ( n350 & n3372 ) | ( ~n778 & n3372 ) ;
  assign n3374 = n778 | n3373 ;
  assign n3375 = ( n192 & ~n334 ) | ( n192 & n3374 ) | ( ~n334 & n3374 ) ;
  assign n3376 = n334 | n3375 ;
  assign n3377 = n156 | n3376 ;
  assign n3393 = ( n405 & ~n493 ) | ( n405 & n628 ) | ( ~n493 & n628 ) ;
  assign n3394 = n493 | n3393 ;
  assign n3395 = n120 | n216 ;
  assign n3396 = ( n3394 & ~n2672 ) | ( n3394 & n3395 ) | ( ~n2672 & n3395 ) ;
  assign n3397 = n2672 | n3396 ;
  assign n3398 = ( n189 & ~n1672 ) | ( n189 & n3397 ) | ( ~n1672 & n3397 ) ;
  assign n3399 = n1672 | n3398 ;
  assign n3378 = x27 | n50 ;
  assign n3379 = ( x27 & ~n3378 ) | ( x27 & n98 ) | ( ~n3378 & n98 ) ;
  assign n3380 = ( n205 & ~n560 ) | ( n205 & n221 ) | ( ~n560 & n221 ) ;
  assign n3381 = n560 | n3380 ;
  assign n3382 = ( n341 & n354 ) | ( n341 & n1060 ) | ( n354 & n1060 ) ;
  assign n3383 = ( n354 & ~n3382 ) | ( n354 & 1'b0 ) | ( ~n3382 & 1'b0 ) ;
  assign n3384 = ( n3159 & ~n3381 ) | ( n3159 & n3383 ) | ( ~n3381 & n3383 ) ;
  assign n3385 = ~n3159 & n3384 ;
  assign n3386 = ( n1955 & ~n953 ) | ( n1955 & n3385 ) | ( ~n953 & n3385 ) ;
  assign n3387 = ~n1955 & n3386 ;
  assign n3388 = ~n58 & n3387 ;
  assign n3389 = ( n3379 & ~n98 ) | ( n3379 & n3388 ) | ( ~n98 & n3388 ) ;
  assign n3390 = ( n236 & ~n256 ) | ( n236 & n3389 ) | ( ~n256 & n3389 ) ;
  assign n3391 = ~n236 & n3390 ;
  assign n3392 = ~n664 & n3391 ;
  assign n3400 = ( n3377 & ~n3399 ) | ( n3377 & n3392 ) | ( ~n3399 & n3392 ) ;
  assign n3401 = ~n3377 & n3400 ;
  assign n3402 = ( n278 & ~n865 ) | ( n278 & n3401 ) | ( ~n865 & n3401 ) ;
  assign n3403 = ~n278 & n3402 ;
  assign n3404 = ( n408 & ~n668 ) | ( n408 & n3403 ) | ( ~n668 & n3403 ) ;
  assign n3405 = ~n408 & n3404 ;
  assign n3406 = ( n224 & ~n241 ) | ( n224 & n3405 ) | ( ~n241 & n3405 ) ;
  assign n3407 = ~n224 & n3406 ;
  assign n3408 = ~n761 & n3407 ;
  assign n3409 = ( n3369 & ~n73 ) | ( n3369 & n3408 ) | ( ~n73 & n3408 ) ;
  assign n3410 = n259 | n345 ;
  assign n3411 = ( n253 & ~n138 ) | ( n253 & n3410 ) | ( ~n138 & n3410 ) ;
  assign n3412 = n138 | n3411 ;
  assign n3413 = ( n343 & n453 ) | ( n343 & n3412 ) | ( n453 & n3412 ) ;
  assign n3414 = ( n343 & ~n3413 ) | ( n343 & 1'b0 ) | ( ~n3413 & 1'b0 ) ;
  assign n3415 = ( n279 & ~n332 ) | ( n279 & n3414 ) | ( ~n332 & n3414 ) ;
  assign n3416 = ~n279 & n3415 ;
  assign n3417 = ~n643 & n3416 ;
  assign n3418 = n415 | n1702 ;
  assign n3419 = n300 | n3418 ;
  assign n3420 = n125 | n376 ;
  assign n3421 = n559 | n3420 ;
  assign n3422 = ( n3419 & ~n3171 ) | ( n3419 & n3421 ) | ( ~n3171 & n3421 ) ;
  assign n3423 = n3171 | n3422 ;
  assign n3424 = ( n905 & ~n72 ) | ( n905 & n3423 ) | ( ~n72 & n3423 ) ;
  assign n3425 = n72 | n3424 ;
  assign n3426 = n137 | n3425 ;
  assign n3427 = ( n38 & ~n57 ) | ( n38 & n119 ) | ( ~n57 & n119 ) ;
  assign n3428 = ~n119 & n3427 ;
  assign n3429 = n2485 | n2703 ;
  assign n3430 = ( n173 & ~n2632 ) | ( n173 & n3429 ) | ( ~n2632 & n3429 ) ;
  assign n3431 = n2632 | n3430 ;
  assign n3432 = ( n2342 & ~n1828 ) | ( n2342 & n3431 ) | ( ~n1828 & n3431 ) ;
  assign n3433 = n1828 | n3432 ;
  assign n3434 = ( n887 & ~n81 ) | ( n887 & n3433 ) | ( ~n81 & n3433 ) ;
  assign n3435 = n81 | n3434 ;
  assign n3436 = ( n3281 & ~n69 ) | ( n3281 & n3435 ) | ( ~n69 & n3435 ) ;
  assign n3437 = n69 | n3436 ;
  assign n3438 = ( n627 & ~n456 ) | ( n627 & n3437 ) | ( ~n456 & n3437 ) ;
  assign n3439 = n456 | n3438 ;
  assign n3440 = ( n38 & ~n3428 ) | ( n38 & n3439 ) | ( ~n3428 & n3439 ) ;
  assign n3441 = ( n123 & ~n1072 ) | ( n123 & n1360 ) | ( ~n1072 & n1360 ) ;
  assign n3442 = n1072 | n3441 ;
  assign n3443 = n257 | n712 ;
  assign n3444 = ( n43 & n484 ) | ( n43 & n3443 ) | ( n484 & n3443 ) ;
  assign n3445 = ( n484 & ~n3444 ) | ( n484 & 1'b0 ) | ( ~n3444 & 1'b0 ) ;
  assign n3446 = ~n3442 & n3445 ;
  assign n3447 = ( n3426 & ~n3440 ) | ( n3426 & n3446 ) | ( ~n3440 & n3446 ) ;
  assign n3448 = ~n3426 & n3447 ;
  assign n3449 = ( n3417 & ~n3409 ) | ( n3417 & n3448 ) | ( ~n3409 & n3448 ) ;
  assign n3450 = ( n654 & n3409 ) | ( n654 & n3449 ) | ( n3409 & n3449 ) ;
  assign n3451 = ~n654 & n3450 ;
  assign n3452 = ( n842 & ~n675 ) | ( n842 & n3451 ) | ( ~n675 & n3451 ) ;
  assign n3453 = ~n842 & n3452 ;
  assign n3454 = n645 &  n3453 ;
  assign n3455 = ( n3367 & ~n60 ) | ( n3367 & n3454 ) | ( ~n60 & n3454 ) ;
  assign n3456 = ( n787 & ~n452 ) | ( n787 & n3455 ) | ( ~n452 & n3455 ) ;
  assign n3457 = ~n787 & n3456 ;
  assign n3458 = ( n3365 & ~n76 ) | ( n3365 & n3457 ) | ( ~n76 & n3457 ) ;
  assign n3459 = ~n630 & n3458 ;
  assign n3460 = ( ~n38 & n3363 ) | ( ~n38 & n3459 ) | ( n3363 & n3459 ) ;
  assign n3461 = ( n35 & ~n55 ) | ( n35 & n79 ) | ( ~n55 & n79 ) ;
  assign n3462 = ( n79 & ~n3461 ) | ( n79 & 1'b0 ) | ( ~n3461 & 1'b0 ) ;
  assign n3474 = n222 | n864 ;
  assign n3475 = ( n3326 & ~n1430 ) | ( n3326 & n3474 ) | ( ~n1430 & n3474 ) ;
  assign n3476 = ( n1430 & ~n3247 ) | ( n1430 & n3475 ) | ( ~n3247 & n3475 ) ;
  assign n3477 = n3247 | n3476 ;
  assign n3478 = n1617 | n3477 ;
  assign n3479 = n245 | n259 ;
  assign n3480 = ( n2253 & ~n761 ) | ( n2253 & n3479 ) | ( ~n761 & n3479 ) ;
  assign n3481 = n761 | n3480 ;
  assign n3482 = n3478 | n3481 ;
  assign n3463 = n416 | n672 ;
  assign n3464 = n155 | n3463 ;
  assign n3465 = ( n717 & n929 ) | ( n717 & n3464 ) | ( n929 & n3464 ) ;
  assign n3466 = ( n337 & ~n3465 ) | ( n337 & n929 ) | ( ~n3465 & n929 ) ;
  assign n3467 = ~n337 & n3466 ;
  assign n3468 = ( n280 & ~n207 ) | ( n280 & n3467 ) | ( ~n207 & n3467 ) ;
  assign n3469 = ~n280 & n3468 ;
  assign n3470 = ( n350 & ~n348 ) | ( n350 & n3469 ) | ( ~n348 & n3469 ) ;
  assign n3471 = ~n350 & n3470 ;
  assign n3472 = ( n167 & ~n534 ) | ( n167 & n3471 ) | ( ~n534 & n3471 ) ;
  assign n3473 = ~n167 & n3472 ;
  assign n3483 = ( n128 & n3482 ) | ( n128 & n3473 ) | ( n3482 & n3473 ) ;
  assign n3484 = ( n2192 & ~n3483 ) | ( n2192 & n3473 ) | ( ~n3483 & n3473 ) ;
  assign n3485 = ~n2192 & n3484 ;
  assign n3486 = ( n1625 & ~n1360 ) | ( n1625 & n3485 ) | ( ~n1360 & n3485 ) ;
  assign n3487 = ~n1625 & n3486 ;
  assign n3488 = ( n3462 & ~n55 ) | ( n3462 & n3487 ) | ( ~n55 & n3487 ) ;
  assign n3489 = ( n3488 & ~n192 ) | ( n3488 & n714 ) | ( ~n192 & n714 ) ;
  assign n3490 = ( n3489 & ~n714 ) | ( n3489 & 1'b0 ) | ( ~n714 & 1'b0 ) ;
  assign n3491 = ( n74 & ~n104 ) | ( n74 & n3490 ) | ( ~n104 & n3490 ) ;
  assign n3492 = ~n74 & n3491 ;
  assign n3493 = ( n875 & ~n1655 ) | ( n875 & 1'b0 ) | ( ~n1655 & 1'b0 ) ;
  assign n3494 = ( n424 & ~n792 ) | ( n424 & n3493 ) | ( ~n792 & n3493 ) ;
  assign n3495 = ~n424 & n3494 ;
  assign n3496 = ~n558 & n3495 ;
  assign n3503 = n409 | n549 ;
  assign n3504 = n205 | n3503 ;
  assign n3505 = ( n1168 & n1687 ) | ( n1168 & n3504 ) | ( n1687 & n3504 ) ;
  assign n3506 = ( n1168 & ~n3505 ) | ( n1168 & 1'b0 ) | ( ~n3505 & 1'b0 ) ;
  assign n3497 = n425 | n789 ;
  assign n3498 = ( n372 & ~n101 ) | ( n372 & n3497 ) | ( ~n101 & n3497 ) ;
  assign n3499 = n101 | n3498 ;
  assign n3500 = ( n485 & ~n353 ) | ( n485 & n3499 ) | ( ~n353 & n3499 ) ;
  assign n3501 = n353 | n3500 ;
  assign n3502 = n630 | n3501 ;
  assign n3507 = ( n3496 & ~n3506 ) | ( n3496 & n3502 ) | ( ~n3506 & n3502 ) ;
  assign n3508 = ( n2784 & ~n3507 ) | ( n2784 & n3496 ) | ( ~n3507 & n3496 ) ;
  assign n3509 = ~n2784 & n3508 ;
  assign n3510 = ( n906 & ~n70 ) | ( n906 & n3509 ) | ( ~n70 & n3509 ) ;
  assign n3511 = ~n906 & n3510 ;
  assign n3512 = ( n451 & ~n412 ) | ( n451 & n3511 ) | ( ~n412 & n3511 ) ;
  assign n3513 = ~n451 & n3512 ;
  assign n3514 = ( n574 & ~n559 ) | ( n574 & n3513 ) | ( ~n559 & n3513 ) ;
  assign n3515 = ~n574 & n3514 ;
  assign n3516 = ~n643 & n3515 ;
  assign n3527 = n252 | n556 ;
  assign n3528 = ~n495 & n644 ;
  assign n3529 = ~n356 & n3528 ;
  assign n3530 = ( n377 & ~n3529 ) | ( n377 & n198 ) | ( ~n3529 & n198 ) ;
  assign n3531 = ( n198 & ~n3530 ) | ( n198 & n2703 ) | ( ~n3530 & n2703 ) ;
  assign n3532 = ~n2703 & n3531 ;
  assign n3533 = ( n2610 & ~n3527 ) | ( n2610 & n3532 ) | ( ~n3527 & n3532 ) ;
  assign n3534 = ~n2610 & n3533 ;
  assign n3517 = n278 | n1960 ;
  assign n3518 = ( n2348 & ~n1703 ) | ( n2348 & n3517 ) | ( ~n1703 & n3517 ) ;
  assign n3519 = n1703 | n3518 ;
  assign n3520 = ( n195 & ~n788 ) | ( n195 & n3519 ) | ( ~n788 & n3519 ) ;
  assign n3521 = n788 | n3520 ;
  assign n3522 = ( n284 & ~n300 ) | ( n284 & n3521 ) | ( ~n300 & n3521 ) ;
  assign n3523 = n300 | n3522 ;
  assign n3524 = ( n628 & ~n93 ) | ( n628 & n3523 ) | ( ~n93 & n3523 ) ;
  assign n3525 = n93 | n3524 ;
  assign n3526 = n666 | n3525 ;
  assign n3535 = ( n3516 & ~n3534 ) | ( n3516 & n3526 ) | ( ~n3534 & n3526 ) ;
  assign n3536 = ( n3516 & ~n3535 ) | ( n3516 & 1'b0 ) | ( ~n3535 & 1'b0 ) ;
  assign n3537 = ( n1796 & n3492 ) | ( n1796 & n3536 ) | ( n3492 & n3536 ) ;
  assign n3538 = ~n1796 & n3537 ;
  assign n3539 = ( n843 & ~n1045 ) | ( n843 & n3538 ) | ( ~n1045 & n3538 ) ;
  assign n3540 = ~n843 & n3539 ;
  assign n3541 = ( n713 & ~n620 ) | ( n713 & n3540 ) | ( ~n620 & n3540 ) ;
  assign n3542 = ~n713 & n3541 ;
  assign n3543 = ( n671 & ~n413 ) | ( n671 & n3542 ) | ( ~n413 & n3542 ) ;
  assign n3544 = ~n671 & n3543 ;
  assign n3545 = ( n3544 & ~n214 ) | ( n3544 & n745 ) | ( ~n214 & n745 ) ;
  assign n3546 = ( n3545 & ~n745 ) | ( n3545 & 1'b0 ) | ( ~n745 & 1'b0 ) ;
  assign n3547 = ~n554 &  n3546 ;
  assign n3602 = ( n3460 & ~n3547 ) | ( n3460 & 1'b0 ) | ( ~n3547 & 1'b0 ) ;
  assign n3552 = n58 | n227 ;
  assign n3553 = ( n888 & ~n3552 ) | ( n888 & 1'b0 ) | ( ~n3552 & 1'b0 ) ;
  assign n3554 = ( n719 & ~n3553 ) | ( n719 & n2316 ) | ( ~n3553 & n2316 ) ;
  assign n3555 = ( n2316 & ~n3554 ) | ( n2316 & 1'b0 ) | ( ~n3554 & 1'b0 ) ;
  assign n3548 = n96 | n2076 ;
  assign n3549 = ( n221 & ~n240 ) | ( n221 & n3548 ) | ( ~n240 & n3548 ) ;
  assign n3550 = n240 | n3549 ;
  assign n3551 = n104 | n3550 ;
  assign n3556 = ( n3137 & ~n3555 ) | ( n3137 & n3551 ) | ( ~n3555 & n3551 ) ;
  assign n3557 = ( n3137 & ~n3556 ) | ( n3137 & 1'b0 ) | ( ~n3556 & 1'b0 ) ;
  assign n3558 = ( n675 & ~n1061 ) | ( n675 & n3557 ) | ( ~n1061 & n3557 ) ;
  assign n3559 = ~n675 & n3558 ;
  assign n3560 = ( n493 & ~n865 ) | ( n493 & n3559 ) | ( ~n865 & n3559 ) ;
  assign n3561 = ~n493 & n3560 ;
  assign n3562 = ( n271 & ~n492 ) | ( n271 & n3561 ) | ( ~n492 & n3561 ) ;
  assign n3563 = ~n271 & n3562 ;
  assign n3564 = ( n336 & ~n3563 ) | ( n336 & n354 ) | ( ~n3563 & n354 ) ;
  assign n3565 = ( n354 & ~n3564 ) | ( n354 & 1'b0 ) | ( ~n3564 & 1'b0 ) ;
  assign n3569 = n155 | n237 ;
  assign n3570 = n285 | n778 ;
  assign n3571 = ( n3304 & ~n3569 ) | ( n3304 & n3570 ) | ( ~n3569 & n3570 ) ;
  assign n3572 = ( n3569 & ~n2540 ) | ( n3569 & n3571 ) | ( ~n2540 & n3571 ) ;
  assign n3573 = n2540 | n3572 ;
  assign n3574 = ( n425 & ~n233 ) | ( n425 & n3573 ) | ( ~n233 & n3573 ) ;
  assign n3575 = n233 | n3574 ;
  assign n3576 = ( n222 & ~n761 ) | ( n222 & n3575 ) | ( ~n761 & n3575 ) ;
  assign n3577 = n761 | n3576 ;
  assign n3578 = ( n270 & ~n239 ) | ( n270 & n3577 ) | ( ~n239 & n3577 ) ;
  assign n3579 = n239 | n3578 ;
  assign n3580 = ( n229 & ~n670 ) | ( n229 & n3579 ) | ( ~n670 & n3579 ) ;
  assign n3581 = n670 | n3580 ;
  assign n3582 = n526 | n2687 ;
  assign n3583 = ( n572 & ~n347 ) | ( n572 & n3582 ) | ( ~n347 & n3582 ) ;
  assign n3584 = n347 | n3583 ;
  assign n3585 = n569 | n676 ;
  assign n3586 = n459 | n3585 ;
  assign n3587 = ( n1434 & ~n3586 ) | ( n1434 & n3115 ) | ( ~n3586 & n3115 ) ;
  assign n3588 = ~n1434 & n3587 ;
  assign n3589 = ~n3584 & n3588 ;
  assign n3590 = ( n3581 & ~n727 ) | ( n3581 & n3589 ) | ( ~n727 & n3589 ) ;
  assign n3591 = ( n3440 & ~n3581 ) | ( n3440 & n3590 ) | ( ~n3581 & n3590 ) ;
  assign n3592 = ( n3591 & ~n3440 ) | ( n3591 & 1'b0 ) | ( ~n3440 & 1'b0 ) ;
  assign n3593 = ( n2128 & ~n866 ) | ( n2128 & n3592 ) | ( ~n866 & n3592 ) ;
  assign n3594 = ~n2128 & n3593 ;
  assign n3566 = n120 | n672 ;
  assign n3567 = ( n478 & ~n560 ) | ( n478 & n3566 ) | ( ~n560 & n3566 ) ;
  assign n3568 = n560 | n3567 ;
  assign n3595 = ( n3565 & ~n3594 ) | ( n3565 & n3568 ) | ( ~n3594 & n3568 ) ;
  assign n3596 = ( n947 & ~n3595 ) | ( n947 & n3565 ) | ( ~n3595 & n3565 ) ;
  assign n3597 = ~n947 & n3596 ;
  assign n3598 = ( n274 & ~n911 ) | ( n274 & n3597 ) | ( ~n911 & n3597 ) ;
  assign n3599 = ~n274 & n3598 ;
  assign n3600 = ( n135 & ~n3599 ) | ( n135 & n623 ) | ( ~n3599 & n623 ) ;
  assign n3601 = n623 &  ~n3600 ;
  assign n3603 = ( n3460 & ~n3602 ) | ( n3460 & n3601 ) | ( ~n3602 & n3601 ) ;
  assign n3604 = ( n3361 & n3460 ) | ( n3361 & n3603 ) | ( n3460 & n3603 ) ;
  assign n3605 = ( n3325 & n3361 ) | ( n3325 & n3604 ) | ( n3361 & n3604 ) ;
  assign n3606 = ( n3325 & ~n3266 ) | ( n3325 & n3605 ) | ( ~n3266 & n3605 ) ;
  assign n3607 = ( n3197 & ~n3266 ) | ( n3197 & n3606 ) | ( ~n3266 & n3606 ) ;
  assign n3608 = ( n3106 & n3197 ) | ( n3106 & n3607 ) | ( n3197 & n3607 ) ;
  assign n3609 = ( n3030 & n3106 ) | ( n3030 & n3608 ) | ( n3106 & n3608 ) ;
  assign n3610 = ( n2995 & n3030 ) | ( n2995 & n3609 ) | ( n3030 & n3609 ) ;
  assign n3611 = ( n2839 & n2995 ) | ( n2839 & n3610 ) | ( n2995 & n3610 ) ;
  assign n3612 = ( n2783 & ~n2839 ) | ( n2783 & n3611 ) | ( ~n2839 & n3611 ) ;
  assign n3613 = ( n2839 & ~n2910 ) | ( n2839 & n3612 ) | ( ~n2910 & n3612 ) ;
  assign n3614 = ( n2751 & n2783 ) | ( n2751 & n3613 ) | ( n2783 & n3613 ) ;
  assign n3615 = ( n2665 & n2751 ) | ( n2665 & n3614 ) | ( n2751 & n3614 ) ;
  assign n3616 = ( n2569 & n2665 ) | ( n2569 & n3615 ) | ( n2665 & n3615 ) ;
  assign n3617 = ( n2483 & n2569 ) | ( n2483 & n3616 ) | ( n2569 & n3616 ) ;
  assign n3618 = ( n2392 & n2483 ) | ( n2392 & n3617 ) | ( n2483 & n3617 ) ;
  assign n3619 = ( n2296 & n2392 ) | ( n2296 & n3618 ) | ( n2392 & n3618 ) ;
  assign n3620 = ( n2178 & n2296 ) | ( n2178 & n3619 ) | ( n2296 & n3619 ) ;
  assign n3621 = ( n2127 & n2178 ) | ( n2127 & n3620 ) | ( n2178 & n3620 ) ;
  assign n3622 = ( n2022 & n2127 ) | ( n2022 & n3621 ) | ( n2127 & n3621 ) ;
  assign n3623 = ( n1940 & n2022 ) | ( n1940 & n3622 ) | ( n2022 & n3622 ) ;
  assign n3624 = ( n1875 & n1940 ) | ( n1875 & n3623 ) | ( n1940 & n3623 ) ;
  assign n3625 = ( n1748 & n1875 ) | ( n1748 & n3624 ) | ( n1875 & n3624 ) ;
  assign n3626 = ( n1671 & n1748 ) | ( n1671 & n3625 ) | ( n1748 & n3625 ) ;
  assign n3627 = ( n1566 & n1671 ) | ( n1566 & n3626 ) | ( n1671 & n3626 ) ;
  assign n3628 = ( n1566 & ~n1483 ) | ( n1566 & n3627 ) | ( ~n1483 & n3627 ) ;
  assign n3629 = ( n1378 & ~n1483 ) | ( n1378 & n3628 ) | ( ~n1483 & n3628 ) ;
  assign n3630 = ( n1378 & ~n1267 ) | ( n1378 & n3629 ) | ( ~n1267 & n3629 ) ;
  assign n3631 = ( n1151 & ~n1267 ) | ( n1151 & n3630 ) | ( ~n1267 & n3630 ) ;
  assign n3632 = ( n1043 & n1151 ) | ( n1043 & n3631 ) | ( n1151 & n3631 ) ;
  assign n3633 = ( n946 & n1043 ) | ( n946 & n3632 ) | ( n1043 & n3632 ) ;
  assign n3634 = ( n863 & n946 ) | ( n863 & n3633 ) | ( n946 & n3633 ) ;
  assign n3635 = ( n702 & n863 ) | ( n702 & n3634 ) | ( n863 & n3634 ) ;
  assign n3636 = ~n702 & n3635 ;
  assign n3637 = ( n599 & ~n3636 ) | ( n599 & n3635 ) | ( ~n3636 & n3635 ) ;
  assign n3638 = n601 | n3637 ;
  assign n3639 = n600 &  n3638 ;
  assign n3640 = ~x29 & n3639 ;
  assign n3641 = ( x29 & ~n3639 ) | ( x29 & 1'b0 ) | ( ~n3639 & 1'b0 ) ;
  assign n3642 = n3640 | n3641 ;
  assign n3645 = n702 | n863 ;
  assign n3646 = n702 &  n863 ;
  assign n3647 = ( n3645 & ~n3646 ) | ( n3645 & 1'b0 ) | ( ~n3646 & 1'b0 ) ;
  assign n3648 = ~n3634 & n3647 ;
  assign n3649 = ( n3634 & ~n3647 ) | ( n3634 & 1'b0 ) | ( ~n3647 & 1'b0 ) ;
  assign n3650 = n3648 | n3649 ;
  assign n3651 = n3644 | n3650 ;
  assign n3652 = x31 &  n50 ;
  assign n3660 = n3652 | n946 ;
  assign n3653 = ~n3643 |  x31 ;
  assign n3654 = n702 | n3653 ;
  assign n3655 = ( x30 & x31 ) | ( x30 & n54 ) | ( x31 & n54 ) ;
  assign n3656 = ( x30 & ~n37 ) | ( x30 & x31 ) | ( ~n37 & x31 ) ;
  assign n3657 = ~n3655 & n3656 ;
  assign n3658 = ~n863 & n3657 ;
  assign n3659 = ( n3654 & ~n3658 ) | ( n3654 & 1'b0 ) | ( ~n3658 & 1'b0 ) ;
  assign n3661 = ( n946 & ~n3660 ) | ( n946 & n3659 ) | ( ~n3660 & n3659 ) ;
  assign n3662 = n3651 &  n3661 ;
  assign n3663 = n271 | n338 ;
  assign n3664 = n217 | n266 ;
  assign n3665 = n256 | n3664 ;
  assign n3666 = ( n159 & ~n3663 ) | ( n159 & n3665 ) | ( ~n3663 & n3665 ) ;
  assign n3667 = ( n3663 & ~n2976 ) | ( n3663 & n3666 ) | ( ~n2976 & n3666 ) ;
  assign n3668 = n2976 | n3667 ;
  assign n3669 = ( n3110 & n3668 ) | ( n3110 & n3041 ) | ( n3668 & n3041 ) ;
  assign n3670 = ( n3041 & ~n3669 ) | ( n3041 & 1'b0 ) | ( ~n3669 & 1'b0 ) ;
  assign n3671 = ( n1567 & ~n1820 ) | ( n1567 & n3670 ) | ( ~n1820 & n3670 ) ;
  assign n3672 = ~n1567 & n3671 ;
  assign n3673 = ( n1490 & ~n461 ) | ( n1490 & n3672 ) | ( ~n461 & n3672 ) ;
  assign n3674 = ~n1490 & n3673 ;
  assign n3675 = ( n235 & ~n3674 ) | ( n235 & n813 ) | ( ~n3674 & n813 ) ;
  assign n3676 = ( n813 & ~n3675 ) | ( n813 & 1'b0 ) | ( ~n3675 & 1'b0 ) ;
  assign n3677 = ( n333 & ~n793 ) | ( n333 & n3676 ) | ( ~n793 & n3676 ) ;
  assign n3678 = ~n333 & n3677 ;
  assign n3679 = ~n137 & n3678 ;
  assign n3680 = ~n558 & n644 ;
  assign n3681 = ~n136 & n3680 ;
  assign n3682 = n142 | n1678 ;
  assign n3683 = ( n1824 & ~n679 ) | ( n1824 & n3682 ) | ( ~n679 & n3682 ) ;
  assign n3684 = n679 | n3683 ;
  assign n3685 = ( n602 & n786 ) | ( n602 & n3684 ) | ( n786 & n3684 ) ;
  assign n3686 = ( n786 & ~n3685 ) | ( n786 & 1'b0 ) | ( ~n3685 & 1'b0 ) ;
  assign n3687 = ( n424 & ~n191 ) | ( n424 & n3686 ) | ( ~n191 & n3686 ) ;
  assign n3688 = ~n424 & n3687 ;
  assign n3689 = ( n230 & ~n556 ) | ( n230 & n3688 ) | ( ~n556 & n3688 ) ;
  assign n3690 = ~n230 & n3689 ;
  assign n3691 = ( n623 & ~n3690 ) | ( n623 & n666 ) | ( ~n3690 & n666 ) ;
  assign n3692 = ( n623 & ~n3691 ) | ( n623 & 1'b0 ) | ( ~n3691 & 1'b0 ) ;
  assign n3693 = n281 | n382 ;
  assign n3694 = n643 | n3693 ;
  assign n3695 = n2090 | n3694 ;
  assign n3696 = ( n811 & ~n1428 ) | ( n811 & n3695 ) | ( ~n1428 & n3695 ) ;
  assign n3697 = n1428 | n3696 ;
  assign n3698 = ( n779 & ~n604 ) | ( n779 & n3697 ) | ( ~n604 & n3697 ) ;
  assign n3699 = n604 | n3698 ;
  assign n3700 = ( n479 & ~n258 ) | ( n479 & n3699 ) | ( ~n258 & n3699 ) ;
  assign n3701 = n258 | n3700 ;
  assign n3702 = ( n372 & ~n277 ) | ( n372 & n3701 ) | ( ~n277 & n3701 ) ;
  assign n3703 = n277 | n3702 ;
  assign n3704 = ( n91 & ~n89 ) | ( n91 & n3703 ) | ( ~n89 & n3703 ) ;
  assign n3705 = n89 | n3704 ;
  assign n3706 = ( n540 & ~n213 ) | ( n540 & n3705 ) | ( ~n213 & n3705 ) ;
  assign n3707 = n213 | n3706 ;
  assign n3708 = ( n354 & ~n3707 ) | ( n354 & 1'b0 ) | ( ~n3707 & 1'b0 ) ;
  assign n3709 = n80 | n99 ;
  assign n3710 = n83 | n3709 ;
  assign n3711 = n1004 | n3710 ;
  assign n3712 = ( n683 & ~n1617 ) | ( n683 & n3711 ) | ( ~n1617 & n3711 ) ;
  assign n3713 = n1617 | n3712 ;
  assign n3714 = ( n1425 & ~n3713 ) | ( n1425 & 1'b0 ) | ( ~n3713 & 1'b0 ) ;
  assign n3715 = ( n3708 & ~n3692 ) | ( n3708 & n3714 ) | ( ~n3692 & n3714 ) ;
  assign n3716 = ( n3692 & ~n3681 ) | ( n3692 & n3715 ) | ( ~n3681 & n3715 ) ;
  assign n3717 = n3681 &  n3716 ;
  assign n3718 = ( n677 & n3679 ) | ( n677 & n3717 ) | ( n3679 & n3717 ) ;
  assign n3719 = ~n677 & n3718 ;
  assign n3720 = ( n65 & ~n647 ) | ( n65 & n3719 ) | ( ~n647 & n3719 ) ;
  assign n3721 = ~n65 & n3720 ;
  assign n3722 = ( n192 & ~n348 ) | ( n192 & n3721 ) | ( ~n348 & n3721 ) ;
  assign n3723 = ~n192 & n3722 ;
  assign n3724 = ( n549 & ~n120 ) | ( n549 & n3723 ) | ( ~n120 & n3723 ) ;
  assign n3725 = ~n549 & n3724 ;
  assign n3726 = ( n454 & ~n526 ) | ( n454 & n3725 ) | ( ~n526 & n3725 ) ;
  assign n3727 = ( n3726 & ~n454 ) | ( n3726 & 1'b0 ) | ( ~n454 & 1'b0 ) ;
  assign n3728 = n260 | n279 ;
  assign n3729 = n347 | n3728 ;
  assign n3730 = ( n223 & ~n3663 ) | ( n223 & n3729 ) | ( ~n3663 & n3729 ) ;
  assign n3731 = n3663 | n3730 ;
  assign n3732 = ( n747 & ~n101 ) | ( n747 & n3731 ) | ( ~n101 & n3731 ) ;
  assign n3733 = n101 | n3732 ;
  assign n3734 = ( n187 & ~n162 ) | ( n187 & n3733 ) | ( ~n162 & n3733 ) ;
  assign n3735 = n162 | n3734 ;
  assign n3736 = ( n88 & ~n95 ) | ( n88 & n3735 ) | ( ~n95 & n3735 ) ;
  assign n3737 = n95 | n3736 ;
  assign n3738 = n196 | n3737 ;
  assign n3739 = n267 | n485 ;
  assign n3740 = ( n43 & ~n300 ) | ( n43 & n3739 ) | ( ~n300 & n3739 ) ;
  assign n3741 = n300 | n3740 ;
  assign n3742 = n669 | n1357 ;
  assign n3743 = ( n234 & ~n3742 ) | ( n234 & n929 ) | ( ~n3742 & n929 ) ;
  assign n3744 = ~n234 & n3743 ;
  assign n3745 = ( n122 & ~n243 ) | ( n122 & n3744 ) | ( ~n243 & n3744 ) ;
  assign n3746 = ~n122 & n3745 ;
  assign n3747 = ( n744 & ~n404 ) | ( n744 & n3746 ) | ( ~n404 & n3746 ) ;
  assign n3748 = ~n744 & n3747 ;
  assign n3749 = ( n148 & ~n139 ) | ( n148 & n3748 ) | ( ~n139 & n3748 ) ;
  assign n3750 = ~n148 & n3749 ;
  assign n3751 = ( n459 & ~n618 ) | ( n459 & n3750 ) | ( ~n618 & n3750 ) ;
  assign n3752 = ~n459 & n3751 ;
  assign n3753 = ~n358 & n3752 ;
  assign n3754 = ( n561 & ~n161 ) | ( n561 & n3753 ) | ( ~n161 & n3753 ) ;
  assign n3755 = ~n561 & n3754 ;
  assign n3756 = ~n617 & n3755 ;
  assign n3757 = ( n2112 & ~n3326 ) | ( n2112 & 1'b0 ) | ( ~n3326 & 1'b0 ) ;
  assign n3758 = ( n2629 & n3756 ) | ( n2629 & n3757 ) | ( n3756 & n3757 ) ;
  assign n3759 = ~n2629 & n3758 ;
  assign n3760 = ( n3738 & ~n3741 ) | ( n3738 & n3759 ) | ( ~n3741 & n3759 ) ;
  assign n3761 = ( n2147 & ~n3760 ) | ( n2147 & n3738 ) | ( ~n3760 & n3738 ) ;
  assign n3762 = ( n2147 & ~n3761 ) | ( n2147 & 1'b0 ) | ( ~n3761 & 1'b0 ) ;
  assign n3763 = ( n238 & ~n171 ) | ( n238 & n3762 ) | ( ~n171 & n3762 ) ;
  assign n3764 = ~n238 & n3763 ;
  assign n3765 = ( n1761 & ~n2191 ) | ( n1761 & n3764 ) | ( ~n2191 & n3764 ) ;
  assign n3766 = ( n3765 & ~n1761 ) | ( n3765 & 1'b0 ) | ( ~n1761 & 1'b0 ) ;
  assign n3767 = ( n912 & ~n1426 ) | ( n912 & n3766 ) | ( ~n1426 & n3766 ) ;
  assign n3768 = ~n912 & n3767 ;
  assign n3769 = ( n124 & ~n194 ) | ( n124 & n3768 ) | ( ~n194 & n3768 ) ;
  assign n3770 = ~n124 & n3769 ;
  assign n3771 = ( n671 & ~n424 ) | ( n671 & n3770 ) | ( ~n424 & n3770 ) ;
  assign n3772 = ~n671 & n3771 ;
  assign n3773 = ( n554 & ~n734 ) | ( n554 & n3772 ) | ( ~n734 & n3772 ) ;
  assign n3774 = ~n554 & n3773 ;
  assign n3775 = ( n628 & ~n353 ) | ( n628 & n3774 ) | ( ~n353 & n3774 ) ;
  assign n3776 = ~n628 & n3775 ;
  assign n3777 = n359 | n424 ;
  assign n3778 = n376 | n493 ;
  assign n3779 = ( n52 & ~n253 ) | ( n52 & n3778 ) | ( ~n253 & n3778 ) ;
  assign n3780 = n253 | n3779 ;
  assign n3781 = ( n711 & ~n239 ) | ( n711 & n3780 ) | ( ~n239 & n3780 ) ;
  assign n3782 = n239 | n3781 ;
  assign n3783 = ( n340 & ~n276 ) | ( n340 & n3782 ) | ( ~n276 & n3782 ) ;
  assign n3784 = n276 | n3783 ;
  assign n3785 = ( n415 & n813 ) | ( n415 & n3710 ) | ( n813 & n3710 ) ;
  assign n3786 = ( n813 & ~n3785 ) | ( n813 & 1'b0 ) | ( ~n3785 & 1'b0 ) ;
  assign n3787 = ( n453 & ~n765 ) | ( n453 & n3786 ) | ( ~n765 & n3786 ) ;
  assign n3788 = ~n453 & n3787 ;
  assign n3801 = ~n257 & n786 ;
  assign n3802 = ~n333 & n3801 ;
  assign n3789 = n338 | n408 ;
  assign n3790 = n93 | n3789 ;
  assign n3791 = n602 | n678 ;
  assign n3792 = n217 | n3791 ;
  assign n3793 = ( n3790 & ~n72 ) | ( n3790 & n3792 ) | ( ~n72 & n3792 ) ;
  assign n3794 = n72 | n3793 ;
  assign n3795 = ( n206 & ~n224 ) | ( n206 & n3794 ) | ( ~n224 & n3794 ) ;
  assign n3796 = n224 | n3795 ;
  assign n3797 = ( n540 & ~n226 ) | ( n540 & n3796 ) | ( ~n226 & n3796 ) ;
  assign n3798 = n226 | n3797 ;
  assign n3799 = ( n617 & ~n459 ) | ( n617 & n3798 ) | ( ~n459 & n3798 ) ;
  assign n3800 = n459 | n3799 ;
  assign n3803 = ( n3788 & ~n3802 ) | ( n3788 & n3800 ) | ( ~n3802 & n3800 ) ;
  assign n3804 = ( n70 & ~n3803 ) | ( n70 & n3788 ) | ( ~n3803 & n3788 ) ;
  assign n3805 = ~n70 & n3804 ;
  assign n3806 = ( n355 & ~n3805 ) | ( n355 & n1490 ) | ( ~n3805 & n1490 ) ;
  assign n3807 = ( n355 & ~n3806 ) | ( n355 & 1'b0 ) | ( ~n3806 & 1'b0 ) ;
  assign n3808 = ( n242 & ~n3479 ) | ( n242 & n3807 ) | ( ~n3479 & n3807 ) ;
  assign n3809 = ~n242 & n3808 ;
  assign n3810 = ( n273 & ~n418 ) | ( n273 & n3809 ) | ( ~n418 & n3809 ) ;
  assign n3811 = ~n273 & n3810 ;
  assign n3812 = ( n299 & ~n123 ) | ( n299 & n3811 ) | ( ~n123 & n3811 ) ;
  assign n3813 = ~n299 & n3812 ;
  assign n3814 = ( n43 & ~n156 ) | ( n43 & n3813 ) | ( ~n156 & n3813 ) ;
  assign n3815 = ~n43 & n3814 ;
  assign n3816 = n1600 | n2515 ;
  assign n3817 = ( n718 & ~n712 ) | ( n718 & n3816 ) | ( ~n712 & n3816 ) ;
  assign n3818 = n712 | n3817 ;
  assign n3819 = ( n191 & ~n222 ) | ( n191 & n3818 ) | ( ~n222 & n3818 ) ;
  assign n3820 = n222 | n3819 ;
  assign n3821 = ( n451 & n524 ) | ( n451 & n3820 ) | ( n524 & n3820 ) ;
  assign n3822 = ( n524 & ~n3821 ) | ( n524 & 1'b0 ) | ( ~n3821 & 1'b0 ) ;
  assign n3823 = ( n268 & ~n569 ) | ( n268 & n3822 ) | ( ~n569 & n3822 ) ;
  assign n3824 = ~n268 & n3823 ;
  assign n3825 = ( n74 & ~n559 ) | ( n74 & n3824 ) | ( ~n559 & n3824 ) ;
  assign n3826 = ~n74 & n3825 ;
  assign n3827 = n234 | n574 ;
  assign n3828 = n169 | n3827 ;
  assign n3829 = ( n1047 & ~n2752 ) | ( n1047 & n3828 ) | ( ~n2752 & n3828 ) ;
  assign n3830 = n2752 | n3829 ;
  assign n3831 = ( n3815 & ~n3826 ) | ( n3815 & n3830 ) | ( ~n3826 & n3830 ) ;
  assign n3832 = ( n3815 & ~n3831 ) | ( n3815 & 1'b0 ) | ( ~n3831 & 1'b0 ) ;
  assign n3833 = ( n2451 & ~n3832 ) | ( n2451 & n3304 ) | ( ~n3832 & n3304 ) ;
  assign n3834 = ( n2451 & ~n3833 ) | ( n2451 & 1'b0 ) | ( ~n3833 & 1'b0 ) ;
  assign n3835 = ( n843 & ~n654 ) | ( n843 & n3834 ) | ( ~n654 & n3834 ) ;
  assign n3836 = ~n843 & n3835 ;
  assign n3837 = ( n1484 & ~n3784 ) | ( n1484 & n3836 ) | ( ~n3784 & n3836 ) ;
  assign n3838 = ~n1484 & n3837 ;
  assign n3839 = ( n673 & ~n3777 ) | ( n673 & n3838 ) | ( ~n3777 & n3838 ) ;
  assign n3840 = ~n673 & n3839 ;
  assign n3841 = ( n62 & ~n275 ) | ( n62 & n3840 ) | ( ~n275 & n3840 ) ;
  assign n3842 = ~n62 & n3841 ;
  assign n3843 = ( n456 & ~n348 ) | ( n456 & n3842 ) | ( ~n348 & n3842 ) ;
  assign n3844 = ~n456 & n3843 ;
  assign n3845 = ( n670 & ~n356 ) | ( n670 & n3844 ) | ( ~n356 & n3844 ) ;
  assign n3846 = ~n670 & n3845 ;
  assign n3873 = n190 | n765 ;
  assign n3874 = ( n540 & ~n347 ) | ( n540 & n3873 ) | ( ~n347 & n3873 ) ;
  assign n3875 = n347 | n3874 ;
  assign n3876 = n570 | n737 ;
  assign n3877 = ( n281 & ~n572 ) | ( n281 & n3876 ) | ( ~n572 & n3876 ) ;
  assign n3878 = n572 | n3877 ;
  assign n3879 = n3875 | n3878 ;
  assign n3880 = ( n1245 & ~n409 ) | ( n1245 & n3879 ) | ( ~n409 & n3879 ) ;
  assign n3881 = n409 | n3880 ;
  assign n3882 = ( n241 & ~n299 ) | ( n241 & n3881 ) | ( ~n299 & n3881 ) ;
  assign n3883 = n299 | n3882 ;
  assign n3884 = ( n212 & ~n252 ) | ( n212 & n3883 ) | ( ~n252 & n3883 ) ;
  assign n3885 = n252 | n3884 ;
  assign n3886 = n332 | n434 ;
  assign n3887 = ( n39 & ~n95 ) | ( n39 & n3886 ) | ( ~n95 & n3886 ) ;
  assign n3888 = n95 | n3887 ;
  assign n3889 = n160 | n556 ;
  assign n3890 = n196 | n456 ;
  assign n3891 = n61 | n3890 ;
  assign n3892 = n240 | n3891 ;
  assign n3893 = n3889 | n3892 ;
  assign n3894 = ( n3492 & ~n3893 ) | ( n3492 & n3888 ) | ( ~n3893 & n3888 ) ;
  assign n3895 = ( n2468 & ~n3888 ) | ( n2468 & n3894 ) | ( ~n3888 & n3894 ) ;
  assign n3896 = ~n2468 & n3895 ;
  assign n3847 = n2348 | n2548 ;
  assign n3848 = ( n349 & ~n244 ) | ( n349 & n3847 ) | ( ~n244 & n3847 ) ;
  assign n3849 = n244 | n3848 ;
  assign n3850 = ( n494 & ~n101 ) | ( n494 & n3849 ) | ( ~n101 & n3849 ) ;
  assign n3851 = n101 | n3850 ;
  assign n3852 = ( n135 & ~n300 ) | ( n135 & n3851 ) | ( ~n300 & n3851 ) ;
  assign n3853 = n300 | n3852 ;
  assign n3854 = n285 | n382 ;
  assign n3855 = n679 | n745 ;
  assign n3856 = n93 | n3855 ;
  assign n3857 = ( n3854 & ~n1729 ) | ( n3854 & n3856 ) | ( ~n1729 & n3856 ) ;
  assign n3858 = n1729 | n3857 ;
  assign n3859 = ( n3853 & ~n794 ) | ( n3853 & n3858 ) | ( ~n794 & n3858 ) ;
  assign n3860 = n794 | n3859 ;
  assign n3861 = ( n1184 & ~n1511 ) | ( n1184 & n3860 ) | ( ~n1511 & n3860 ) ;
  assign n3862 = n1511 | n3861 ;
  assign n3863 = ( n1427 & ~n238 ) | ( n1427 & n3862 ) | ( ~n238 & n3862 ) ;
  assign n3864 = n238 | n3863 ;
  assign n3865 = ( n260 & ~n157 ) | ( n260 & n3864 ) | ( ~n157 & n3864 ) ;
  assign n3866 = n157 | n3865 ;
  assign n3867 = ( n793 & ~n226 ) | ( n793 & n3866 ) | ( ~n226 & n3866 ) ;
  assign n3868 = n226 | n3867 ;
  assign n3869 = ( n404 & n3868 ) | ( n404 & n524 ) | ( n3868 & n524 ) ;
  assign n3870 = ( n524 & ~n3869 ) | ( n524 & 1'b0 ) | ( ~n3869 & 1'b0 ) ;
  assign n3871 = ( n162 & ~n646 ) | ( n162 & n3870 ) | ( ~n646 & n3870 ) ;
  assign n3872 = ~n162 & n3871 ;
  assign n3897 = ( n3885 & ~n3896 ) | ( n3885 & n3872 ) | ( ~n3896 & n3872 ) ;
  assign n3898 = ( n1385 & ~n3897 ) | ( n1385 & n3872 ) | ( ~n3897 & n3872 ) ;
  assign n3899 = ~n1385 & n3898 ;
  assign n3900 = ( n1244 & ~n3213 ) | ( n1244 & n3899 ) | ( ~n3213 & n3899 ) ;
  assign n3901 = ~n1244 & n3900 ;
  assign n3902 = ( n1152 & ~n357 ) | ( n1152 & n3901 ) | ( ~n357 & n3901 ) ;
  assign n3903 = ~n1152 & n3902 ;
  assign n3904 = ( n234 & ~n775 ) | ( n234 & n3903 ) | ( ~n775 & n3903 ) ;
  assign n3905 = ~n234 & n3904 ;
  assign n3906 = ( n558 & ~n561 ) | ( n558 & n3905 ) | ( ~n561 & n3905 ) ;
  assign n3907 = ~n558 & n3906 ;
  assign n3908 = ( x26 & n3846 ) | ( x26 & n3907 ) | ( n3846 & n3907 ) ;
  assign n3909 = n863 | n946 ;
  assign n3910 = n863 &  n946 ;
  assign n3911 = ( n3909 & ~n3910 ) | ( n3909 & 1'b0 ) | ( ~n3910 & 1'b0 ) ;
  assign n3912 = ~n3633 & n3911 ;
  assign n3913 = ( n3633 & ~n3911 ) | ( n3633 & 1'b0 ) | ( ~n3911 & 1'b0 ) ;
  assign n3914 = n3912 | n3913 ;
  assign n3915 = n3644 | n3914 ;
  assign n3919 = n946 | n3657 ;
  assign n3916 = n863 | n3653 ;
  assign n3917 = ~n1043 & n3652 ;
  assign n3918 = ( n3916 & ~n3917 ) | ( n3916 & 1'b0 ) | ( ~n3917 & 1'b0 ) ;
  assign n3920 = ( n946 & ~n3919 ) | ( n946 & n3918 ) | ( ~n3919 & n3918 ) ;
  assign n3921 = n3915 &  n3920 ;
  assign n3922 = ( n3908 & ~n3727 ) | ( n3908 & n3921 ) | ( ~n3727 & n3921 ) ;
  assign n3923 = ( n3727 & ~n3776 ) | ( n3727 & n3922 ) | ( ~n3776 & n3922 ) ;
  assign n3924 = ( n3727 & ~n3922 ) | ( n3727 & n3776 ) | ( ~n3922 & n3776 ) ;
  assign n3925 = ( n3923 & ~n3727 ) | ( n3923 & n3924 ) | ( ~n3727 & n3924 ) ;
  assign n3926 = ( n3642 & ~n3662 ) | ( n3642 & n3925 ) | ( ~n3662 & n3925 ) ;
  assign n3927 = ( n3662 & ~n3642 ) | ( n3662 & n3925 ) | ( ~n3642 & n3925 ) ;
  assign n3928 = ( n3926 & ~n3925 ) | ( n3926 & n3927 ) | ( ~n3925 & n3927 ) ;
  assign n3947 = n1043 | n1151 ;
  assign n3948 = n1043 &  n1151 ;
  assign n3949 = ( n3947 & ~n3948 ) | ( n3947 & 1'b0 ) | ( ~n3948 & 1'b0 ) ;
  assign n3950 = ~n3631 & n3949 ;
  assign n3951 = ( n3631 & ~n3949 ) | ( n3631 & 1'b0 ) | ( ~n3949 & 1'b0 ) ;
  assign n3952 = n3950 | n3951 ;
  assign n3953 = n3644 | n3952 ;
  assign n3954 = n1043 | n3653 ;
  assign n3955 = ~n1151 & n3657 ;
  assign n3956 = ( n3954 & ~n3955 ) | ( n3954 & 1'b0 ) | ( ~n3955 & 1'b0 ) ;
  assign n3957 = ( n1267 & ~n3652 ) | ( n1267 & 1'b0 ) | ( ~n3652 & 1'b0 ) ;
  assign n3958 = ( n3956 & ~n1267 ) | ( n3956 & n3957 ) | ( ~n1267 & n3957 ) ;
  assign n3959 = n3953 &  n3958 ;
  assign n3960 = n65 | n101 ;
  assign n3961 = n559 | n3960 ;
  assign n3962 = ( n654 & ~n668 ) | ( n654 & n3961 ) | ( ~n668 & n3961 ) ;
  assign n3963 = ( n668 & n1701 ) | ( n668 & n3962 ) | ( n1701 & n3962 ) ;
  assign n3964 = ( n1701 & ~n3963 ) | ( n1701 & 1'b0 ) | ( ~n3963 & 1'b0 ) ;
  assign n3965 = ( n362 & ~n373 ) | ( n362 & n3964 ) | ( ~n373 & n3964 ) ;
  assign n3966 = ~n362 & n3965 ;
  assign n3967 = ( n118 & ~n80 ) | ( n118 & n3966 ) | ( ~n80 & n3966 ) ;
  assign n3968 = ~n118 & n3967 ;
  assign n3969 = ( n236 & ~n137 ) | ( n236 & n3968 ) | ( ~n137 & n3968 ) ;
  assign n3970 = ~n236 & n3969 ;
  assign n3971 = ~n431 & n3970 ;
  assign n3972 = n415 | n571 ;
  assign n3973 = n478 | n3972 ;
  assign n3974 = ( n2996 & ~n260 ) | ( n2996 & n3973 ) | ( ~n260 & n3973 ) ;
  assign n3975 = n260 | n3974 ;
  assign n3976 = ( n69 & ~n333 ) | ( n69 & n3975 ) | ( ~n333 & n3975 ) ;
  assign n3977 = n333 | n3976 ;
  assign n3978 = ( n720 & ~n276 ) | ( n720 & n3977 ) | ( ~n276 & n3977 ) ;
  assign n3979 = n276 | n3978 ;
  assign n3980 = n106 | n235 ;
  assign n3981 = ( n718 & n786 ) | ( n718 & n3980 ) | ( n786 & n3980 ) ;
  assign n3982 = ( n786 & ~n3981 ) | ( n786 & 1'b0 ) | ( ~n3981 & 1'b0 ) ;
  assign n3983 = ( n95 & ~n99 ) | ( n95 & n3982 ) | ( ~n99 & n3982 ) ;
  assign n3984 = ~n95 & n3983 ;
  assign n3985 = n150 | n212 ;
  assign n3986 = n225 | n3985 ;
  assign n3987 = ( n665 & ~n2395 ) | ( n665 & n3986 ) | ( ~n2395 & n3986 ) ;
  assign n3988 = ( n2395 & ~n1653 ) | ( n2395 & n3987 ) | ( ~n1653 & n3987 ) ;
  assign n3989 = n1653 | n3988 ;
  assign n3990 = ( n575 & ~n1072 ) | ( n575 & n3989 ) | ( ~n1072 & n3989 ) ;
  assign n3991 = n1072 | n3990 ;
  assign n3992 = ( n2187 & ~n165 ) | ( n2187 & n3991 ) | ( ~n165 & n3991 ) ;
  assign n3993 = n165 | n3992 ;
  assign n3994 = ( n568 & ~n104 ) | ( n568 & n3993 ) | ( ~n104 & n3993 ) ;
  assign n3995 = n104 | n3994 ;
  assign n3996 = n492 | n3995 ;
  assign n3997 = n187 | n418 ;
  assign n3998 = n237 | n3997 ;
  assign n3999 = n2431 | n3998 ;
  assign n4000 = ( n3984 & n3996 ) | ( n3984 & n3999 ) | ( n3996 & n3999 ) ;
  assign n4001 = ( n3979 & ~n4000 ) | ( n3979 & n3984 ) | ( ~n4000 & n3984 ) ;
  assign n4002 = ~n3979 & n4001 ;
  assign n4003 = ( n244 & n624 ) | ( n244 & n4002 ) | ( n624 & n4002 ) ;
  assign n4004 = ~n244 & n4003 ;
  assign n4005 = ( n349 & ~n676 ) | ( n349 & n4004 ) | ( ~n676 & n4004 ) ;
  assign n4006 = ~n349 & n4005 ;
  assign n4007 = ( n273 & ~n372 ) | ( n273 & n4006 ) | ( ~n372 & n4006 ) ;
  assign n4008 = ~n273 & n4007 ;
  assign n4009 = ( n226 & ~n909 ) | ( n226 & n4008 ) | ( ~n909 & n4008 ) ;
  assign n4010 = ~n226 & n4009 ;
  assign n4011 = ( n74 & ~n88 ) | ( n74 & n4010 ) | ( ~n88 & n4010 ) ;
  assign n4012 = ~n74 & n4011 ;
  assign n4013 = ( n141 & ~n432 ) | ( n141 & n4012 ) | ( ~n432 & n4012 ) ;
  assign n4014 = ~n141 & n4013 ;
  assign n4015 = n105 | n232 ;
  assign n4016 = n167 | n4015 ;
  assign n4017 = ( n3854 & ~n535 ) | ( n3854 & n4016 ) | ( ~n535 & n4016 ) ;
  assign n4018 = n535 | n4017 ;
  assign n4019 = ( n3971 & ~n4014 ) | ( n3971 & n4018 ) | ( ~n4014 & n4018 ) ;
  assign n4020 = ( n3971 & ~n4019 ) | ( n3971 & 1'b0 ) | ( ~n4019 & 1'b0 ) ;
  assign n4021 = ( n842 & ~n886 ) | ( n842 & n4020 ) | ( ~n886 & n4020 ) ;
  assign n4022 = ~n842 & n4021 ;
  assign n4023 = ( n477 & ~n2576 ) | ( n477 & n4022 ) | ( ~n2576 & n4022 ) ;
  assign n4024 = ~n477 & n4023 ;
  assign n4025 = ( n343 & ~n4024 ) | ( n343 & n671 ) | ( ~n4024 & n671 ) ;
  assign n4026 = ( n343 & ~n4025 ) | ( n343 & 1'b0 ) | ( ~n4025 & 1'b0 ) ;
  assign n4027 = ( n281 & ~n631 ) | ( n281 & n4026 ) | ( ~n631 & n4026 ) ;
  assign n4028 = ~n281 & n4027 ;
  assign n4029 = ( n3959 & ~n3846 ) | ( n3959 & n4028 ) | ( ~n3846 & n4028 ) ;
  assign n4030 = ( n3846 & ~x26 ) | ( n3846 & n3907 ) | ( ~x26 & n3907 ) ;
  assign n4031 = ( x26 & ~n3907 ) | ( x26 & n3846 ) | ( ~n3907 & n3846 ) ;
  assign n4032 = ( n4030 & ~n3846 ) | ( n4030 & n4031 ) | ( ~n3846 & n4031 ) ;
  assign n4033 = n946 | n1043 ;
  assign n4034 = n946 &  n1043 ;
  assign n4035 = ( n4033 & ~n4034 ) | ( n4033 & 1'b0 ) | ( ~n4034 & 1'b0 ) ;
  assign n4036 = ~n3632 & n4035 ;
  assign n4037 = ( n3632 & ~n4035 ) | ( n3632 & 1'b0 ) | ( ~n4035 & 1'b0 ) ;
  assign n4038 = n4036 | n4037 ;
  assign n4039 = n3644 | n4038 ;
  assign n4040 = ~n1151 & n3652 ;
  assign n4041 = ~n1043 & n3657 ;
  assign n4042 = n4040 | n4041 ;
  assign n4043 = ~n946 & n3653 ;
  assign n4044 = ( n946 & ~n4042 ) | ( n946 & n4043 ) | ( ~n4042 & n4043 ) ;
  assign n4045 = n4039 &  n4044 ;
  assign n4443 = ( n4029 & ~n4032 ) | ( n4029 & n4045 ) | ( ~n4032 & n4045 ) ;
  assign n4444 = ( n4029 & ~n4045 ) | ( n4029 & n4032 ) | ( ~n4045 & n4032 ) ;
  assign n4445 = ( n4443 & ~n4029 ) | ( n4443 & n4444 ) | ( ~n4029 & n4444 ) ;
  assign n4054 = ( n3846 & ~n3959 ) | ( n3846 & n4028 ) | ( ~n3959 & n4028 ) ;
  assign n4055 = ( n4029 & ~n4028 ) | ( n4029 & n4054 ) | ( ~n4028 & n4054 ) ;
  assign n4056 = ~n1151 & n1267 ;
  assign n4057 = ( n1151 & ~n1267 ) | ( n1151 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n4058 = n4056 | n4057 ;
  assign n4059 = n3630 | n4058 ;
  assign n4060 = n3630 &  n4058 ;
  assign n4061 = ( n4059 & ~n4060 ) | ( n4059 & 1'b0 ) | ( ~n4060 & 1'b0 ) ;
  assign n4062 = ~n3644 & n4061 ;
  assign n4063 = n1151 | n3653 ;
  assign n4064 = ~n1378 & n3652 ;
  assign n4065 = ( n4063 & ~n4064 ) | ( n4063 & 1'b0 ) | ( ~n4064 & 1'b0 ) ;
  assign n4066 = ( n1267 & ~n3657 ) | ( n1267 & 1'b0 ) | ( ~n3657 & 1'b0 ) ;
  assign n4067 = ( n4065 & ~n1267 ) | ( n4065 & n4066 ) | ( ~n1267 & n4066 ) ;
  assign n4068 = ~n4062 & n4067 ;
  assign n4069 = n126 | n195 ;
  assign n4070 = ( n216 & ~n765 ) | ( n216 & n4069 ) | ( ~n765 & n4069 ) ;
  assign n4071 = n765 | n4070 ;
  assign n4072 = ( n221 & ~n451 ) | ( n221 & n4071 ) | ( ~n451 & n4071 ) ;
  assign n4073 = n451 | n4072 ;
  assign n4074 = n167 | n4073 ;
  assign n4115 = n120 | n797 ;
  assign n4116 = ( n572 & ~n228 ) | ( n572 & n4115 ) | ( ~n228 & n4115 ) ;
  assign n4117 = n228 | n4116 ;
  assign n4118 = n225 | n4117 ;
  assign n4119 = n43 | n2309 ;
  assign n4120 = n135 | n4119 ;
  assign n4121 = ( n3229 & ~n1754 ) | ( n3229 & n4120 ) | ( ~n1754 & n4120 ) ;
  assign n4122 = n1754 | n4121 ;
  assign n4123 = ( n4118 & ~n2262 ) | ( n4118 & n4122 ) | ( ~n2262 & n4122 ) ;
  assign n4124 = n2262 | n4123 ;
  assign n4075 = n274 | n647 ;
  assign n4076 = n788 | n1289 ;
  assign n4077 = ( n718 & ~n415 ) | ( n718 & n4076 ) | ( ~n415 & n4076 ) ;
  assign n4078 = n415 | n4077 ;
  assign n4079 = ( n490 & ~n122 ) | ( n490 & n4078 ) | ( ~n122 & n4078 ) ;
  assign n4080 = n122 | n4079 ;
  assign n4081 = ( n424 & ~n205 ) | ( n424 & n4080 ) | ( ~n205 & n4080 ) ;
  assign n4082 = n205 | n4081 ;
  assign n4083 = n664 | n4082 ;
  assign n4084 = ( n193 & n624 ) | ( n193 & n3889 ) | ( n624 & n3889 ) ;
  assign n4085 = ( n624 & ~n4084 ) | ( n624 & 1'b0 ) | ( ~n4084 & 1'b0 ) ;
  assign n4086 = ( n778 & ~n674 ) | ( n778 & n4085 ) | ( ~n674 & n4085 ) ;
  assign n4087 = ~n778 & n4086 ;
  assign n4088 = ( n74 & ~n476 ) | ( n74 & n4087 ) | ( ~n476 & n4087 ) ;
  assign n4089 = ~n74 & n4088 ;
  assign n4090 = ( n484 & ~n744 ) | ( n484 & 1'b0 ) | ( ~n744 & 1'b0 ) ;
  assign n4091 = n1399 | n2378 ;
  assign n4092 = ( n1282 & n4090 ) | ( n1282 & n4091 ) | ( n4090 & n4091 ) ;
  assign n4093 = ( n4090 & ~n4092 ) | ( n4090 & 1'b0 ) | ( ~n4092 & 1'b0 ) ;
  assign n4094 = ( n234 & ~n812 ) | ( n234 & n4093 ) | ( ~n812 & n4093 ) ;
  assign n4095 = ~n234 & n4094 ;
  assign n4096 = ( n475 & ~n714 ) | ( n475 & n4095 ) | ( ~n714 & n4095 ) ;
  assign n4097 = ~n475 & n4096 ;
  assign n4098 = ( n905 & ~n132 ) | ( n905 & n4097 ) | ( ~n132 & n4097 ) ;
  assign n4099 = ~n905 & n4098 ;
  assign n4100 = ( n354 & ~n4099 ) | ( n354 & n406 ) | ( ~n4099 & n406 ) ;
  assign n4101 = ( n354 & ~n4100 ) | ( n354 & 1'b0 ) | ( ~n4100 & 1'b0 ) ;
  assign n4102 = ~n410 & n4101 ;
  assign n4103 = ( n4089 & ~n3417 ) | ( n4089 & n4102 ) | ( ~n3417 & n4102 ) ;
  assign n4104 = n3417 &  n4103 ;
  assign n4105 = ( n1495 & ~n4083 ) | ( n1495 & n4104 ) | ( ~n4083 & n4104 ) ;
  assign n4106 = ~n1495 & n4105 ;
  assign n4107 = ( n4075 & ~n268 ) | ( n4075 & n4106 ) | ( ~n268 & n4106 ) ;
  assign n4108 = ( n813 & ~n4107 ) | ( n813 & n4075 ) | ( ~n4107 & n4075 ) ;
  assign n4109 = ( n813 & ~n4108 ) | ( n813 & 1'b0 ) | ( ~n4108 & 1'b0 ) ;
  assign n4110 = ( n554 & ~n89 ) | ( n554 & n4109 ) | ( ~n89 & n4109 ) ;
  assign n4111 = ~n554 & n4110 ;
  assign n4112 = ( n129 & ~n49 ) | ( n129 & n4111 ) | ( ~n49 & n4111 ) ;
  assign n4113 = ~n129 & n4112 ;
  assign n4114 = ~n666 & n4113 ;
  assign n4125 = ( n4074 & ~n4124 ) | ( n4074 & n4114 ) | ( ~n4124 & n4114 ) ;
  assign n4126 = ( n2840 & ~n4074 ) | ( n2840 & n4125 ) | ( ~n4074 & n4125 ) ;
  assign n4127 = ~n2840 & n4126 ;
  assign n4128 = ( n163 & ~n238 ) | ( n163 & n4127 ) | ( ~n238 & n4127 ) ;
  assign n4129 = ~n163 & n4128 ;
  assign n4130 = ( n493 & ~n194 ) | ( n493 & n4129 ) | ( ~n194 & n4129 ) ;
  assign n4131 = ~n493 & n4130 ;
  assign n4132 = ( n761 & n786 ) | ( n761 & n4131 ) | ( n786 & n4131 ) ;
  assign n4133 = ~n761 & n4132 ;
  assign n4134 = ( n165 & ~n281 ) | ( n165 & n4133 ) | ( ~n281 & n4133 ) ;
  assign n4135 = ~n165 & n4134 ;
  assign n4136 = n413 | n1428 ;
  assign n4137 = ( n431 & ~n124 ) | ( n431 & n4136 ) | ( ~n124 & n4136 ) ;
  assign n4138 = n124 | n4137 ;
  assign n4139 = n233 | n1454 ;
  assign n4140 = ( n424 & ~n190 ) | ( n424 & n4139 ) | ( ~n190 & n4139 ) ;
  assign n4141 = n190 | n4140 ;
  assign n4142 = ( n3370 & ~n4138 ) | ( n3370 & n4141 ) | ( ~n4138 & n4141 ) ;
  assign n4143 = ( n4138 & ~n668 ) | ( n4138 & n4142 ) | ( ~n668 & n4142 ) ;
  assign n4144 = n668 | n4143 ;
  assign n4145 = ( n475 & ~n273 ) | ( n475 & n4144 ) | ( ~n273 & n4144 ) ;
  assign n4146 = n273 | n4145 ;
  assign n4147 = n160 | n4146 ;
  assign n4148 = n104 | n276 ;
  assign n4149 = ( n478 & ~n225 ) | ( n478 & n4148 ) | ( ~n225 & n4148 ) ;
  assign n4150 = n225 | n4149 ;
  assign n4151 = n526 | n778 ;
  assign n4152 = n212 | n4151 ;
  assign n4153 = ( n3802 & ~n4152 ) | ( n3802 & 1'b0 ) | ( ~n4152 & 1'b0 ) ;
  assign n4154 = ( n1600 & ~n1809 ) | ( n1600 & n4153 ) | ( ~n1809 & n4153 ) ;
  assign n4155 = ~n1600 & n4154 ;
  assign n4156 = ( n128 & ~n4150 ) | ( n128 & n4155 ) | ( ~n4150 & n4155 ) ;
  assign n4157 = ~n128 & n4156 ;
  assign n4158 = ( n1060 & ~n1195 ) | ( n1060 & n4157 ) | ( ~n1195 & n4157 ) ;
  assign n4159 = ~n1060 & n4158 ;
  assign n4160 = ( n885 & ~n495 ) | ( n885 & n4159 ) | ( ~n495 & n4159 ) ;
  assign n4161 = ~n885 & n4160 ;
  assign n4162 = ( n49 & ~n531 ) | ( n49 & n4161 ) | ( ~n531 & n4161 ) ;
  assign n4163 = ~n49 & n4162 ;
  assign n4164 = ( n239 & ~n240 ) | ( n239 & n4163 ) | ( ~n240 & n4163 ) ;
  assign n4165 = ~n239 & n4164 ;
  assign n4166 = ~n336 & n4165 ;
  assign n4174 = n374 | n417 ;
  assign n4175 = ( n410 & ~n117 ) | ( n410 & n4174 ) | ( ~n117 & n4174 ) ;
  assign n4176 = n117 | n4175 ;
  assign n4198 = n1497 | n1753 ;
  assign n4177 = n620 | n2034 ;
  assign n4178 = ( n217 & ~n376 ) | ( n217 & n4177 ) | ( ~n376 & n4177 ) ;
  assign n4179 = n376 | n4178 ;
  assign n4180 = ( n187 & ~n284 ) | ( n187 & n4179 ) | ( ~n284 & n4179 ) ;
  assign n4181 = n284 | n4180 ;
  assign n4182 = ( n2548 & ~n4181 ) | ( n2548 & n3878 ) | ( ~n4181 & n3878 ) ;
  assign n4183 = ( n4182 & ~n2411 ) | ( n4182 & n4181 ) | ( ~n2411 & n4181 ) ;
  assign n4184 = n4183 | n2411 ;
  assign n4185 = ( n1433 & ~n1828 ) | ( n1433 & n4184 ) | ( ~n1828 & n4184 ) ;
  assign n4186 = n1828 | n4185 ;
  assign n4187 = ( n2192 & ~n1807 ) | ( n2192 & n4186 ) | ( ~n1807 & n4186 ) ;
  assign n4188 = n1807 | n4187 ;
  assign n4189 = ( n2784 & ~n461 ) | ( n2784 & n4188 ) | ( ~n461 & n4188 ) ;
  assign n4190 = n461 | n4189 ;
  assign n4191 = ( n194 & ~n362 ) | ( n194 & n4190 ) | ( ~n362 & n4190 ) ;
  assign n4192 = n362 | n4191 ;
  assign n4193 = ( n672 & ~n230 ) | ( n672 & n4192 ) | ( ~n230 & n4192 ) ;
  assign n4194 = n230 | n4193 ;
  assign n4195 = ( n99 & ~n411 ) | ( n99 & n4194 ) | ( ~n411 & n4194 ) ;
  assign n4196 = n411 | n4195 ;
  assign n4197 = n664 | n4196 ;
  assign n4199 = ( n4198 & ~n4176 ) | ( n4198 & n4197 ) | ( ~n4176 & n4197 ) ;
  assign n4200 = ( n4176 & ~n2108 ) | ( n4176 & n4199 ) | ( ~n2108 & n4199 ) ;
  assign n4201 = n2108 | n4200 ;
  assign n4167 = ( n223 & ~n61 ) | ( n223 & n2462 ) | ( ~n61 & n2462 ) ;
  assign n4168 = n61 | n4167 ;
  assign n4169 = ( n792 & ~n243 ) | ( n792 & n4168 ) | ( ~n243 & n4168 ) ;
  assign n4170 = n243 | n4169 ;
  assign n4171 = ( n80 & ~n149 ) | ( n80 & n4170 ) | ( ~n149 & n4170 ) ;
  assign n4172 = n149 | n4171 ;
  assign n4173 = n141 | n4172 ;
  assign n4202 = ( n4166 & n4201 ) | ( n4166 & n4173 ) | ( n4201 & n4173 ) ;
  assign n4203 = ( n4166 & ~n4202 ) | ( n4166 & 1'b0 ) | ( ~n4202 & 1'b0 ) ;
  assign n4204 = ( n414 & ~n4147 ) | ( n414 & n4203 ) | ( ~n4147 & n4203 ) ;
  assign n4205 = ~n414 & n4204 ;
  assign n4206 = ( n234 & ~n260 ) | ( n234 & n4205 ) | ( ~n260 & n4205 ) ;
  assign n4207 = ~n234 & n4206 ;
  assign n4208 = ( n722 & ~n490 ) | ( n722 & n4207 ) | ( ~n490 & n4207 ) ;
  assign n4209 = ~n722 & n4208 ;
  assign n4210 = ( n905 & ~n630 ) | ( n905 & n4209 ) | ( ~n630 & n4209 ) ;
  assign n4211 = ~n905 & n4210 ;
  assign n4212 = ( n140 & ~n476 ) | ( n140 & n4211 ) | ( ~n476 & n4211 ) ;
  assign n4213 = ~n140 & n4212 ;
  assign n4214 = ~n432 & n4213 ;
  assign n4215 = ( x23 & n4135 ) | ( x23 & n4214 ) | ( n4135 & n4214 ) ;
  assign n4216 = ( n4068 & ~n3846 ) | ( n4068 & n4215 ) | ( ~n3846 & n4215 ) ;
  assign n4217 = ( n3846 & ~n4215 ) | ( n3846 & n4068 ) | ( ~n4215 & n4068 ) ;
  assign n4218 = ( n3846 & ~n4068 ) | ( n3846 & n4215 ) | ( ~n4068 & n4215 ) ;
  assign n4219 = ( n4217 & ~n3846 ) | ( n4217 & n4218 ) | ( ~n3846 & n4218 ) ;
  assign n3939 = ~n515 |  n521 ;
  assign n4434 = ~n946 & n3939 ;
  assign n4430 = ~n521 |  n518 ;
  assign n4431 = n863 | n4430 ;
  assign n4432 = n523 | n1043 ;
  assign n4433 = n4431 &  n4432 ;
  assign n4435 = ( n946 & n4434 ) | ( n946 & n4433 ) | ( n4434 & n4433 ) ;
  assign n4436 = ( n3914 & ~n601 ) | ( n3914 & n4435 ) | ( ~n601 & n4435 ) ;
  assign n4437 = ~n3914 & n4436 ;
  assign n4438 = ( x29 & ~n4435 ) | ( x29 & n4437 ) | ( ~n4435 & n4437 ) ;
  assign n4439 = ( n4435 & ~x29 ) | ( n4435 & n4437 ) | ( ~x29 & n4437 ) ;
  assign n4440 = ( n4438 & ~n4437 ) | ( n4438 & n4439 ) | ( ~n4437 & n4439 ) ;
  assign n4220 = n765 | n3481 ;
  assign n4221 = ( n905 & ~n734 ) | ( n905 & n4220 ) | ( ~n734 & n4220 ) ;
  assign n4222 = n734 | n4221 ;
  assign n4223 = ( n554 & ~n205 ) | ( n554 & n4222 ) | ( ~n205 & n4222 ) ;
  assign n4224 = n205 | n4223 ;
  assign n4225 = ( n618 & ~n643 ) | ( n618 & n4224 ) | ( ~n643 & n4224 ) ;
  assign n4226 = n643 | n4225 ;
  assign n4227 = n433 | n490 ;
  assign n4228 = n123 | n244 ;
  assign n4229 = n222 | n679 ;
  assign n4230 = ( n343 & ~n4229 ) | ( n343 & 1'b0 ) | ( ~n4229 & 1'b0 ) ;
  assign n4231 = ( n4227 & ~n4228 ) | ( n4227 & n4230 ) | ( ~n4228 & n4230 ) ;
  assign n4232 = ~n4227 & n4231 ;
  assign n4233 = ( n889 & ~n998 ) | ( n889 & n4232 ) | ( ~n998 & n4232 ) ;
  assign n4234 = ( n2666 & ~n889 ) | ( n2666 & n4233 ) | ( ~n889 & n4233 ) ;
  assign n4235 = ~n2666 & n4234 ;
  assign n4236 = ( n4235 & ~n620 ) | ( n4235 & n4226 ) | ( ~n620 & n4226 ) ;
  assign n4237 = ( n1511 & ~n4226 ) | ( n1511 & n4236 ) | ( ~n4226 & n4236 ) ;
  assign n4238 = ~n1511 & n4237 ;
  assign n4239 = ( n788 & ~n948 ) | ( n788 & n4238 ) | ( ~n948 & n4238 ) ;
  assign n4240 = ~n788 & n4239 ;
  assign n4241 = ( n4240 & ~n235 ) | ( n4240 & n569 ) | ( ~n235 & n569 ) ;
  assign n4242 = ( n4241 & ~n569 ) | ( n4241 & 1'b0 ) | ( ~n569 & 1'b0 ) ;
  assign n4243 = n258 | n797 ;
  assign n4244 = n494 | n4243 ;
  assign n4245 = ( n69 & ~n362 ) | ( n69 & n4244 ) | ( ~n362 & n4244 ) ;
  assign n4246 = n362 | n4245 ;
  assign n4247 = ( n404 & n623 ) | ( n404 & n4246 ) | ( n623 & n4246 ) ;
  assign n4248 = ( n623 & ~n4247 ) | ( n623 & 1'b0 ) | ( ~n4247 & 1'b0 ) ;
  assign n4249 = ( n276 & ~n135 ) | ( n276 & n4248 ) | ( ~n135 & n4248 ) ;
  assign n4250 = ~n276 & n4249 ;
  assign n4251 = n127 | n887 ;
  assign n4252 = ( n351 & ~n280 ) | ( n351 & n4251 ) | ( ~n280 & n4251 ) ;
  assign n4253 = n280 | n4252 ;
  assign n4254 = ( n1547 & ~n1657 ) | ( n1547 & 1'b0 ) | ( ~n1657 & 1'b0 ) ;
  assign n4255 = ( n4253 & ~n2358 ) | ( n4253 & n4254 ) | ( ~n2358 & n4254 ) ;
  assign n4256 = ( n1617 & ~n4253 ) | ( n1617 & n4255 ) | ( ~n4253 & n4255 ) ;
  assign n4257 = ~n1617 & n4256 ;
  assign n4258 = n1917 &  n4257 ;
  assign n4259 = ( n1360 & ~n4258 ) | ( n1360 & n4250 ) | ( ~n4258 & n4250 ) ;
  assign n4260 = ( n3129 & ~n4250 ) | ( n3129 & n4259 ) | ( ~n4250 & n4259 ) ;
  assign n4261 = ( n3129 & ~n4260 ) | ( n3129 & 1'b0 ) | ( ~n4260 & 1'b0 ) ;
  assign n4262 = ( n416 & n4242 ) | ( n416 & n4261 ) | ( n4242 & n4261 ) ;
  assign n4263 = ~n416 & n4262 ;
  assign n4264 = ( n674 & ~n345 ) | ( n674 & n4263 ) | ( ~n345 & n4263 ) ;
  assign n4265 = ~n674 & n4264 ;
  assign n4266 = ( n217 & ~n793 ) | ( n217 & n4265 ) | ( ~n793 & n4265 ) ;
  assign n4267 = ~n217 & n4266 ;
  assign n4268 = ~n560 & n4267 ;
  assign n4291 = n1618 | n4244 ;
  assign n4282 = ( n1279 & n3665 ) | ( n1279 & n1754 ) | ( n3665 & n1754 ) ;
  assign n4283 = ( n1279 & ~n4282 ) | ( n1279 & 1'b0 ) | ( ~n4282 & 1'b0 ) ;
  assign n4284 = ( n280 & ~n127 ) | ( n280 & n4283 ) | ( ~n127 & n4283 ) ;
  assign n4285 = ~n280 & n4284 ;
  assign n4286 = ( n4285 & ~n602 ) | ( n4285 & n737 ) | ( ~n602 & n737 ) ;
  assign n4287 = ( n4286 & ~n737 ) | ( n4286 & 1'b0 ) | ( ~n737 & 1'b0 ) ;
  assign n4288 = ( n417 & ~n540 ) | ( n417 & n4287 ) | ( ~n540 & n4287 ) ;
  assign n4289 = ~n417 & n4288 ;
  assign n4290 = ~n166 & n4289 ;
  assign n4292 = ( n866 & ~n4291 ) | ( n866 & n4290 ) | ( ~n4291 & n4290 ) ;
  assign n4293 = ~n866 & n4292 ;
  assign n4294 = ( n2702 & ~n654 ) | ( n2702 & n4293 ) | ( ~n654 & n4293 ) ;
  assign n4295 = ~n2702 & n4294 ;
  assign n4296 = ( n813 & ~n4295 ) | ( n813 & n2757 ) | ( ~n4295 & n2757 ) ;
  assign n4297 = ( n813 & ~n4296 ) | ( n813 & 1'b0 ) | ( ~n4296 & 1'b0 ) ;
  assign n4298 = ( n761 & ~n168 ) | ( n761 & n4297 ) | ( ~n168 & n4297 ) ;
  assign n4299 = ~n761 & n4298 ;
  assign n4300 = ( n453 & ~n226 ) | ( n453 & n4299 ) | ( ~n226 & n4299 ) ;
  assign n4301 = ~n453 & n4300 ;
  assign n4302 = ( n4301 & ~n91 ) | ( n4301 & n454 ) | ( ~n91 & n454 ) ;
  assign n4303 = ( n4302 & ~n454 ) | ( n4302 & 1'b0 ) | ( ~n454 & 1'b0 ) ;
  assign n4304 = ~n646 & n4303 ;
  assign n4323 = ( n791 & ~n1585 ) | ( n791 & n1885 ) | ( ~n1585 & n1885 ) ;
  assign n4324 = n1585 | n4323 ;
  assign n4325 = ( n463 & ~n385 ) | ( n463 & n4324 ) | ( ~n385 & n4324 ) ;
  assign n4326 = n385 | n4325 ;
  assign n4327 = ( n2403 & ~n2081 ) | ( n2403 & n4326 ) | ( ~n2081 & n4326 ) ;
  assign n4328 = n2081 | n4327 ;
  assign n4305 = n106 | n363 ;
  assign n4306 = ( n679 & ~n678 ) | ( n679 & n4305 ) | ( ~n678 & n4305 ) ;
  assign n4307 = n678 | n4306 ;
  assign n4308 = ( n221 & n484 ) | ( n221 & n4307 ) | ( n484 & n4307 ) ;
  assign n4309 = ( n484 & ~n4308 ) | ( n484 & 1'b0 ) | ( ~n4308 & 1'b0 ) ;
  assign n4310 = n765 | n3158 ;
  assign n4311 = ( n2266 & ~n1004 ) | ( n2266 & n4310 ) | ( ~n1004 & n4310 ) ;
  assign n4312 = ( n1071 & ~n4310 ) | ( n1071 & n4311 ) | ( ~n4310 & n4311 ) ;
  assign n4313 = ~n1071 & n4312 ;
  assign n4314 = ( n1045 & n4309 ) | ( n1045 & n4313 ) | ( n4309 & n4313 ) ;
  assign n4315 = ~n1045 & n4314 ;
  assign n4316 = ( n2666 & ~n3568 ) | ( n2666 & n4315 ) | ( ~n3568 & n4315 ) ;
  assign n4317 = ~n2666 & n4316 ;
  assign n4318 = ( n716 & ~n238 ) | ( n716 & n4317 ) | ( ~n238 & n4317 ) ;
  assign n4319 = ~n716 & n4318 ;
  assign n4320 = ( n72 & ~n4319 ) | ( n72 & n343 ) | ( ~n4319 & n343 ) ;
  assign n4321 = ( n343 & ~n4320 ) | ( n343 & 1'b0 ) | ( ~n4320 & 1'b0 ) ;
  assign n4322 = ~n93 & n4321 ;
  assign n4329 = ( n1627 & ~n4328 ) | ( n1627 & n4322 ) | ( ~n4328 & n4322 ) ;
  assign n4330 = ~n1627 & n4329 ;
  assign n4331 = ( n2784 & n4304 ) | ( n2784 & n4330 ) | ( n4304 & n4330 ) ;
  assign n4332 = ~n2784 & n4331 ;
  assign n4333 = ( n335 & ~n70 ) | ( n335 & n4332 ) | ( ~n70 & n4332 ) ;
  assign n4334 = ~n335 & n4333 ;
  assign n4335 = ( n216 & ~n260 ) | ( n216 & n4334 ) | ( ~n260 & n4334 ) ;
  assign n4336 = ~n216 & n4335 ;
  assign n4337 = ( n187 & ~n549 ) | ( n187 & n4336 ) | ( ~n549 & n4336 ) ;
  assign n4338 = ~n187 & n4337 ;
  assign n4339 = ( n160 & ~n141 ) | ( n160 & n4338 ) | ( ~n141 & n4338 ) ;
  assign n4340 = ~n160 & n4339 ;
  assign n4341 = n137 | n910 ;
  assign n4342 = n135 | n4341 ;
  assign n4343 = ( n414 & ~n225 ) | ( n414 & n631 ) | ( ~n225 & n631 ) ;
  assign n4344 = n225 | n4343 ;
  assign n4345 = ( n254 & ~n4342 ) | ( n254 & n4344 ) | ( ~n4342 & n4344 ) ;
  assign n4346 = ( n4342 & ~n3159 ) | ( n4342 & n4345 ) | ( ~n3159 & n4345 ) ;
  assign n4347 = n3159 | n4346 ;
  assign n4348 = ( n887 & ~n530 ) | ( n887 & n4347 ) | ( ~n530 & n4347 ) ;
  assign n4349 = n530 | n4348 ;
  assign n4350 = ( n2091 & ~n2029 ) | ( n2091 & n4349 ) | ( ~n2029 & n4349 ) ;
  assign n4351 = n2029 | n4350 ;
  assign n4352 = ( n339 & ~n381 ) | ( n339 & n4351 ) | ( ~n381 & n4351 ) ;
  assign n4353 = ( n381 & ~n416 ) | ( n381 & n4352 ) | ( ~n416 & n4352 ) ;
  assign n4354 = n416 | n4353 ;
  assign n4355 = ( n335 & n4354 ) | ( n335 & n813 ) | ( n4354 & n813 ) ;
  assign n4356 = ( n813 & ~n4355 ) | ( n813 & 1'b0 ) | ( ~n4355 & 1'b0 ) ;
  assign n4357 = ( n676 & ~n490 ) | ( n676 & n4356 ) | ( ~n490 & n4356 ) ;
  assign n4358 = ~n676 & n4357 ;
  assign n4359 = ~n191 & n4358 ;
  assign n4360 = n974 | n1626 ;
  assign n4361 = ( n61 & ~n4360 ) | ( n61 & n525 ) | ( ~n4360 & n525 ) ;
  assign n4362 = ~n61 & n4361 ;
  assign n4363 = ( n217 & ~n406 ) | ( n217 & n4362 ) | ( ~n406 & n4362 ) ;
  assign n4364 = ~n217 & n4363 ;
  assign n4365 = ( n160 & ~n118 ) | ( n160 & n4364 ) | ( ~n118 & n4364 ) ;
  assign n4366 = ~n160 & n4365 ;
  assign n4367 = ( n236 & ~n627 ) | ( n236 & n4366 ) | ( ~n627 & n4366 ) ;
  assign n4368 = ~n236 & n4367 ;
  assign n4369 = ( n670 & ~n285 ) | ( n670 & n4368 ) | ( ~n285 & n4368 ) ;
  assign n4370 = ~n670 & n4369 ;
  assign n4371 = n425 | n1625 ;
  assign n4372 = n150 | n362 ;
  assign n4373 = n245 | n4372 ;
  assign n4374 = ( n1437 & n4371 ) | ( n1437 & n4373 ) | ( n4371 & n4373 ) ;
  assign n4375 = ( n1437 & ~n4374 ) | ( n1437 & 1'b0 ) | ( ~n4374 & 1'b0 ) ;
  assign n4376 = ( n1427 & ~n4375 ) | ( n1427 & n4370 ) | ( ~n4375 & n4370 ) ;
  assign n4377 = ( n2467 & ~n4370 ) | ( n2467 & n4376 ) | ( ~n4370 & n4376 ) ;
  assign n4378 = ( n2467 & ~n4377 ) | ( n2467 & 1'b0 ) | ( ~n4377 & 1'b0 ) ;
  assign n4379 = ( n1762 & ~n2191 ) | ( n1762 & n4378 ) | ( ~n2191 & n4378 ) ;
  assign n4380 = ~n1762 & n4379 ;
  assign n4381 = ( n775 & ~n721 ) | ( n775 & n4380 ) | ( ~n721 & n4380 ) ;
  assign n4382 = ~n775 & n4381 ;
  assign n4383 = ( n151 & ~n417 ) | ( n151 & n4382 ) | ( ~n417 & n4382 ) ;
  assign n4384 = ~n151 & n4383 ;
  assign n4385 = ( n259 & ~n157 ) | ( n259 & n430 ) | ( ~n157 & n430 ) ;
  assign n4386 = n157 | n4385 ;
  assign n4387 = ( n258 & ~n712 ) | ( n258 & n4386 ) | ( ~n712 & n4386 ) ;
  assign n4388 = n712 | n4387 ;
  assign n4389 = ( n52 & ~n231 ) | ( n52 & n4388 ) | ( ~n231 & n4388 ) ;
  assign n4390 = n231 | n4389 ;
  assign n4391 = ( n485 & ~n456 ) | ( n485 & n4390 ) | ( ~n456 & n4390 ) ;
  assign n4392 = n456 | n4391 ;
  assign n4393 = ( n4392 & ~n161 ) | ( n4392 & n266 ) | ( ~n161 & n266 ) ;
  assign n4394 = n161 | n4393 ;
  assign n4395 = ( n603 & ~n129 ) | ( n603 & n4394 ) | ( ~n129 & n4394 ) ;
  assign n4396 = n129 | n4395 ;
  assign n4397 = n433 | n4396 ;
  assign n4398 = ( n1129 & n4397 ) | ( n1129 & n1289 ) | ( n4397 & n1289 ) ;
  assign n4399 = ( n3144 & ~n4398 ) | ( n3144 & n1129 ) | ( ~n4398 & n1129 ) ;
  assign n4400 = ( n4399 & ~n3144 ) | ( n4399 & 1'b0 ) | ( ~n3144 & 1'b0 ) ;
  assign n4401 = ( n4384 & ~n4359 ) | ( n4384 & n4400 ) | ( ~n4359 & n4400 ) ;
  assign n4402 = n4359 &  n4401 ;
  assign n4403 = ( n1484 & ~n115 ) | ( n1484 & n4402 ) | ( ~n115 & n4402 ) ;
  assign n4404 = ~n1484 & n4403 ;
  assign n4405 = ( n1678 & ~n1185 ) | ( n1678 & n4404 ) | ( ~n1185 & n4404 ) ;
  assign n4406 = ~n1678 & n4405 ;
  assign n4407 = ( n166 & ~n679 ) | ( n166 & n4406 ) | ( ~n679 & n4406 ) ;
  assign n4408 = ~n166 & n4407 ;
  assign n4409 = ( n617 & ~n347 ) | ( n617 & n4408 ) | ( ~n347 & n4408 ) ;
  assign n4410 = ~n617 & n4409 ;
  assign n4411 = ( x20 & n4340 ) | ( x20 & n4410 ) | ( n4340 & n4410 ) ;
  assign n4270 = n1483 &  n1566 ;
  assign n4269 = ( n1483 & ~n1566 ) | ( n1483 & 1'b0 ) | ( ~n1566 & 1'b0 ) ;
  assign n4271 = ( n1566 & ~n4270 ) | ( n1566 & n4269 ) | ( ~n4270 & n4269 ) ;
  assign n4272 = n3627 | n4271 ;
  assign n4273 = n3627 &  n4271 ;
  assign n4274 = ( n4272 & ~n4273 ) | ( n4272 & 1'b0 ) | ( ~n4273 & 1'b0 ) ;
  assign n4280 = n4274 | n3644 ;
  assign n4275 = ( n1483 & ~n3653 ) | ( n1483 & 1'b0 ) | ( ~n3653 & 1'b0 ) ;
  assign n4276 = ~n1671 & n3652 ;
  assign n4277 = ~n1566 & n3657 ;
  assign n4278 = n4276 | n4277 ;
  assign n4279 = n4275 | n4278 ;
  assign n4281 = ( n4280 & ~n3644 ) | ( n4280 & n4279 ) | ( ~n3644 & n4279 ) ;
  assign n4412 = ( n4268 & ~n4411 ) | ( n4268 & n4281 ) | ( ~n4411 & n4281 ) ;
  assign n4413 = ( n4135 & ~n4268 ) | ( n4135 & n4412 ) | ( ~n4268 & n4412 ) ;
  assign n4414 = ( x23 & ~n4135 ) | ( x23 & n4214 ) | ( ~n4135 & n4214 ) ;
  assign n4415 = ( n4135 & ~n4215 ) | ( n4135 & n4414 ) | ( ~n4215 & n4414 ) ;
  assign n4417 = ( n1267 & ~n1378 ) | ( n1267 & 1'b0 ) | ( ~n1378 & 1'b0 ) ;
  assign n4418 = ~n1267 & n1378 ;
  assign n4419 = n4417 | n4418 ;
  assign n4420 = n3629 | n4419 ;
  assign n4421 = n3629 &  n4419 ;
  assign n4422 = ( n4420 & ~n4421 ) | ( n4420 & 1'b0 ) | ( ~n4421 & 1'b0 ) ;
  assign n4427 = n4422 | n3644 ;
  assign n4425 = ( n1483 & ~n3652 ) | ( n1483 & 1'b0 ) | ( ~n3652 & 1'b0 ) ;
  assign n4416 = ( n1267 & ~n3653 ) | ( n1267 & 1'b0 ) | ( ~n3653 & 1'b0 ) ;
  assign n4423 = ~n1378 & n3657 ;
  assign n4424 = n4416 | n4423 ;
  assign n4426 = ( n1483 & ~n4425 ) | ( n1483 & n4424 ) | ( ~n4425 & n4424 ) ;
  assign n4428 = ( n4427 & ~n3644 ) | ( n4427 & n4426 ) | ( ~n3644 & n4426 ) ;
  assign n4429 = ( n4413 & ~n4415 ) | ( n4413 & n4428 ) | ( ~n4415 & n4428 ) ;
  assign n4441 = ( n4219 & ~n4440 ) | ( n4219 & n4429 ) | ( ~n4440 & n4429 ) ;
  assign n4442 = ( n4055 & ~n4216 ) | ( n4055 & n4441 ) | ( ~n4216 & n4441 ) ;
  assign n4449 = ~n523 & n863 ;
  assign n4446 = n599 | n4430 ;
  assign n4447 = n702 | n3939 ;
  assign n4448 = n4446 &  n4447 ;
  assign n4450 = ( n523 & n4449 ) | ( n523 & n4448 ) | ( n4449 & n4448 ) ;
  assign n3932 = n599 | n702 ;
  assign n3933 = ~n599 & n702 ;
  assign n3934 = ( n3932 & ~n702 ) | ( n3932 & n3933 ) | ( ~n702 & n3933 ) ;
  assign n3935 = ~n3635 & n3934 ;
  assign n4451 = ( n3635 & ~n3934 ) | ( n3635 & 1'b0 ) | ( ~n3934 & 1'b0 ) ;
  assign n4452 = n3935 | n4451 ;
  assign n4453 = n601 | n4452 ;
  assign n4454 = n4450 &  n4453 ;
  assign n4455 = x29 &  n4454 ;
  assign n4456 = x29 | n4454 ;
  assign n4457 = ~n4455 & n4456 ;
  assign n4458 = ( n4445 & ~n4442 ) | ( n4445 & n4457 ) | ( ~n4442 & n4457 ) ;
  assign n3936 = n3935 &  n599 ;
  assign n3937 = ( n3936 & ~n599 ) | ( n3936 & n3637 ) | ( ~n599 & n3637 ) ;
  assign n3942 = n3937 | n601 ;
  assign n3938 = n523 | n702 ;
  assign n3940 = n599 | n3939 ;
  assign n3941 = n3938 &  n3940 ;
  assign n3943 = ( n601 & ~n3942 ) | ( n601 & n3941 ) | ( ~n3942 & n3941 ) ;
  assign n4046 = ( n4029 & n4032 ) | ( n4029 & n4045 ) | ( n4032 & n4045 ) ;
  assign n3929 = ( n3727 & ~n3908 ) | ( n3727 & n3921 ) | ( ~n3908 & n3921 ) ;
  assign n3930 = ( n3727 & ~n3921 ) | ( n3727 & n3908 ) | ( ~n3921 & n3908 ) ;
  assign n3931 = ( n3929 & ~n3727 ) | ( n3929 & n3930 ) | ( ~n3727 & n3930 ) ;
  assign n4048 = ~x29 & n3931 ;
  assign n4049 = x29 | n3931 ;
  assign n4050 = ( n4048 & ~n3931 ) | ( n4048 & n4049 ) | ( ~n3931 & n4049 ) ;
  assign n4051 = ( n3943 & ~n4046 ) | ( n3943 & n4050 ) | ( ~n4046 & n4050 ) ;
  assign n4052 = ( n4046 & ~n3943 ) | ( n4046 & n4050 ) | ( ~n3943 & n4050 ) ;
  assign n4053 = ( n4051 & ~n4050 ) | ( n4051 & n4052 ) | ( ~n4050 & n4052 ) ;
  assign n4465 = ~n523 & n946 ;
  assign n4462 = n702 | n4430 ;
  assign n4463 = n863 | n3939 ;
  assign n4464 = n4462 &  n4463 ;
  assign n4466 = ( n523 & n4465 ) | ( n523 & n4464 ) | ( n4465 & n4464 ) ;
  assign n4467 = n601 | n3650 ;
  assign n4468 = n4466 &  n4467 ;
  assign n4469 = x29 &  n4468 ;
  assign n4470 = x29 | n4468 ;
  assign n4471 = ~n4469 & n4470 ;
  assign n4472 = ( x23 & ~x24 ) | ( x23 & 1'b0 ) | ( ~x24 & 1'b0 ) ;
  assign n4473 = ~x23 & x24 ;
  assign n4474 = n4472 | n4473 ;
  assign n4475 = ( x25 & ~x26 ) | ( x25 & 1'b0 ) | ( ~x26 & 1'b0 ) ;
  assign n4476 = ~x25 & x26 ;
  assign n4477 = n4475 | n4476 ;
  assign n4478 = ~n4474 | ~n4477 ;
  assign n4479 = n3637 | n4478 ;
  assign n4481 = ~n4474 & n4477 ;
  assign n4480 = ~n34 & n78 ;
  assign n4482 = ~n4481 |  n4480 ;
  assign n4483 = n599 | n4482 ;
  assign n4484 = n4479 &  n4483 ;
  assign n4485 = ~x26 & n4484 ;
  assign n4486 = ( x26 & ~n4484 ) | ( x26 & 1'b0 ) | ( ~n4484 & 1'b0 ) ;
  assign n4487 = n4485 | n4486 ;
  assign n4488 = ( n4055 & ~n4441 ) | ( n4055 & n4216 ) | ( ~n4441 & n4216 ) ;
  assign n4489 = ( n4216 & ~n4055 ) | ( n4216 & n4441 ) | ( ~n4055 & n4441 ) ;
  assign n4490 = ( n4488 & ~n4216 ) | ( n4488 & n4489 ) | ( ~n4216 & n4489 ) ;
  assign n4491 = ( n4471 & n4487 ) | ( n4471 & n4490 ) | ( n4487 & n4490 ) ;
  assign n4459 = ( n4442 & n4445 ) | ( n4442 & n4457 ) | ( n4445 & n4457 ) ;
  assign n4460 = ( n4442 & ~n4445 ) | ( n4442 & n4457 ) | ( ~n4445 & n4457 ) ;
  assign n4461 = ( n4445 & ~n4459 ) | ( n4445 & n4460 ) | ( ~n4459 & n4460 ) ;
  assign n4492 = ( n4471 & ~n4487 ) | ( n4471 & n4490 ) | ( ~n4487 & n4490 ) ;
  assign n4493 = ( n4487 & ~n4491 ) | ( n4487 & n4492 ) | ( ~n4491 & n4492 ) ;
  assign n4494 = n702 | n4482 ;
  assign n4495 = ~n4480 |  n4474 ;
  assign n4496 = n599 | n4495 ;
  assign n4497 = n4494 &  n4496 ;
  assign n4498 = n3937 &  n4478 ;
  assign n4499 = ( n4497 & ~n3937 ) | ( n4497 & n4498 ) | ( ~n3937 & n4498 ) ;
  assign n4500 = x26 | n4499 ;
  assign n4501 = ( x26 & ~n4499 ) | ( x26 & 1'b0 ) | ( ~n4499 & 1'b0 ) ;
  assign n4502 = ( n4500 & ~x26 ) | ( n4500 & n4501 ) | ( ~x26 & n4501 ) ;
  assign n4503 = ( n4413 & ~n4428 ) | ( n4413 & n4415 ) | ( ~n4428 & n4415 ) ;
  assign n4504 = ( n4415 & ~n4413 ) | ( n4415 & n4428 ) | ( ~n4413 & n4428 ) ;
  assign n4505 = ( n4503 & ~n4415 ) | ( n4503 & n4504 ) | ( ~n4415 & n4504 ) ;
  assign n4506 = n127 | n193 ;
  assign n4507 = ( n253 & ~n105 ) | ( n253 & n4506 ) | ( ~n105 & n4506 ) ;
  assign n4508 = n105 | n4507 ;
  assign n4509 = ( n123 & ~n714 ) | ( n123 & n4508 ) | ( ~n714 & n4508 ) ;
  assign n4510 = n714 | n4509 ;
  assign n4511 = ( n911 & ~n628 ) | ( n911 & n4510 ) | ( ~n628 & n4510 ) ;
  assign n4512 = n628 | n4511 ;
  assign n4513 = n670 | n4512 ;
  assign n4514 = ( n645 & ~n800 ) | ( n645 & 1'b0 ) | ( ~n800 & 1'b0 ) ;
  assign n4515 = ( n348 & ~n540 ) | ( n348 & n4514 ) | ( ~n540 & n4514 ) ;
  assign n4516 = ~n348 & n4515 ;
  assign n4517 = ( n417 & ~n80 ) | ( n417 & n4516 ) | ( ~n80 & n4516 ) ;
  assign n4518 = ~n417 & n4517 ;
  assign n4519 = ~n104 & n4518 ;
  assign n4520 = ( n1362 & ~n3694 ) | ( n1362 & n4519 ) | ( ~n3694 & n4519 ) ;
  assign n4521 = ( n2427 & ~n1362 ) | ( n2427 & n4520 ) | ( ~n1362 & n4520 ) ;
  assign n4522 = ~n2427 & n4521 ;
  assign n4523 = ( n886 & ~n4513 ) | ( n886 & n4522 ) | ( ~n4513 & n4522 ) ;
  assign n4524 = ~n886 & n4523 ;
  assign n4525 = ( n96 & ~n1580 ) | ( n96 & n4524 ) | ( ~n1580 & n4524 ) ;
  assign n4526 = ~n96 & n4525 ;
  assign n4527 = ( n1625 & ~n1762 ) | ( n1625 & n4526 ) | ( ~n1762 & n4526 ) ;
  assign n4528 = ~n1625 & n4527 ;
  assign n4529 = ( n574 & ~n99 ) | ( n574 & n4528 ) | ( ~n99 & n4528 ) ;
  assign n4530 = ~n574 & n4529 ;
  assign n4531 = ~n431 & n4530 ;
  assign n4532 = ~n676 & n2318 ;
  assign n4533 = ~n118 & n4532 ;
  assign n4534 = n812 | n3570 ;
  assign n4535 = ( n678 & ~n275 ) | ( n678 & n4534 ) | ( ~n275 & n4534 ) ;
  assign n4536 = n275 | n4535 ;
  assign n4537 = ( n490 & ~n494 ) | ( n490 & n4536 ) | ( ~n494 & n4536 ) ;
  assign n4538 = n494 | n4537 ;
  assign n4539 = ( n524 & n266 ) | ( n524 & n4538 ) | ( n266 & n4538 ) ;
  assign n4540 = ( n524 & ~n4539 ) | ( n524 & 1'b0 ) | ( ~n4539 & 1'b0 ) ;
  assign n4541 = n277 | n528 ;
  assign n4542 = ( n646 & ~n65 ) | ( n646 & n4541 ) | ( ~n65 & n4541 ) ;
  assign n4543 = n65 | n4542 ;
  assign n4544 = n337 | n2029 ;
  assign n4545 = n236 | n4544 ;
  assign n4546 = ( n4543 & ~n1075 ) | ( n4543 & n4545 ) | ( ~n1075 & n4545 ) ;
  assign n4547 = ( n1075 & ~n1388 ) | ( n1075 & n4546 ) | ( ~n1388 & n4546 ) ;
  assign n4548 = n1388 | n4547 ;
  assign n4549 = ( n4533 & ~n4540 ) | ( n4533 & n4548 ) | ( ~n4540 & n4548 ) ;
  assign n4550 = ( n1963 & ~n4549 ) | ( n1963 & n4533 ) | ( ~n4549 & n4533 ) ;
  assign n4551 = ~n1963 & n4550 ;
  assign n4552 = ( n1093 & ~n1808 ) | ( n1093 & n4551 ) | ( ~n1808 & n4551 ) ;
  assign n4553 = ( n4552 & ~n1093 ) | ( n4552 & 1'b0 ) | ( ~n1093 & 1'b0 ) ;
  assign n4554 = ( n674 & ~n797 ) | ( n674 & n4553 ) | ( ~n797 & n4553 ) ;
  assign n4555 = ~n674 & n4554 ;
  assign n4556 = ( n241 & ~n569 ) | ( n241 & n4555 ) | ( ~n569 & n4555 ) ;
  assign n4557 = ~n241 & n4556 ;
  assign n4558 = ( n433 & ~n410 ) | ( n433 & n4557 ) | ( ~n410 & n4557 ) ;
  assign n4559 = ~n433 & n4558 ;
  assign n4560 = n69 | n232 ;
  assign n4561 = n534 | n4560 ;
  assign n4562 = ( n2034 & ~n4561 ) | ( n2034 & n2853 ) | ( ~n4561 & n2853 ) ;
  assign n4563 = ~n2034 & n4562 ;
  assign n4564 = ( n1631 & ~n3066 ) | ( n1631 & n4563 ) | ( ~n3066 & n4563 ) ;
  assign n4565 = ~n1631 & n4564 ;
  assign n4566 = ( n4559 & ~n4531 ) | ( n4559 & n4565 ) | ( ~n4531 & n4565 ) ;
  assign n4567 = ( n1001 & n4531 ) | ( n1001 & n4566 ) | ( n4531 & n4566 ) ;
  assign n4568 = ~n1001 & n4567 ;
  assign n4569 = ( n416 & n4090 ) | ( n416 & n4568 ) | ( n4090 & n4568 ) ;
  assign n4570 = ~n416 & n4569 ;
  assign n4571 = ( n720 & ~n477 ) | ( n720 & n4570 ) | ( ~n477 & n4570 ) ;
  assign n4572 = ~n720 & n4571 ;
  assign n4573 = ( n617 & ~n272 ) | ( n617 & n4572 ) | ( ~n272 & n4572 ) ;
  assign n4574 = ~n617 & n4573 ;
  assign n4575 = n1671 | n1748 ;
  assign n4576 = ( n1671 & ~n1748 ) | ( n1671 & 1'b0 ) | ( ~n1748 & 1'b0 ) ;
  assign n4577 = ( n4575 & ~n1671 ) | ( n4575 & n4576 ) | ( ~n1671 & n4576 ) ;
  assign n4578 = ~n3625 & n4577 ;
  assign n4579 = ( n3625 & ~n4577 ) | ( n3625 & 1'b0 ) | ( ~n4577 & 1'b0 ) ;
  assign n4580 = n4578 | n4579 ;
  assign n4581 = n3644 | n4580 ;
  assign n4585 = n1875 | n3652 ;
  assign n4582 = n1671 | n3653 ;
  assign n4583 = ~n1748 & n3657 ;
  assign n4584 = ( n4582 & ~n4583 ) | ( n4582 & 1'b0 ) | ( ~n4583 & 1'b0 ) ;
  assign n4586 = ( n1875 & ~n4585 ) | ( n1875 & n4584 ) | ( ~n4585 & n4584 ) ;
  assign n4587 = n4581 &  n4586 ;
  assign n4588 = ( n4574 & ~n4340 ) | ( n4574 & n4587 ) | ( ~n4340 & n4587 ) ;
  assign n4589 = ( n4340 & ~x20 ) | ( n4340 & n4410 ) | ( ~x20 & n4410 ) ;
  assign n4590 = ( x20 & ~n4410 ) | ( x20 & n4340 ) | ( ~n4410 & n4340 ) ;
  assign n4591 = ( n4589 & ~n4340 ) | ( n4589 & n4590 ) | ( ~n4340 & n4590 ) ;
  assign n4592 = n1566 | n1671 ;
  assign n4593 = ( n1566 & ~n1671 ) | ( n1566 & 1'b0 ) | ( ~n1671 & 1'b0 ) ;
  assign n4594 = ( n4592 & ~n1566 ) | ( n4592 & n4593 ) | ( ~n1566 & n4593 ) ;
  assign n4595 = ~n3626 & n4594 ;
  assign n4596 = ( n3626 & ~n4594 ) | ( n3626 & 1'b0 ) | ( ~n4594 & 1'b0 ) ;
  assign n4597 = n4595 | n4596 ;
  assign n4598 = n3644 | n4597 ;
  assign n4599 = ~n1748 & n3652 ;
  assign n4600 = ~n1671 & n3657 ;
  assign n4601 = n4599 | n4600 ;
  assign n4602 = ~n1566 & n3653 ;
  assign n4603 = ( n1566 & ~n4601 ) | ( n1566 & n4602 ) | ( ~n4601 & n4602 ) ;
  assign n4604 = n4598 &  n4603 ;
  assign n4605 = ( n4588 & n4591 ) | ( n4588 & n4604 ) | ( n4591 & n4604 ) ;
  assign n4606 = n4268 | n4411 ;
  assign n4607 = ( n4268 & ~n4411 ) | ( n4268 & 1'b0 ) | ( ~n4411 & 1'b0 ) ;
  assign n4608 = ( n4606 & ~n4268 ) | ( n4606 & n4607 ) | ( ~n4268 & n4607 ) ;
  assign n4609 = ( n4605 & ~n4281 ) | ( n4605 & n4608 ) | ( ~n4281 & n4608 ) ;
  assign n4610 = ( n4281 & ~n4608 ) | ( n4281 & n4605 ) | ( ~n4608 & n4605 ) ;
  assign n4611 = n4609 | n4610 ;
  assign n4617 = n4061 | n601 ;
  assign n4612 = n1151 | n4430 ;
  assign n4613 = n523 | n1378 ;
  assign n4614 = n4612 &  n4613 ;
  assign n4615 = n1267 &  n3939 ;
  assign n4616 = ( n4614 & ~n1267 ) | ( n4614 & n4615 ) | ( ~n1267 & n4615 ) ;
  assign n4618 = ( n601 & ~n4617 ) | ( n601 & n4616 ) | ( ~n4617 & n4616 ) ;
  assign n4620 = ( n4281 & n4605 ) | ( n4281 & n4608 ) | ( n4605 & n4608 ) ;
  assign n4621 = ( n4608 & ~n4620 ) | ( n4608 & n4610 ) | ( ~n4620 & n4610 ) ;
  assign n4622 = ( n4618 & ~x29 ) | ( n4618 & n4621 ) | ( ~x29 & n4621 ) ;
  assign n4619 = ~x29 & n4618 ;
  assign n4623 = ( n4611 & ~n4622 ) | ( n4611 & n4619 ) | ( ~n4622 & n4619 ) ;
  assign n4625 = ( n4135 & n4268 ) | ( n4135 & n4412 ) | ( n4268 & n4412 ) ;
  assign n4624 = ( n4135 & ~n4412 ) | ( n4135 & n4268 ) | ( ~n4412 & n4268 ) ;
  assign n4626 = ( n4412 & ~n4625 ) | ( n4412 & n4624 ) | ( ~n4625 & n4624 ) ;
  assign n4627 = n1483 &  n3657 ;
  assign n4628 = ~n1566 & n3652 ;
  assign n4629 = ~n1378 & n1483 ;
  assign n4630 = ( n1378 & ~n1483 ) | ( n1378 & 1'b0 ) | ( ~n1483 & 1'b0 ) ;
  assign n4631 = n4629 | n4630 ;
  assign n4632 = n3628 &  n4631 ;
  assign n4633 = ( n3628 & ~n3644 ) | ( n3628 & n4631 ) | ( ~n3644 & n4631 ) ;
  assign n4634 = ( n4628 & ~n4632 ) | ( n4628 & n4633 ) | ( ~n4632 & n4633 ) ;
  assign n4635 = n4627 | n4634 ;
  assign n4636 = ~n1378 & n3653 ;
  assign n4637 = ( n1378 & ~n4635 ) | ( n1378 & n4636 ) | ( ~n4635 & n4636 ) ;
  assign n4638 = ( n4623 & n4626 ) | ( n4623 & n4637 ) | ( n4626 & n4637 ) ;
  assign n4642 = ~n946 & n4430 ;
  assign n4639 = n523 | n1151 ;
  assign n4640 = n1043 | n3939 ;
  assign n4641 = n4639 &  n4640 ;
  assign n4643 = ( n946 & n4642 ) | ( n946 & n4641 ) | ( n4642 & n4641 ) ;
  assign n4644 = n601 | n4038 ;
  assign n4645 = n4643 &  n4644 ;
  assign n4646 = x29 &  n4645 ;
  assign n4647 = x29 | n4645 ;
  assign n4648 = ~n4646 & n4647 ;
  assign n4649 = ( n4505 & n4638 ) | ( n4505 & n4648 ) | ( n4638 & n4648 ) ;
  assign n4651 = ( n4219 & n4429 ) | ( n4219 & n4440 ) | ( n4429 & n4440 ) ;
  assign n4650 = ( n4219 & ~n4429 ) | ( n4219 & n4440 ) | ( ~n4429 & n4440 ) ;
  assign n4652 = ( n4429 & ~n4651 ) | ( n4429 & n4650 ) | ( ~n4651 & n4650 ) ;
  assign n4653 = ( n4502 & n4649 ) | ( n4502 & n4652 ) | ( n4649 & n4652 ) ;
  assign n4654 = ~n523 & n1483 ;
  assign n4655 = n1378 | n3939 ;
  assign n4656 = ~n4654 & n4655 ;
  assign n4657 = n1267 &  n4430 ;
  assign n4658 = ( n4656 & ~n1267 ) | ( n4656 & n4657 ) | ( ~n1267 & n4657 ) ;
  assign n4659 = ( n601 & n4422 ) | ( n601 & n4658 ) | ( n4422 & n4658 ) ;
  assign n4660 = ~n601 & n4659 ;
  assign n4661 = ( x29 & ~n4658 ) | ( x29 & n4660 ) | ( ~n4658 & n4660 ) ;
  assign n4662 = ( n4658 & ~x29 ) | ( n4658 & n4660 ) | ( ~x29 & n4660 ) ;
  assign n4663 = ( n4661 & ~n4660 ) | ( n4661 & n4662 ) | ( ~n4660 & n4662 ) ;
  assign n4664 = ( n4588 & ~n4591 ) | ( n4588 & n4604 ) | ( ~n4591 & n4604 ) ;
  assign n4665 = ( n4588 & ~n4604 ) | ( n4588 & n4591 ) | ( ~n4604 & n4591 ) ;
  assign n4666 = ( n4664 & ~n4588 ) | ( n4664 & n4665 ) | ( ~n4588 & n4665 ) ;
  assign n4670 = n680 | n1496 ;
  assign n4671 = ( n3031 & ~n1271 ) | ( n3031 & n4670 ) | ( ~n1271 & n4670 ) ;
  assign n4672 = n1271 | n4671 ;
  assign n4673 = ( n428 & ~n1384 ) | ( n428 & n4672 ) | ( ~n1384 & n4672 ) ;
  assign n4674 = n1384 | n4673 ;
  assign n4675 = ( n1877 & ~n4674 ) | ( n1877 & n3050 ) | ( ~n4674 & n3050 ) ;
  assign n4676 = ~n1877 & n4675 ;
  assign n4677 = ( n904 & ~n1122 ) | ( n904 & n4676 ) | ( ~n1122 & n4676 ) ;
  assign n4678 = n1122 &  n4677 ;
  assign n4679 = ( n2128 & ~n3303 ) | ( n2128 & n4678 ) | ( ~n3303 & n4678 ) ;
  assign n4680 = ~n2128 & n4679 ;
  assign n4681 = ( n383 & ~n1625 ) | ( n383 & n4680 ) | ( ~n1625 & n4680 ) ;
  assign n4682 = ( n775 & ~n383 ) | ( n775 & n4681 ) | ( ~n383 & n4681 ) ;
  assign n4683 = ~n775 & n4682 ;
  assign n4684 = ( n255 & ~n734 ) | ( n255 & n4683 ) | ( ~n734 & n4683 ) ;
  assign n4685 = ~n255 & n4684 ;
  assign n4686 = ~n492 & n4685 ;
  assign n4687 = n2091 | n2666 ;
  assign n4688 = ( n351 & ~n72 ) | ( n351 & n4687 ) | ( ~n72 & n4687 ) ;
  assign n4689 = n72 | n4688 ;
  assign n4690 = n382 | n2036 ;
  assign n4691 = ( n452 & ~n561 ) | ( n452 & n4690 ) | ( ~n561 & n4690 ) ;
  assign n4692 = n561 | n4691 ;
  assign n4693 = ( n80 & ~n571 ) | ( n80 & n4692 ) | ( ~n571 & n4692 ) ;
  assign n4694 = n571 | n4693 ;
  assign n4695 = n459 | n4694 ;
  assign n4696 = n372 | n1107 ;
  assign n4697 = n451 | n4696 ;
  assign n4698 = ( n1073 & ~n4697 ) | ( n1073 & n1829 ) | ( ~n4697 & n1829 ) ;
  assign n4699 = ~n1829 & n4698 ;
  assign n4700 = ~n2593 & n4699 ;
  assign n4701 = ( n4689 & ~n4695 ) | ( n4689 & n4700 ) | ( ~n4695 & n4700 ) ;
  assign n4702 = ( n1044 & ~n4689 ) | ( n1044 & n4701 ) | ( ~n4689 & n4701 ) ;
  assign n4703 = ( n4702 & ~n1044 ) | ( n4702 & 1'b0 ) | ( ~n1044 & 1'b0 ) ;
  assign n4704 = ( n948 & n2190 ) | ( n948 & n4703 ) | ( n2190 & n4703 ) ;
  assign n4705 = ~n948 & n4704 ;
  assign n4706 = ( n124 & ~n105 ) | ( n124 & n4705 ) | ( ~n105 & n4705 ) ;
  assign n4707 = ~n124 & n4706 ;
  assign n4708 = ( n272 & ~n52 ) | ( n272 & n4707 ) | ( ~n52 & n4707 ) ;
  assign n4709 = ~n272 & n4708 ;
  assign n4710 = ( n123 & ~n384 ) | ( n123 & n4709 ) | ( ~n384 & n4709 ) ;
  assign n4711 = ~n123 & n4710 ;
  assign n4712 = ( n492 & ~n4711 ) | ( n492 & n623 ) | ( ~n4711 & n623 ) ;
  assign n4713 = ( n623 & ~n4712 ) | ( n623 & 1'b0 ) | ( ~n4712 & 1'b0 ) ;
  assign n4714 = n221 | n224 ;
  assign n4715 = ( n229 & ~n433 ) | ( n229 & n4714 ) | ( ~n433 & n4714 ) ;
  assign n4716 = n433 | n4715 ;
  assign n4717 = n357 | n403 ;
  assign n4718 = n239 | n4717 ;
  assign n4719 = ( n4716 & ~n3171 ) | ( n4716 & n4718 ) | ( ~n3171 & n4718 ) ;
  assign n4720 = n3171 | n4719 ;
  assign n4721 = ( n4713 & ~n1352 ) | ( n4713 & n4720 ) | ( ~n1352 & n4720 ) ;
  assign n4722 = ( n764 & ~n4721 ) | ( n764 & n4713 ) | ( ~n4721 & n4713 ) ;
  assign n4723 = ~n764 & n4722 ;
  assign n4724 = ( n1493 & ~n1808 ) | ( n1493 & n4723 ) | ( ~n1808 & n4723 ) ;
  assign n4725 = ~n1493 & n4724 ;
  assign n4726 = ( n527 & ~n479 ) | ( n527 & n4725 ) | ( ~n479 & n4725 ) ;
  assign n4727 = ~n527 & n4726 ;
  assign n4728 = ( n277 & ~n69 ) | ( n277 & n4727 ) | ( ~n69 & n4727 ) ;
  assign n4729 = ~n277 & n4728 ;
  assign n4730 = ( n775 & ~n793 ) | ( n775 & n4729 ) | ( ~n793 & n4729 ) ;
  assign n4731 = ~n775 & n4730 ;
  assign n4732 = ( n187 & ~n2428 ) | ( n187 & n4731 ) | ( ~n2428 & n4731 ) ;
  assign n4733 = ~n187 & n4732 ;
  assign n4734 = ( n269 & ~n534 ) | ( n269 & n4733 ) | ( ~n534 & n4733 ) ;
  assign n4735 = ~n269 & n4734 ;
  assign n4736 = ~n169 & n4735 ;
  assign n4737 = ( x17 & n4686 ) | ( x17 & n4736 ) | ( n4686 & n4736 ) ;
  assign n4738 = n1748 | n1875 ;
  assign n4739 = ( n1748 & ~n1875 ) | ( n1748 & 1'b0 ) | ( ~n1875 & 1'b0 ) ;
  assign n4740 = ( n4738 & ~n1748 ) | ( n4738 & n4739 ) | ( ~n1748 & n4739 ) ;
  assign n4741 = ~n3624 & n4740 ;
  assign n4742 = ( n3624 & ~n4740 ) | ( n3624 & 1'b0 ) | ( ~n4740 & 1'b0 ) ;
  assign n4743 = n4741 | n4742 ;
  assign n4744 = n3644 | n4743 ;
  assign n4745 = ~n1940 & n3652 ;
  assign n4746 = ~n1875 & n3657 ;
  assign n4747 = n4745 | n4746 ;
  assign n4748 = ~n1748 & n3653 ;
  assign n4749 = ( n1748 & ~n4747 ) | ( n1748 & n4748 ) | ( ~n4747 & n4748 ) ;
  assign n4750 = n4744 &  n4749 ;
  assign n4751 = ( n4737 & ~n4340 ) | ( n4737 & n4750 ) | ( ~n4340 & n4750 ) ;
  assign n4667 = ( n4340 & ~n4574 ) | ( n4340 & n4587 ) | ( ~n4574 & n4587 ) ;
  assign n4668 = ( n4340 & ~n4587 ) | ( n4340 & n4574 ) | ( ~n4587 & n4574 ) ;
  assign n4669 = ( n4667 & ~n4340 ) | ( n4667 & n4668 ) | ( ~n4340 & n4668 ) ;
  assign n4951 = n4274 | n601 ;
  assign n4946 = n523 | n1671 ;
  assign n4947 = n1566 | n3939 ;
  assign n4948 = n4946 &  n4947 ;
  assign n4949 = n1483 &  n4430 ;
  assign n4950 = ( n4948 & ~n1483 ) | ( n4948 & n4949 ) | ( ~n1483 & n4949 ) ;
  assign n4952 = ( n601 & ~n4951 ) | ( n601 & n4950 ) | ( ~n4951 & n4950 ) ;
  assign n4953 = ~x29 & n4952 ;
  assign n4752 = ( n4340 & ~n4737 ) | ( n4340 & n4750 ) | ( ~n4737 & n4750 ) ;
  assign n4753 = ( n4340 & ~n4750 ) | ( n4340 & n4737 ) | ( ~n4750 & n4737 ) ;
  assign n4754 = ( n4752 & ~n4340 ) | ( n4752 & n4753 ) | ( ~n4340 & n4753 ) ;
  assign n4755 = ( x17 & ~n4686 ) | ( x17 & n4736 ) | ( ~n4686 & n4736 ) ;
  assign n4756 = ( n4686 & ~n4737 ) | ( n4686 & n4755 ) | ( ~n4737 & n4755 ) ;
  assign n4766 = ~n1875 & n3653 ;
  assign n4757 = ~n1940 & n3657 ;
  assign n4759 = n1875 | n1940 ;
  assign n4760 = ( n1875 & ~n1940 ) | ( n1875 & 1'b0 ) | ( ~n1940 & 1'b0 ) ;
  assign n4761 = ( n4759 & ~n1875 ) | ( n4759 & n4760 ) | ( ~n1875 & n4760 ) ;
  assign n4762 = ( n3623 & ~n4761 ) | ( n3623 & 1'b0 ) | ( ~n4761 & 1'b0 ) ;
  assign n4758 = ~n2022 & n3652 ;
  assign n4763 = ( n3644 & ~n3623 ) | ( n3644 & n4761 ) | ( ~n3623 & n4761 ) ;
  assign n4764 = ( n4762 & ~n4758 ) | ( n4762 & n4763 ) | ( ~n4758 & n4763 ) ;
  assign n4765 = ~n4757 & n4764 ;
  assign n4767 = ( n1875 & n4766 ) | ( n1875 & n4765 ) | ( n4766 & n4765 ) ;
  assign n4768 = n1232 | n3307 ;
  assign n4769 = ( n1385 & ~n1955 ) | ( n1385 & n4768 ) | ( ~n1955 & n4768 ) ;
  assign n4770 = n1955 | n4769 ;
  assign n4771 = ( n83 & n4770 ) | ( n83 & n354 ) | ( n4770 & n354 ) ;
  assign n4772 = ( n354 & ~n4771 ) | ( n354 & 1'b0 ) | ( ~n4771 & 1'b0 ) ;
  assign n4773 = ~n212 & n4772 ;
  assign n4774 = n139 | n3267 ;
  assign n4775 = n336 | n4774 ;
  assign n4776 = ( n535 & ~n1810 ) | ( n535 & n4775 ) | ( ~n1810 & n4775 ) ;
  assign n4777 = n1810 | n4776 ;
  assign n4778 = ( n929 & ~n4777 ) | ( n929 & n2804 ) | ( ~n4777 & n2804 ) ;
  assign n4779 = ~n2804 & n4778 ;
  assign n4780 = ( n124 & ~n1152 ) | ( n124 & n4779 ) | ( ~n1152 & n4779 ) ;
  assign n4781 = ~n124 & n4780 ;
  assign n4782 = ( n58 & ~n674 ) | ( n58 & n4781 ) | ( ~n674 & n4781 ) ;
  assign n4783 = ~n58 & n4782 ;
  assign n4784 = ( n720 & ~n911 ) | ( n720 & n4783 ) | ( ~n911 & n4783 ) ;
  assign n4785 = ~n720 & n4784 ;
  assign n4786 = ( n151 & ~n268 ) | ( n151 & n4785 ) | ( ~n268 & n4785 ) ;
  assign n4787 = ~n151 & n4786 ;
  assign n4788 = ~n572 & n4787 ;
  assign n4789 = n1635 | n3070 ;
  assign n4790 = ( n3304 & ~n3142 ) | ( n3304 & n4789 ) | ( ~n3142 & n4789 ) ;
  assign n4791 = n3142 | n4790 ;
  assign n4792 = ( n3679 & ~n4788 ) | ( n3679 & n4791 ) | ( ~n4788 & n4791 ) ;
  assign n4793 = ( n3679 & ~n4792 ) | ( n3679 & 1'b0 ) | ( ~n4792 & 1'b0 ) ;
  assign n4794 = ( n171 & n4773 ) | ( n171 & n4793 ) | ( n4773 & n4793 ) ;
  assign n4795 = ~n171 & n4794 ;
  assign n4796 = ( n2666 & ~n3551 ) | ( n2666 & n4795 ) | ( ~n3551 & n4795 ) ;
  assign n4797 = ~n2666 & n4796 ;
  assign n4798 = ( n345 & ~n216 ) | ( n345 & n4797 ) | ( ~n216 & n4797 ) ;
  assign n4799 = ~n345 & n4798 ;
  assign n4800 = ( n453 & ~n269 ) | ( n453 & n4799 ) | ( ~n269 & n4799 ) ;
  assign n4801 = ~n453 & n4800 ;
  assign n4802 = ( n382 & ~n559 ) | ( n382 & n4801 ) | ( ~n559 & n4801 ) ;
  assign n4803 = ~n382 & n4802 ;
  assign n4804 = ( n478 & ~n646 ) | ( n478 & n4803 ) | ( ~n646 & n4803 ) ;
  assign n4805 = ~n478 & n4804 ;
  assign n4806 = ( n358 & ~n229 ) | ( n358 & n4805 ) | ( ~n229 & n4805 ) ;
  assign n4807 = ~n358 & n4806 ;
  assign n4808 = n735 | n796 ;
  assign n4809 = ( n258 & ~n1496 ) | ( n258 & n4808 ) | ( ~n1496 & n4808 ) ;
  assign n4810 = n1496 | n4809 ;
  assign n4811 = ( n338 & ~n372 ) | ( n338 & n4810 ) | ( ~n372 & n4810 ) ;
  assign n4812 = n372 | n4811 ;
  assign n4813 = n39 | n4812 ;
  assign n4814 = n362 | n711 ;
  assign n4815 = ( n411 & ~n187 ) | ( n411 & n4814 ) | ( ~n187 & n4814 ) ;
  assign n4816 = n187 | n4815 ;
  assign n4817 = ( n336 & ~n454 ) | ( n336 & n4816 ) | ( ~n454 & n4816 ) ;
  assign n4818 = n454 | n4817 ;
  assign n4819 = n2864 | n3552 ;
  assign n4820 = ( n4773 & n4818 ) | ( n4773 & n4819 ) | ( n4818 & n4819 ) ;
  assign n4821 = ( n4773 & ~n4820 ) | ( n4773 & 1'b0 ) | ( ~n4820 & 1'b0 ) ;
  assign n4822 = ( n1045 & ~n4813 ) | ( n1045 & n4821 ) | ( ~n4813 & n4821 ) ;
  assign n4823 = ~n1045 & n4822 ;
  assign n4824 = ( n1808 & ~n70 ) | ( n1808 & n4823 ) | ( ~n70 & n4823 ) ;
  assign n4825 = ~n1808 & n4824 ;
  assign n4826 = ( n208 & ~n101 ) | ( n208 & n4825 ) | ( ~n101 & n4825 ) ;
  assign n4827 = ~n208 & n4826 ;
  assign n4828 = ( n456 & ~n745 ) | ( n456 & n4827 ) | ( ~n745 & n4827 ) ;
  assign n4829 = ~n456 & n4828 ;
  assign n4830 = ( n80 & ~n4829 ) | ( n80 & n623 ) | ( ~n4829 & n623 ) ;
  assign n4831 = ( n623 & ~n4830 ) | ( n623 & 1'b0 ) | ( ~n4830 & 1'b0 ) ;
  assign n4832 = ~n630 & n4831 ;
  assign n4842 = n348 | n720 ;
  assign n4840 = ( n524 & ~n788 ) | ( n524 & 1'b0 ) | ( ~n788 & 1'b0 ) ;
  assign n4841 = ~n334 & n4840 ;
  assign n4843 = ( n4310 & ~n4842 ) | ( n4310 & n4841 ) | ( ~n4842 & n4841 ) ;
  assign n4844 = ( n4843 & ~n4310 ) | ( n4843 & 1'b0 ) | ( ~n4310 & 1'b0 ) ;
  assign n4833 = ( n410 & ~n554 ) | ( n410 & n792 ) | ( ~n554 & n792 ) ;
  assign n4834 = n554 | n4833 ;
  assign n4835 = n3171 | n4834 ;
  assign n4836 = ( n495 & ~n415 ) | ( n495 & n4835 ) | ( ~n415 & n4835 ) ;
  assign n4837 = n415 | n4836 ;
  assign n4838 = ( n340 & ~n490 ) | ( n340 & n4837 ) | ( ~n490 & n4837 ) ;
  assign n4839 = n490 | n4838 ;
  assign n4845 = ( n929 & ~n4844 ) | ( n929 & n4839 ) | ( ~n4844 & n4839 ) ;
  assign n4846 = ( n929 & ~n4845 ) | ( n929 & 1'b0 ) | ( ~n4845 & 1'b0 ) ;
  assign n4847 = ( n3011 & ~n298 ) | ( n3011 & n4846 ) | ( ~n298 & n4846 ) ;
  assign n4848 = ( n186 & ~n3011 ) | ( n186 & n4847 ) | ( ~n3011 & n4847 ) ;
  assign n4849 = ~n186 & n4848 ;
  assign n4850 = ( n4832 & n1044 ) | ( n4832 & n4849 ) | ( n1044 & n4849 ) ;
  assign n4851 = ~n1044 & n4850 ;
  assign n4852 = ( n761 & ~n1061 ) | ( n761 & n4851 ) | ( ~n1061 & n4851 ) ;
  assign n4853 = ~n761 & n4852 ;
  assign n4854 = ( n356 & ~n384 ) | ( n356 & n4853 ) | ( ~n384 & n4853 ) ;
  assign n4855 = ~n356 & n4854 ;
  assign n4856 = ( n459 & ~n353 ) | ( n459 & n4855 ) | ( ~n353 & n4855 ) ;
  assign n4857 = ~n459 & n4856 ;
  assign n4858 = ~n433 & n4857 ;
  assign n4859 = n260 | n568 ;
  assign n4860 = n2087 | n3146 ;
  assign n4861 = ( n4859 & ~n479 ) | ( n4859 & n4860 ) | ( ~n479 & n4860 ) ;
  assign n4862 = n479 | n4861 ;
  assign n4863 = ( n676 & ~n234 ) | ( n676 & n4862 ) | ( ~n234 & n4862 ) ;
  assign n4864 = n234 | n4863 ;
  assign n4865 = ( n207 & ~n217 ) | ( n207 & n4864 ) | ( ~n217 & n4864 ) ;
  assign n4866 = n217 | n4865 ;
  assign n4867 = ( n197 & ~n4866 ) | ( n197 & n349 ) | ( ~n4866 & n349 ) ;
  assign n4868 = ~n349 & n4867 ;
  assign n4874 = ~n1797 & n4519 ;
  assign n4875 = ( n1279 & ~n4874 ) | ( n1279 & n3113 ) | ( ~n4874 & n3113 ) ;
  assign n4876 = ( n1279 & ~n4875 ) | ( n1279 & 1'b0 ) | ( ~n4875 & 1'b0 ) ;
  assign n4877 = ( n605 & ~n1244 ) | ( n605 & n4876 ) | ( ~n1244 & n4876 ) ;
  assign n4878 = ~n605 & n4877 ;
  assign n4879 = ( n434 & ~n912 ) | ( n434 & n4878 ) | ( ~n912 & n4878 ) ;
  assign n4880 = ~n434 & n4879 ;
  assign n4881 = ( n672 & ~n235 ) | ( n672 & n4880 ) | ( ~n235 & n4880 ) ;
  assign n4882 = ~n672 & n4881 ;
  assign n4883 = ( n245 & ~n415 ) | ( n245 & n4882 ) | ( ~n415 & n4882 ) ;
  assign n4884 = ~n245 & n4883 ;
  assign n4885 = ( n272 & ~n494 ) | ( n272 & n4884 ) | ( ~n494 & n4884 ) ;
  assign n4886 = ~n272 & n4885 ;
  assign n4887 = ( n457 & ~n237 ) | ( n457 & n4886 ) | ( ~n237 & n4886 ) ;
  assign n4888 = ~n457 & n4887 ;
  assign n4889 = ( n129 & ~n240 ) | ( n129 & n4888 ) | ( ~n240 & n4888 ) ;
  assign n4890 = ~n129 & n4889 ;
  assign n4891 = ~n375 & n3043 ;
  assign n4892 = ( n1233 & ~n4718 ) | ( n1233 & n4891 ) | ( ~n4718 & n4891 ) ;
  assign n4893 = ~n1233 & n4892 ;
  assign n4894 = ( n3890 & ~n3527 ) | ( n3890 & n4893 ) | ( ~n3527 & n4893 ) ;
  assign n4895 = ( n493 & ~n3890 ) | ( n493 & n4894 ) | ( ~n3890 & n4894 ) ;
  assign n4896 = ~n493 & n4895 ;
  assign n4897 = ( n244 & ~n232 ) | ( n244 & n4896 ) | ( ~n232 & n4896 ) ;
  assign n4898 = ~n244 & n4897 ;
  assign n4899 = n2206 | n4775 ;
  assign n4900 = ( n4898 & n1059 ) | ( n4898 & n4899 ) | ( n1059 & n4899 ) ;
  assign n4901 = ( n1585 & ~n4900 ) | ( n1585 & n4898 ) | ( ~n4900 & n4898 ) ;
  assign n4902 = ~n1585 & n4901 ;
  assign n4903 = ( n345 & ~n2462 ) | ( n345 & n4902 ) | ( ~n2462 & n4902 ) ;
  assign n4904 = ~n345 & n4903 ;
  assign n4905 = ( n4904 & ~n712 ) | ( n4904 & n745 ) | ( ~n712 & n745 ) ;
  assign n4906 = ( n4905 & ~n745 ) | ( n4905 & 1'b0 ) | ( ~n745 & 1'b0 ) ;
  assign n4907 = ( n460 & ~n452 ) | ( n460 & n4906 ) | ( ~n452 & n4906 ) ;
  assign n4908 = ~n460 & n4907 ;
  assign n4909 = ( n169 & ~n141 ) | ( n169 & n4908 ) | ( ~n141 & n4908 ) ;
  assign n4910 = ~n169 & n4909 ;
  assign n4911 = ~n347 & n4910 ;
  assign n4912 = n562 | n1076 ;
  assign n4913 = ( n2279 & ~n1993 ) | ( n2279 & n4912 ) | ( ~n1993 & n4912 ) ;
  assign n4914 = n1993 | n4913 ;
  assign n4915 = ( n4890 & ~n4911 ) | ( n4890 & n4914 ) | ( ~n4911 & n4914 ) ;
  assign n4916 = ( n577 & ~n4915 ) | ( n577 & n4890 ) | ( ~n4915 & n4890 ) ;
  assign n4917 = ~n577 & n4916 ;
  assign n4869 = n127 | n2578 ;
  assign n4870 = ( n216 & ~n243 ) | ( n216 & n4869 ) | ( ~n243 & n4869 ) ;
  assign n4871 = n243 | n4870 ;
  assign n4872 = ( n351 & ~n83 ) | ( n351 & n4871 ) | ( ~n83 & n4871 ) ;
  assign n4873 = n83 | n4872 ;
  assign n4918 = ( n4868 & ~n4917 ) | ( n4868 & n4873 ) | ( ~n4917 & n4873 ) ;
  assign n4919 = ( n1807 & ~n4918 ) | ( n1807 & n4868 ) | ( ~n4918 & n4868 ) ;
  assign n4920 = ~n1807 & n4919 ;
  assign n4921 = ( n1511 & ~n866 ) | ( n1511 & n4920 ) | ( ~n866 & n4920 ) ;
  assign n4922 = ~n1511 & n4921 ;
  assign n4923 = ( n157 & ~n69 ) | ( n157 & n4922 ) | ( ~n69 & n4922 ) ;
  assign n4924 = ~n157 & n4923 ;
  assign n4925 = ( n359 & ~n569 ) | ( n359 & n4924 ) | ( ~n569 & n4924 ) ;
  assign n4926 = ~n359 & n4925 ;
  assign n4927 = ~n643 & n4926 ;
  assign n4928 = ( x14 & n4858 ) | ( x14 & n4927 ) | ( n4858 & n4927 ) ;
  assign n4929 = n2022 | n2127 ;
  assign n4930 = ( n2022 & ~n2127 ) | ( n2022 & 1'b0 ) | ( ~n2127 & 1'b0 ) ;
  assign n4931 = ( n4929 & ~n2022 ) | ( n4929 & n4930 ) | ( ~n2022 & n4930 ) ;
  assign n4932 = ~n3621 & n4931 ;
  assign n4933 = ( n3621 & ~n4931 ) | ( n3621 & 1'b0 ) | ( ~n4931 & 1'b0 ) ;
  assign n4934 = n4932 | n4933 ;
  assign n4935 = n3644 | n4934 ;
  assign n4936 = ~n2178 & n3652 ;
  assign n4937 = ~n2127 & n3657 ;
  assign n4938 = n4936 | n4937 ;
  assign n4939 = ~n2022 & n3653 ;
  assign n4940 = ( n2022 & ~n4938 ) | ( n2022 & n4939 ) | ( ~n4938 & n4939 ) ;
  assign n4941 = n4935 &  n4940 ;
  assign n4942 = ( n4928 & ~n4807 ) | ( n4928 & n4941 ) | ( ~n4807 & n4941 ) ;
  assign n4943 = ( n4807 & ~n4686 ) | ( n4807 & n4942 ) | ( ~n4686 & n4942 ) ;
  assign n4944 = ( n4756 & n4767 ) | ( n4756 & n4943 ) | ( n4767 & n4943 ) ;
  assign n4945 = ( n4754 & ~n4944 ) | ( n4754 & 1'b0 ) | ( ~n4944 & 1'b0 ) ;
  assign n4954 = ~n4754 & n4944 ;
  assign n4955 = ( x29 & ~n4952 ) | ( x29 & n4954 ) | ( ~n4952 & n4954 ) ;
  assign n4956 = ( n4953 & ~n4945 ) | ( n4953 & n4955 ) | ( ~n4945 & n4955 ) ;
  assign n4957 = ( n4751 & ~n4669 ) | ( n4751 & n4956 ) | ( ~n4669 & n4956 ) ;
  assign n4958 = ( n4663 & n4666 ) | ( n4663 & n4957 ) | ( n4666 & n4957 ) ;
  assign n4960 = ( x29 & n4618 ) | ( x29 & n4621 ) | ( n4618 & n4621 ) ;
  assign n4959 = ( x29 & ~n4621 ) | ( x29 & n4618 ) | ( ~n4621 & n4618 ) ;
  assign n4961 = ( n4621 & ~n4960 ) | ( n4621 & n4959 ) | ( ~n4960 & n4959 ) ;
  assign n4966 = ~n946 & n4495 ;
  assign n4962 = ~n4474 |  n4477 ;
  assign n4963 = n863 | n4962 ;
  assign n4964 = n1043 | n4482 ;
  assign n4965 = n4963 &  n4964 ;
  assign n4967 = ( n946 & n4966 ) | ( n946 & n4965 ) | ( n4966 & n4965 ) ;
  assign n4968 = ( n4478 & ~n3914 ) | ( n4478 & n4967 ) | ( ~n3914 & n4967 ) ;
  assign n4969 = ~n4478 & n4968 ;
  assign n4970 = ( x26 & ~n4967 ) | ( x26 & n4969 ) | ( ~n4967 & n4969 ) ;
  assign n4971 = ( n4967 & ~x26 ) | ( n4967 & n4969 ) | ( ~x26 & n4969 ) ;
  assign n4972 = ( n4970 & ~n4969 ) | ( n4970 & n4971 ) | ( ~n4969 & n4971 ) ;
  assign n4973 = ( n4958 & n4961 ) | ( n4958 & n4972 ) | ( n4961 & n4972 ) ;
  assign n4977 = n1267 | n523 ;
  assign n4974 = n1043 | n4430 ;
  assign n4975 = n1151 | n3939 ;
  assign n4976 = n4974 &  n4975 ;
  assign n4978 = ( n523 & ~n4977 ) | ( n523 & n4976 ) | ( ~n4977 & n4976 ) ;
  assign n4979 = ( n601 & ~n3952 ) | ( n601 & n4978 ) | ( ~n3952 & n4978 ) ;
  assign n4980 = ~n601 & n4979 ;
  assign n4981 = ( x29 & ~n4978 ) | ( x29 & n4980 ) | ( ~n4978 & n4980 ) ;
  assign n4982 = ( n4978 & ~x29 ) | ( n4978 & n4980 ) | ( ~x29 & n4980 ) ;
  assign n4983 = ( n4981 & ~n4980 ) | ( n4981 & n4982 ) | ( ~n4980 & n4982 ) ;
  assign n4984 = ( n4626 & ~n4623 ) | ( n4626 & n4637 ) | ( ~n4623 & n4637 ) ;
  assign n4985 = ( n4623 & ~n4637 ) | ( n4623 & n4626 ) | ( ~n4637 & n4626 ) ;
  assign n4986 = ( n4984 & ~n4626 ) | ( n4984 & n4985 ) | ( ~n4626 & n4985 ) ;
  assign n4990 = ~n946 & n4482 ;
  assign n4987 = n702 | n4962 ;
  assign n4988 = n863 | n4495 ;
  assign n4989 = n4987 &  n4988 ;
  assign n4991 = ( n946 & n4990 ) | ( n946 & n4989 ) | ( n4990 & n4989 ) ;
  assign n4992 = ( n3650 & ~n4478 ) | ( n3650 & n4991 ) | ( ~n4478 & n4991 ) ;
  assign n4993 = ~n3650 & n4992 ;
  assign n4994 = ( x26 & ~n4991 ) | ( x26 & n4993 ) | ( ~n4991 & n4993 ) ;
  assign n4995 = ( n4991 & ~x26 ) | ( n4991 & n4993 ) | ( ~x26 & n4993 ) ;
  assign n4996 = ( n4994 & ~n4993 ) | ( n4994 & n4995 ) | ( ~n4993 & n4995 ) ;
  assign n4997 = ( n4983 & ~n4986 ) | ( n4983 & n4996 ) | ( ~n4986 & n4996 ) ;
  assign n4998 = ( n4983 & ~n4996 ) | ( n4983 & n4986 ) | ( ~n4996 & n4986 ) ;
  assign n4999 = ( n4997 & ~n4983 ) | ( n4997 & n4998 ) | ( ~n4983 & n4998 ) ;
  assign n5003 = ( x20 & ~x21 ) | ( x20 & 1'b0 ) | ( ~x21 & 1'b0 ) ;
  assign n5004 = ~x20 & x21 ;
  assign n5005 = n5003 | n5004 ;
  assign n5006 = ~x22 & x23 ;
  assign n5007 = ( x22 & ~x23 ) | ( x22 & 1'b0 ) | ( ~x23 & 1'b0 ) ;
  assign n5008 = n5006 | n5007 ;
  assign n5012 = ~n5005 | ~n5008 ;
  assign n5000 = ~x21 & x22 ;
  assign n5001 = ( x21 & ~x22 ) | ( x21 & 1'b0 ) | ( ~x22 & 1'b0 ) ;
  assign n5002 = n5000 | n5001 ;
  assign n5009 = ( n5002 & ~n5005 ) | ( n5002 & n5008 ) | ( ~n5005 & n5008 ) ;
  assign n5010 = ~n5009 |  n5002 ;
  assign n5011 = n599 | n5010 ;
  assign n5013 = ( n3637 & ~n5012 ) | ( n3637 & n5011 ) | ( ~n5012 & n5011 ) ;
  assign n5014 = ~n3637 & n5013 ;
  assign n5016 = ( x23 & n5011 ) | ( x23 & n5014 ) | ( n5011 & n5014 ) ;
  assign n5015 = ( x23 & ~n5014 ) | ( x23 & n5011 ) | ( ~n5014 & n5011 ) ;
  assign n5017 = ( n5014 & ~n5016 ) | ( n5014 & n5015 ) | ( ~n5016 & n5015 ) ;
  assign n5018 = ( n4973 & ~n4999 ) | ( n4973 & n5017 ) | ( ~n4999 & n5017 ) ;
  assign n5019 = ( n4973 & ~n5017 ) | ( n4973 & n4999 ) | ( ~n5017 & n4999 ) ;
  assign n5020 = ( n5018 & ~n4973 ) | ( n5018 & n5019 ) | ( ~n4973 & n5019 ) ;
  assign n5021 = ( n4666 & ~n4663 ) | ( n4666 & n4957 ) | ( ~n4663 & n4957 ) ;
  assign n5022 = ( n4663 & ~n4957 ) | ( n4663 & n4666 ) | ( ~n4957 & n4666 ) ;
  assign n5023 = ( n5021 & ~n4666 ) | ( n5021 & n5022 ) | ( ~n4666 & n5022 ) ;
  assign n5027 = ~n946 & n4962 ;
  assign n5024 = n1151 | n4482 ;
  assign n5025 = n1043 | n4495 ;
  assign n5026 = n5024 &  n5025 ;
  assign n5028 = ( n946 & n5027 ) | ( n946 & n5026 ) | ( n5027 & n5026 ) ;
  assign n5029 = ( n4478 & ~n4038 ) | ( n4478 & n5028 ) | ( ~n4038 & n5028 ) ;
  assign n5030 = ~n4478 & n5029 ;
  assign n5031 = ( x26 & ~n5028 ) | ( x26 & n5030 ) | ( ~n5028 & n5030 ) ;
  assign n5032 = ( n5028 & ~x26 ) | ( n5028 & n5030 ) | ( ~x26 & n5030 ) ;
  assign n5033 = ( n5031 & ~n5030 ) | ( n5031 & n5032 ) | ( ~n5030 & n5032 ) ;
  assign n5049 = n1043 | n4962 ;
  assign n5050 = n1151 | n4495 ;
  assign n5051 = n5049 &  n5050 ;
  assign n5052 = n1267 &  n4482 ;
  assign n5053 = ( n5051 & ~n1267 ) | ( n5051 & n5052 ) | ( ~n1267 & n5052 ) ;
  assign n5054 = n3952 | n4478 ;
  assign n5055 = n5053 &  n5054 ;
  assign n5056 = ~x26 & n5055 ;
  assign n5037 = n3628 | n4631 ;
  assign n5038 = ~n4632 & n5037 ;
  assign n5044 = n601 | n5038 ;
  assign n5039 = n1378 | n4430 ;
  assign n5040 = n523 | n1566 ;
  assign n5041 = n5039 &  n5040 ;
  assign n5042 = n1483 &  n3939 ;
  assign n5043 = ( n5041 & ~n1483 ) | ( n5041 & n5042 ) | ( ~n1483 & n5042 ) ;
  assign n5045 = ( n601 & ~n5044 ) | ( n601 & n5043 ) | ( ~n5044 & n5043 ) ;
  assign n5034 = ( n4669 & n4751 ) | ( n4669 & n4956 ) | ( n4751 & n4956 ) ;
  assign n5035 = ( n4669 & ~n4751 ) | ( n4669 & n4956 ) | ( ~n4751 & n4956 ) ;
  assign n5036 = ( n4751 & ~n5034 ) | ( n4751 & n5035 ) | ( ~n5034 & n5035 ) ;
  assign n5046 = ( x29 & ~n5045 ) | ( x29 & n5036 ) | ( ~n5045 & n5036 ) ;
  assign n5047 = ( n5036 & ~x29 ) | ( n5036 & n5045 ) | ( ~x29 & n5045 ) ;
  assign n5048 = n5046 &  n5047 ;
  assign n5058 = ( x29 & n5036 ) | ( x29 & n5045 ) | ( n5036 & n5045 ) ;
  assign n5057 = ( x29 & ~n5036 ) | ( x29 & n5045 ) | ( ~n5036 & n5045 ) ;
  assign n5059 = ( n5036 & ~n5058 ) | ( n5036 & n5057 ) | ( ~n5058 & n5057 ) ;
  assign n5060 = ( x26 & ~n5055 ) | ( x26 & n5059 ) | ( ~n5055 & n5059 ) ;
  assign n5061 = ( n5056 & ~n5048 ) | ( n5056 & n5060 ) | ( ~n5048 & n5060 ) ;
  assign n5062 = ( n5023 & n5033 ) | ( n5023 & n5061 ) | ( n5033 & n5061 ) ;
  assign n5063 = ( n4958 & ~n4972 ) | ( n4958 & n4961 ) | ( ~n4972 & n4961 ) ;
  assign n5064 = ( n4961 & ~n4958 ) | ( n4961 & n4972 ) | ( ~n4958 & n4972 ) ;
  assign n5065 = ( n5063 & ~n4961 ) | ( n5063 & n5064 ) | ( ~n4961 & n5064 ) ;
  assign n5066 = n702 | n5010 ;
  assign n5067 = ~n5002 |  n5005 ;
  assign n5068 = n599 | n5067 ;
  assign n5069 = n5066 &  n5068 ;
  assign n5070 = ( n3937 & ~n5012 ) | ( n3937 & 1'b0 ) | ( ~n5012 & 1'b0 ) ;
  assign n5071 = ( n5069 & ~n5070 ) | ( n5069 & 1'b0 ) | ( ~n5070 & 1'b0 ) ;
  assign n5072 = x23 | n5071 ;
  assign n5073 = x23 &  n5071 ;
  assign n5074 = ( n5072 & ~n5073 ) | ( n5072 & 1'b0 ) | ( ~n5073 & 1'b0 ) ;
  assign n5075 = ( n5062 & n5065 ) | ( n5062 & n5074 ) | ( n5065 & n5074 ) ;
  assign n5081 = ~n2022 & n3657 ;
  assign n5083 = n1940 | n2022 ;
  assign n5084 = ( n1940 & ~n2022 ) | ( n1940 & 1'b0 ) | ( ~n2022 & 1'b0 ) ;
  assign n5085 = ( n5083 & ~n1940 ) | ( n5083 & n5084 ) | ( ~n1940 & n5084 ) ;
  assign n5086 = ( n3622 & ~n5085 ) | ( n3622 & 1'b0 ) | ( ~n5085 & 1'b0 ) ;
  assign n5082 = ~n2127 & n3652 ;
  assign n5087 = ( n3644 & ~n3622 ) | ( n3644 & n5085 ) | ( ~n3622 & n5085 ) ;
  assign n5088 = ( n5086 & ~n5082 ) | ( n5086 & n5087 ) | ( ~n5082 & n5087 ) ;
  assign n5089 = ~n5081 & n5088 ;
  assign n5090 = ~n1940 & n3653 ;
  assign n5091 = ( n1940 & n5089 ) | ( n1940 & n5090 ) | ( n5089 & n5090 ) ;
  assign n5079 = ( n4686 & n4807 ) | ( n4686 & n4942 ) | ( n4807 & n4942 ) ;
  assign n5078 = ( n4686 & ~n4807 ) | ( n4686 & n4942 ) | ( ~n4807 & n4942 ) ;
  assign n5080 = ( n4807 & ~n5079 ) | ( n4807 & n5078 ) | ( ~n5079 & n5078 ) ;
  assign n5095 = ~n523 & n1875 ;
  assign n5092 = n1671 | n4430 ;
  assign n5093 = n1748 | n3939 ;
  assign n5094 = n5092 &  n5093 ;
  assign n5096 = ( n523 & n5095 ) | ( n523 & n5094 ) | ( n5095 & n5094 ) ;
  assign n5097 = n601 | n4580 ;
  assign n5098 = n5096 &  n5097 ;
  assign n5099 = x29 &  n5098 ;
  assign n5100 = x29 | n5098 ;
  assign n5101 = ~n5099 & n5100 ;
  assign n5102 = ( n5091 & ~n5080 ) | ( n5091 & n5101 ) | ( ~n5080 & n5101 ) ;
  assign n5103 = ( n4767 & ~n4756 ) | ( n4767 & n4943 ) | ( ~n4756 & n4943 ) ;
  assign n5104 = ( n4756 & ~n4943 ) | ( n4756 & n4767 ) | ( ~n4943 & n4767 ) ;
  assign n5105 = ( n5103 & ~n4767 ) | ( n5103 & n5104 ) | ( ~n4767 & n5104 ) ;
  assign n5106 = n5102 | n5105 ;
  assign n5110 = ~n1566 & n4430 ;
  assign n5107 = n523 | n1748 ;
  assign n5108 = n1671 | n3939 ;
  assign n5109 = n5107 &  n5108 ;
  assign n5111 = ( n1566 & n5110 ) | ( n1566 & n5109 ) | ( n5110 & n5109 ) ;
  assign n5112 = n601 | n4597 ;
  assign n5113 = n5111 &  n5112 ;
  assign n5114 = ( x29 & ~n5113 ) | ( x29 & 1'b0 ) | ( ~n5113 & 1'b0 ) ;
  assign n5115 = n5102 &  n5105 ;
  assign n5116 = ( n5113 & ~x29 ) | ( n5113 & n5115 ) | ( ~x29 & n5115 ) ;
  assign n5117 = ( n5106 & n5114 ) | ( n5106 & n5116 ) | ( n5114 & n5116 ) ;
  assign n5118 = n4945 | n4954 ;
  assign n5119 = ( n4952 & ~x29 ) | ( n4952 & n5118 ) | ( ~x29 & n5118 ) ;
  assign n5120 = ( x29 & ~n5118 ) | ( x29 & n4952 ) | ( ~n5118 & n4952 ) ;
  assign n5121 = ( n5119 & ~n4952 ) | ( n5119 & n5120 ) | ( ~n4952 & n5120 ) ;
  assign n5123 = n1151 | n4962 ;
  assign n5124 = n1378 | n4482 ;
  assign n5125 = n5123 &  n5124 ;
  assign n5126 = n1267 &  n4495 ;
  assign n5127 = ( n5125 & ~n1267 ) | ( n5125 & n5126 ) | ( ~n1267 & n5126 ) ;
  assign n5128 = ( n4061 & ~n4478 ) | ( n4061 & 1'b0 ) | ( ~n4478 & 1'b0 ) ;
  assign n5129 = ( n5127 & ~n5128 ) | ( n5127 & 1'b0 ) | ( ~n5128 & 1'b0 ) ;
  assign n5131 = x26 | n5129 ;
  assign n5132 = x26 &  n5129 ;
  assign n5133 = ( n5131 & ~n5132 ) | ( n5131 & 1'b0 ) | ( ~n5132 & 1'b0 ) ;
  assign n5134 = ( n5117 & ~n5121 ) | ( n5117 & n5133 ) | ( ~n5121 & n5133 ) ;
  assign n5076 = ( x26 & n5055 ) | ( x26 & n5059 ) | ( n5055 & n5059 ) ;
  assign n5077 = ( n5055 & ~n5076 ) | ( n5055 & n5060 ) | ( ~n5076 & n5060 ) ;
  assign n5139 = ~n946 & n5010 ;
  assign n5135 = ~n5005 |  n5008 ;
  assign n5136 = n702 | n5135 ;
  assign n5137 = n863 | n5067 ;
  assign n5138 = n5136 &  n5137 ;
  assign n5140 = ( n946 & n5139 ) | ( n946 & n5138 ) | ( n5139 & n5138 ) ;
  assign n5141 = n3650 | n5012 ;
  assign n5142 = n5140 &  n5141 ;
  assign n5143 = x23 &  n5142 ;
  assign n5144 = x23 | n5142 ;
  assign n5145 = ~n5143 & n5144 ;
  assign n5146 = ( n5134 & ~n5077 ) | ( n5134 & n5145 ) | ( ~n5077 & n5145 ) ;
  assign n5150 = ~n863 & n5010 ;
  assign n5147 = n599 | n5135 ;
  assign n5148 = n702 | n5067 ;
  assign n5149 = n5147 &  n5148 ;
  assign n5151 = ( n863 & n5150 ) | ( n863 & n5149 ) | ( n5150 & n5149 ) ;
  assign n5152 = ( n5012 & ~n4452 ) | ( n5012 & n5151 ) | ( ~n4452 & n5151 ) ;
  assign n5153 = ~n5012 & n5152 ;
  assign n5154 = ( x23 & ~n5151 ) | ( x23 & n5153 ) | ( ~n5151 & n5153 ) ;
  assign n5155 = ( n5151 & ~x23 ) | ( n5151 & n5153 ) | ( ~x23 & n5153 ) ;
  assign n5156 = ( n5154 & ~n5153 ) | ( n5154 & n5155 ) | ( ~n5153 & n5155 ) ;
  assign n5157 = ( n5023 & ~n5033 ) | ( n5023 & n5061 ) | ( ~n5033 & n5061 ) ;
  assign n5158 = ( n5033 & ~n5062 ) | ( n5033 & n5157 ) | ( ~n5062 & n5157 ) ;
  assign n5159 = ( n5146 & n5156 ) | ( n5146 & n5158 ) | ( n5156 & n5158 ) ;
  assign n5160 = ~x23 & n5062 ;
  assign n5161 = x23 | n5062 ;
  assign n5162 = ( n5160 & ~n5062 ) | ( n5160 & n5161 ) | ( ~n5062 & n5161 ) ;
  assign n5163 = ( n5071 & ~n5065 ) | ( n5071 & n5162 ) | ( ~n5065 & n5162 ) ;
  assign n5164 = ( n5065 & ~n5071 ) | ( n5065 & n5162 ) | ( ~n5071 & n5162 ) ;
  assign n5165 = ( n5163 & ~n5162 ) | ( n5163 & n5164 ) | ( ~n5162 & n5164 ) ;
  assign n5166 = ( n5156 & ~n5146 ) | ( n5156 & n5158 ) | ( ~n5146 & n5158 ) ;
  assign n5167 = ( n5146 & ~n5158 ) | ( n5146 & n5156 ) | ( ~n5158 & n5156 ) ;
  assign n5168 = ( n5166 & ~n5156 ) | ( n5166 & n5167 ) | ( ~n5156 & n5167 ) ;
  assign n5321 = ~n946 & n5067 ;
  assign n5318 = n863 | n5135 ;
  assign n5319 = n1043 | n5010 ;
  assign n5320 = n5318 &  n5319 ;
  assign n5322 = ( n946 & n5321 ) | ( n946 & n5320 ) | ( n5321 & n5320 ) ;
  assign n5323 = n3914 | n5012 ;
  assign n5324 = n5322 &  n5323 ;
  assign n5325 = ( x23 & ~n5324 ) | ( x23 & 1'b0 ) | ( ~n5324 & 1'b0 ) ;
  assign n5122 = ~n5117 & n5121 ;
  assign n5130 = ( n5117 & ~n5121 ) | ( n5117 & 1'b0 ) | ( ~n5121 & 1'b0 ) ;
  assign n5169 = n5122 | n5130 ;
  assign n5170 = ( x26 & ~n5169 ) | ( x26 & n5129 ) | ( ~n5169 & n5129 ) ;
  assign n5171 = ( n5129 & ~x26 ) | ( n5129 & n5169 ) | ( ~x26 & n5169 ) ;
  assign n5172 = ( n5170 & ~n5129 ) | ( n5170 & n5171 ) | ( ~n5129 & n5171 ) ;
  assign n5173 = ( n5106 & ~n5115 ) | ( n5106 & 1'b0 ) | ( ~n5115 & 1'b0 ) ;
  assign n5175 = ( x29 & n5113 ) | ( x29 & n5173 ) | ( n5113 & n5173 ) ;
  assign n5174 = ( x29 & ~n5113 ) | ( x29 & n5173 ) | ( ~n5113 & n5173 ) ;
  assign n5176 = ( n5113 & ~n5175 ) | ( n5113 & n5174 ) | ( ~n5175 & n5174 ) ;
  assign n5177 = ( n1483 & ~n4482 ) | ( n1483 & 1'b0 ) | ( ~n4482 & 1'b0 ) ;
  assign n5178 = n1378 | n4495 ;
  assign n5179 = ~n5177 & n5178 ;
  assign n5180 = n1267 &  n4962 ;
  assign n5181 = ( n5179 & ~n1267 ) | ( n5179 & n5180 ) | ( ~n1267 & n5180 ) ;
  assign n5182 = ( n4422 & ~n5181 ) | ( n4422 & n4478 ) | ( ~n5181 & n4478 ) ;
  assign n5183 = ( n4422 & ~n5182 ) | ( n4422 & 1'b0 ) | ( ~n5182 & 1'b0 ) ;
  assign n5184 = ( x26 & ~n5181 ) | ( x26 & n5183 ) | ( ~n5181 & n5183 ) ;
  assign n5185 = ( n5181 & ~x26 ) | ( n5181 & n5183 ) | ( ~x26 & n5183 ) ;
  assign n5186 = ( n5184 & ~n5183 ) | ( n5184 & n5185 ) | ( ~n5183 & n5185 ) ;
  assign n5305 = n1378 | n4962 ;
  assign n5306 = n1566 | n4482 ;
  assign n5307 = n5305 &  n5306 ;
  assign n5308 = n1483 &  n4495 ;
  assign n5309 = ( n5307 & ~n1483 ) | ( n5307 & n5308 ) | ( ~n1483 & n5308 ) ;
  assign n5310 = ~n4478 & n5038 ;
  assign n5311 = ( n5309 & ~n5310 ) | ( n5309 & 1'b0 ) | ( ~n5310 & 1'b0 ) ;
  assign n5312 = ( x26 & ~n5311 ) | ( x26 & 1'b0 ) | ( ~n5311 & 1'b0 ) ;
  assign n5187 = ( n5080 & n5091 ) | ( n5080 & n5101 ) | ( n5091 & n5101 ) ;
  assign n5188 = ( n5080 & ~n5091 ) | ( n5080 & n5101 ) | ( ~n5091 & n5101 ) ;
  assign n5189 = ( n5091 & ~n5187 ) | ( n5091 & n5188 ) | ( ~n5187 & n5188 ) ;
  assign n5298 = ~n601 & n4743 ;
  assign n5293 = n523 | n1940 ;
  assign n5294 = n1875 | n3939 ;
  assign n5295 = n5293 &  n5294 ;
  assign n5296 = ~n1748 & n4430 ;
  assign n5297 = ( n1748 & n5295 ) | ( n1748 & n5296 ) | ( n5295 & n5296 ) ;
  assign n5299 = ( n601 & n5298 ) | ( n601 & n5297 ) | ( n5298 & n5297 ) ;
  assign n5300 = ~x29 & n5299 ;
  assign n5190 = ( n4807 & ~n4928 ) | ( n4807 & n4941 ) | ( ~n4928 & n4941 ) ;
  assign n5191 = ( n4807 & ~n4941 ) | ( n4807 & n4928 ) | ( ~n4941 & n4928 ) ;
  assign n5192 = ( n5190 & ~n4807 ) | ( n5190 & n5191 ) | ( ~n4807 & n5191 ) ;
  assign n5193 = ( x14 & ~n4858 ) | ( x14 & n4927 ) | ( ~n4858 & n4927 ) ;
  assign n5194 = ( n4858 & ~n4928 ) | ( n4858 & n5193 ) | ( ~n4928 & n5193 ) ;
  assign n5195 = n117 | n1305 ;
  assign n5196 = n229 | n5195 ;
  assign n5197 = ( n220 & ~n5196 ) | ( n220 & n1047 ) | ( ~n5196 & n1047 ) ;
  assign n5198 = ( n1489 & n5196 ) | ( n1489 & n5197 ) | ( n5196 & n5197 ) ;
  assign n5199 = ( n1489 & ~n5198 ) | ( n1489 & 1'b0 ) | ( ~n5198 & 1'b0 ) ;
  assign n5200 = ( n1883 & ~n1107 ) | ( n1883 & n5199 ) | ( ~n1107 & n5199 ) ;
  assign n5201 = ~n1883 & n5200 ;
  assign n5202 = ( n4090 & n665 ) | ( n4090 & n5201 ) | ( n665 & n5201 ) ;
  assign n5203 = ~n665 & n5202 ;
  assign n5204 = ( n2702 & ~n865 ) | ( n2702 & n5203 ) | ( ~n865 & n5203 ) ;
  assign n5205 = ~n2702 & n5204 ;
  assign n5206 = ( n493 & ~n383 ) | ( n493 & n5205 ) | ( ~n383 & n5205 ) ;
  assign n5207 = ~n493 & n5206 ;
  assign n5208 = ( n255 & ~n403 ) | ( n255 & n5207 ) | ( ~n403 & n5207 ) ;
  assign n5209 = ~n255 & n5208 ;
  assign n5210 = ~n167 & n5209 ;
  assign n5221 = n3370 | n3586 ;
  assign n5217 = ~n125 & n644 ;
  assign n5218 = ( n405 & ~n5217 ) | ( n405 & n623 ) | ( ~n5217 & n623 ) ;
  assign n5219 = ( n623 & ~n5218 ) | ( n623 & 1'b0 ) | ( ~n5218 & 1'b0 ) ;
  assign n5220 = ~n353 & n5219 ;
  assign n5222 = ( n779 & ~n5221 ) | ( n779 & n5220 ) | ( ~n5221 & n5220 ) ;
  assign n5223 = ~n779 & n5222 ;
  assign n5224 = ( n477 & ~n425 ) | ( n477 & n5223 ) | ( ~n425 & n5223 ) ;
  assign n5225 = ~n477 & n5224 ;
  assign n5226 = ( n162 & ~n737 ) | ( n162 & n5225 ) | ( ~n737 & n5225 ) ;
  assign n5227 = ~n162 & n5226 ;
  assign n5228 = ~n574 & n5227 ;
  assign n5229 = n555 | n3890 ;
  assign n5230 = n348 | n5229 ;
  assign n5231 = ( n3875 & ~n1513 ) | ( n3875 & n5230 ) | ( ~n1513 & n5230 ) ;
  assign n5232 = n1513 | n5231 ;
  assign n5233 = n1585 | n5232 ;
  assign n5234 = ( n3777 & ~n3979 ) | ( n3777 & n5233 ) | ( ~n3979 & n5233 ) ;
  assign n5235 = ( n3979 & ~n81 ) | ( n3979 & n5234 ) | ( ~n81 & n5234 ) ;
  assign n5236 = n81 | n5235 ;
  assign n5237 = ( n5236 & ~n335 ) | ( n5236 & n1380 ) | ( ~n335 & n1380 ) ;
  assign n5238 = n335 | n5237 ;
  assign n5239 = ( n814 & ~n362 ) | ( n814 & n5238 ) | ( ~n362 & n5238 ) ;
  assign n5240 = n362 | n5239 ;
  assign n5241 = ( n257 & ~n193 ) | ( n257 & n5240 ) | ( ~n193 & n5240 ) ;
  assign n5242 = n193 | n5241 ;
  assign n5243 = ( n451 & ~n796 ) | ( n451 & n5242 ) | ( ~n796 & n5242 ) ;
  assign n5244 = n796 | n5243 ;
  assign n5245 = ( n266 & n343 ) | ( n266 & n5244 ) | ( n343 & n5244 ) ;
  assign n5246 = ( n343 & ~n5245 ) | ( n343 & 1'b0 ) | ( ~n5245 & 1'b0 ) ;
  assign n5247 = n139 | n206 ;
  assign n5248 = ( n2891 & ~n5247 ) | ( n2891 & 1'b0 ) | ( ~n5247 & 1'b0 ) ;
  assign n5249 = ( n5246 & ~n5228 ) | ( n5246 & n5248 ) | ( ~n5228 & n5248 ) ;
  assign n5250 = ( n1224 & n5228 ) | ( n1224 & n5249 ) | ( n5228 & n5249 ) ;
  assign n5251 = ~n1224 & n5250 ;
  assign n5211 = n259 | n4228 ;
  assign n5212 = ( n797 & ~n275 ) | ( n797 & n5211 ) | ( ~n275 & n5211 ) ;
  assign n5213 = n275 | n5212 ;
  assign n5214 = ( n239 & ~n602 ) | ( n239 & n5213 ) | ( ~n602 & n5213 ) ;
  assign n5215 = n602 | n5214 ;
  assign n5216 = n646 | n5215 ;
  assign n5252 = ( n5210 & ~n5251 ) | ( n5210 & n5216 ) | ( ~n5251 & n5216 ) ;
  assign n5253 = ( n1278 & ~n5252 ) | ( n1278 & n5210 ) | ( ~n5252 & n5210 ) ;
  assign n5254 = ~n1278 & n5253 ;
  assign n5255 = ( n5254 & ~n102 ) | ( n5254 & n1580 ) | ( ~n102 & n1580 ) ;
  assign n5256 = ( n5255 & ~n1580 ) | ( n5255 & 1'b0 ) | ( ~n1580 & 1'b0 ) ;
  assign n5257 = ( n230 & ~n235 ) | ( n230 & n5256 ) | ( ~n235 & n5256 ) ;
  assign n5258 = ~n230 & n5257 ;
  assign n5259 = ( n74 & ~n136 ) | ( n74 & n5258 ) | ( ~n136 & n5258 ) ;
  assign n5260 = ~n74 & n5259 ;
  assign n5261 = ( n627 & ~n279 ) | ( n627 & n5260 ) | ( ~n279 & n5260 ) ;
  assign n5262 = ~n627 & n5261 ;
  assign n5263 = ~n141 & n5262 ;
  assign n5264 = n2178 | n2296 ;
  assign n5265 = ( n2178 & ~n2296 ) | ( n2178 & 1'b0 ) | ( ~n2296 & 1'b0 ) ;
  assign n5266 = ( n5264 & ~n2178 ) | ( n5264 & n5265 ) | ( ~n2178 & n5265 ) ;
  assign n5267 = ~n3619 & n5266 ;
  assign n5268 = ( n3619 & ~n5266 ) | ( n3619 & 1'b0 ) | ( ~n5266 & 1'b0 ) ;
  assign n5269 = n5267 | n5268 ;
  assign n5270 = n3644 | n5269 ;
  assign n5271 = ~n2392 & n3652 ;
  assign n5272 = ~n2296 & n3657 ;
  assign n5273 = n5271 | n5272 ;
  assign n5274 = ~n2178 & n3653 ;
  assign n5275 = ( n2178 & ~n5273 ) | ( n2178 & n5274 ) | ( ~n5273 & n5274 ) ;
  assign n5276 = n5270 &  n5275 ;
  assign n5277 = ( n5263 & ~n4858 ) | ( n5263 & n5276 ) | ( ~n4858 & n5276 ) ;
  assign n5278 = n2127 | n2178 ;
  assign n5279 = ( n2127 & ~n2178 ) | ( n2127 & 1'b0 ) | ( ~n2178 & 1'b0 ) ;
  assign n5280 = ( n5278 & ~n2127 ) | ( n5278 & n5279 ) | ( ~n2127 & n5279 ) ;
  assign n5281 = ~n3620 & n5280 ;
  assign n5282 = ( n3620 & ~n5280 ) | ( n3620 & 1'b0 ) | ( ~n5280 & 1'b0 ) ;
  assign n5283 = n5281 | n5282 ;
  assign n5284 = n3644 | n5283 ;
  assign n5285 = n2296 &  n3652 ;
  assign n5286 = n2127 | n3653 ;
  assign n5287 = ~n2178 & n3657 ;
  assign n5288 = ( n5286 & ~n5287 ) | ( n5286 & 1'b0 ) | ( ~n5287 & 1'b0 ) ;
  assign n5289 = ( n5285 & ~n3652 ) | ( n5285 & n5288 ) | ( ~n3652 & n5288 ) ;
  assign n5290 = n5284 &  n5289 ;
  assign n5291 = ( n5194 & n5277 ) | ( n5194 & n5290 ) | ( n5277 & n5290 ) ;
  assign n5292 = ( n5192 & ~n5291 ) | ( n5192 & 1'b0 ) | ( ~n5291 & 1'b0 ) ;
  assign n5301 = ~n5192 & n5291 ;
  assign n5302 = ( x29 & ~n5299 ) | ( x29 & n5301 ) | ( ~n5299 & n5301 ) ;
  assign n5303 = ( n5300 & ~n5292 ) | ( n5300 & n5302 ) | ( ~n5292 & n5302 ) ;
  assign n5304 = ( n5189 & ~n5303 ) | ( n5189 & 1'b0 ) | ( ~n5303 & 1'b0 ) ;
  assign n5313 = ~n5189 & n5303 ;
  assign n5314 = ( n5311 & ~x26 ) | ( n5311 & n5313 ) | ( ~x26 & n5313 ) ;
  assign n5315 = ( n5312 & ~n5304 ) | ( n5312 & n5314 ) | ( ~n5304 & n5314 ) ;
  assign n5316 = ( n5176 & n5186 ) | ( n5176 & n5315 ) | ( n5186 & n5315 ) ;
  assign n5317 = ( n5172 & ~n5316 ) | ( n5172 & 1'b0 ) | ( ~n5316 & 1'b0 ) ;
  assign n5326 = ~n5172 & n5316 ;
  assign n5327 = ( n5324 & ~x23 ) | ( n5324 & n5326 ) | ( ~x23 & n5326 ) ;
  assign n5328 = ( n5325 & ~n5317 ) | ( n5325 & n5327 ) | ( ~n5317 & n5327 ) ;
  assign n5347 = ( n5077 & n5134 ) | ( n5077 & n5145 ) | ( n5134 & n5145 ) ;
  assign n5348 = ( n5077 & ~n5134 ) | ( n5077 & n5145 ) | ( ~n5134 & n5145 ) ;
  assign n5349 = ( n5134 & ~n5347 ) | ( n5134 & n5348 ) | ( ~n5347 & n5348 ) ;
  assign n5329 = ~x18 & x19 ;
  assign n5330 = ( x18 & ~x19 ) | ( x18 & 1'b0 ) | ( ~x19 & 1'b0 ) ;
  assign n5331 = n5329 | n5330 ;
  assign n5335 = ( x17 & ~x18 ) | ( x17 & 1'b0 ) | ( ~x18 & 1'b0 ) ;
  assign n5336 = ~x17 & x18 ;
  assign n5337 = n5335 | n5336 ;
  assign n5332 = ( x19 & ~x20 ) | ( x19 & 1'b0 ) | ( ~x20 & 1'b0 ) ;
  assign n5333 = ~x19 & x20 ;
  assign n5334 = n5332 | n5333 ;
  assign n5338 = ( n5331 & ~n5337 ) | ( n5331 & n5334 ) | ( ~n5337 & n5334 ) ;
  assign n5339 = ~n5331 & n5338 ;
  assign n5340 = ~n599 & n5339 ;
  assign n5341 = ~n5334 | ~n5337 ;
  assign n5342 = ( n5340 & ~n3637 ) | ( n5340 & n5341 ) | ( ~n3637 & n5341 ) ;
  assign n5343 = n3637 | n5342 ;
  assign n5344 = ( x20 & ~n5340 ) | ( x20 & n5343 ) | ( ~n5340 & n5343 ) ;
  assign n5345 = ( n5340 & ~x20 ) | ( n5340 & n5343 ) | ( ~x20 & n5343 ) ;
  assign n5346 = ( n5344 & ~n5343 ) | ( n5344 & n5345 ) | ( ~n5343 & n5345 ) ;
  assign n5350 = ( n5328 & ~n5349 ) | ( n5328 & n5346 ) | ( ~n5349 & n5346 ) ;
  assign n5760 = ~n702 & n5339 ;
  assign n5761 = ~n5331 |  n5337 ;
  assign n5762 = n599 | n5761 ;
  assign n5763 = ~n5760 & n5762 ;
  assign n5764 = ( n3937 & ~n5341 ) | ( n3937 & 1'b0 ) | ( ~n5341 & 1'b0 ) ;
  assign n5765 = ( n5763 & ~n5764 ) | ( n5763 & 1'b0 ) | ( ~n5764 & 1'b0 ) ;
  assign n5766 = ( x20 & ~n5765 ) | ( x20 & 1'b0 ) | ( ~n5765 & 1'b0 ) ;
  assign n5354 = n5317 | n5326 ;
  assign n5355 = ( x23 & ~n5354 ) | ( x23 & n5324 ) | ( ~n5354 & n5324 ) ;
  assign n5356 = ( n5324 & ~x23 ) | ( n5324 & n5354 ) | ( ~x23 & n5354 ) ;
  assign n5357 = ( n5355 & ~n5324 ) | ( n5355 & n5356 ) | ( ~n5324 & n5356 ) ;
  assign n5361 = ~n946 & n5135 ;
  assign n5358 = n1151 | n5010 ;
  assign n5359 = n1043 | n5067 ;
  assign n5360 = n5358 &  n5359 ;
  assign n5362 = ( n946 & n5361 ) | ( n946 & n5360 ) | ( n5361 & n5360 ) ;
  assign n5363 = n4038 | n5012 ;
  assign n5364 = n5362 &  n5363 ;
  assign n5365 = x23 &  n5364 ;
  assign n5366 = x23 | n5364 ;
  assign n5367 = ~n5365 & n5366 ;
  assign n5368 = ( n5186 & ~n5176 ) | ( n5186 & n5315 ) | ( ~n5176 & n5315 ) ;
  assign n5369 = ( n5176 & ~n5315 ) | ( n5176 & n5186 ) | ( ~n5315 & n5186 ) ;
  assign n5370 = ( n5368 & ~n5186 ) | ( n5368 & n5369 ) | ( ~n5186 & n5369 ) ;
  assign n5747 = n1043 | n5135 ;
  assign n5748 = n1151 | n5067 ;
  assign n5749 = n5747 &  n5748 ;
  assign n5750 = n1267 &  n5010 ;
  assign n5751 = ( n5749 & ~n1267 ) | ( n5749 & n5750 ) | ( ~n1267 & n5750 ) ;
  assign n5752 = n3952 | n5012 ;
  assign n5753 = n5751 &  n5752 ;
  assign n5754 = ( x23 & ~n5753 ) | ( x23 & 1'b0 ) | ( ~n5753 & 1'b0 ) ;
  assign n5371 = n5304 | n5313 ;
  assign n5372 = ( x26 & ~n5371 ) | ( x26 & n5311 ) | ( ~n5371 & n5311 ) ;
  assign n5373 = ( n5311 & ~x26 ) | ( n5311 & n5371 ) | ( ~x26 & n5371 ) ;
  assign n5374 = ( n5372 & ~n5311 ) | ( n5372 & n5373 ) | ( ~n5311 & n5373 ) ;
  assign n5735 = n1671 | n4482 ;
  assign n5736 = n1566 | n4495 ;
  assign n5737 = n5735 &  n5736 ;
  assign n5738 = n1483 &  n4962 ;
  assign n5739 = ( n5737 & ~n1483 ) | ( n5737 & n5738 ) | ( ~n1483 & n5738 ) ;
  assign n5740 = ( n4274 & ~n4478 ) | ( n4274 & 1'b0 ) | ( ~n4478 & 1'b0 ) ;
  assign n5741 = ( n5739 & ~n5740 ) | ( n5739 & 1'b0 ) | ( ~n5740 & 1'b0 ) ;
  assign n5742 = ( x26 & ~n5741 ) | ( x26 & 1'b0 ) | ( ~n5741 & 1'b0 ) ;
  assign n5378 = ~n1875 & n4430 ;
  assign n5375 = n523 | n2022 ;
  assign n5376 = n1940 | n3939 ;
  assign n5377 = n5375 &  n5376 ;
  assign n5379 = ( n1875 & n5378 ) | ( n1875 & n5377 ) | ( n5378 & n5377 ) ;
  assign n5380 = ~n3623 & n4761 ;
  assign n5381 = n4762 | n5380 ;
  assign n5382 = n601 | n5381 ;
  assign n5383 = n5379 &  n5382 ;
  assign n5384 = x29 &  n5383 ;
  assign n5385 = x29 | n5383 ;
  assign n5386 = ~n5384 & n5385 ;
  assign n5387 = ( n5194 & ~n5277 ) | ( n5194 & n5290 ) | ( ~n5277 & n5290 ) ;
  assign n5388 = ( n5194 & ~n5290 ) | ( n5194 & n5277 ) | ( ~n5290 & n5277 ) ;
  assign n5389 = ( n5387 & ~n5194 ) | ( n5387 & n5388 ) | ( ~n5194 & n5388 ) ;
  assign n5392 = n408 | n2610 ;
  assign n5393 = ( n49 & ~n273 ) | ( n49 & n5392 ) | ( ~n273 & n5392 ) ;
  assign n5394 = n273 | n5393 ;
  assign n5395 = ( n252 & ~n300 ) | ( n252 & n5394 ) | ( ~n300 & n5394 ) ;
  assign n5396 = n300 | n5395 ;
  assign n5397 = n617 | n5396 ;
  assign n5398 = n454 | n485 ;
  assign n5399 = n88 | n5398 ;
  assign n5400 = n2264 | n2735 ;
  assign n5401 = ( n5399 & ~n1828 ) | ( n5399 & n5400 ) | ( ~n1828 & n5400 ) ;
  assign n5402 = n1828 | n5401 ;
  assign n5403 = ( n5397 & ~n414 ) | ( n5397 & n5402 ) | ( ~n414 & n5402 ) ;
  assign n5404 = n414 | n5403 ;
  assign n5405 = ( n275 & ~n280 ) | ( n275 & n5404 ) | ( ~n280 & n5404 ) ;
  assign n5406 = n280 | n5405 ;
  assign n5407 = ( n793 & ~n372 ) | ( n793 & n5406 ) | ( ~n372 & n5406 ) ;
  assign n5408 = n372 | n5407 ;
  assign n5409 = ( n132 & ~n737 ) | ( n132 & n5408 ) | ( ~n737 & n5408 ) ;
  assign n5410 = n737 | n5409 ;
  assign n5411 = ( n384 & ~n431 ) | ( n384 & n5410 ) | ( ~n431 & n5410 ) ;
  assign n5412 = n431 | n5411 ;
  assign n5413 = n239 | n718 ;
  assign n5414 = ( n1130 & ~n4859 ) | ( n1130 & n5413 ) | ( ~n4859 & n5413 ) ;
  assign n5415 = ( n4859 & ~n3328 ) | ( n4859 & n5414 ) | ( ~n3328 & n5414 ) ;
  assign n5416 = n3328 | n5415 ;
  assign n5417 = ( n884 & ~n713 ) | ( n884 & n5416 ) | ( ~n713 & n5416 ) ;
  assign n5418 = n713 | n5417 ;
  assign n5419 = ( n70 & ~n101 ) | ( n70 & n5418 ) | ( ~n101 & n5418 ) ;
  assign n5420 = n101 | n5419 ;
  assign n5421 = ( n403 & ~n909 ) | ( n403 & n5420 ) | ( ~n909 & n5420 ) ;
  assign n5422 = n909 | n5421 ;
  assign n5423 = ( n336 & ~n342 ) | ( n336 & n5422 ) | ( ~n342 & n5422 ) ;
  assign n5424 = n342 | n5423 ;
  assign n5425 = n130 | n812 ;
  assign n5426 = n279 | n5425 ;
  assign n5427 = n188 | n478 ;
  assign n5428 = n86 | n5427 ;
  assign n5429 = ( n195 & ~n675 ) | ( n195 & n3213 ) | ( ~n675 & n3213 ) ;
  assign n5430 = n675 | n5429 ;
  assign n5431 = n1829 | n5430 ;
  assign n5432 = ( n5428 & ~n5426 ) | ( n5428 & n5431 ) | ( ~n5426 & n5431 ) ;
  assign n5433 = ( n5426 & ~n3663 ) | ( n5426 & n5432 ) | ( ~n3663 & n5432 ) ;
  assign n5434 = n3663 | n5433 ;
  assign n5435 = ( n4839 & ~n2514 ) | ( n4839 & n5434 ) | ( ~n2514 & n5434 ) ;
  assign n5436 = n2514 | n5435 ;
  assign n5437 = ( n1453 & ~n5436 ) | ( n1453 & 1'b0 ) | ( ~n5436 & 1'b0 ) ;
  assign n5438 = ( n5412 & ~n5424 ) | ( n5412 & n5437 ) | ( ~n5424 & n5437 ) ;
  assign n5439 = ( n258 & ~n5412 ) | ( n258 & n5438 ) | ( ~n5412 & n5438 ) ;
  assign n5440 = ~n258 & n5439 ;
  assign n5441 = ( n169 & ~n52 ) | ( n169 & n5440 ) | ( ~n52 & n5440 ) ;
  assign n5442 = ~n169 & n5441 ;
  assign n5443 = ~n351 & n5442 ;
  assign n5444 = n415 | n789 ;
  assign n5445 = ( n351 & ~n279 ) | ( n351 & n5444 ) | ( ~n279 & n5444 ) ;
  assign n5446 = n279 | n5445 ;
  assign n5447 = n3395 | n4228 ;
  assign n5448 = ( n5446 & ~n1678 ) | ( n5446 & n5447 ) | ( ~n1678 & n5447 ) ;
  assign n5449 = n1678 | n5448 ;
  assign n5450 = ( n5449 & ~n187 ) | ( n5449 & n1884 ) | ( ~n187 & n1884 ) ;
  assign n5451 = n187 | n5450 ;
  assign n5452 = ( n451 & ~n299 ) | ( n451 & n5451 ) | ( ~n299 & n5451 ) ;
  assign n5453 = n299 | n5452 ;
  assign n5455 = n194 | n800 ;
  assign n5456 = n372 | n5455 ;
  assign n5454 = n236 | n531 ;
  assign n5457 = ( n2188 & n5456 ) | ( n2188 & n5454 ) | ( n5456 & n5454 ) ;
  assign n5458 = ( n2188 & ~n5457 ) | ( n2188 & 1'b0 ) | ( ~n5457 & 1'b0 ) ;
  assign n5459 = ( n1710 & ~n5453 ) | ( n1710 & n5458 ) | ( ~n5453 & n5458 ) ;
  assign n5460 = ~n1710 & n5459 ;
  assign n5461 = ( n2576 & ~n2577 ) | ( n2576 & n5460 ) | ( ~n2577 & n5460 ) ;
  assign n5462 = ~n2576 & n5461 ;
  assign n5463 = ( n673 & ~n479 ) | ( n673 & n5462 ) | ( ~n479 & n5462 ) ;
  assign n5464 = ~n673 & n5463 ;
  assign n5465 = ( n493 & ~n259 ) | ( n493 & n5464 ) | ( ~n259 & n5464 ) ;
  assign n5466 = ~n493 & n5465 ;
  assign n5467 = ( n429 & ~n359 ) | ( n429 & n5466 ) | ( ~n359 & n5466 ) ;
  assign n5468 = ~n429 & n5467 ;
  assign n5469 = ( n253 & ~n221 ) | ( n253 & n5468 ) | ( ~n221 & n5468 ) ;
  assign n5470 = ~n253 & n5469 ;
  assign n5471 = ( n617 & ~n571 ) | ( n617 & n5470 ) | ( ~n571 & n5470 ) ;
  assign n5472 = ~n617 & n5471 ;
  assign n5473 = n1963 | n2061 ;
  assign n5474 = ( n1796 & ~n5473 ) | ( n1796 & n4102 ) | ( ~n5473 & n4102 ) ;
  assign n5475 = ~n1796 & n5474 ;
  assign n5476 = ( n4290 & n1828 ) | ( n4290 & n5475 ) | ( n1828 & n5475 ) ;
  assign n5477 = ~n1828 & n5476 ;
  assign n5478 = ( n575 & ~n3741 ) | ( n575 & n5477 ) | ( ~n3741 & n5477 ) ;
  assign n5479 = ~n575 & n5478 ;
  assign n5480 = ( n5424 & n5472 ) | ( n5424 & n5479 ) | ( n5472 & n5479 ) ;
  assign n5481 = ~n5424 & n5480 ;
  assign n5482 = ( n62 & ~n1454 ) | ( n62 & n5481 ) | ( ~n1454 & n5481 ) ;
  assign n5483 = ~n62 & n5482 ;
  assign n5484 = ( n208 & ~n409 ) | ( n208 & n5483 ) | ( ~n409 & n5483 ) ;
  assign n5485 = ~n208 & n5484 ;
  assign n5486 = ( n418 & ~n272 ) | ( n418 & n5485 ) | ( ~n272 & n5485 ) ;
  assign n5487 = ~n418 & n5486 ;
  assign n5488 = ( n255 & ~n411 ) | ( n255 & n5487 ) | ( ~n411 & n5487 ) ;
  assign n5489 = ~n255 & n5488 ;
  assign n5490 = ( n334 & ~n80 ) | ( n334 & n5489 ) | ( ~n80 & n5489 ) ;
  assign n5491 = ~n334 & n5490 ;
  assign n5492 = ( n5491 & ~n432 ) | ( n5491 & n663 ) | ( ~n432 & n663 ) ;
  assign n5493 = ( n5492 & ~n663 ) | ( n5492 & 1'b0 ) | ( ~n663 & 1'b0 ) ;
  assign n5494 = ( x11 & n5443 ) | ( x11 & n5493 ) | ( n5443 & n5493 ) ;
  assign n5495 = n2296 | n2392 ;
  assign n5496 = ( n2296 & ~n2392 ) | ( n2296 & 1'b0 ) | ( ~n2392 & 1'b0 ) ;
  assign n5497 = ( n5495 & ~n2296 ) | ( n5495 & n5496 ) | ( ~n2296 & n5496 ) ;
  assign n5498 = ~n3618 & n5497 ;
  assign n5499 = ( n3618 & ~n5497 ) | ( n3618 & 1'b0 ) | ( ~n5497 & 1'b0 ) ;
  assign n5500 = n5498 | n5499 ;
  assign n5501 = n3644 | n5500 ;
  assign n5502 = ~n2483 & n3652 ;
  assign n5503 = ~n2392 & n3657 ;
  assign n5504 = n5502 | n5503 ;
  assign n5505 = ~n2296 & n3653 ;
  assign n5506 = ( n2296 & ~n5504 ) | ( n2296 & n5505 ) | ( ~n5504 & n5505 ) ;
  assign n5507 = n5501 &  n5506 ;
  assign n5508 = ( n5494 & ~n4858 ) | ( n5494 & n5507 ) | ( ~n4858 & n5507 ) ;
  assign n5390 = ( n4858 & ~n5263 ) | ( n4858 & n5276 ) | ( ~n5263 & n5276 ) ;
  assign n5391 = ( n5277 & ~n5276 ) | ( n5277 & n5390 ) | ( ~n5276 & n5390 ) ;
  assign n5722 = ~n601 & n4934 ;
  assign n5717 = n523 | n2178 ;
  assign n5718 = n2127 | n3939 ;
  assign n5719 = n5717 &  n5718 ;
  assign n5720 = ~n2022 & n4430 ;
  assign n5721 = ( n2022 & n5719 ) | ( n2022 & n5720 ) | ( n5719 & n5720 ) ;
  assign n5723 = ( n601 & n5722 ) | ( n601 & n5721 ) | ( n5722 & n5721 ) ;
  assign n5724 = ~x29 & n5723 ;
  assign n5509 = ( n4858 & ~n5494 ) | ( n4858 & n5507 ) | ( ~n5494 & n5507 ) ;
  assign n5510 = ( n4858 & ~n5507 ) | ( n4858 & n5494 ) | ( ~n5507 & n5494 ) ;
  assign n5511 = ( n5509 & ~n4858 ) | ( n5509 & n5510 ) | ( ~n4858 & n5510 ) ;
  assign n5512 = ( n5443 & ~x11 ) | ( n5443 & n5493 ) | ( ~x11 & n5493 ) ;
  assign n5513 = ( x11 & ~n5443 ) | ( x11 & n5493 ) | ( ~n5443 & n5493 ) ;
  assign n5514 = ( n5512 & ~n5493 ) | ( n5512 & n5513 ) | ( ~n5493 & n5513 ) ;
  assign n5524 = ~n2392 & n3653 ;
  assign n5515 = ~n2483 & n3657 ;
  assign n5517 = n2392 | n2483 ;
  assign n5518 = ( n2392 & ~n2483 ) | ( n2392 & 1'b0 ) | ( ~n2483 & 1'b0 ) ;
  assign n5519 = ( n5517 & ~n2392 ) | ( n5517 & n5518 ) | ( ~n2392 & n5518 ) ;
  assign n5520 = ( n3617 & ~n5519 ) | ( n3617 & 1'b0 ) | ( ~n5519 & 1'b0 ) ;
  assign n5516 = ~n2569 & n3652 ;
  assign n5521 = ( n3644 & ~n3617 ) | ( n3644 & n5519 ) | ( ~n3617 & n5519 ) ;
  assign n5522 = ( n5520 & ~n5516 ) | ( n5520 & n5521 ) | ( ~n5516 & n5521 ) ;
  assign n5523 = ~n5515 & n5522 ;
  assign n5525 = ( n2392 & n5524 ) | ( n2392 & n5523 ) | ( n5524 & n5523 ) ;
  assign n5526 = n58 | n2128 ;
  assign n5527 = ( n190 & ~n457 ) | ( n190 & n5526 ) | ( ~n457 & n5526 ) ;
  assign n5528 = n457 | n5527 ;
  assign n5529 = n117 | n5528 ;
  assign n5530 = n39 | n2427 ;
  assign n5531 = n670 | n5530 ;
  assign n5532 = n224 | n1244 ;
  assign n5533 = n167 | n5532 ;
  assign n5534 = ( n5531 & ~n1907 ) | ( n5531 & n5533 ) | ( ~n1907 & n5533 ) ;
  assign n5535 = n1907 | n5534 ;
  assign n5536 = ( n4089 & ~n5535 ) | ( n4089 & n5529 ) | ( ~n5535 & n5529 ) ;
  assign n5537 = ( n2539 & ~n5529 ) | ( n2539 & n5536 ) | ( ~n5529 & n5536 ) ;
  assign n5538 = ( n5537 & ~n2539 ) | ( n5537 & 1'b0 ) | ( ~n2539 & 1'b0 ) ;
  assign n5539 = ( n2492 & ~n2840 ) | ( n2492 & n5538 ) | ( ~n2840 & n5538 ) ;
  assign n5540 = ~n2492 & n5539 ;
  assign n5541 = ( n1794 & ~n5540 ) | ( n1794 & n3281 ) | ( ~n5540 & n3281 ) ;
  assign n5542 = ( n1794 & ~n5541 ) | ( n1794 & 1'b0 ) | ( ~n5541 & 1'b0 ) ;
  assign n5543 = ( n721 & ~n195 ) | ( n721 & n5542 ) | ( ~n195 & n5542 ) ;
  assign n5544 = ~n721 & n5543 ;
  assign n5545 = ( n5544 & ~n485 ) | ( n5544 & n737 ) | ( ~n485 & n737 ) ;
  assign n5546 = ( n5545 & ~n737 ) | ( n5545 & 1'b0 ) | ( ~n737 & 1'b0 ) ;
  assign n5547 = ( n405 & ~n568 ) | ( n405 & n5546 ) | ( ~n568 & n5546 ) ;
  assign n5548 = ~n405 & n5547 ;
  assign n5549 = ~n252 & n5548 ;
  assign n5550 = n52 | n679 ;
  assign n5551 = n337 | n602 ;
  assign n5552 = n226 | n5551 ;
  assign n5553 = ( n3093 & ~n1885 ) | ( n3093 & n5552 ) | ( ~n1885 & n5552 ) ;
  assign n5554 = n1885 | n5553 ;
  assign n5555 = ( n4873 & ~n1627 ) | ( n4873 & n5554 ) | ( ~n1627 & n5554 ) ;
  assign n5556 = n1627 | n5555 ;
  assign n5557 = ( n1703 & ~n673 ) | ( n1703 & n5556 ) | ( ~n673 & n5556 ) ;
  assign n5558 = n673 | n5557 ;
  assign n5559 = ( n414 & ~n722 ) | ( n414 & n5558 ) | ( ~n722 & n5558 ) ;
  assign n5560 = n722 | n5559 ;
  assign n5561 = ( n271 & ~n744 ) | ( n271 & n5560 ) | ( ~n744 & n5560 ) ;
  assign n5562 = n744 | n5561 ;
  assign n5563 = ( n452 & ~n911 ) | ( n452 & n5562 ) | ( ~n911 & n5562 ) ;
  assign n5564 = n911 | n5563 ;
  assign n5565 = ( n228 & n623 ) | ( n228 & n5564 ) | ( n623 & n5564 ) ;
  assign n5566 = ( n623 & ~n5565 ) | ( n623 & 1'b0 ) | ( ~n5565 & 1'b0 ) ;
  assign n5567 = ~n285 & n5566 ;
  assign n5568 = ( n60 & ~n103 ) | ( n60 & n63 ) | ( ~n103 & n63 ) ;
  assign n5569 = ~n63 & n5568 ;
  assign n5570 = ( n60 & ~n5569 ) | ( n60 & n4152 ) | ( ~n5569 & n4152 ) ;
  assign n5571 = ( n126 & ~n534 ) | ( n126 & n5570 ) | ( ~n534 & n5570 ) ;
  assign n5572 = ( n534 & ~n796 ) | ( n534 & n5571 ) | ( ~n796 & n5571 ) ;
  assign n5573 = n796 | n5572 ;
  assign n5574 = ( n74 & ~n5573 ) | ( n74 & n197 ) | ( ~n5573 & n197 ) ;
  assign n5575 = ~n74 & n5574 ;
  assign n5576 = ~n666 & n5575 ;
  assign n5583 = ( n746 & ~n1284 ) | ( n746 & n283 ) | ( ~n1284 & n283 ) ;
  assign n5584 = n1284 | n5583 ;
  assign n5585 = ( n1959 & ~n5584 ) | ( n1959 & n2084 ) | ( ~n5584 & n2084 ) ;
  assign n5586 = ~n1959 & n5585 ;
  assign n5577 = ( n568 & ~n269 ) | ( n568 & n3069 ) | ( ~n269 & n3069 ) ;
  assign n5578 = n269 | n5577 ;
  assign n5579 = ( n240 & ~n540 ) | ( n240 & n5578 ) | ( ~n540 & n5578 ) ;
  assign n5580 = ( n540 & ~n332 ) | ( n540 & n5579 ) | ( ~n332 & n5579 ) ;
  assign n5581 = n332 | n5580 ;
  assign n5582 = n229 | n5581 ;
  assign n5587 = ( n5576 & ~n5586 ) | ( n5576 & n5582 ) | ( ~n5586 & n5582 ) ;
  assign n5588 = ( n61 & ~n5587 ) | ( n61 & n5576 ) | ( ~n5587 & n5576 ) ;
  assign n5589 = ~n61 & n5588 ;
  assign n5590 = ( n242 & ~n191 ) | ( n242 & n5589 ) | ( ~n191 & n5589 ) ;
  assign n5591 = ( n161 & ~n242 ) | ( n161 & n5590 ) | ( ~n242 & n5590 ) ;
  assign n5592 = ~n161 & n5591 ;
  assign n5593 = ( n484 & ~n5592 ) | ( n484 & n618 ) | ( ~n5592 & n618 ) ;
  assign n5594 = ( n484 & ~n5593 ) | ( n484 & 1'b0 ) | ( ~n5593 & 1'b0 ) ;
  assign n5595 = ( n492 & ~n476 ) | ( n492 & n5594 ) | ( ~n476 & n5594 ) ;
  assign n5596 = ( n631 & ~n492 ) | ( n631 & n5595 ) | ( ~n492 & n5595 ) ;
  assign n5597 = ~n631 & n5596 ;
  assign n5603 = n719 | n2626 ;
  assign n5604 = ( n676 & ~n234 ) | ( n676 & n5603 ) | ( ~n234 & n5603 ) ;
  assign n5605 = n234 | n5604 ;
  assign n5606 = ( n123 & ~n714 ) | ( n123 & n5605 ) | ( ~n714 & n5605 ) ;
  assign n5607 = n714 | n5606 ;
  assign n5608 = n617 | n5607 ;
  assign n5609 = n1430 | n2044 ;
  assign n5610 = ( n455 & ~n619 ) | ( n455 & n5609 ) | ( ~n619 & n5609 ) ;
  assign n5611 = n619 | n5610 ;
  assign n5612 = ( n150 & ~n267 ) | ( n150 & n5611 ) | ( ~n267 & n5611 ) ;
  assign n5613 = n267 | n5612 ;
  assign n5614 = ( n137 & ~n300 ) | ( n137 & n5613 ) | ( ~n300 & n5613 ) ;
  assign n5615 = n300 | n5614 ;
  assign n5616 = ( n256 & ~n664 ) | ( n256 & n5615 ) | ( ~n664 & n5615 ) ;
  assign n5617 = n664 | n5616 ;
  assign n5618 = n1689 | n5456 ;
  assign n5619 = ( n5617 & ~n5608 ) | ( n5617 & n5618 ) | ( ~n5608 & n5618 ) ;
  assign n5620 = ( n5608 & ~n2701 ) | ( n5608 & n5619 ) | ( ~n2701 & n5619 ) ;
  assign n5621 = n2701 | n5620 ;
  assign n5598 = n106 | n493 ;
  assign n5599 = n255 | n5598 ;
  assign n5600 = ( n3222 & ~n425 ) | ( n3222 & n5599 ) | ( ~n425 & n5599 ) ;
  assign n5601 = n425 | n5600 ;
  assign n5602 = n775 | n5601 ;
  assign n5622 = ( n5597 & n5621 ) | ( n5597 & n5602 ) | ( n5621 & n5602 ) ;
  assign n5623 = ( n5567 & ~n5597 ) | ( n5567 & n5622 ) | ( ~n5597 & n5622 ) ;
  assign n5624 = ( n5567 & ~n5623 ) | ( n5567 & 1'b0 ) | ( ~n5623 & 1'b0 ) ;
  assign n5625 = ( n5550 & ~n257 ) | ( n5550 & n5624 ) | ( ~n257 & n5624 ) ;
  assign n5626 = ( n130 & ~n5550 ) | ( n130 & n5625 ) | ( ~n5550 & n5625 ) ;
  assign n5627 = ~n130 & n5626 ;
  assign n5628 = ( n558 & ~n169 ) | ( n558 & n5627 ) | ( ~n169 & n5627 ) ;
  assign n5629 = ~n558 & n5628 ;
  assign n5630 = ( n5629 & ~n646 ) | ( n5629 & n663 ) | ( ~n646 & n663 ) ;
  assign n5631 = ( n5630 & ~n663 ) | ( n5630 & 1'b0 ) | ( ~n663 & 1'b0 ) ;
  assign n5632 = ~n432 & n5631 ;
  assign n5633 = n412 | n947 ;
  assign n5634 = ( n765 & ~n560 ) | ( n765 & n5633 ) | ( ~n560 & n5633 ) ;
  assign n5635 = n560 | n5634 ;
  assign n5636 = ( n347 & ~n433 ) | ( n347 & n5635 ) | ( ~n433 & n5635 ) ;
  assign n5637 = n433 | n5636 ;
  assign n5638 = n998 | n3228 ;
  assign n5639 = ( n1325 & ~n408 ) | ( n1325 & n5638 ) | ( ~n408 & n5638 ) ;
  assign n5640 = n408 | n5639 ;
  assign n5641 = ( n672 & ~n245 ) | ( n672 & n5640 ) | ( ~n245 & n5640 ) ;
  assign n5642 = n245 | n5641 ;
  assign n5643 = ( n206 & ~n58 ) | ( n206 & n5642 ) | ( ~n58 & n5642 ) ;
  assign n5644 = n58 | n5643 ;
  assign n5645 = ( n343 & n492 ) | ( n343 & n5644 ) | ( n492 & n5644 ) ;
  assign n5646 = ( n343 & ~n5645 ) | ( n343 & 1'b0 ) | ( ~n5645 & 1'b0 ) ;
  assign n5647 = ~n212 & n5646 ;
  assign n5648 = ~n188 & n624 ;
  assign n5649 = ~n39 & n5648 ;
  assign n5650 = ( n1284 & ~n4545 ) | ( n1284 & n5649 ) | ( ~n4545 & n5649 ) ;
  assign n5651 = ~n1284 & n5650 ;
  assign n5652 = ( n5637 & n5647 ) | ( n5637 & n5651 ) | ( n5647 & n5651 ) ;
  assign n5653 = ( n1060 & ~n5637 ) | ( n1060 & n5652 ) | ( ~n5637 & n5652 ) ;
  assign n5654 = ~n1060 & n5653 ;
  assign n5655 = ( n1001 & ~n570 ) | ( n1001 & n5654 ) | ( ~n570 & n5654 ) ;
  assign n5656 = ~n1001 & n5655 ;
  assign n5657 = ( n1678 & ~n2484 ) | ( n1678 & n5656 ) | ( ~n2484 & n5656 ) ;
  assign n5658 = ~n1678 & n5657 ;
  assign n5659 = ( n671 & ~n260 ) | ( n671 & n5658 ) | ( ~n260 & n5658 ) ;
  assign n5660 = ~n671 & n5659 ;
  assign n5661 = ( n572 & ~n268 ) | ( n572 & n5660 ) | ( ~n268 & n5660 ) ;
  assign n5662 = ~n572 & n5661 ;
  assign n5663 = ( n148 & ~n88 ) | ( n148 & n5662 ) | ( ~n88 & n5662 ) ;
  assign n5664 = ~n148 & n5663 ;
  assign n5665 = n1010 | n2508 ;
  assign n5666 = ( n2062 & ~n530 ) | ( n2062 & n5665 ) | ( ~n530 & n5665 ) ;
  assign n5667 = n530 | n5666 ;
  assign n5668 = ( n124 & ~n457 ) | ( n124 & n5667 ) | ( ~n457 & n5667 ) ;
  assign n5669 = n457 | n5668 ;
  assign n5670 = ( n101 & ~n226 ) | ( n101 & n5669 ) | ( ~n226 & n5669 ) ;
  assign n5671 = n226 | n5670 ;
  assign n5672 = ( n404 & ~n571 ) | ( n404 & n5671 ) | ( ~n571 & n5671 ) ;
  assign n5673 = n571 | n5672 ;
  assign n5674 = n356 | n5673 ;
  assign n5675 = n275 | n716 ;
  assign n5676 = ( n235 & ~n208 ) | ( n235 & n5675 ) | ( ~n208 & n5675 ) ;
  assign n5677 = n208 | n5676 ;
  assign n5678 = ( n137 & ~n403 ) | ( n137 & n5677 ) | ( ~n403 & n5677 ) ;
  assign n5679 = n403 | n5678 ;
  assign n5680 = ( n117 & ~n129 ) | ( n117 & n5679 ) | ( ~n129 & n5679 ) ;
  assign n5681 = n129 | n5680 ;
  assign n5682 = n166 | n5681 ;
  assign n5683 = n3421 | n4543 ;
  assign n5684 = ( n4531 & ~n5683 ) | ( n4531 & n5682 ) | ( ~n5683 & n5682 ) ;
  assign n5685 = ( n843 & ~n5682 ) | ( n843 & n5684 ) | ( ~n5682 & n5684 ) ;
  assign n5686 = ~n843 & n5685 ;
  assign n5687 = ( n5674 & ~n677 ) | ( n5674 & n5686 ) | ( ~n677 & n5686 ) ;
  assign n5688 = ( n1046 & ~n5674 ) | ( n1046 & n5687 ) | ( ~n5674 & n5687 ) ;
  assign n5689 = ~n1046 & n5688 ;
  assign n5690 = ( n1279 & ~n5664 ) | ( n1279 & n5689 ) | ( ~n5664 & n5689 ) ;
  assign n5691 = ( n5664 & ~n355 ) | ( n5664 & n5690 ) | ( ~n355 & n5690 ) ;
  assign n5692 = n355 &  n5691 ;
  assign n5693 = ( n359 & ~n372 ) | ( n359 & n5692 ) | ( ~n372 & n5692 ) ;
  assign n5694 = ~n359 & n5693 ;
  assign n5695 = ( n460 & ~n485 ) | ( n460 & n5694 ) | ( ~n485 & n5694 ) ;
  assign n5696 = ~n460 & n5695 ;
  assign n5697 = ( n432 & ~n5696 ) | ( n432 & n524 ) | ( ~n5696 & n524 ) ;
  assign n5698 = ( n524 & ~n5697 ) | ( n524 & 1'b0 ) | ( ~n5697 & 1'b0 ) ;
  assign n5699 = ( x8 & n5632 ) | ( x8 & n5698 ) | ( n5632 & n5698 ) ;
  assign n5700 = n2569 | n2665 ;
  assign n5701 = ( n2569 & ~n2665 ) | ( n2569 & 1'b0 ) | ( ~n2665 & 1'b0 ) ;
  assign n5702 = ( n5700 & ~n2569 ) | ( n5700 & n5701 ) | ( ~n2569 & n5701 ) ;
  assign n5703 = ~n3615 & n5702 ;
  assign n5704 = ( n3615 & ~n5702 ) | ( n3615 & 1'b0 ) | ( ~n5702 & 1'b0 ) ;
  assign n5705 = n5703 | n5704 ;
  assign n5706 = n3644 | n5705 ;
  assign n5707 = n2751 &  n3652 ;
  assign n5708 = n2569 | n3653 ;
  assign n5709 = ~n2665 & n3657 ;
  assign n5710 = ( n5708 & ~n5709 ) | ( n5708 & 1'b0 ) | ( ~n5709 & 1'b0 ) ;
  assign n5711 = ( n5707 & ~n3652 ) | ( n5707 & n5710 ) | ( ~n3652 & n5710 ) ;
  assign n5712 = n5706 &  n5711 ;
  assign n5713 = ( n5699 & ~n5443 ) | ( n5699 & n5712 ) | ( ~n5443 & n5712 ) ;
  assign n5714 = ( n5549 & ~n5443 ) | ( n5549 & n5713 ) | ( ~n5443 & n5713 ) ;
  assign n5715 = ( n5514 & n5525 ) | ( n5514 & n5714 ) | ( n5525 & n5714 ) ;
  assign n5716 = ( n5511 & ~n5715 ) | ( n5511 & 1'b0 ) | ( ~n5715 & 1'b0 ) ;
  assign n5725 = ~n5511 & n5715 ;
  assign n5726 = ( x29 & ~n5723 ) | ( x29 & n5725 ) | ( ~n5723 & n5725 ) ;
  assign n5727 = ( n5724 & ~n5716 ) | ( n5724 & n5726 ) | ( ~n5716 & n5726 ) ;
  assign n5728 = ( n5508 & ~n5391 ) | ( n5508 & n5727 ) | ( ~n5391 & n5727 ) ;
  assign n5729 = ( n5386 & n5389 ) | ( n5386 & n5728 ) | ( n5389 & n5728 ) ;
  assign n5730 = n5292 | n5301 ;
  assign n5731 = ( n5299 & ~x29 ) | ( n5299 & n5730 ) | ( ~x29 & n5730 ) ;
  assign n5732 = ( x29 & ~n5730 ) | ( x29 & n5299 ) | ( ~n5730 & n5299 ) ;
  assign n5733 = ( n5731 & ~n5299 ) | ( n5731 & n5732 ) | ( ~n5299 & n5732 ) ;
  assign n5734 = ~n5729 & n5733 ;
  assign n5743 = ( n5729 & ~n5733 ) | ( n5729 & 1'b0 ) | ( ~n5733 & 1'b0 ) ;
  assign n5744 = ( n5741 & ~x26 ) | ( n5741 & n5743 ) | ( ~x26 & n5743 ) ;
  assign n5745 = ( n5742 & ~n5734 ) | ( n5742 & n5744 ) | ( ~n5734 & n5744 ) ;
  assign n5746 = ( n5374 & ~n5745 ) | ( n5374 & 1'b0 ) | ( ~n5745 & 1'b0 ) ;
  assign n5755 = ~n5374 & n5745 ;
  assign n5756 = ( n5753 & ~x23 ) | ( n5753 & n5755 ) | ( ~x23 & n5755 ) ;
  assign n5757 = ( n5754 & ~n5746 ) | ( n5754 & n5756 ) | ( ~n5746 & n5756 ) ;
  assign n5758 = ( n5367 & n5370 ) | ( n5367 & n5757 ) | ( n5370 & n5757 ) ;
  assign n5759 = ( n5357 & ~n5758 ) | ( n5357 & 1'b0 ) | ( ~n5758 & 1'b0 ) ;
  assign n5767 = ~n5357 & n5758 ;
  assign n5768 = ( n5765 & ~x20 ) | ( n5765 & n5767 ) | ( ~x20 & n5767 ) ;
  assign n5769 = ( n5766 & ~n5759 ) | ( n5766 & n5768 ) | ( ~n5759 & n5768 ) ;
  assign n5352 = ( n5328 & n5346 ) | ( n5328 & n5349 ) | ( n5346 & n5349 ) ;
  assign n5351 = ( n5328 & ~n5346 ) | ( n5328 & n5349 ) | ( ~n5346 & n5349 ) ;
  assign n5353 = ( n5346 & ~n5352 ) | ( n5346 & n5351 ) | ( ~n5352 & n5351 ) ;
  assign n5825 = n1151 | n5135 ;
  assign n5826 = n1378 | n5010 ;
  assign n5827 = n5825 &  n5826 ;
  assign n5828 = n1267 &  n5067 ;
  assign n5829 = ( n5827 & ~n1267 ) | ( n5827 & n5828 ) | ( ~n1267 & n5828 ) ;
  assign n5830 = ( n4061 & ~n5012 ) | ( n4061 & 1'b0 ) | ( ~n5012 & 1'b0 ) ;
  assign n5831 = ( n5829 & ~n5830 ) | ( n5829 & 1'b0 ) | ( ~n5830 & 1'b0 ) ;
  assign n5832 = ( x23 & ~n5831 ) | ( x23 & 1'b0 ) | ( ~n5831 & 1'b0 ) ;
  assign n5778 = n5734 | n5743 ;
  assign n5779 = ( x26 & ~n5778 ) | ( x26 & n5741 ) | ( ~n5778 & n5741 ) ;
  assign n5780 = ( n5741 & ~x26 ) | ( n5741 & n5778 ) | ( ~x26 & n5778 ) ;
  assign n5781 = ( n5779 & ~n5741 ) | ( n5779 & n5780 ) | ( ~n5741 & n5780 ) ;
  assign n5782 = ( n5389 & ~n5386 ) | ( n5389 & n5728 ) | ( ~n5386 & n5728 ) ;
  assign n5783 = ( n5386 & ~n5728 ) | ( n5386 & n5389 ) | ( ~n5728 & n5389 ) ;
  assign n5784 = ( n5782 & ~n5389 ) | ( n5782 & n5783 ) | ( ~n5389 & n5783 ) ;
  assign n5788 = ~n1566 & n4962 ;
  assign n5785 = n1748 | n4482 ;
  assign n5786 = n1671 | n4495 ;
  assign n5787 = n5785 &  n5786 ;
  assign n5789 = ( n1566 & n5788 ) | ( n1566 & n5787 ) | ( n5788 & n5787 ) ;
  assign n5790 = ( n4478 & ~n4597 ) | ( n4478 & n5789 ) | ( ~n4597 & n5789 ) ;
  assign n5791 = ~n4478 & n5790 ;
  assign n5792 = ( x26 & ~n5789 ) | ( x26 & n5791 ) | ( ~n5789 & n5791 ) ;
  assign n5793 = ( n5789 & ~x26 ) | ( n5789 & n5791 ) | ( ~x26 & n5791 ) ;
  assign n5794 = ( n5792 & ~n5791 ) | ( n5792 & n5793 ) | ( ~n5791 & n5793 ) ;
  assign n5813 = ~n1875 & n4482 ;
  assign n5810 = n1671 | n4962 ;
  assign n5811 = n1748 | n4495 ;
  assign n5812 = n5810 &  n5811 ;
  assign n5814 = ( n1875 & n5813 ) | ( n1875 & n5812 ) | ( n5813 & n5812 ) ;
  assign n5815 = n4478 | n4580 ;
  assign n5816 = n5814 &  n5815 ;
  assign n5817 = ~x26 & n5816 ;
  assign n5798 = ~n3622 & n5085 ;
  assign n5799 = n5086 | n5798 ;
  assign n5805 = ~n601 & n5799 ;
  assign n5800 = n523 | n2127 ;
  assign n5801 = n2022 | n3939 ;
  assign n5802 = n5800 &  n5801 ;
  assign n5803 = ~n1940 & n4430 ;
  assign n5804 = ( n1940 & n5802 ) | ( n1940 & n5803 ) | ( n5802 & n5803 ) ;
  assign n5806 = ( n601 & n5805 ) | ( n601 & n5804 ) | ( n5805 & n5804 ) ;
  assign n5795 = ( n5391 & n5508 ) | ( n5391 & n5727 ) | ( n5508 & n5727 ) ;
  assign n5796 = ( n5391 & ~n5508 ) | ( n5391 & n5727 ) | ( ~n5508 & n5727 ) ;
  assign n5797 = ( n5508 & ~n5795 ) | ( n5508 & n5796 ) | ( ~n5795 & n5796 ) ;
  assign n5807 = ( x29 & ~n5806 ) | ( x29 & n5797 ) | ( ~n5806 & n5797 ) ;
  assign n5808 = ( n5797 & ~x29 ) | ( n5797 & n5806 ) | ( ~x29 & n5806 ) ;
  assign n5809 = n5807 &  n5808 ;
  assign n5819 = ( x29 & n5797 ) | ( x29 & n5806 ) | ( n5797 & n5806 ) ;
  assign n5818 = ( x29 & ~n5797 ) | ( x29 & n5806 ) | ( ~n5797 & n5806 ) ;
  assign n5820 = ( n5797 & ~n5819 ) | ( n5797 & n5818 ) | ( ~n5819 & n5818 ) ;
  assign n5821 = ( x26 & ~n5816 ) | ( x26 & n5820 ) | ( ~n5816 & n5820 ) ;
  assign n5822 = ( n5817 & ~n5809 ) | ( n5817 & n5821 ) | ( ~n5809 & n5821 ) ;
  assign n5823 = ( n5784 & n5794 ) | ( n5784 & n5822 ) | ( n5794 & n5822 ) ;
  assign n5824 = ( n5781 & ~n5823 ) | ( n5781 & 1'b0 ) | ( ~n5823 & 1'b0 ) ;
  assign n5833 = ~n5781 & n5823 ;
  assign n5834 = ( n5831 & ~x23 ) | ( n5831 & n5833 ) | ( ~x23 & n5833 ) ;
  assign n5835 = ( n5832 & ~n5824 ) | ( n5832 & n5834 ) | ( ~n5824 & n5834 ) ;
  assign n5774 = n5746 | n5755 ;
  assign n5775 = ( x23 & ~n5774 ) | ( x23 & n5753 ) | ( ~n5774 & n5753 ) ;
  assign n5776 = ( n5753 & ~x23 ) | ( n5753 & n5774 ) | ( ~x23 & n5774 ) ;
  assign n5777 = ( n5775 & ~n5753 ) | ( n5775 & n5776 ) | ( ~n5753 & n5776 ) ;
  assign n5836 = n946 &  n5339 ;
  assign n5837 = ~n5337 |  n5334 ;
  assign n5838 = n702 | n5837 ;
  assign n5839 = n863 | n5761 ;
  assign n5840 = n5838 &  n5839 ;
  assign n5841 = ( n5836 & ~n5339 ) | ( n5836 & n5840 ) | ( ~n5339 & n5840 ) ;
  assign n5842 = n3650 | n5341 ;
  assign n5843 = n5841 &  n5842 ;
  assign n5844 = x20 &  n5843 ;
  assign n5845 = x20 | n5843 ;
  assign n5846 = ~n5844 & n5845 ;
  assign n5847 = ( n5835 & ~n5777 ) | ( n5835 & n5846 ) | ( ~n5777 & n5846 ) ;
  assign n5848 = n863 &  n5339 ;
  assign n5849 = n599 | n5837 ;
  assign n5850 = n702 | n5761 ;
  assign n5851 = n5849 &  n5850 ;
  assign n5852 = ( n5848 & ~n5339 ) | ( n5848 & n5851 ) | ( ~n5339 & n5851 ) ;
  assign n5853 = ( n5341 & ~n4452 ) | ( n5341 & n5852 ) | ( ~n4452 & n5852 ) ;
  assign n5854 = ~n5341 & n5853 ;
  assign n5855 = ( x20 & ~n5852 ) | ( x20 & n5854 ) | ( ~n5852 & n5854 ) ;
  assign n5856 = ( n5852 & ~x20 ) | ( n5852 & n5854 ) | ( ~x20 & n5854 ) ;
  assign n5857 = ( n5855 & ~n5854 ) | ( n5855 & n5856 ) | ( ~n5854 & n5856 ) ;
  assign n5858 = ( n5367 & ~n5757 ) | ( n5367 & n5370 ) | ( ~n5757 & n5370 ) ;
  assign n5859 = ( n5370 & ~n5367 ) | ( n5370 & n5757 ) | ( ~n5367 & n5757 ) ;
  assign n5860 = ( n5858 & ~n5370 ) | ( n5858 & n5859 ) | ( ~n5370 & n5859 ) ;
  assign n5861 = ( n5847 & n5857 ) | ( n5847 & n5860 ) | ( n5857 & n5860 ) ;
  assign n5770 = n5759 | n5767 ;
  assign n5771 = ( x20 & ~n5770 ) | ( x20 & n5765 ) | ( ~n5770 & n5765 ) ;
  assign n5772 = ( n5765 & ~x20 ) | ( n5765 & n5770 ) | ( ~x20 & n5770 ) ;
  assign n5773 = ( n5771 & ~n5765 ) | ( n5771 & n5772 ) | ( ~n5765 & n5772 ) ;
  assign n5866 = ( n1483 & ~n5010 ) | ( n1483 & 1'b0 ) | ( ~n5010 & 1'b0 ) ;
  assign n5867 = n1378 | n5067 ;
  assign n5868 = ~n5866 & n5867 ;
  assign n5869 = n1267 &  n5135 ;
  assign n5870 = ( n5868 & ~n1267 ) | ( n5868 & n5869 ) | ( ~n1267 & n5869 ) ;
  assign n5871 = ( n4422 & ~n5012 ) | ( n4422 & 1'b0 ) | ( ~n5012 & 1'b0 ) ;
  assign n5872 = ( n5870 & ~n5871 ) | ( n5870 & 1'b0 ) | ( ~n5871 & 1'b0 ) ;
  assign n5873 = x23 &  n5872 ;
  assign n5874 = x23 | n5872 ;
  assign n5875 = ~n5873 & n5874 ;
  assign n5876 = ( n5784 & ~n5794 ) | ( n5784 & n5822 ) | ( ~n5794 & n5822 ) ;
  assign n5877 = ( n5794 & ~n5823 ) | ( n5794 & n5876 ) | ( ~n5823 & n5876 ) ;
  assign n5937 = n1378 | n5135 ;
  assign n5938 = n1566 | n5010 ;
  assign n5939 = n5937 &  n5938 ;
  assign n5940 = n1483 &  n5067 ;
  assign n5941 = ( n5939 & ~n1483 ) | ( n5939 & n5940 ) | ( ~n1483 & n5940 ) ;
  assign n5942 = ~n5012 & n5038 ;
  assign n5943 = ( n5941 & ~n5942 ) | ( n5941 & 1'b0 ) | ( ~n5942 & 1'b0 ) ;
  assign n5944 = ( x23 & ~n5943 ) | ( x23 & 1'b0 ) | ( ~n5943 & 1'b0 ) ;
  assign n5878 = ( x26 & n5816 ) | ( x26 & n5820 ) | ( n5816 & n5820 ) ;
  assign n5879 = ( n5816 & ~n5878 ) | ( n5816 & n5821 ) | ( ~n5878 & n5821 ) ;
  assign n5882 = ~n2569 & n3657 ;
  assign n5884 = n2483 | n2569 ;
  assign n5885 = ( n2483 & ~n2569 ) | ( n2483 & 1'b0 ) | ( ~n2569 & 1'b0 ) ;
  assign n5886 = ( n5884 & ~n2483 ) | ( n5884 & n5885 ) | ( ~n2483 & n5885 ) ;
  assign n5887 = ( n3616 & ~n5886 ) | ( n3616 & 1'b0 ) | ( ~n5886 & 1'b0 ) ;
  assign n5883 = ~n2665 & n3652 ;
  assign n5888 = ( n3644 & ~n3616 ) | ( n3644 & n5886 ) | ( ~n3616 & n5886 ) ;
  assign n5889 = ( n5887 & ~n5883 ) | ( n5887 & n5888 ) | ( ~n5883 & n5888 ) ;
  assign n5890 = ~n5882 & n5889 ;
  assign n5891 = ~n2483 & n3653 ;
  assign n5892 = ( n2483 & n5890 ) | ( n2483 & n5891 ) | ( n5890 & n5891 ) ;
  assign n5880 = ( n5443 & ~n5549 ) | ( n5443 & n5713 ) | ( ~n5549 & n5713 ) ;
  assign n5881 = ( n5714 & ~n5713 ) | ( n5714 & n5880 ) | ( ~n5713 & n5880 ) ;
  assign n5896 = ~n2178 & n4430 ;
  assign n5893 = n523 | n2392 ;
  assign n5894 = n2296 | n3939 ;
  assign n5895 = n5893 &  n5894 ;
  assign n5897 = ( n2178 & n5896 ) | ( n2178 & n5895 ) | ( n5896 & n5895 ) ;
  assign n5898 = n601 | n5269 ;
  assign n5899 = n5897 &  n5898 ;
  assign n5900 = x29 &  n5899 ;
  assign n5901 = x29 | n5899 ;
  assign n5902 = ~n5900 & n5901 ;
  assign n5903 = ( n5892 & ~n5881 ) | ( n5892 & n5902 ) | ( ~n5881 & n5902 ) ;
  assign n5904 = ( n5525 & ~n5514 ) | ( n5525 & n5714 ) | ( ~n5514 & n5714 ) ;
  assign n5905 = ( n5514 & ~n5714 ) | ( n5514 & n5525 ) | ( ~n5714 & n5525 ) ;
  assign n5906 = ( n5904 & ~n5525 ) | ( n5904 & n5905 ) | ( ~n5525 & n5905 ) ;
  assign n5907 = n5903 | n5906 ;
  assign n5911 = ~n523 & n2296 ;
  assign n5908 = n2127 | n4430 ;
  assign n5909 = n2178 | n3939 ;
  assign n5910 = n5908 &  n5909 ;
  assign n5912 = ( n523 & n5911 ) | ( n523 & n5910 ) | ( n5911 & n5910 ) ;
  assign n5913 = n601 | n5283 ;
  assign n5914 = n5912 &  n5913 ;
  assign n5915 = ( x29 & ~n5914 ) | ( x29 & 1'b0 ) | ( ~n5914 & 1'b0 ) ;
  assign n5916 = n5903 &  n5906 ;
  assign n5917 = ( n5914 & ~x29 ) | ( n5914 & n5916 ) | ( ~x29 & n5916 ) ;
  assign n5918 = ( n5907 & n5915 ) | ( n5907 & n5917 ) | ( n5915 & n5917 ) ;
  assign n5919 = n5716 | n5725 ;
  assign n5920 = ( n5723 & ~x29 ) | ( n5723 & n5919 ) | ( ~x29 & n5919 ) ;
  assign n5921 = ( x29 & ~n5919 ) | ( x29 & n5723 ) | ( ~n5919 & n5723 ) ;
  assign n5922 = ( n5920 & ~n5723 ) | ( n5920 & n5921 ) | ( ~n5723 & n5921 ) ;
  assign n5924 = n1940 | n4482 ;
  assign n5925 = n1875 | n4495 ;
  assign n5926 = n5924 &  n5925 ;
  assign n5927 = ~n1748 & n4962 ;
  assign n5928 = ( n1748 & n5926 ) | ( n1748 & n5927 ) | ( n5926 & n5927 ) ;
  assign n5929 = n4478 | n4743 ;
  assign n5930 = n5928 &  n5929 ;
  assign n5932 = ( x26 & ~n5930 ) | ( x26 & 1'b0 ) | ( ~n5930 & 1'b0 ) ;
  assign n5933 = ~x26 & n5930 ;
  assign n5934 = n5932 | n5933 ;
  assign n5935 = ( n5918 & ~n5922 ) | ( n5918 & n5934 ) | ( ~n5922 & n5934 ) ;
  assign n5936 = ( n5879 & ~n5935 ) | ( n5879 & 1'b0 ) | ( ~n5935 & 1'b0 ) ;
  assign n5945 = ~n5879 & n5935 ;
  assign n5946 = ( n5943 & ~x23 ) | ( n5943 & n5945 ) | ( ~x23 & n5945 ) ;
  assign n5947 = ( n5944 & ~n5936 ) | ( n5944 & n5946 ) | ( ~n5936 & n5946 ) ;
  assign n5948 = ( n5875 & n5877 ) | ( n5875 & n5947 ) | ( n5877 & n5947 ) ;
  assign n5862 = n5824 | n5833 ;
  assign n5863 = ( x23 & ~n5862 ) | ( x23 & n5831 ) | ( ~n5862 & n5831 ) ;
  assign n5864 = ( n5831 & ~x23 ) | ( n5831 & n5862 ) | ( ~x23 & n5862 ) ;
  assign n5865 = ( n5863 & ~n5831 ) | ( n5863 & n5864 ) | ( ~n5831 & n5864 ) ;
  assign n5952 = ~n946 & n5761 ;
  assign n5949 = n863 | n5837 ;
  assign n5950 = ~n1043 & n5339 ;
  assign n5951 = ( n5949 & ~n5950 ) | ( n5949 & 1'b0 ) | ( ~n5950 & 1'b0 ) ;
  assign n5953 = ( n946 & n5952 ) | ( n946 & n5951 ) | ( n5952 & n5951 ) ;
  assign n5954 = n3914 | n5341 ;
  assign n5955 = n5953 &  n5954 ;
  assign n5956 = x20 &  n5955 ;
  assign n5957 = x20 | n5955 ;
  assign n5958 = ~n5956 & n5957 ;
  assign n5959 = ( n5948 & ~n5865 ) | ( n5948 & n5958 ) | ( ~n5865 & n5958 ) ;
  assign n5978 = ( n5777 & n5835 ) | ( n5777 & n5846 ) | ( n5835 & n5846 ) ;
  assign n5979 = ( n5777 & ~n5835 ) | ( n5777 & n5846 ) | ( ~n5835 & n5846 ) ;
  assign n5980 = ( n5835 & ~n5978 ) | ( n5835 & n5979 ) | ( ~n5978 & n5979 ) ;
  assign n5963 = ( x14 & ~x15 ) | ( x14 & 1'b0 ) | ( ~x15 & 1'b0 ) ;
  assign n5964 = ~x14 & x15 ;
  assign n5965 = n5963 | n5964 ;
  assign n5966 = ( x16 & ~x17 ) | ( x16 & 1'b0 ) | ( ~x17 & 1'b0 ) ;
  assign n5967 = ~x16 & x17 ;
  assign n5968 = n5966 | n5967 ;
  assign n5972 = ~n5965 | ~n5968 ;
  assign n5960 = ~x15 & x16 ;
  assign n5961 = ( x15 & ~x16 ) | ( x15 & 1'b0 ) | ( ~x16 & 1'b0 ) ;
  assign n5962 = n5960 | n5961 ;
  assign n5969 = ( n5962 & ~n5965 ) | ( n5962 & n5968 ) | ( ~n5965 & n5968 ) ;
  assign n5970 = ~n5969 |  n5962 ;
  assign n5971 = n599 | n5970 ;
  assign n5973 = ( n3637 & ~n5972 ) | ( n3637 & n5971 ) | ( ~n5972 & n5971 ) ;
  assign n5974 = ~n3637 & n5973 ;
  assign n5976 = ( x17 & n5971 ) | ( x17 & n5974 ) | ( n5971 & n5974 ) ;
  assign n5975 = ( x17 & ~n5974 ) | ( x17 & n5971 ) | ( ~n5974 & n5971 ) ;
  assign n5977 = ( n5974 & ~n5976 ) | ( n5974 & n5975 ) | ( ~n5976 & n5975 ) ;
  assign n5981 = ( n5959 & ~n5980 ) | ( n5959 & n5977 ) | ( ~n5980 & n5977 ) ;
  assign n5982 = ( n5847 & ~n5857 ) | ( n5847 & n5860 ) | ( ~n5857 & n5860 ) ;
  assign n5983 = ( n5857 & ~n5861 ) | ( n5857 & n5982 ) | ( ~n5861 & n5982 ) ;
  assign n6169 = n702 | n5970 ;
  assign n6170 = ~n5962 |  n5965 ;
  assign n6171 = n599 | n6170 ;
  assign n6172 = n6169 &  n6171 ;
  assign n6173 = ( n3937 & ~n5972 ) | ( n3937 & 1'b0 ) | ( ~n5972 & 1'b0 ) ;
  assign n6174 = ( n6172 & ~n6173 ) | ( n6172 & 1'b0 ) | ( ~n6173 & 1'b0 ) ;
  assign n6175 = ( x17 & ~n6174 ) | ( x17 & 1'b0 ) | ( ~n6174 & 1'b0 ) ;
  assign n5990 = ( n5875 & ~n5947 ) | ( n5875 & n5877 ) | ( ~n5947 & n5877 ) ;
  assign n5991 = ( n5877 & ~n5875 ) | ( n5877 & n5947 ) | ( ~n5875 & n5947 ) ;
  assign n5992 = ( n5990 & ~n5877 ) | ( n5990 & n5991 ) | ( ~n5877 & n5991 ) ;
  assign n5996 = ~n946 & n5837 ;
  assign n5993 = ~n1151 & n5339 ;
  assign n5994 = n1043 | n5761 ;
  assign n5995 = ~n5993 & n5994 ;
  assign n5997 = ( n946 & n5996 ) | ( n946 & n5995 ) | ( n5996 & n5995 ) ;
  assign n5998 = ( n5341 & ~n4038 ) | ( n5341 & n5997 ) | ( ~n4038 & n5997 ) ;
  assign n5999 = ~n5341 & n5998 ;
  assign n6000 = ( x20 & ~n5997 ) | ( x20 & n5999 ) | ( ~n5997 & n5999 ) ;
  assign n6001 = ( n5997 & ~x20 ) | ( n5997 & n5999 ) | ( ~x20 & n5999 ) ;
  assign n6002 = ( n6000 & ~n5999 ) | ( n6000 & n6001 ) | ( ~n5999 & n6001 ) ;
  assign n6143 = n1671 | n5010 ;
  assign n6144 = n1566 | n5067 ;
  assign n6145 = n6143 &  n6144 ;
  assign n6146 = n1483 &  n5135 ;
  assign n6147 = ( n6145 & ~n1483 ) | ( n6145 & n6146 ) | ( ~n1483 & n6146 ) ;
  assign n6148 = ( n4274 & ~n5012 ) | ( n4274 & 1'b0 ) | ( ~n5012 & 1'b0 ) ;
  assign n6149 = ( n6147 & ~n6148 ) | ( n6147 & 1'b0 ) | ( ~n6148 & 1'b0 ) ;
  assign n6150 = ( x23 & ~n6149 ) | ( x23 & 1'b0 ) | ( ~n6149 & 1'b0 ) ;
  assign n5923 = ~n5918 & n5922 ;
  assign n5931 = ( n5918 & ~n5922 ) | ( n5918 & 1'b0 ) | ( ~n5922 & 1'b0 ) ;
  assign n6007 = n5923 | n5931 ;
  assign n6008 = ( x26 & ~n6007 ) | ( x26 & n5930 ) | ( ~n6007 & n5930 ) ;
  assign n6009 = ( n5930 & ~x26 ) | ( n5930 & n6007 ) | ( ~x26 & n6007 ) ;
  assign n6010 = ( n6008 & ~n5930 ) | ( n6008 & n6009 ) | ( ~n5930 & n6009 ) ;
  assign n6011 = ( n5907 & ~n5916 ) | ( n5907 & 1'b0 ) | ( ~n5916 & 1'b0 ) ;
  assign n6013 = ( x29 & n5914 ) | ( x29 & n6011 ) | ( n5914 & n6011 ) ;
  assign n6012 = ( x29 & ~n5914 ) | ( x29 & n6011 ) | ( ~n5914 & n6011 ) ;
  assign n6014 = ( n5914 & ~n6013 ) | ( n5914 & n6012 ) | ( ~n6013 & n6012 ) ;
  assign n6018 = ~n1875 & n4962 ;
  assign n6015 = n2022 | n4482 ;
  assign n6016 = n1940 | n4495 ;
  assign n6017 = n6015 &  n6016 ;
  assign n6019 = ( n1875 & n6018 ) | ( n1875 & n6017 ) | ( n6018 & n6017 ) ;
  assign n6020 = ( n5381 & ~n4478 ) | ( n5381 & n6019 ) | ( ~n4478 & n6019 ) ;
  assign n6021 = ~n5381 & n6020 ;
  assign n6022 = ( x26 & ~n6019 ) | ( x26 & n6021 ) | ( ~n6019 & n6021 ) ;
  assign n6023 = ( n6019 & ~x26 ) | ( n6019 & n6021 ) | ( ~x26 & n6021 ) ;
  assign n6024 = ( n6022 & ~n6021 ) | ( n6022 & n6023 ) | ( ~n6021 & n6023 ) ;
  assign n6130 = n2127 | n4482 ;
  assign n6131 = n2022 | n4495 ;
  assign n6132 = n6130 &  n6131 ;
  assign n6133 = ~n1940 & n4962 ;
  assign n6134 = ( n1940 & n6132 ) | ( n1940 & n6133 ) | ( n6132 & n6133 ) ;
  assign n6135 = n4478 | n5799 ;
  assign n6136 = n6134 &  n6135 ;
  assign n6137 = ( x26 & ~n6136 ) | ( x26 & 1'b0 ) | ( ~n6136 & 1'b0 ) ;
  assign n6025 = ( n5881 & n5892 ) | ( n5881 & n5902 ) | ( n5892 & n5902 ) ;
  assign n6026 = ( n5881 & ~n5892 ) | ( n5881 & n5902 ) | ( ~n5892 & n5902 ) ;
  assign n6027 = ( n5892 & ~n6025 ) | ( n5892 & n6026 ) | ( ~n6025 & n6026 ) ;
  assign n6036 = ~n601 & n5500 ;
  assign n6034 = ~n2296 & n4430 ;
  assign n6031 = n523 | n2483 ;
  assign n6032 = n2392 | n3939 ;
  assign n6033 = n6031 &  n6032 ;
  assign n6035 = ( n2296 & n6034 ) | ( n2296 & n6033 ) | ( n6034 & n6033 ) ;
  assign n6037 = ( n601 & n6036 ) | ( n601 & n6035 ) | ( n6036 & n6035 ) ;
  assign n6038 = x29 &  n6037 ;
  assign n6039 = x29 | n6037 ;
  assign n6040 = ~n6038 & n6039 ;
  assign n6028 = ( n5443 & ~n5699 ) | ( n5443 & n5712 ) | ( ~n5699 & n5712 ) ;
  assign n6029 = ( n5443 & ~n5712 ) | ( n5443 & n5699 ) | ( ~n5712 & n5699 ) ;
  assign n6030 = ( n6028 & ~n5443 ) | ( n6028 & n6029 ) | ( ~n5443 & n6029 ) ;
  assign n6041 = ( n5632 & ~x8 ) | ( n5632 & n5698 ) | ( ~x8 & n5698 ) ;
  assign n6042 = ( x8 & ~n5632 ) | ( x8 & n5698 ) | ( ~n5632 & n5698 ) ;
  assign n6043 = ( n6041 & ~n5698 ) | ( n6041 & n6042 ) | ( ~n5698 & n6042 ) ;
  assign n6044 = n620 | n1268 ;
  assign n6045 = n460 | n6044 ;
  assign n6046 = ( n4120 & ~n1227 ) | ( n4120 & n6045 ) | ( ~n1227 & n6045 ) ;
  assign n6047 = n1227 | n6046 ;
  assign n6048 = ( n254 & ~n2346 ) | ( n254 & n6047 ) | ( ~n2346 & n6047 ) ;
  assign n6049 = n2346 | n6048 ;
  assign n6050 = ( n2484 & ~n1955 ) | ( n2484 & n6049 ) | ( ~n1955 & n6049 ) ;
  assign n6051 = n1955 | n6050 ;
  assign n6052 = ( n206 & ~n814 ) | ( n206 & n6051 ) | ( ~n814 & n6051 ) ;
  assign n6053 = n814 | n6052 ;
  assign n6054 = ( n221 & ~n405 ) | ( n221 & n6053 ) | ( ~n405 & n6053 ) ;
  assign n6055 = n405 | n6054 ;
  assign n6056 = ( n666 & ~n212 ) | ( n666 & n6055 ) | ( ~n212 & n6055 ) ;
  assign n6057 = n212 | n6056 ;
  assign n6058 = n243 | n408 ;
  assign n6059 = n226 | n6058 ;
  assign n6060 = ( n5637 & ~n1704 ) | ( n5637 & n6059 ) | ( ~n1704 & n6059 ) ;
  assign n6061 = n1704 | n6060 ;
  assign n6062 = ( n6061 & ~n1841 ) | ( n6061 & n5608 ) | ( ~n1841 & n5608 ) ;
  assign n6063 = n6062 | n1841 ;
  assign n6064 = ( n4384 & ~n6063 ) | ( n4384 & n6057 ) | ( ~n6063 & n6057 ) ;
  assign n6065 = ( n887 & ~n6057 ) | ( n887 & n6064 ) | ( ~n6057 & n6064 ) ;
  assign n6066 = ~n887 & n6065 ;
  assign n6067 = ( n458 & ~n477 ) | ( n458 & n6066 ) | ( ~n477 & n6066 ) ;
  assign n6068 = ~n458 & n6067 ;
  assign n6069 = ( n58 & ~n277 ) | ( n58 & n6068 ) | ( ~n277 & n6068 ) ;
  assign n6070 = ~n58 & n6069 ;
  assign n6071 = ( n168 & ~n905 ) | ( n168 & n6070 ) | ( ~n905 & n6070 ) ;
  assign n6072 = ~n168 & n6071 ;
  assign n6073 = ( n569 & ~n6072 ) | ( n569 & n484 ) | ( ~n6072 & n484 ) ;
  assign n6074 = ( n484 & ~n6073 ) | ( n484 & 1'b0 ) | ( ~n6073 & 1'b0 ) ;
  assign n6075 = ( n279 & ~n237 ) | ( n279 & n6074 ) | ( ~n237 & n6074 ) ;
  assign n6076 = ~n279 & n6075 ;
  assign n6077 = n1363 | n2412 ;
  assign n6078 = ( n120 & ~n157 ) | ( n120 & n6077 ) | ( ~n157 & n6077 ) ;
  assign n6079 = n157 | n6078 ;
  assign n6080 = ( n405 & ~n190 ) | ( n405 & n6079 ) | ( ~n190 & n6079 ) ;
  assign n6081 = n190 | n6080 ;
  assign n6082 = n646 | n6081 ;
  assign n6083 = ( n3815 & ~n4911 ) | ( n3815 & n3986 ) | ( ~n4911 & n3986 ) ;
  assign n6084 = ( n1464 & ~n6083 ) | ( n1464 & n3815 ) | ( ~n6083 & n3815 ) ;
  assign n6085 = ( n6084 & ~n1464 ) | ( n6084 & 1'b0 ) | ( ~n1464 & 1'b0 ) ;
  assign n6086 = ( n6082 & ~n1360 ) | ( n6082 & n6085 ) | ( ~n1360 & n6085 ) ;
  assign n6087 = ( n1702 & ~n6082 ) | ( n1702 & n6086 ) | ( ~n6082 & n6086 ) ;
  assign n6088 = ~n1702 & n6087 ;
  assign n6089 = ( n864 & ~n1397 ) | ( n864 & n6088 ) | ( ~n1397 & n6088 ) ;
  assign n6090 = ~n864 & n6089 ;
  assign n6091 = ( n679 & ~n194 ) | ( n679 & n6090 ) | ( ~n194 & n6090 ) ;
  assign n6092 = ~n679 & n6091 ;
  assign n6093 = ( n475 & ~n373 ) | ( n475 & n6092 ) | ( ~n373 & n6092 ) ;
  assign n6094 = ~n475 & n6093 ;
  assign n6095 = ( n162 & ~n214 ) | ( n162 & n6094 ) | ( ~n214 & n6094 ) ;
  assign n6096 = ~n162 & n6095 ;
  assign n6097 = ( n664 & ~n618 ) | ( n664 & n6096 ) | ( ~n618 & n6096 ) ;
  assign n6098 = ~n664 & n6097 ;
  assign n6099 = ~n431 & n6098 ;
  assign n6100 = ( x2 & x5 ) | ( x2 & n6099 ) | ( x5 & n6099 ) ;
  assign n6101 = ( n2783 & ~n2839 ) | ( n2783 & n2910 ) | ( ~n2839 & n2910 ) ;
  assign n6102 = ( n3611 & ~n2910 ) | ( n3611 & n6101 ) | ( ~n2910 & n6101 ) ;
  assign n6103 = ( n2839 & ~n3611 ) | ( n2839 & n6101 ) | ( ~n3611 & n6101 ) ;
  assign n6104 = ( n6102 & ~n2783 ) | ( n6102 & n6103 ) | ( ~n2783 & n6103 ) ;
  assign n6105 = ~n3644 & n6104 ;
  assign n6109 = ~n3657 & n2910 ;
  assign n6106 = n2783 | n3653 ;
  assign n6107 = ~n2839 & n3652 ;
  assign n6108 = ( n6106 & ~n6107 ) | ( n6106 & 1'b0 ) | ( ~n6107 & 1'b0 ) ;
  assign n6110 = ( n6109 & ~n2910 ) | ( n6109 & n6108 ) | ( ~n2910 & n6108 ) ;
  assign n6111 = ~n6105 & n6110 ;
  assign n6112 = ( n6100 & ~n5632 ) | ( n6100 & n6111 ) | ( ~n5632 & n6111 ) ;
  assign n6113 = ( n6076 & ~n5632 ) | ( n6076 & n6112 ) | ( ~n5632 & n6112 ) ;
  assign n6114 = n2665 | n2751 ;
  assign n6115 = ( n2665 & ~n2751 ) | ( n2665 & 1'b0 ) | ( ~n2751 & 1'b0 ) ;
  assign n6116 = ( n6114 & ~n2665 ) | ( n6114 & n6115 ) | ( ~n2665 & n6115 ) ;
  assign n6117 = ~n3614 & n6116 ;
  assign n6118 = ( n3614 & ~n6116 ) | ( n3614 & 1'b0 ) | ( ~n6116 & 1'b0 ) ;
  assign n6119 = n6117 | n6118 ;
  assign n6120 = n3644 | n6119 ;
  assign n6121 = n2751 &  n3657 ;
  assign n6122 = n2665 | n3653 ;
  assign n6123 = ~n2783 & n3652 ;
  assign n6124 = ( n6122 & ~n6123 ) | ( n6122 & 1'b0 ) | ( ~n6123 & 1'b0 ) ;
  assign n6125 = ( n6121 & ~n3657 ) | ( n6121 & n6124 ) | ( ~n3657 & n6124 ) ;
  assign n6126 = n6120 &  n6125 ;
  assign n6127 = ( n6043 & n6113 ) | ( n6043 & n6126 ) | ( n6113 & n6126 ) ;
  assign n6128 = ( n6040 & ~n6030 ) | ( n6040 & n6127 ) | ( ~n6030 & n6127 ) ;
  assign n6129 = ( n6027 & ~n6128 ) | ( n6027 & 1'b0 ) | ( ~n6128 & 1'b0 ) ;
  assign n6138 = ~n6027 & n6128 ;
  assign n6139 = ( n6136 & ~x26 ) | ( n6136 & n6138 ) | ( ~x26 & n6138 ) ;
  assign n6140 = ( n6137 & ~n6129 ) | ( n6137 & n6139 ) | ( ~n6129 & n6139 ) ;
  assign n6141 = ( n6014 & n6024 ) | ( n6014 & n6140 ) | ( n6024 & n6140 ) ;
  assign n6142 = ( n6010 & ~n6141 ) | ( n6010 & 1'b0 ) | ( ~n6141 & 1'b0 ) ;
  assign n6151 = ~n6010 & n6141 ;
  assign n6152 = ( n6149 & ~x23 ) | ( n6149 & n6151 ) | ( ~x23 & n6151 ) ;
  assign n6153 = ( n6150 & ~n6142 ) | ( n6150 & n6152 ) | ( ~n6142 & n6152 ) ;
  assign n6003 = n5936 | n5945 ;
  assign n6004 = ( x23 & ~n6003 ) | ( x23 & n5943 ) | ( ~n6003 & n5943 ) ;
  assign n6005 = ( n5943 & ~x23 ) | ( n5943 & n6003 ) | ( ~x23 & n6003 ) ;
  assign n6006 = ( n6004 & ~n5943 ) | ( n6004 & n6005 ) | ( ~n5943 & n6005 ) ;
  assign n6157 = ~n5339 & n1267 ;
  assign n6154 = n1043 | n5837 ;
  assign n6155 = n1151 | n5761 ;
  assign n6156 = n6154 &  n6155 ;
  assign n6158 = ( n6157 & ~n1267 ) | ( n6157 & n6156 ) | ( ~n1267 & n6156 ) ;
  assign n6159 = n3952 | n5341 ;
  assign n6160 = n6158 &  n6159 ;
  assign n6161 = x20 &  n6160 ;
  assign n6162 = x20 | n6160 ;
  assign n6163 = ~n6161 & n6162 ;
  assign n6164 = ( n6153 & ~n6006 ) | ( n6153 & n6163 ) | ( ~n6006 & n6163 ) ;
  assign n6165 = ( n5992 & n6002 ) | ( n5992 & n6164 ) | ( n6002 & n6164 ) ;
  assign n5987 = ( n5865 & ~n5948 ) | ( n5865 & 1'b0 ) | ( ~n5948 & 1'b0 ) ;
  assign n5988 = ~n5865 & n5948 ;
  assign n5989 = n5987 | n5988 ;
  assign n6166 = ( n5958 & ~n6165 ) | ( n5958 & n5989 ) | ( ~n6165 & n5989 ) ;
  assign n6167 = ( n5958 & n5989 ) | ( n5958 & n6165 ) | ( n5989 & n6165 ) ;
  assign n6168 = ( n6166 & ~n6167 ) | ( n6166 & 1'b0 ) | ( ~n6167 & 1'b0 ) ;
  assign n6176 = ( n5989 & ~n5958 ) | ( n5989 & n6165 ) | ( ~n5958 & n6165 ) ;
  assign n6177 = ( n5958 & ~n6167 ) | ( n5958 & n6176 ) | ( ~n6167 & n6176 ) ;
  assign n6178 = ( n6174 & ~x17 ) | ( n6174 & n6177 ) | ( ~x17 & n6177 ) ;
  assign n6179 = ( n6175 & ~n6168 ) | ( n6175 & n6178 ) | ( ~n6168 & n6178 ) ;
  assign n5985 = ( n5959 & n5977 ) | ( n5959 & n5980 ) | ( n5977 & n5980 ) ;
  assign n5984 = ( n5959 & ~n5977 ) | ( n5959 & n5980 ) | ( ~n5977 & n5980 ) ;
  assign n5986 = ( n5977 & ~n5985 ) | ( n5977 & n5984 ) | ( ~n5985 & n5984 ) ;
  assign n6399 = ~n946 & n5970 ;
  assign n6395 = ~n5965 |  n5968 ;
  assign n6396 = n702 | n6395 ;
  assign n6397 = n863 | n6170 ;
  assign n6398 = n6396 &  n6397 ;
  assign n6400 = ( n946 & n6399 ) | ( n946 & n6398 ) | ( n6399 & n6398 ) ;
  assign n6401 = n3650 | n5972 ;
  assign n6402 = n6400 &  n6401 ;
  assign n6403 = ( x17 & ~n6402 ) | ( x17 & 1'b0 ) | ( ~n6402 & 1'b0 ) ;
  assign n6182 = ( n6006 & n6153 ) | ( n6006 & n6163 ) | ( n6153 & n6163 ) ;
  assign n6183 = ( n6006 & ~n6153 ) | ( n6006 & n6163 ) | ( ~n6153 & n6163 ) ;
  assign n6184 = ( n6153 & ~n6182 ) | ( n6153 & n6183 ) | ( ~n6182 & n6183 ) ;
  assign n6192 = ~n1566 & n5135 ;
  assign n6189 = n1748 | n5010 ;
  assign n6190 = n1671 | n5067 ;
  assign n6191 = n6189 &  n6190 ;
  assign n6193 = ( n1566 & n6192 ) | ( n1566 & n6191 ) | ( n6192 & n6191 ) ;
  assign n6194 = n4597 | n5012 ;
  assign n6195 = n6193 &  n6194 ;
  assign n6196 = x23 &  n6195 ;
  assign n6197 = x23 | n6195 ;
  assign n6198 = ~n6196 & n6197 ;
  assign n6199 = ( n6024 & ~n6014 ) | ( n6024 & n6140 ) | ( ~n6014 & n6140 ) ;
  assign n6200 = ( n6014 & ~n6140 ) | ( n6014 & n6024 ) | ( ~n6140 & n6024 ) ;
  assign n6201 = ( n6199 & ~n6024 ) | ( n6199 & n6200 ) | ( ~n6024 & n6200 ) ;
  assign n6360 = n2178 | n4482 ;
  assign n6361 = n2127 | n4495 ;
  assign n6362 = n6360 &  n6361 ;
  assign n6363 = ~n2022 & n4962 ;
  assign n6364 = ( n2022 & n6362 ) | ( n2022 & n6363 ) | ( n6362 & n6363 ) ;
  assign n6365 = n4478 | n4934 ;
  assign n6366 = n6364 &  n6365 ;
  assign n6367 = ( x26 & ~n6366 ) | ( x26 & 1'b0 ) | ( ~n6366 & 1'b0 ) ;
  assign n6209 = ~n2392 & n4430 ;
  assign n6206 = n523 | n2569 ;
  assign n6207 = n2483 | n3939 ;
  assign n6208 = n6206 &  n6207 ;
  assign n6210 = ( n2392 & n6209 ) | ( n2392 & n6208 ) | ( n6209 & n6208 ) ;
  assign n6211 = ~n3617 & n5519 ;
  assign n6212 = n5520 | n6211 ;
  assign n6213 = n601 | n6212 ;
  assign n6214 = n6210 &  n6213 ;
  assign n6215 = x29 &  n6214 ;
  assign n6216 = x29 | n6214 ;
  assign n6217 = ~n6215 & n6216 ;
  assign n6218 = ( n6043 & ~n6113 ) | ( n6043 & n6126 ) | ( ~n6113 & n6126 ) ;
  assign n6219 = ( n6043 & ~n6126 ) | ( n6043 & n6113 ) | ( ~n6126 & n6113 ) ;
  assign n6220 = ( n6218 & ~n6043 ) | ( n6218 & n6219 ) | ( ~n6043 & n6219 ) ;
  assign n6225 = ( n2751 & ~n2783 ) | ( n2751 & n3613 ) | ( ~n2783 & n3613 ) ;
  assign n6226 = ( n2783 & ~n3614 ) | ( n2783 & n6225 ) | ( ~n3614 & n6225 ) ;
  assign n6231 = ~n3644 & n6226 ;
  assign n6229 = ~n3652 & n2910 ;
  assign n6224 = n2751 | n3653 ;
  assign n6227 = ~n2783 & n3657 ;
  assign n6228 = ( n6224 & ~n6227 ) | ( n6224 & 1'b0 ) | ( ~n6227 & 1'b0 ) ;
  assign n6230 = ( n6229 & ~n2910 ) | ( n6229 & n6228 ) | ( ~n2910 & n6228 ) ;
  assign n6232 = ( n3644 & n6231 ) | ( n3644 & n6230 ) | ( n6231 & n6230 ) ;
  assign n6222 = ( n5632 & n6076 ) | ( n5632 & n6112 ) | ( n6076 & n6112 ) ;
  assign n6221 = ( n5632 & ~n6076 ) | ( n5632 & n6112 ) | ( ~n6076 & n6112 ) ;
  assign n6223 = ( n6076 & ~n6222 ) | ( n6076 & n6221 ) | ( ~n6222 & n6221 ) ;
  assign n6345 = ~n601 & n5705 ;
  assign n6343 = ~n523 & n2751 ;
  assign n6340 = n2569 | n4430 ;
  assign n6341 = n2665 | n3939 ;
  assign n6342 = n6340 &  n6341 ;
  assign n6344 = ( n523 & n6343 ) | ( n523 & n6342 ) | ( n6343 & n6342 ) ;
  assign n6346 = ( n601 & n6345 ) | ( n601 & n6344 ) | ( n6345 & n6344 ) ;
  assign n6347 = ~x29 & n6346 ;
  assign n6233 = ( n5632 & ~n6100 ) | ( n5632 & n6111 ) | ( ~n6100 & n6111 ) ;
  assign n6234 = ( n5632 & ~n6111 ) | ( n5632 & n6100 ) | ( ~n6111 & n6100 ) ;
  assign n6235 = ( n6233 & ~n5632 ) | ( n6233 & n6234 ) | ( ~n5632 & n6234 ) ;
  assign n6236 = ( n875 & ~n3570 ) | ( n875 & 1'b0 ) | ( ~n3570 & 1'b0 ) ;
  assign n6237 = ( n150 & ~n975 ) | ( n150 & n6236 ) | ( ~n975 & n6236 ) ;
  assign n6238 = ~n150 & n6237 ;
  assign n6239 = ( n89 & ~n1208 ) | ( n89 & n6238 ) | ( ~n1208 & n6238 ) ;
  assign n6240 = ~n89 & n6239 ;
  assign n6241 = ~n670 & n6240 ;
  assign n6242 = n4842 | n5533 ;
  assign n6243 = ( n5446 & ~n2033 ) | ( n5446 & n6242 ) | ( ~n2033 & n6242 ) ;
  assign n6244 = n2033 | n6243 ;
  assign n6245 = ( n6241 & n1243 ) | ( n6241 & n6244 ) | ( n1243 & n6244 ) ;
  assign n6246 = ( n2957 & ~n6245 ) | ( n2957 & n6241 ) | ( ~n6245 & n6241 ) ;
  assign n6247 = ( n6246 & ~n2957 ) | ( n6246 & 1'b0 ) | ( ~n2957 & 1'b0 ) ;
  assign n6248 = ( n251 & n3241 ) | ( n251 & n6247 ) | ( n3241 & n6247 ) ;
  assign n6249 = ( n1270 & ~n251 ) | ( n1270 & n6248 ) | ( ~n251 & n6248 ) ;
  assign n6250 = ~n1270 & n6249 ;
  assign n6251 = ( n790 & ~n3777 ) | ( n790 & n6250 ) | ( ~n3777 & n6250 ) ;
  assign n6252 = ~n790 & n6251 ;
  assign n6253 = ( n74 & ~n88 ) | ( n74 & n6252 ) | ( ~n88 & n6252 ) ;
  assign n6254 = ~n74 & n6253 ;
  assign n6255 = ( n664 & ~n93 ) | ( n664 & n6254 ) | ( ~n93 & n6254 ) ;
  assign n6256 = ~n664 & n6255 ;
  assign n6257 = ~n385 & n4090 ;
  assign n6258 = ~n790 & n6257 ;
  assign n6259 = ( n1168 & ~n6258 ) | ( n1168 & n5247 ) | ( ~n6258 & n5247 ) ;
  assign n6260 = ( n1168 & ~n6259 ) | ( n1168 & 1'b0 ) | ( ~n6259 & 1'b0 ) ;
  assign n6261 = ~n1531 & n6260 ;
  assign n6262 = n3826 &  n6261 ;
  assign n6263 = ( n6262 & ~n1433 ) | ( n6262 & n4813 ) | ( ~n1433 & n4813 ) ;
  assign n6264 = ( n3409 & ~n6263 ) | ( n3409 & n4813 ) | ( ~n6263 & n4813 ) ;
  assign n6265 = ( n3409 & ~n6264 ) | ( n3409 & 1'b0 ) | ( ~n6264 & 1'b0 ) ;
  assign n6266 = ( n527 & ~n573 ) | ( n527 & n6265 ) | ( ~n573 & n6265 ) ;
  assign n6267 = ~n527 & n6266 ;
  assign n6268 = ( n1580 & ~n1762 ) | ( n1580 & n6267 ) | ( ~n1762 & n6267 ) ;
  assign n6269 = ( n6268 & ~n1580 ) | ( n6268 & 1'b0 ) | ( ~n1580 & 1'b0 ) ;
  assign n6270 = ( n122 & ~n2308 ) | ( n122 & n6269 ) | ( ~n2308 & n6269 ) ;
  assign n6271 = ~n122 & n6270 ;
  assign n6272 = ( n162 & ~n266 ) | ( n162 & n6271 ) | ( ~n266 & n6271 ) ;
  assign n6273 = ~n162 & n6272 ;
  assign n6274 = ( n603 & ~n229 ) | ( n603 & n6273 ) | ( ~n229 & n6273 ) ;
  assign n6275 = ~n603 & n6274 ;
  assign n6276 = ~n212 & n6275 ;
  assign n6277 = n3381 | n5531 ;
  assign n6278 = ( n5602 & ~n3854 ) | ( n5602 & n6277 ) | ( ~n3854 & n6277 ) ;
  assign n6279 = ( n3854 & ~n2358 ) | ( n3854 & n6278 ) | ( ~n2358 & n6278 ) ;
  assign n6280 = n2358 | n6279 ;
  assign n6281 = ( n1283 & ~n1270 ) | ( n1283 & n6280 ) | ( ~n1270 & n6280 ) ;
  assign n6282 = n1270 | n6281 ;
  assign n6283 = ( n675 & ~n527 ) | ( n675 & n6282 ) | ( ~n527 & n6282 ) ;
  assign n6284 = n527 | n6283 ;
  assign n6285 = ( n258 & ~n65 ) | ( n258 & n6284 ) | ( ~n65 & n6284 ) ;
  assign n6286 = n65 | n6285 ;
  assign n6287 = ( n765 & ~n744 ) | ( n765 & n6286 ) | ( ~n744 & n6286 ) ;
  assign n6288 = n744 | n6287 ;
  assign n6289 = n99 | n6288 ;
  assign n6290 = n195 | n434 ;
  assign n6291 = ( n559 & ~n165 ) | ( n559 & n6290 ) | ( ~n165 & n6290 ) ;
  assign n6292 = n165 | n6291 ;
  assign n6293 = ( n384 & ~n631 ) | ( n384 & n6292 ) | ( ~n631 & n6292 ) ;
  assign n6294 = n631 | n6293 ;
  assign n6295 = ( n3892 & ~n3070 ) | ( n3892 & n4808 ) | ( ~n3070 & n4808 ) ;
  assign n6296 = n3070 | n6295 ;
  assign n6297 = ( n3527 & ~n6294 ) | ( n3527 & n6296 ) | ( ~n6294 & n6296 ) ;
  assign n6298 = ( n3473 & n6297 ) | ( n3473 & n6294 ) | ( n6297 & n6294 ) ;
  assign n6299 = ( n3473 & ~n6298 ) | ( n3473 & 1'b0 ) | ( ~n6298 & 1'b0 ) ;
  assign n6300 = ( n6289 & ~n3853 ) | ( n6289 & n6299 ) | ( ~n3853 & n6299 ) ;
  assign n6301 = ( n215 & ~n6289 ) | ( n215 & n6300 ) | ( ~n6289 & n6300 ) ;
  assign n6302 = ~n215 & n6301 ;
  assign n6303 = ( n2227 & ~n6302 ) | ( n2227 & n3777 ) | ( ~n6302 & n3777 ) ;
  assign n6304 = ( n2227 & ~n6303 ) | ( n2227 & 1'b0 ) | ( ~n6303 & 1'b0 ) ;
  assign n6305 = ( n169 & ~n117 ) | ( n169 & n6304 ) | ( ~n117 & n6304 ) ;
  assign n6306 = ~n169 & n6305 ;
  assign n6307 = ( n6306 & ~n229 ) | ( n6306 & n643 ) | ( ~n229 & n643 ) ;
  assign n6308 = ( n6307 & ~n643 ) | ( n6307 & 1'b0 ) | ( ~n643 & 1'b0 ) ;
  assign n6309 = n3030 | n3106 ;
  assign n6310 = ( n3030 & ~n3106 ) | ( n3030 & 1'b0 ) | ( ~n3106 & 1'b0 ) ;
  assign n6311 = ( n6309 & ~n3030 ) | ( n6309 & n6310 ) | ( ~n3030 & n6310 ) ;
  assign n6312 = ~n3608 & n6311 ;
  assign n6313 = ( n3608 & ~n6311 ) | ( n3608 & 1'b0 ) | ( ~n6311 & 1'b0 ) ;
  assign n6314 = n6312 | n6313 ;
  assign n6315 = n3644 | n6314 ;
  assign n6316 = ~n3197 & n3652 ;
  assign n6317 = ~n3106 & n3657 ;
  assign n6318 = n6316 | n6317 ;
  assign n6319 = ~n3030 & n3653 ;
  assign n6320 = ( n3030 & ~n6318 ) | ( n3030 & n6319 ) | ( ~n6318 & n6319 ) ;
  assign n6321 = n6315 &  n6320 ;
  assign n6322 = ( n6308 & ~x2 ) | ( n6308 & n6321 ) | ( ~x2 & n6321 ) ;
  assign n6323 = ( n6276 & ~x2 ) | ( n6276 & n6322 ) | ( ~x2 & n6322 ) ;
  assign n6324 = ( n6256 & ~x2 ) | ( n6256 & n6323 ) | ( ~x2 & n6323 ) ;
  assign n6328 = ( n2839 & n2910 ) | ( n2839 & n3611 ) | ( n2910 & n3611 ) ;
  assign n6329 = ( n2839 & ~n3611 ) | ( n2839 & n2910 ) | ( ~n3611 & n2910 ) ;
  assign n6330 = ( n3611 & ~n6328 ) | ( n3611 & n6329 ) | ( ~n6328 & n6329 ) ;
  assign n6331 = ~n3644 & n6330 ;
  assign n6335 = n2910 &  n3653 ;
  assign n6332 = ~n2995 & n3652 ;
  assign n6333 = ~n2839 & n3657 ;
  assign n6334 = n6332 | n6333 ;
  assign n6336 = ( n2910 & ~n6335 ) | ( n2910 & n6334 ) | ( ~n6335 & n6334 ) ;
  assign n6337 = n6331 | n6336 ;
  assign n6325 = ( x2 & ~x5 ) | ( x2 & n6099 ) | ( ~x5 & n6099 ) ;
  assign n6326 = ( x2 & ~n6099 ) | ( x2 & x5 ) | ( ~n6099 & x5 ) ;
  assign n6327 = ( n6325 & ~x2 ) | ( n6325 & n6326 ) | ( ~x2 & n6326 ) ;
  assign n6338 = ( n6324 & ~n6337 ) | ( n6324 & n6327 ) | ( ~n6337 & n6327 ) ;
  assign n6339 = ( n6235 & ~n6338 ) | ( n6235 & 1'b0 ) | ( ~n6338 & 1'b0 ) ;
  assign n6348 = ~n6235 & n6338 ;
  assign n6349 = ( x29 & ~n6346 ) | ( x29 & n6348 ) | ( ~n6346 & n6348 ) ;
  assign n6350 = ( n6347 & ~n6339 ) | ( n6347 & n6349 ) | ( ~n6339 & n6349 ) ;
  assign n6351 = ( n6232 & ~n6223 ) | ( n6232 & n6350 ) | ( ~n6223 & n6350 ) ;
  assign n6352 = ( n6217 & n6220 ) | ( n6217 & n6351 ) | ( n6220 & n6351 ) ;
  assign n6353 = ~x29 & n6030 ;
  assign n6354 = x29 | n6030 ;
  assign n6355 = ( n6353 & ~n6030 ) | ( n6353 & n6354 ) | ( ~n6030 & n6354 ) ;
  assign n6357 = ( n6037 & n6127 ) | ( n6037 & n6355 ) | ( n6127 & n6355 ) ;
  assign n6356 = ( n6037 & ~n6355 ) | ( n6037 & n6127 ) | ( ~n6355 & n6127 ) ;
  assign n6358 = ( n6355 & ~n6357 ) | ( n6355 & n6356 ) | ( ~n6357 & n6356 ) ;
  assign n6359 = ~n6352 & n6358 ;
  assign n6368 = ( n6352 & ~n6358 ) | ( n6352 & 1'b0 ) | ( ~n6358 & 1'b0 ) ;
  assign n6369 = ( n6366 & ~x26 ) | ( n6366 & n6368 ) | ( ~x26 & n6368 ) ;
  assign n6370 = ( n6367 & ~n6359 ) | ( n6367 & n6369 ) | ( ~n6359 & n6369 ) ;
  assign n6202 = n6129 | n6138 ;
  assign n6203 = ( x26 & ~n6202 ) | ( x26 & n6136 ) | ( ~n6202 & n6136 ) ;
  assign n6204 = ( n6136 & ~x26 ) | ( n6136 & n6202 ) | ( ~x26 & n6202 ) ;
  assign n6205 = ( n6203 & ~n6136 ) | ( n6203 & n6204 ) | ( ~n6136 & n6204 ) ;
  assign n6374 = ~n1875 & n5010 ;
  assign n6371 = n1671 | n5135 ;
  assign n6372 = n1748 | n5067 ;
  assign n6373 = n6371 &  n6372 ;
  assign n6375 = ( n1875 & n6374 ) | ( n1875 & n6373 ) | ( n6374 & n6373 ) ;
  assign n6376 = n4580 | n5012 ;
  assign n6377 = n6375 &  n6376 ;
  assign n6378 = x23 &  n6377 ;
  assign n6379 = x23 | n6377 ;
  assign n6380 = ~n6378 & n6379 ;
  assign n6381 = ( n6370 & ~n6205 ) | ( n6370 & n6380 ) | ( ~n6205 & n6380 ) ;
  assign n6382 = ( n6198 & n6201 ) | ( n6198 & n6381 ) | ( n6201 & n6381 ) ;
  assign n6185 = n6142 | n6151 ;
  assign n6186 = ( x23 & ~n6185 ) | ( x23 & n6149 ) | ( ~n6185 & n6149 ) ;
  assign n6187 = ( n6149 & ~x23 ) | ( n6149 & n6185 ) | ( ~x23 & n6185 ) ;
  assign n6188 = ( n6186 & ~n6149 ) | ( n6186 & n6187 ) | ( ~n6149 & n6187 ) ;
  assign n6383 = n1151 | n5837 ;
  assign n6384 = ~n1378 & n5339 ;
  assign n6385 = ( n6383 & ~n6384 ) | ( n6383 & 1'b0 ) | ( ~n6384 & 1'b0 ) ;
  assign n6386 = n1267 &  n5761 ;
  assign n6387 = ( n6385 & ~n1267 ) | ( n6385 & n6386 ) | ( ~n1267 & n6386 ) ;
  assign n6388 = ( n4061 & ~n5341 ) | ( n4061 & 1'b0 ) | ( ~n5341 & 1'b0 ) ;
  assign n6389 = ( n6387 & ~n6388 ) | ( n6387 & 1'b0 ) | ( ~n6388 & 1'b0 ) ;
  assign n6390 = x20 &  n6389 ;
  assign n6391 = x20 | n6389 ;
  assign n6392 = ~n6390 & n6391 ;
  assign n6393 = ( n6382 & ~n6188 ) | ( n6382 & n6392 ) | ( ~n6188 & n6392 ) ;
  assign n6394 = ( n6184 & ~n6393 ) | ( n6184 & 1'b0 ) | ( ~n6393 & 1'b0 ) ;
  assign n6404 = ~n6184 & n6393 ;
  assign n6405 = ( n6402 & ~x17 ) | ( n6402 & n6404 ) | ( ~x17 & n6404 ) ;
  assign n6406 = ( n6403 & ~n6394 ) | ( n6403 & n6405 ) | ( ~n6394 & n6405 ) ;
  assign n6410 = ~n863 & n5970 ;
  assign n6407 = n599 | n6395 ;
  assign n6408 = n702 | n6170 ;
  assign n6409 = n6407 &  n6408 ;
  assign n6411 = ( n863 & n6410 ) | ( n863 & n6409 ) | ( n6410 & n6409 ) ;
  assign n6412 = ( n5972 & ~n4452 ) | ( n5972 & n6411 ) | ( ~n4452 & n6411 ) ;
  assign n6413 = ~n5972 & n6412 ;
  assign n6414 = ( x17 & ~n6411 ) | ( x17 & n6413 ) | ( ~n6411 & n6413 ) ;
  assign n6415 = ( n6411 & ~x17 ) | ( n6411 & n6413 ) | ( ~x17 & n6413 ) ;
  assign n6416 = ( n6414 & ~n6413 ) | ( n6414 & n6415 ) | ( ~n6413 & n6415 ) ;
  assign n6417 = ( n5992 & ~n6002 ) | ( n5992 & n6164 ) | ( ~n6002 & n6164 ) ;
  assign n6418 = ( n6002 & ~n6165 ) | ( n6002 & n6417 ) | ( ~n6165 & n6417 ) ;
  assign n6419 = ( n6406 & n6416 ) | ( n6406 & n6418 ) | ( n6416 & n6418 ) ;
  assign n6180 = ( x17 & n6174 ) | ( x17 & n6177 ) | ( n6174 & n6177 ) ;
  assign n6181 = ( x17 & ~n6180 ) | ( x17 & n6178 ) | ( ~n6180 & n6178 ) ;
  assign n6512 = ~n946 & n6170 ;
  assign n6509 = n863 | n6395 ;
  assign n6510 = n1043 | n5970 ;
  assign n6511 = n6509 &  n6510 ;
  assign n6513 = ( n946 & n6512 ) | ( n946 & n6511 ) | ( n6512 & n6511 ) ;
  assign n6514 = n3914 | n5972 ;
  assign n6515 = n6513 &  n6514 ;
  assign n6516 = ( x17 & ~n6515 ) | ( x17 & 1'b0 ) | ( ~n6515 & 1'b0 ) ;
  assign n6420 = ( n6188 & n6382 ) | ( n6188 & n6392 ) | ( n6382 & n6392 ) ;
  assign n6421 = ( n6188 & ~n6382 ) | ( n6188 & n6392 ) | ( ~n6382 & n6392 ) ;
  assign n6422 = ( n6382 & ~n6420 ) | ( n6382 & n6421 ) | ( ~n6420 & n6421 ) ;
  assign n6423 = ( n6198 & ~n6381 ) | ( n6198 & n6201 ) | ( ~n6381 & n6201 ) ;
  assign n6424 = ( n6201 & ~n6198 ) | ( n6201 & n6381 ) | ( ~n6198 & n6381 ) ;
  assign n6425 = ( n6423 & ~n6201 ) | ( n6423 & n6424 ) | ( ~n6201 & n6424 ) ;
  assign n6426 = n1483 &  n5339 ;
  assign n6427 = n1378 | n5761 ;
  assign n6428 = ~n6426 & n6427 ;
  assign n6429 = n1267 &  n5837 ;
  assign n6430 = ( n6428 & ~n1267 ) | ( n6428 & n6429 ) | ( ~n1267 & n6429 ) ;
  assign n6431 = ( n4422 & n5341 ) | ( n4422 & n6430 ) | ( n5341 & n6430 ) ;
  assign n6432 = ~n5341 & n6431 ;
  assign n6433 = ( x20 & ~n6430 ) | ( x20 & n6432 ) | ( ~n6430 & n6432 ) ;
  assign n6434 = ( n6430 & ~x20 ) | ( n6430 & n6432 ) | ( ~x20 & n6432 ) ;
  assign n6435 = ( n6433 & ~n6432 ) | ( n6433 & n6434 ) | ( ~n6432 & n6434 ) ;
  assign n6485 = n1940 | n5010 ;
  assign n6486 = n1875 | n5067 ;
  assign n6487 = n6485 &  n6486 ;
  assign n6488 = ~n1748 & n5135 ;
  assign n6489 = ( n1748 & n6487 ) | ( n1748 & n6488 ) | ( n6487 & n6488 ) ;
  assign n6490 = n4743 | n5012 ;
  assign n6491 = n6489 &  n6490 ;
  assign n6492 = ( x23 & ~n6491 ) | ( x23 & 1'b0 ) | ( ~n6491 & 1'b0 ) ;
  assign n6439 = n6359 | n6368 ;
  assign n6440 = ( x26 & ~n6439 ) | ( x26 & n6366 ) | ( ~n6439 & n6366 ) ;
  assign n6441 = ( n6366 & ~x26 ) | ( n6366 & n6439 ) | ( ~x26 & n6439 ) ;
  assign n6442 = ( n6440 & ~n6366 ) | ( n6440 & n6441 ) | ( ~n6366 & n6441 ) ;
  assign n6443 = ( n6220 & ~n6217 ) | ( n6220 & n6351 ) | ( ~n6217 & n6351 ) ;
  assign n6444 = ( n6217 & ~n6351 ) | ( n6217 & n6220 ) | ( ~n6351 & n6220 ) ;
  assign n6445 = ( n6443 & ~n6220 ) | ( n6443 & n6444 ) | ( ~n6220 & n6444 ) ;
  assign n6449 = ~n2296 & n4482 ;
  assign n6446 = n2127 | n4962 ;
  assign n6447 = n2178 | n4495 ;
  assign n6448 = n6446 &  n6447 ;
  assign n6450 = ( n2296 & n6449 ) | ( n2296 & n6448 ) | ( n6449 & n6448 ) ;
  assign n6451 = ( n5283 & ~n4478 ) | ( n5283 & n6450 ) | ( ~n4478 & n6450 ) ;
  assign n6452 = ~n5283 & n6451 ;
  assign n6453 = ( x26 & ~n6450 ) | ( x26 & n6452 ) | ( ~n6450 & n6452 ) ;
  assign n6454 = ( n6450 & ~x26 ) | ( n6450 & n6452 ) | ( ~x26 & n6452 ) ;
  assign n6455 = ( n6453 & ~n6452 ) | ( n6453 & n6454 ) | ( ~n6452 & n6454 ) ;
  assign n6475 = ~n2178 & n4962 ;
  assign n6472 = n2392 | n4482 ;
  assign n6473 = n2296 | n4495 ;
  assign n6474 = n6472 &  n6473 ;
  assign n6476 = ( n2178 & n6475 ) | ( n2178 & n6474 ) | ( n6475 & n6474 ) ;
  assign n6477 = n4478 | n5269 ;
  assign n6478 = n6476 &  n6477 ;
  assign n6479 = ( x26 & ~n6478 ) | ( x26 & 1'b0 ) | ( ~n6478 & 1'b0 ) ;
  assign n6456 = ( n6223 & n6232 ) | ( n6223 & n6350 ) | ( n6232 & n6350 ) ;
  assign n6457 = ( n6223 & ~n6350 ) | ( n6223 & n6232 ) | ( ~n6350 & n6232 ) ;
  assign n6458 = ( n6350 & ~n6456 ) | ( n6350 & n6457 ) | ( ~n6456 & n6457 ) ;
  assign n6462 = ~n523 & n2665 ;
  assign n6459 = n2483 | n4430 ;
  assign n6460 = n2569 | n3939 ;
  assign n6461 = n6459 &  n6460 ;
  assign n6463 = ( n523 & n6462 ) | ( n523 & n6461 ) | ( n6462 & n6461 ) ;
  assign n6464 = ~n3616 & n5886 ;
  assign n6465 = n5887 | n6464 ;
  assign n6466 = ( n6463 & ~n601 ) | ( n6463 & n6465 ) | ( ~n601 & n6465 ) ;
  assign n6467 = ~n6465 & n6466 ;
  assign n6468 = ( x29 & ~n6463 ) | ( x29 & n6467 ) | ( ~n6463 & n6467 ) ;
  assign n6469 = ( n6463 & ~x29 ) | ( n6463 & n6467 ) | ( ~x29 & n6467 ) ;
  assign n6470 = ( n6468 & ~n6467 ) | ( n6468 & n6469 ) | ( ~n6467 & n6469 ) ;
  assign n6471 = ( n6458 & ~n6470 ) | ( n6458 & 1'b0 ) | ( ~n6470 & 1'b0 ) ;
  assign n6480 = ~n6458 & n6470 ;
  assign n6481 = ( n6478 & ~x26 ) | ( n6478 & n6480 ) | ( ~x26 & n6480 ) ;
  assign n6482 = ( n6479 & ~n6471 ) | ( n6479 & n6481 ) | ( ~n6471 & n6481 ) ;
  assign n6483 = ( n6445 & n6455 ) | ( n6445 & n6482 ) | ( n6455 & n6482 ) ;
  assign n6484 = ( n6442 & ~n6483 ) | ( n6442 & 1'b0 ) | ( ~n6483 & 1'b0 ) ;
  assign n6493 = ~n6442 & n6483 ;
  assign n6494 = ( n6491 & ~x23 ) | ( n6491 & n6493 ) | ( ~x23 & n6493 ) ;
  assign n6495 = ( n6492 & ~n6484 ) | ( n6492 & n6494 ) | ( ~n6484 & n6494 ) ;
  assign n6436 = ( n6205 & n6370 ) | ( n6205 & n6380 ) | ( n6370 & n6380 ) ;
  assign n6437 = ( n6205 & ~n6370 ) | ( n6205 & n6380 ) | ( ~n6370 & n6380 ) ;
  assign n6438 = ( n6370 & ~n6436 ) | ( n6370 & n6437 ) | ( ~n6436 & n6437 ) ;
  assign n6496 = n1378 | n5837 ;
  assign n6497 = ~n1566 & n5339 ;
  assign n6498 = ( n6496 & ~n6497 ) | ( n6496 & 1'b0 ) | ( ~n6497 & 1'b0 ) ;
  assign n6499 = n1483 &  n5761 ;
  assign n6500 = ( n6498 & ~n1483 ) | ( n6498 & n6499 ) | ( ~n1483 & n6499 ) ;
  assign n6501 = ( n5038 & ~n5341 ) | ( n5038 & 1'b0 ) | ( ~n5341 & 1'b0 ) ;
  assign n6502 = ( n6500 & ~n6501 ) | ( n6500 & 1'b0 ) | ( ~n6501 & 1'b0 ) ;
  assign n6503 = x20 &  n6502 ;
  assign n6504 = x20 | n6502 ;
  assign n6505 = ~n6503 & n6504 ;
  assign n6506 = ( n6495 & ~n6438 ) | ( n6495 & n6505 ) | ( ~n6438 & n6505 ) ;
  assign n6507 = ( n6425 & n6435 ) | ( n6425 & n6506 ) | ( n6435 & n6506 ) ;
  assign n6508 = ( n6422 & ~n6507 ) | ( n6422 & 1'b0 ) | ( ~n6507 & 1'b0 ) ;
  assign n6517 = ~n6422 & n6507 ;
  assign n6518 = ( n6515 & ~x17 ) | ( n6515 & n6517 ) | ( ~x17 & n6517 ) ;
  assign n6519 = ( n6516 & ~n6508 ) | ( n6516 & n6518 ) | ( ~n6508 & n6518 ) ;
  assign n6538 = n6394 | n6404 ;
  assign n6539 = ( x17 & ~n6538 ) | ( x17 & n6402 ) | ( ~n6538 & n6402 ) ;
  assign n6540 = ( n6402 & ~x17 ) | ( n6402 & n6538 ) | ( ~x17 & n6538 ) ;
  assign n6541 = ( n6539 & ~n6402 ) | ( n6539 & n6540 ) | ( ~n6402 & n6540 ) ;
  assign n6523 = ( x11 & ~x12 ) | ( x11 & 1'b0 ) | ( ~x12 & 1'b0 ) ;
  assign n6524 = ~x11 & x12 ;
  assign n6525 = n6523 | n6524 ;
  assign n6526 = ( x13 & ~x14 ) | ( x13 & 1'b0 ) | ( ~x14 & 1'b0 ) ;
  assign n6527 = ~x13 & x14 ;
  assign n6528 = n6526 | n6527 ;
  assign n6532 = ~n6525 | ~n6528 ;
  assign n6529 = ~n6525 & n6528 ;
  assign n6520 = ~x12 & x13 ;
  assign n6521 = ( x12 & ~x13 ) | ( x12 & 1'b0 ) | ( ~x13 & 1'b0 ) ;
  assign n6522 = n6520 | n6521 ;
  assign n6530 = ~n6529 |  n6522 ;
  assign n6531 = n599 | n6530 ;
  assign n6533 = ( n6531 & ~n3637 ) | ( n6531 & n6532 ) | ( ~n3637 & n6532 ) ;
  assign n6534 = ~n6532 & n6533 ;
  assign n6536 = ( x14 & n6531 ) | ( x14 & n6534 ) | ( n6531 & n6534 ) ;
  assign n6535 = ( x14 & ~n6534 ) | ( x14 & n6531 ) | ( ~n6534 & n6531 ) ;
  assign n6537 = ( n6534 & ~n6536 ) | ( n6534 & n6535 ) | ( ~n6536 & n6535 ) ;
  assign n6542 = ( n6519 & ~n6541 ) | ( n6519 & n6537 ) | ( ~n6541 & n6537 ) ;
  assign n6543 = ( n6406 & ~n6416 ) | ( n6406 & n6418 ) | ( ~n6416 & n6418 ) ;
  assign n6544 = ( n6416 & ~n6419 ) | ( n6416 & n6543 ) | ( ~n6419 & n6543 ) ;
  assign n6551 = ~n946 & n6395 ;
  assign n6548 = n1151 | n5970 ;
  assign n6549 = n1043 | n6170 ;
  assign n6550 = n6548 &  n6549 ;
  assign n6552 = ( n946 & n6551 ) | ( n946 & n6550 ) | ( n6551 & n6550 ) ;
  assign n6553 = n4038 | n5972 ;
  assign n6554 = n6552 &  n6553 ;
  assign n6555 = x17 &  n6554 ;
  assign n6556 = x17 | n6554 ;
  assign n6557 = ~n6555 & n6556 ;
  assign n6558 = ( n6425 & ~n6435 ) | ( n6425 & n6506 ) | ( ~n6435 & n6506 ) ;
  assign n6559 = ( n6435 & ~n6507 ) | ( n6435 & n6558 ) | ( ~n6507 & n6558 ) ;
  assign n6570 = ~n1875 & n5135 ;
  assign n6567 = n2022 | n5010 ;
  assign n6568 = n1940 | n5067 ;
  assign n6569 = n6567 &  n6568 ;
  assign n6571 = ( n1875 & n6570 ) | ( n1875 & n6569 ) | ( n6570 & n6569 ) ;
  assign n6572 = n5012 | n5381 ;
  assign n6573 = n6571 &  n6572 ;
  assign n6574 = x23 &  n6573 ;
  assign n6575 = x23 | n6573 ;
  assign n6576 = ~n6574 & n6575 ;
  assign n6577 = ( n6445 & ~n6455 ) | ( n6445 & n6482 ) | ( ~n6455 & n6482 ) ;
  assign n6578 = ( n6455 & ~n6483 ) | ( n6455 & n6577 ) | ( ~n6483 & n6577 ) ;
  assign n6596 = ~n2839 & n3653 ;
  assign n6587 = ~n2995 & n3657 ;
  assign n6589 = n2839 | n2995 ;
  assign n6590 = ( n2839 & ~n2995 ) | ( n2839 & 1'b0 ) | ( ~n2995 & 1'b0 ) ;
  assign n6591 = ( n6589 & ~n2839 ) | ( n6589 & n6590 ) | ( ~n2839 & n6590 ) ;
  assign n6592 = ( n3610 & ~n6591 ) | ( n3610 & 1'b0 ) | ( ~n6591 & 1'b0 ) ;
  assign n6588 = ~n3030 & n3652 ;
  assign n6593 = ( n3644 & ~n3610 ) | ( n3644 & n6591 ) | ( ~n3610 & n6591 ) ;
  assign n6594 = ( n6592 & ~n6588 ) | ( n6592 & n6593 ) | ( ~n6588 & n6593 ) ;
  assign n6595 = ~n6587 & n6594 ;
  assign n6597 = ( n2839 & n6596 ) | ( n2839 & n6595 ) | ( n6596 & n6595 ) ;
  assign n6585 = ( x2 & ~n6323 ) | ( x2 & n6256 ) | ( ~n6323 & n6256 ) ;
  assign n6586 = ( n6324 & ~n6256 ) | ( n6324 & n6585 ) | ( ~n6256 & n6585 ) ;
  assign n6600 = ~n3030 & n3657 ;
  assign n6602 = n2995 | n3030 ;
  assign n6603 = ( n2995 & ~n3030 ) | ( n2995 & 1'b0 ) | ( ~n3030 & 1'b0 ) ;
  assign n6604 = ( n6602 & ~n2995 ) | ( n6602 & n6603 ) | ( ~n2995 & n6603 ) ;
  assign n6605 = ( n3609 & ~n6604 ) | ( n3609 & 1'b0 ) | ( ~n6604 & 1'b0 ) ;
  assign n6601 = ~n3106 & n3652 ;
  assign n6606 = ( n3644 & ~n3609 ) | ( n3644 & n6604 ) | ( ~n3609 & n6604 ) ;
  assign n6607 = ( n6605 & ~n6601 ) | ( n6605 & n6606 ) | ( ~n6601 & n6606 ) ;
  assign n6608 = ~n6600 & n6607 ;
  assign n6609 = ~n2995 & n3653 ;
  assign n6610 = ( n2995 & n6608 ) | ( n2995 & n6609 ) | ( n6608 & n6609 ) ;
  assign n6598 = ( x2 & ~n6276 ) | ( x2 & n6322 ) | ( ~n6276 & n6322 ) ;
  assign n6599 = ( n6323 & ~n6322 ) | ( n6323 & n6598 ) | ( ~n6322 & n6598 ) ;
  assign n6614 = n3395 | n4859 ;
  assign n6615 = ( n5247 & ~n4818 ) | ( n5247 & n6614 ) | ( ~n4818 & n6614 ) ;
  assign n6616 = n4818 | n6615 ;
  assign n6617 = ( n2696 & ~n794 ) | ( n2696 & n6616 ) | ( ~n794 & n6616 ) ;
  assign n6618 = n794 | n6617 ;
  assign n6619 = ( n2091 & ~n1883 ) | ( n2091 & n6618 ) | ( ~n1883 & n6618 ) ;
  assign n6620 = n1883 | n6619 ;
  assign n6621 = ( n766 & ~n62 ) | ( n766 & n6620 ) | ( ~n62 & n6620 ) ;
  assign n6622 = n62 | n6621 ;
  assign n6623 = ( n259 & ~n138 ) | ( n259 & n6622 ) | ( ~n138 & n6622 ) ;
  assign n6624 = n138 | n6623 ;
  assign n6625 = ( n207 & ~n406 ) | ( n207 & n6624 ) | ( ~n406 & n6624 ) ;
  assign n6626 = n406 | n6625 ;
  assign n6627 = n266 | n6626 ;
  assign n6628 = n778 | n5550 ;
  assign n6629 = ( n666 & ~n165 ) | ( n666 & n6628 ) | ( ~n165 & n6628 ) ;
  assign n6630 = n165 | n6629 ;
  assign n6631 = ( n148 & ~n124 ) | ( n148 & n787 ) | ( ~n124 & n787 ) ;
  assign n6632 = n124 | n6631 ;
  assign n6633 = n670 | n6632 ;
  assign n6634 = n1363 | n3790 ;
  assign n6635 = ( n6633 & ~n1729 ) | ( n6633 & n6634 ) | ( ~n1729 & n6634 ) ;
  assign n6636 = n1729 | n6635 ;
  assign n6637 = ( n6630 & ~n2610 ) | ( n6630 & n6636 ) | ( ~n2610 & n6636 ) ;
  assign n6638 = n2610 | n6637 ;
  assign n6639 = ( n4898 & ~n4890 ) | ( n4898 & n6638 ) | ( ~n4890 & n6638 ) ;
  assign n6640 = ( n4898 & ~n6639 ) | ( n4898 & 1'b0 ) | ( ~n6639 & 1'b0 ) ;
  assign n6641 = ( n527 & ~n6627 ) | ( n527 & n6640 ) | ( ~n6627 & n6640 ) ;
  assign n6642 = ~n527 & n6641 ;
  assign n6643 = ( n1762 & ~n777 ) | ( n1762 & n6642 ) | ( ~n777 & n6642 ) ;
  assign n6644 = ~n1762 & n6643 ;
  assign n6645 = ( n231 & ~n6644 ) | ( n231 & n813 ) | ( ~n6644 & n813 ) ;
  assign n6646 = ( n813 & ~n6645 ) | ( n813 & 1'b0 ) | ( ~n6645 & 1'b0 ) ;
  assign n6647 = ( n118 & ~n267 ) | ( n118 & n6646 ) | ( ~n267 & n6646 ) ;
  assign n6648 = ~n118 & n6647 ;
  assign n6649 = ~n77 & n6648 ;
  assign n6659 = ~n3106 & n3653 ;
  assign n6650 = ~n3197 & n3657 ;
  assign n6652 = n3106 | n3197 ;
  assign n6653 = ( n3106 & ~n3197 ) | ( n3106 & 1'b0 ) | ( ~n3197 & 1'b0 ) ;
  assign n6654 = ( n6652 & ~n3106 ) | ( n6652 & n6653 ) | ( ~n3106 & n6653 ) ;
  assign n6655 = ( n3607 & ~n6654 ) | ( n3607 & 1'b0 ) | ( ~n6654 & 1'b0 ) ;
  assign n6651 = n3266 &  n3652 ;
  assign n6656 = ( n3644 & ~n3607 ) | ( n3644 & n6654 ) | ( ~n3607 & n6654 ) ;
  assign n6657 = ( n6655 & ~n6651 ) | ( n6655 & n6656 ) | ( ~n6651 & n6656 ) ;
  assign n6658 = ~n6650 & n6657 ;
  assign n6660 = ( n3106 & n6659 ) | ( n3106 & n6658 ) | ( n6659 & n6658 ) ;
  assign n6661 = n208 | n271 ;
  assign n6662 = n256 | n6661 ;
  assign n6663 = ( n6662 & ~n577 ) | ( n6662 & n5399 ) | ( ~n577 & n5399 ) ;
  assign n6664 = n577 | n6663 ;
  assign n6665 = ( n4695 & ~n1356 ) | ( n4695 & n6664 ) | ( ~n1356 & n6664 ) ;
  assign n6666 = n1356 | n6665 ;
  assign n6667 = ( n355 & n6666 ) | ( n355 & n865 ) | ( n6666 & n865 ) ;
  assign n6668 = ( n355 & ~n6667 ) | ( n355 & 1'b0 ) | ( ~n6667 & 1'b0 ) ;
  assign n6669 = ( n797 & ~n235 ) | ( n797 & n6668 ) | ( ~n235 & n6668 ) ;
  assign n6670 = ~n797 & n6669 ;
  assign n6671 = ( n457 & ~n333 ) | ( n457 & n6670 ) | ( ~n333 & n6670 ) ;
  assign n6672 = ~n457 & n6671 ;
  assign n6673 = ( n117 & ~n270 ) | ( n117 & n6672 ) | ( ~n270 & n6672 ) ;
  assign n6674 = ~n117 & n6673 ;
  assign n6675 = ~n664 & n6674 ;
  assign n6680 = n337 | n671 ;
  assign n6681 = n373 | n6680 ;
  assign n6682 = n1076 | n2633 ;
  assign n6683 = ( n1326 & ~n6681 ) | ( n1326 & n6682 ) | ( ~n6681 & n6682 ) ;
  assign n6684 = ( n6681 & ~n2593 ) | ( n6681 & n6683 ) | ( ~n2593 & n6683 ) ;
  assign n6685 = n2593 | n6684 ;
  assign n6676 = n718 | n1580 ;
  assign n6677 = ( n206 & ~n267 ) | ( n206 & n6676 ) | ( ~n267 & n6676 ) ;
  assign n6678 = n267 | n6677 ;
  assign n6679 = n628 | n6678 ;
  assign n6686 = ( n6685 & ~n1877 ) | ( n6685 & n6679 ) | ( ~n1877 & n6679 ) ;
  assign n6687 = n1877 | n6686 ;
  assign n6688 = ( n2610 & ~n3890 ) | ( n2610 & n6687 ) | ( ~n3890 & n6687 ) ;
  assign n6689 = ( n3890 & ~n1510 ) | ( n3890 & n6688 ) | ( ~n1510 & n6688 ) ;
  assign n6690 = n1510 | n6689 ;
  assign n6691 = ( n6675 & ~n6690 ) | ( n6675 & n5453 ) | ( ~n6690 & n5453 ) ;
  assign n6692 = ~n5453 & n6691 ;
  assign n6693 = ( n1581 & ~n555 ) | ( n1581 & n6692 ) | ( ~n555 & n6692 ) ;
  assign n6694 = ~n1581 & n6693 ;
  assign n6695 = ( n376 & ~n6694 ) | ( n376 & n786 ) | ( ~n6694 & n786 ) ;
  assign n6696 = ( n786 & ~n6695 ) | ( n786 & 1'b0 ) | ( ~n6695 & 1'b0 ) ;
  assign n6697 = ( n484 & ~n6696 ) | ( n484 & n765 ) | ( ~n6696 & n765 ) ;
  assign n6698 = ( n484 & ~n6697 ) | ( n484 & 1'b0 ) | ( ~n6697 & 1'b0 ) ;
  assign n6699 = ( n43 & ~n6698 ) | ( n43 & n623 ) | ( ~n6698 & n623 ) ;
  assign n6700 = ( n623 & ~n6699 ) | ( n623 & 1'b0 ) | ( ~n6699 & 1'b0 ) ;
  assign n6701 = n3266 &  n3657 ;
  assign n6702 = ~n3325 & n3652 ;
  assign n6704 = n3197 &  n3266 ;
  assign n6703 = ~n3197 & n3266 ;
  assign n6705 = ( n3197 & ~n6704 ) | ( n3197 & n6703 ) | ( ~n6704 & n6703 ) ;
  assign n6706 = n3606 &  n6705 ;
  assign n6707 = ( n3606 & ~n3644 ) | ( n3606 & n6705 ) | ( ~n3644 & n6705 ) ;
  assign n6708 = ( n6702 & ~n6706 ) | ( n6702 & n6707 ) | ( ~n6706 & n6707 ) ;
  assign n6709 = n6701 | n6708 ;
  assign n6710 = ~n3197 & n3653 ;
  assign n6711 = ( n3197 & ~n6709 ) | ( n3197 & n6710 ) | ( ~n6709 & n6710 ) ;
  assign n6715 = n602 | n906 ;
  assign n6716 = ( n342 & ~n271 ) | ( n342 & n6715 ) | ( ~n271 & n6715 ) ;
  assign n6717 = n271 | n6716 ;
  assign n6712 = n258 | n885 ;
  assign n6713 = ( n531 & ~n643 ) | ( n531 & n6712 ) | ( ~n643 & n6712 ) ;
  assign n6714 = n643 | n6713 ;
  assign n6718 = n2346 | n2494 ;
  assign n6719 = ( n6717 & ~n6714 ) | ( n6717 & n6718 ) | ( ~n6714 & n6718 ) ;
  assign n6720 = ( n6719 & ~n5529 ) | ( n6719 & n6714 ) | ( ~n5529 & n6714 ) ;
  assign n6721 = n5529 | n6720 ;
  assign n6722 = ( n412 & ~n6721 ) | ( n412 & n645 ) | ( ~n6721 & n645 ) ;
  assign n6723 = ~n412 & n6722 ;
  assign n6724 = ( n245 & ~n812 ) | ( n245 & n6723 ) | ( ~n812 & n6723 ) ;
  assign n6725 = ~n245 & n6724 ;
  assign n6726 = ( n277 & ~n270 ) | ( n277 & n6725 ) | ( ~n270 & n6725 ) ;
  assign n6727 = ~n277 & n6726 ;
  assign n6728 = ( n406 & ~n451 ) | ( n406 & n6727 ) | ( ~n451 & n6727 ) ;
  assign n6729 = ~n406 & n6728 ;
  assign n6730 = ( n228 & ~n80 ) | ( n228 & n6729 ) | ( ~n80 & n6729 ) ;
  assign n6731 = ~n228 & n6730 ;
  assign n6732 = ~n137 & n6731 ;
  assign n6733 = n125 | n3011 ;
  assign n6734 = ( n130 & ~n775 ) | ( n130 & n6733 ) | ( ~n775 & n6733 ) ;
  assign n6735 = n775 | n6734 ;
  assign n6736 = n1153 | n2412 ;
  assign n6737 = ( n1008 & ~n6735 ) | ( n1008 & n6736 ) | ( ~n6735 & n6736 ) ;
  assign n6738 = ( n6735 & ~n3180 ) | ( n6735 & n6737 ) | ( ~n3180 & n6737 ) ;
  assign n6739 = n6738 | n3180 ;
  assign n6740 = ( n5597 & ~n6739 ) | ( n5597 & 1'b0 ) | ( ~n6739 & 1'b0 ) ;
  assign n6741 = ( n371 & ~n6732 ) | ( n371 & n6740 ) | ( ~n6732 & n6740 ) ;
  assign n6742 = ( n674 & n6732 ) | ( n674 & n6741 ) | ( n6732 & n6741 ) ;
  assign n6743 = ~n674 & n6742 ;
  assign n6744 = ( n424 & ~n485 ) | ( n424 & n6743 ) | ( ~n485 & n6743 ) ;
  assign n6745 = ~n424 & n6744 ;
  assign n6746 = ( n236 & ~n6745 ) | ( n236 & n343 ) | ( ~n6745 & n343 ) ;
  assign n6747 = ( n343 & ~n6746 ) | ( n343 & 1'b0 ) | ( ~n6746 & 1'b0 ) ;
  assign n6748 = ~n77 & n6747 ;
  assign n6758 = n3266 &  n3653 ;
  assign n6749 = ~n3325 & n3657 ;
  assign n6750 = ~n3361 & n3652 ;
  assign n6751 = ( n3266 & ~n3325 ) | ( n3266 & 1'b0 ) | ( ~n3325 & 1'b0 ) ;
  assign n6752 = ~n3266 & n3325 ;
  assign n6753 = n6751 | n6752 ;
  assign n6754 = n3605 &  n6753 ;
  assign n6755 = ( n3605 & ~n3644 ) | ( n3605 & n6753 ) | ( ~n3644 & n6753 ) ;
  assign n6756 = ( n6750 & ~n6754 ) | ( n6750 & n6755 ) | ( ~n6754 & n6755 ) ;
  assign n6757 = n6749 | n6756 ;
  assign n6759 = ( n3266 & ~n6758 ) | ( n3266 & n6757 ) | ( ~n6758 & n6757 ) ;
  assign n6760 = n1196 | n4561 ;
  assign n6761 = ( n795 & ~n607 ) | ( n795 & n6760 ) | ( ~n607 & n6760 ) ;
  assign n6762 = n607 | n6761 ;
  assign n6763 = ( n2427 & ~n124 ) | ( n2427 & n6762 ) | ( ~n124 & n6762 ) ;
  assign n6764 = n124 | n6763 ;
  assign n6765 = ( n345 & ~n429 ) | ( n345 & n6764 ) | ( ~n429 & n6764 ) ;
  assign n6766 = n429 | n6765 ;
  assign n6767 = ( n372 & ~n602 ) | ( n372 & n6766 ) | ( ~n602 & n6766 ) ;
  assign n6768 = n602 | n6767 ;
  assign n6769 = ( n338 & ~n334 ) | ( n338 & n6768 ) | ( ~n334 & n6768 ) ;
  assign n6770 = n334 | n6769 ;
  assign n6771 = n166 | n787 ;
  assign n6772 = n39 | n6771 ;
  assign n6773 = ( n605 & ~n572 ) | ( n605 & n6772 ) | ( ~n572 & n6772 ) ;
  assign n6774 = n572 | n6773 ;
  assign n6775 = n617 | n6774 ;
  assign n6776 = n573 | n800 ;
  assign n6777 = n213 | n6776 ;
  assign n6778 = ( n4808 & ~n2485 ) | ( n4808 & n6777 ) | ( ~n2485 & n6777 ) ;
  assign n6779 = n2485 | n6778 ;
  assign n6780 = ( n6775 & ~n4150 ) | ( n6775 & n6779 ) | ( ~n4150 & n6779 ) ;
  assign n6781 = ( n3087 & n6780 ) | ( n3087 & n4150 ) | ( n6780 & n4150 ) ;
  assign n6782 = ( n3087 & ~n6781 ) | ( n3087 & 1'b0 ) | ( ~n6781 & 1'b0 ) ;
  assign n6783 = ( n1820 & ~n6770 ) | ( n1820 & n6782 ) | ( ~n6770 & n6782 ) ;
  assign n6784 = ~n1820 & n6783 ;
  assign n6785 = ( n647 & ~n654 ) | ( n647 & n6784 ) | ( ~n654 & n6784 ) ;
  assign n6786 = ~n647 & n6785 ;
  assign n6787 = ( n912 & ~n948 ) | ( n912 & n6786 ) | ( ~n948 & n6786 ) ;
  assign n6788 = ~n912 & n6787 ;
  assign n6789 = ( n344 & n674 ) | ( n344 & n6788 ) | ( n674 & n6788 ) ;
  assign n6790 = ~n674 & n6789 ;
  assign n6791 = ( n6790 & ~n404 ) | ( n6790 & n714 ) | ( ~n404 & n714 ) ;
  assign n6792 = ( n6791 & ~n714 ) | ( n6791 & 1'b0 ) | ( ~n714 & 1'b0 ) ;
  assign n6793 = ( n192 & ~n6792 ) | ( n192 & n644 ) | ( ~n6792 & n644 ) ;
  assign n6794 = ( n644 & ~n6793 ) | ( n644 & 1'b0 ) | ( ~n6793 & 1'b0 ) ;
  assign n6795 = ~n618 & n6794 ;
  assign n6796 = ~n3361 & n3657 ;
  assign n6798 = n3325 | n3361 ;
  assign n6799 = ( n3325 & ~n3361 ) | ( n3325 & 1'b0 ) | ( ~n3361 & 1'b0 ) ;
  assign n6800 = ( n6798 & ~n3325 ) | ( n6798 & n6799 ) | ( ~n3325 & n6799 ) ;
  assign n6801 = ( n3604 & ~n6800 ) | ( n3604 & 1'b0 ) | ( ~n6800 & 1'b0 ) ;
  assign n6797 = ~n3460 & n3652 ;
  assign n6802 = ( n3644 & ~n3604 ) | ( n3644 & n6800 ) | ( ~n3604 & n6800 ) ;
  assign n6803 = ( n6801 & ~n6797 ) | ( n6801 & n6802 ) | ( ~n6797 & n6802 ) ;
  assign n6804 = ~n6796 & n6803 ;
  assign n6805 = ~n3325 & n3653 ;
  assign n6806 = ( n3325 & n6804 ) | ( n3325 & n6805 ) | ( n6804 & n6805 ) ;
  assign n6807 = n374 | n1063 ;
  assign n6808 = ( n793 & ~n217 ) | ( n793 & n6807 ) | ( ~n217 & n6807 ) ;
  assign n6809 = n217 | n6808 ;
  assign n6810 = ( n269 & ~n226 ) | ( n269 & n6809 ) | ( ~n226 & n6809 ) ;
  assign n6811 = n226 | n6810 ;
  assign n6819 = n556 | n1225 ;
  assign n6820 = n169 | n6819 ;
  assign n6821 = n193 | n2958 ;
  assign n6822 = ( n3222 & ~n6820 ) | ( n3222 & n6821 ) | ( ~n6820 & n6821 ) ;
  assign n6823 = ( n6820 & ~n1885 ) | ( n6820 & n6822 ) | ( ~n1885 & n6822 ) ;
  assign n6824 = n1885 | n6823 ;
  assign n6825 = ( n2395 & ~n530 ) | ( n2395 & n6824 ) | ( ~n530 & n6824 ) ;
  assign n6826 = n530 | n6825 ;
  assign n6812 = n1062 | n2521 ;
  assign n6813 = ( n884 & ~n887 ) | ( n884 & n6812 ) | ( ~n887 & n6812 ) ;
  assign n6814 = n887 | n6813 ;
  assign n6815 = ( n197 & n348 ) | ( n197 & n6814 ) | ( n348 & n6814 ) ;
  assign n6816 = ( n197 & ~n6815 ) | ( n197 & 1'b0 ) | ( ~n6815 & 1'b0 ) ;
  assign n6817 = ( n332 & ~n410 ) | ( n332 & n6816 ) | ( ~n410 & n6816 ) ;
  assign n6818 = ~n332 & n6817 ;
  assign n6827 = ( n647 & ~n6826 ) | ( n647 & n6818 ) | ( ~n6826 & n6818 ) ;
  assign n6828 = ~n647 & n6827 ;
  assign n6829 = ( n1490 & ~n1824 ) | ( n1490 & n6828 ) | ( ~n1824 & n6828 ) ;
  assign n6830 = ~n1490 & n6829 ;
  assign n6831 = ( n787 & ~n52 ) | ( n787 & n6830 ) | ( ~n52 & n6830 ) ;
  assign n6832 = ~n787 & n6831 ;
  assign n6833 = ( n80 & ~n6832 ) | ( n80 & n524 ) | ( ~n6832 & n524 ) ;
  assign n6834 = ( n524 & ~n6833 ) | ( n524 & 1'b0 ) | ( ~n6833 & 1'b0 ) ;
  assign n6835 = ( n631 & ~n256 ) | ( n631 & n6834 ) | ( ~n256 & n6834 ) ;
  assign n6836 = ~n631 & n6835 ;
  assign n6837 = n461 | n720 ;
  assign n6838 = n299 | n6837 ;
  assign n6839 = ( n2519 & ~n2164 ) | ( n2519 & n6838 ) | ( ~n2164 & n6838 ) ;
  assign n6840 = n2164 | n6839 ;
  assign n6841 = n3426 | n6840 ;
  assign n6842 = ( n2374 & ~n6841 ) | ( n2374 & 1'b0 ) | ( ~n6841 & 1'b0 ) ;
  assign n6843 = ( n3681 & ~n6836 ) | ( n3681 & n6842 ) | ( ~n6836 & n6842 ) ;
  assign n6844 = ( n1325 & n6836 ) | ( n1325 & n6843 ) | ( n6836 & n6843 ) ;
  assign n6845 = ~n1325 & n6844 ;
  assign n6846 = ( n214 & ~n6811 ) | ( n214 & n6845 ) | ( ~n6811 & n6845 ) ;
  assign n6847 = ~n214 & n6846 ;
  assign n6848 = ( n228 & ~n99 ) | ( n228 & n6847 ) | ( ~n99 & n6847 ) ;
  assign n6849 = ~n228 & n6848 ;
  assign n6850 = ( n351 & ~n492 ) | ( n351 & n6849 ) | ( ~n492 & n6849 ) ;
  assign n6851 = ~n351 & n6850 ;
  assign n6852 = ~n666 & n6851 ;
  assign n6853 = n1063 | n3569 ;
  assign n6854 = ( n260 & ~n61 ) | ( n260 & n6853 ) | ( ~n61 & n6853 ) ;
  assign n6855 = n61 | n6854 ;
  assign n6856 = ( n569 & ~n132 ) | ( n569 & n6855 ) | ( ~n132 & n6855 ) ;
  assign n6857 = n132 | n6856 ;
  assign n6858 = ( n630 & ~n214 ) | ( n630 & n6857 ) | ( ~n214 & n6857 ) ;
  assign n6859 = n214 | n6858 ;
  assign n6860 = n156 | n4075 ;
  assign n6861 = n410 | n6860 ;
  assign n6862 = n491 | n1356 ;
  assign n6863 = ( n4713 & n6861 ) | ( n4713 & n6862 ) | ( n6861 & n6862 ) ;
  assign n6864 = ( n4713 & ~n6863 ) | ( n4713 & 1'b0 ) | ( ~n6863 & 1'b0 ) ;
  assign n6865 = ( n6859 & ~n6864 ) | ( n6859 & n4166 ) | ( ~n6864 & n4166 ) ;
  assign n6866 = ( n2971 & ~n4166 ) | ( n2971 & n6865 ) | ( ~n4166 & n6865 ) ;
  assign n6867 = ( n2971 & ~n6866 ) | ( n2971 & 1'b0 ) | ( ~n6866 & 1'b0 ) ;
  assign n6868 = ( n1626 & ~n2577 ) | ( n1626 & n6867 ) | ( ~n2577 & n6867 ) ;
  assign n6869 = ~n1626 & n6868 ;
  assign n6870 = ( n1428 & ~n1876 ) | ( n1428 & n6869 ) | ( ~n1876 & n6869 ) ;
  assign n6871 = ~n1428 & n6870 ;
  assign n6872 = ( n339 & ~n1426 ) | ( n339 & n6871 ) | ( ~n1426 & n6871 ) ;
  assign n6873 = ~n339 & n6872 ;
  assign n6874 = ( n157 & ~n243 ) | ( n157 & n6873 ) | ( ~n243 & n6873 ) ;
  assign n6875 = ~n157 & n6874 ;
  assign n6876 = ( n138 & ~n415 ) | ( n138 & n6875 ) | ( ~n415 & n6875 ) ;
  assign n6877 = ~n138 & n6876 ;
  assign n6878 = ( n217 & ~n424 ) | ( n217 & n6877 ) | ( ~n424 & n6877 ) ;
  assign n6879 = ~n217 & n6878 ;
  assign n6880 = ( n162 & ~n270 ) | ( n162 & n6879 ) | ( ~n270 & n6879 ) ;
  assign n6881 = ~n162 & n6880 ;
  assign n6883 = ( n3547 & ~n3601 ) | ( n3547 & 1'b0 ) | ( ~n3601 & 1'b0 ) ;
  assign n6884 = n3460 &  n6883 ;
  assign n6885 = n3460 | n6883 ;
  assign n6886 = ~n6884 & n6885 ;
  assign n6891 = ~n3644 & n6886 ;
  assign n6882 = n3460 | n3653 ;
  assign n6887 = ~n3601 & n3657 ;
  assign n6888 = ~n3547 & n3652 ;
  assign n6889 = n6887 | n6888 ;
  assign n6890 = ( n6882 & ~n6889 ) | ( n6882 & 1'b0 ) | ( ~n6889 & 1'b0 ) ;
  assign n6892 = ( n3644 & n6891 ) | ( n3644 & n6890 ) | ( n6891 & n6890 ) ;
  assign n6893 = n6881 | n6892 ;
  assign n6894 = ( n3361 & ~n3460 ) | ( n3361 & n3603 ) | ( ~n3460 & n3603 ) ;
  assign n6895 = ( n3460 & ~n3604 ) | ( n3460 & n6894 ) | ( ~n3604 & n6894 ) ;
  assign n6896 = n3644 | n6895 ;
  assign n6897 = n3460 &  n3657 ;
  assign n6898 = n3361 | n3653 ;
  assign n6899 = ~n3601 & n3652 ;
  assign n6900 = ( n6898 & ~n6899 ) | ( n6898 & 1'b0 ) | ( ~n6899 & 1'b0 ) ;
  assign n6901 = ( n6897 & ~n3657 ) | ( n6897 & n6900 ) | ( ~n3657 & n6900 ) ;
  assign n6902 = n6896 &  n6901 ;
  assign n6903 = ( n6852 & n6893 ) | ( n6852 & n6902 ) | ( n6893 & n6902 ) ;
  assign n6904 = ( n6795 & n6806 ) | ( n6795 & n6903 ) | ( n6806 & n6903 ) ;
  assign n6905 = ( n6748 & ~n6759 ) | ( n6748 & n6904 ) | ( ~n6759 & n6904 ) ;
  assign n6906 = ( n6700 & n6711 ) | ( n6700 & n6905 ) | ( n6711 & n6905 ) ;
  assign n6907 = ( n6649 & n6660 ) | ( n6649 & n6906 ) | ( n6660 & n6906 ) ;
  assign n6611 = ( x2 & ~n6308 ) | ( x2 & n6321 ) | ( ~n6308 & n6321 ) ;
  assign n6612 = ( x2 & ~n6321 ) | ( x2 & n6308 ) | ( ~n6321 & n6308 ) ;
  assign n6613 = ( n6611 & ~x2 ) | ( n6611 & n6612 ) | ( ~x2 & n6612 ) ;
  assign n6908 = n523 | n2995 ;
  assign n6909 = n2839 | n3939 ;
  assign n6910 = n6908 &  n6909 ;
  assign n6911 = n2910 &  n4430 ;
  assign n6912 = ( n6910 & ~n2910 ) | ( n6910 & n6911 ) | ( ~n2910 & n6911 ) ;
  assign n6913 = ( n601 & ~n6912 ) | ( n601 & n6330 ) | ( ~n6912 & n6330 ) ;
  assign n6914 = ( n6330 & ~n6913 ) | ( n6330 & 1'b0 ) | ( ~n6913 & 1'b0 ) ;
  assign n6915 = ( x29 & ~n6912 ) | ( x29 & n6914 ) | ( ~n6912 & n6914 ) ;
  assign n6916 = ( n6912 & ~x29 ) | ( n6912 & n6914 ) | ( ~x29 & n6914 ) ;
  assign n6917 = ( n6915 & ~n6914 ) | ( n6915 & n6916 ) | ( ~n6914 & n6916 ) ;
  assign n6918 = ( n6907 & ~n6613 ) | ( n6907 & n6917 ) | ( ~n6613 & n6917 ) ;
  assign n6919 = ( n6610 & ~n6599 ) | ( n6610 & n6918 ) | ( ~n6599 & n6918 ) ;
  assign n6920 = ( n6597 & ~n6586 ) | ( n6597 & n6919 ) | ( ~n6586 & n6919 ) ;
  assign n6583 = ( n6324 & ~n6327 ) | ( n6324 & n6337 ) | ( ~n6327 & n6337 ) ;
  assign n6584 = ( n6338 & ~n6324 ) | ( n6338 & n6583 ) | ( ~n6324 & n6583 ) ;
  assign n6924 = ~n2751 & n3939 ;
  assign n6921 = n2665 | n4430 ;
  assign n6922 = n523 | n2783 ;
  assign n6923 = n6921 &  n6922 ;
  assign n6925 = ( n2751 & n6924 ) | ( n2751 & n6923 ) | ( n6924 & n6923 ) ;
  assign n6926 = n601 | n6119 ;
  assign n6927 = n6925 &  n6926 ;
  assign n6928 = x29 &  n6927 ;
  assign n6929 = x29 | n6927 ;
  assign n6930 = ~n6928 & n6929 ;
  assign n6931 = ( n6920 & ~n6584 ) | ( n6920 & n6930 ) | ( ~n6584 & n6930 ) ;
  assign n6932 = n6339 | n6348 ;
  assign n6933 = ( n6346 & ~x29 ) | ( n6346 & n6932 ) | ( ~x29 & n6932 ) ;
  assign n6934 = ( x29 & ~n6932 ) | ( x29 & n6346 ) | ( ~n6932 & n6346 ) ;
  assign n6935 = ( n6933 & ~n6346 ) | ( n6933 & n6934 ) | ( ~n6346 & n6934 ) ;
  assign n6939 = ~n2296 & n4962 ;
  assign n6936 = n2483 | n4482 ;
  assign n6937 = n2392 | n4495 ;
  assign n6938 = n6936 &  n6937 ;
  assign n6940 = ( n2296 & n6939 ) | ( n2296 & n6938 ) | ( n6939 & n6938 ) ;
  assign n6941 = n4478 | n5500 ;
  assign n6942 = n6940 &  n6941 ;
  assign n6943 = x26 &  n6942 ;
  assign n6944 = x26 | n6942 ;
  assign n6945 = ~n6943 & n6944 ;
  assign n6946 = ( n6931 & ~n6935 ) | ( n6931 & n6945 ) | ( ~n6935 & n6945 ) ;
  assign n6579 = n6471 | n6480 ;
  assign n6580 = ( x26 & ~n6579 ) | ( x26 & n6478 ) | ( ~n6579 & n6478 ) ;
  assign n6581 = ( n6478 & ~x26 ) | ( n6478 & n6579 ) | ( ~x26 & n6579 ) ;
  assign n6582 = ( n6580 & ~n6478 ) | ( n6580 & n6581 ) | ( ~n6478 & n6581 ) ;
  assign n6947 = n2127 | n5010 ;
  assign n6948 = n2022 | n5067 ;
  assign n6949 = n6947 &  n6948 ;
  assign n6950 = ~n1940 & n5135 ;
  assign n6951 = ( n1940 & n6949 ) | ( n1940 & n6950 ) | ( n6949 & n6950 ) ;
  assign n6952 = n5012 | n5799 ;
  assign n6953 = n6951 &  n6952 ;
  assign n6954 = x23 &  n6953 ;
  assign n6955 = x23 | n6953 ;
  assign n6956 = ~n6954 & n6955 ;
  assign n6957 = ( n6946 & ~n6582 ) | ( n6946 & n6956 ) | ( ~n6582 & n6956 ) ;
  assign n6958 = ( n6576 & n6578 ) | ( n6576 & n6957 ) | ( n6578 & n6957 ) ;
  assign n6563 = n6484 | n6493 ;
  assign n6564 = ( x23 & ~n6563 ) | ( x23 & n6491 ) | ( ~n6563 & n6491 ) ;
  assign n6565 = ( n6491 & ~x23 ) | ( n6491 & n6563 ) | ( ~x23 & n6563 ) ;
  assign n6566 = ( n6564 & ~n6491 ) | ( n6564 & n6565 ) | ( ~n6491 & n6565 ) ;
  assign n6959 = ~n1671 & n5339 ;
  assign n6960 = n1566 | n5761 ;
  assign n6961 = ~n6959 & n6960 ;
  assign n6962 = n1483 &  n5837 ;
  assign n6963 = ( n6961 & ~n1483 ) | ( n6961 & n6962 ) | ( ~n1483 & n6962 ) ;
  assign n6964 = ( n4274 & ~n5341 ) | ( n4274 & 1'b0 ) | ( ~n5341 & 1'b0 ) ;
  assign n6965 = ( n6963 & ~n6964 ) | ( n6963 & 1'b0 ) | ( ~n6964 & 1'b0 ) ;
  assign n6966 = x20 &  n6965 ;
  assign n6967 = x20 | n6965 ;
  assign n6968 = ~n6966 & n6967 ;
  assign n6969 = ( n6958 & ~n6566 ) | ( n6958 & n6968 ) | ( ~n6566 & n6968 ) ;
  assign n6560 = ( n6438 & n6495 ) | ( n6438 & n6505 ) | ( n6495 & n6505 ) ;
  assign n6561 = ( n6438 & ~n6495 ) | ( n6438 & n6505 ) | ( ~n6495 & n6505 ) ;
  assign n6562 = ( n6495 & ~n6560 ) | ( n6495 & n6561 ) | ( ~n6560 & n6561 ) ;
  assign n6970 = n1043 | n6395 ;
  assign n6971 = n1151 | n6170 ;
  assign n6972 = n6970 &  n6971 ;
  assign n6973 = n1267 &  n5970 ;
  assign n6974 = ( n6972 & ~n1267 ) | ( n6972 & n6973 ) | ( ~n1267 & n6973 ) ;
  assign n6975 = n3952 | n5972 ;
  assign n6976 = n6974 &  n6975 ;
  assign n6977 = x17 &  n6976 ;
  assign n6978 = x17 | n6976 ;
  assign n6979 = ~n6977 & n6978 ;
  assign n6980 = ( n6969 & ~n6562 ) | ( n6969 & n6979 ) | ( ~n6562 & n6979 ) ;
  assign n6981 = ( n6557 & n6559 ) | ( n6557 & n6980 ) | ( n6559 & n6980 ) ;
  assign n6991 = n6508 | n6517 ;
  assign n6992 = ( x17 & ~n6991 ) | ( x17 & n6515 ) | ( ~n6991 & n6515 ) ;
  assign n6993 = ( n6515 & ~x17 ) | ( n6515 & n6991 ) | ( ~x17 & n6991 ) ;
  assign n6994 = ( n6992 & ~n6515 ) | ( n6992 & n6993 ) | ( ~n6515 & n6993 ) ;
  assign n6982 = n702 | n6530 ;
  assign n6983 = ~n6522 |  n6525 ;
  assign n6984 = n599 | n6983 ;
  assign n6985 = n6982 &  n6984 ;
  assign n6986 = ( n3937 & n6532 ) | ( n3937 & n6985 ) | ( n6532 & n6985 ) ;
  assign n6987 = ~n6532 & n6986 ;
  assign n6988 = ( x14 & ~n6985 ) | ( x14 & n6987 ) | ( ~n6985 & n6987 ) ;
  assign n6989 = ( n6985 & ~x14 ) | ( n6985 & n6987 ) | ( ~x14 & n6987 ) ;
  assign n6990 = ( n6988 & ~n6987 ) | ( n6988 & n6989 ) | ( ~n6987 & n6989 ) ;
  assign n6995 = ( n6981 & ~n6994 ) | ( n6981 & n6990 ) | ( ~n6994 & n6990 ) ;
  assign n6546 = ( n6519 & n6537 ) | ( n6519 & n6541 ) | ( n6537 & n6541 ) ;
  assign n6545 = ( n6519 & ~n6537 ) | ( n6519 & n6541 ) | ( ~n6537 & n6541 ) ;
  assign n6547 = ( n6537 & ~n6546 ) | ( n6537 & n6545 ) | ( ~n6546 & n6545 ) ;
  assign n7101 = ~n946 & n6530 ;
  assign n7097 = ~n6525 |  n6528 ;
  assign n7098 = n702 | n7097 ;
  assign n7099 = n863 | n6983 ;
  assign n7100 = n7098 &  n7099 ;
  assign n7102 = ( n946 & n7101 ) | ( n946 & n7100 ) | ( n7101 & n7100 ) ;
  assign n7103 = n3650 | n6532 ;
  assign n7104 = n7102 &  n7103 ;
  assign n7105 = ( x14 & ~n7104 ) | ( x14 & 1'b0 ) | ( ~n7104 & 1'b0 ) ;
  assign n6996 = ( n6562 & n6969 ) | ( n6562 & n6979 ) | ( n6969 & n6979 ) ;
  assign n6997 = ( n6562 & ~n6969 ) | ( n6562 & n6979 ) | ( ~n6969 & n6979 ) ;
  assign n6998 = ( n6969 & ~n6996 ) | ( n6969 & n6997 ) | ( ~n6996 & n6997 ) ;
  assign n7002 = ( n6576 & ~n6957 ) | ( n6576 & n6578 ) | ( ~n6957 & n6578 ) ;
  assign n7003 = ( n6578 & ~n6576 ) | ( n6578 & n6957 ) | ( ~n6576 & n6957 ) ;
  assign n7004 = ( n7002 & ~n6578 ) | ( n7002 & n7003 ) | ( ~n6578 & n7003 ) ;
  assign n7008 = ~n1566 & n5837 ;
  assign n7005 = ~n1748 & n5339 ;
  assign n7006 = n1671 | n5761 ;
  assign n7007 = ~n7005 & n7006 ;
  assign n7009 = ( n1566 & n7008 ) | ( n1566 & n7007 ) | ( n7008 & n7007 ) ;
  assign n7010 = ( n5341 & ~n4597 ) | ( n5341 & n7009 ) | ( ~n4597 & n7009 ) ;
  assign n7011 = ~n5341 & n7010 ;
  assign n7012 = ( x20 & ~n7009 ) | ( x20 & n7011 ) | ( ~n7009 & n7011 ) ;
  assign n7013 = ( n7009 & ~x20 ) | ( n7009 & n7011 ) | ( ~x20 & n7011 ) ;
  assign n7014 = ( n7012 & ~n7011 ) | ( n7012 & n7013 ) | ( ~n7011 & n7013 ) ;
  assign n7030 = ~n2392 & n4962 ;
  assign n7027 = n2569 | n4482 ;
  assign n7028 = n2483 | n4495 ;
  assign n7029 = n7027 &  n7028 ;
  assign n7031 = ( n2392 & n7030 ) | ( n2392 & n7029 ) | ( n7030 & n7029 ) ;
  assign n7032 = ( n6212 & ~n4478 ) | ( n6212 & n7031 ) | ( ~n4478 & n7031 ) ;
  assign n7033 = ~n6212 & n7032 ;
  assign n7034 = ( x26 & ~n7031 ) | ( x26 & n7033 ) | ( ~n7031 & n7033 ) ;
  assign n7035 = ( n7031 & ~x26 ) | ( n7031 & n7033 ) | ( ~x26 & n7033 ) ;
  assign n7036 = ( n7034 & ~n7033 ) | ( n7034 & n7035 ) | ( ~n7033 & n7035 ) ;
  assign n7024 = ( n6584 & n6920 ) | ( n6584 & n6930 ) | ( n6920 & n6930 ) ;
  assign n7025 = ( n6584 & ~n6920 ) | ( n6584 & n6930 ) | ( ~n6920 & n6930 ) ;
  assign n7026 = ( n6920 & ~n7024 ) | ( n6920 & n7025 ) | ( ~n7024 & n7025 ) ;
  assign n7043 = n2910 | n523 ;
  assign n7040 = n2751 | n4430 ;
  assign n7041 = n2783 | n3939 ;
  assign n7042 = n7040 &  n7041 ;
  assign n7044 = ( n523 & ~n7043 ) | ( n523 & n7042 ) | ( ~n7043 & n7042 ) ;
  assign n7045 = ( n6226 & ~n601 ) | ( n6226 & n7044 ) | ( ~n601 & n7044 ) ;
  assign n7046 = ~n6226 & n7045 ;
  assign n7047 = ( x29 & ~n7044 ) | ( x29 & n7046 ) | ( ~n7044 & n7046 ) ;
  assign n7048 = ( n7044 & ~x29 ) | ( n7044 & n7046 ) | ( ~x29 & n7046 ) ;
  assign n7049 = ( n7047 & ~n7046 ) | ( n7047 & n7048 ) | ( ~n7046 & n7048 ) ;
  assign n7037 = ( n6586 & n6597 ) | ( n6586 & n6919 ) | ( n6597 & n6919 ) ;
  assign n7038 = ( n6586 & ~n6597 ) | ( n6586 & n6919 ) | ( ~n6597 & n6919 ) ;
  assign n7039 = ( n6597 & ~n7037 ) | ( n6597 & n7038 ) | ( ~n7037 & n7038 ) ;
  assign n7053 = ~n2665 & n4482 ;
  assign n7050 = n2483 | n4962 ;
  assign n7051 = n2569 | n4495 ;
  assign n7052 = n7050 &  n7051 ;
  assign n7054 = ( n2665 & n7053 ) | ( n2665 & n7052 ) | ( n7053 & n7052 ) ;
  assign n7055 = n4478 | n6465 ;
  assign n7056 = n7054 &  n7055 ;
  assign n7057 = x26 &  n7056 ;
  assign n7058 = x26 | n7056 ;
  assign n7059 = ~n7057 & n7058 ;
  assign n7060 = ( n7049 & ~n7039 ) | ( n7049 & n7059 ) | ( ~n7039 & n7059 ) ;
  assign n7061 = ( n7036 & ~n7026 ) | ( n7036 & n7060 ) | ( ~n7026 & n7060 ) ;
  assign n7018 = ~n6931 & n6935 ;
  assign n7019 = ( n6931 & ~n6935 ) | ( n6931 & 1'b0 ) | ( ~n6935 & 1'b0 ) ;
  assign n7020 = n7018 | n7019 ;
  assign n7022 = ( x26 & n6942 ) | ( x26 & n7020 ) | ( n6942 & n7020 ) ;
  assign n7021 = ( n6942 & ~x26 ) | ( n6942 & n7020 ) | ( ~x26 & n7020 ) ;
  assign n7023 = ( x26 & ~n7022 ) | ( x26 & n7021 ) | ( ~n7022 & n7021 ) ;
  assign n7062 = n2178 | n5010 ;
  assign n7063 = n2127 | n5067 ;
  assign n7064 = n7062 &  n7063 ;
  assign n7065 = ~n2022 & n5135 ;
  assign n7066 = ( n2022 & n7064 ) | ( n2022 & n7065 ) | ( n7064 & n7065 ) ;
  assign n7067 = n4934 | n5012 ;
  assign n7068 = n7066 &  n7067 ;
  assign n7069 = x23 &  n7068 ;
  assign n7070 = x23 | n7068 ;
  assign n7071 = ~n7069 & n7070 ;
  assign n7072 = ( n7061 & ~n7023 ) | ( n7061 & n7071 ) | ( ~n7023 & n7071 ) ;
  assign n7015 = ( n6582 & n6946 ) | ( n6582 & n6956 ) | ( n6946 & n6956 ) ;
  assign n7016 = ( n6582 & ~n6946 ) | ( n6582 & n6956 ) | ( ~n6946 & n6956 ) ;
  assign n7017 = ( n6946 & ~n7015 ) | ( n6946 & n7016 ) | ( ~n7015 & n7016 ) ;
  assign n7073 = n1875 &  n5339 ;
  assign n7074 = n1671 | n5837 ;
  assign n7075 = n1748 | n5761 ;
  assign n7076 = n7074 &  n7075 ;
  assign n7077 = ( n7073 & ~n5339 ) | ( n7073 & n7076 ) | ( ~n5339 & n7076 ) ;
  assign n7078 = n4580 | n5341 ;
  assign n7079 = n7077 &  n7078 ;
  assign n7080 = x20 &  n7079 ;
  assign n7081 = x20 | n7079 ;
  assign n7082 = ~n7080 & n7081 ;
  assign n7083 = ( n7072 & ~n7017 ) | ( n7072 & n7082 ) | ( ~n7017 & n7082 ) ;
  assign n7084 = ( n7004 & n7014 ) | ( n7004 & n7083 ) | ( n7014 & n7083 ) ;
  assign n6999 = ( n6566 & n6958 ) | ( n6566 & n6968 ) | ( n6958 & n6968 ) ;
  assign n7000 = ( n6566 & ~n6958 ) | ( n6566 & n6968 ) | ( ~n6958 & n6968 ) ;
  assign n7001 = ( n6958 & ~n6999 ) | ( n6958 & n7000 ) | ( ~n6999 & n7000 ) ;
  assign n7085 = n1151 | n6395 ;
  assign n7086 = n1378 | n5970 ;
  assign n7087 = n7085 &  n7086 ;
  assign n7088 = n1267 &  n6170 ;
  assign n7089 = ( n7087 & ~n1267 ) | ( n7087 & n7088 ) | ( ~n1267 & n7088 ) ;
  assign n7090 = ( n4061 & ~n5972 ) | ( n4061 & 1'b0 ) | ( ~n5972 & 1'b0 ) ;
  assign n7091 = ( n7089 & ~n7090 ) | ( n7089 & 1'b0 ) | ( ~n7090 & 1'b0 ) ;
  assign n7092 = x17 &  n7091 ;
  assign n7093 = x17 | n7091 ;
  assign n7094 = ~n7092 & n7093 ;
  assign n7095 = ( n7084 & ~n7001 ) | ( n7084 & n7094 ) | ( ~n7001 & n7094 ) ;
  assign n7096 = ( n6998 & ~n7095 ) | ( n6998 & 1'b0 ) | ( ~n7095 & 1'b0 ) ;
  assign n7106 = ~n6998 & n7095 ;
  assign n7107 = ( n7104 & ~x14 ) | ( n7104 & n7106 ) | ( ~x14 & n7106 ) ;
  assign n7108 = ( n7105 & ~n7096 ) | ( n7105 & n7107 ) | ( ~n7096 & n7107 ) ;
  assign n7112 = ~n863 & n6530 ;
  assign n7109 = n599 | n7097 ;
  assign n7110 = n702 | n6983 ;
  assign n7111 = n7109 &  n7110 ;
  assign n7113 = ( n863 & n7112 ) | ( n863 & n7111 ) | ( n7112 & n7111 ) ;
  assign n7114 = ( n6532 & ~n4452 ) | ( n6532 & n7113 ) | ( ~n4452 & n7113 ) ;
  assign n7115 = ~n6532 & n7114 ;
  assign n7116 = ( x14 & ~n7113 ) | ( x14 & n7115 ) | ( ~n7113 & n7115 ) ;
  assign n7117 = ( n7113 & ~x14 ) | ( n7113 & n7115 ) | ( ~x14 & n7115 ) ;
  assign n7118 = ( n7116 & ~n7115 ) | ( n7116 & n7117 ) | ( ~n7115 & n7117 ) ;
  assign n7119 = ( n6557 & ~n6980 ) | ( n6557 & n6559 ) | ( ~n6980 & n6559 ) ;
  assign n7120 = ( n6559 & ~n6557 ) | ( n6559 & n6980 ) | ( ~n6557 & n6980 ) ;
  assign n7121 = ( n7119 & ~n6559 ) | ( n7119 & n7120 ) | ( ~n6559 & n7120 ) ;
  assign n7122 = ( n7108 & n7118 ) | ( n7108 & n7121 ) | ( n7118 & n7121 ) ;
  assign n7124 = ( n6981 & n6990 ) | ( n6981 & n6994 ) | ( n6990 & n6994 ) ;
  assign n7123 = ( n6981 & ~n6990 ) | ( n6981 & n6994 ) | ( ~n6990 & n6994 ) ;
  assign n7125 = ( n6990 & ~n7124 ) | ( n6990 & n7123 ) | ( ~n7124 & n7123 ) ;
  assign n7235 = ~n946 & n6983 ;
  assign n7232 = n863 | n7097 ;
  assign n7233 = n1043 | n6530 ;
  assign n7234 = n7232 &  n7233 ;
  assign n7236 = ( n946 & n7235 ) | ( n946 & n7234 ) | ( n7235 & n7234 ) ;
  assign n7237 = n3914 | n6532 ;
  assign n7238 = n7236 &  n7237 ;
  assign n7239 = ( x14 & ~n7238 ) | ( x14 & 1'b0 ) | ( ~n7238 & 1'b0 ) ;
  assign n7126 = ( n7001 & n7084 ) | ( n7001 & n7094 ) | ( n7084 & n7094 ) ;
  assign n7127 = ( n7001 & ~n7084 ) | ( n7001 & n7094 ) | ( ~n7084 & n7094 ) ;
  assign n7128 = ( n7084 & ~n7126 ) | ( n7084 & n7127 ) | ( ~n7126 & n7127 ) ;
  assign n7129 = ( n1483 & ~n5970 ) | ( n1483 & 1'b0 ) | ( ~n5970 & 1'b0 ) ;
  assign n7130 = n1378 | n6170 ;
  assign n7131 = ~n7129 & n7130 ;
  assign n7132 = n1267 &  n6395 ;
  assign n7133 = ( n7131 & ~n1267 ) | ( n7131 & n7132 ) | ( ~n1267 & n7132 ) ;
  assign n7134 = ( n4422 & ~n5972 ) | ( n4422 & 1'b0 ) | ( ~n5972 & 1'b0 ) ;
  assign n7135 = ( n7133 & ~n7134 ) | ( n7133 & 1'b0 ) | ( ~n7134 & 1'b0 ) ;
  assign n7136 = x17 &  n7135 ;
  assign n7137 = x17 | n7135 ;
  assign n7138 = ~n7136 & n7137 ;
  assign n7139 = ( n7004 & ~n7014 ) | ( n7004 & n7083 ) | ( ~n7014 & n7083 ) ;
  assign n7140 = ( n7014 & ~n7084 ) | ( n7014 & n7139 ) | ( ~n7084 & n7139 ) ;
  assign n7153 = ~n2296 & n5010 ;
  assign n7150 = n2127 | n5135 ;
  assign n7151 = n2178 | n5067 ;
  assign n7152 = n7150 &  n7151 ;
  assign n7154 = ( n2296 & n7153 ) | ( n2296 & n7152 ) | ( n7153 & n7152 ) ;
  assign n7155 = n5012 | n5283 ;
  assign n7156 = n7154 &  n7155 ;
  assign n7157 = x23 &  n7156 ;
  assign n7158 = x23 | n7156 ;
  assign n7159 = ~n7157 & n7158 ;
  assign n7160 = ( n7026 & n7036 ) | ( n7026 & n7060 ) | ( n7036 & n7060 ) ;
  assign n7161 = ( n7026 & ~n7036 ) | ( n7026 & n7060 ) | ( ~n7036 & n7060 ) ;
  assign n7162 = ( n7036 & ~n7160 ) | ( n7036 & n7161 ) | ( ~n7160 & n7161 ) ;
  assign n7175 = n2783 | n4430 ;
  assign n7176 = n523 | n2839 ;
  assign n7177 = n7175 &  n7176 ;
  assign n7178 = n2910 &  n3939 ;
  assign n7179 = ( n7177 & ~n2910 ) | ( n7177 & n7178 ) | ( ~n2910 & n7178 ) ;
  assign n7180 = ( n601 & ~n7179 ) | ( n601 & n6104 ) | ( ~n7179 & n6104 ) ;
  assign n7181 = ( n6104 & ~n7180 ) | ( n6104 & 1'b0 ) | ( ~n7180 & 1'b0 ) ;
  assign n7182 = ( x29 & ~n7179 ) | ( x29 & n7181 ) | ( ~n7179 & n7181 ) ;
  assign n7183 = ( n7179 & ~x29 ) | ( n7179 & n7181 ) | ( ~x29 & n7181 ) ;
  assign n7184 = ( n7182 & ~n7181 ) | ( n7182 & n7183 ) | ( ~n7181 & n7183 ) ;
  assign n7172 = ( n6599 & n6610 ) | ( n6599 & n6918 ) | ( n6610 & n6918 ) ;
  assign n7173 = ( n6599 & ~n6610 ) | ( n6599 & n6918 ) | ( ~n6610 & n6918 ) ;
  assign n7174 = ( n6610 & ~n7172 ) | ( n6610 & n7173 ) | ( ~n7172 & n7173 ) ;
  assign n7188 = ~n2751 & n4482 ;
  assign n7185 = n2569 | n4962 ;
  assign n7186 = n2665 | n4495 ;
  assign n7187 = n7185 &  n7186 ;
  assign n7189 = ( n2751 & n7188 ) | ( n2751 & n7187 ) | ( n7188 & n7187 ) ;
  assign n7190 = ( n5705 & ~n4478 ) | ( n5705 & n7189 ) | ( ~n4478 & n7189 ) ;
  assign n7191 = ~n5705 & n7190 ;
  assign n7192 = ( x26 & ~n7189 ) | ( x26 & n7191 ) | ( ~n7189 & n7191 ) ;
  assign n7193 = ( n7189 & ~x26 ) | ( n7189 & n7191 ) | ( ~x26 & n7191 ) ;
  assign n7194 = ( n7192 & ~n7191 ) | ( n7192 & n7193 ) | ( ~n7191 & n7193 ) ;
  assign n7195 = ( n7184 & ~n7174 ) | ( n7184 & n7194 ) | ( ~n7174 & n7194 ) ;
  assign n7164 = n6586 &  n6597 ;
  assign n7163 = ( n6586 & ~n6597 ) | ( n6586 & 1'b0 ) | ( ~n6597 & 1'b0 ) ;
  assign n7165 = ( n6597 & ~n7164 ) | ( n6597 & n7163 ) | ( ~n7164 & n7163 ) ;
  assign n7166 = ( n7049 & ~n6919 ) | ( n7049 & n7165 ) | ( ~n6919 & n7165 ) ;
  assign n7167 = ( n6919 & ~n7049 ) | ( n6919 & n7165 ) | ( ~n7049 & n7165 ) ;
  assign n7168 = ( n7166 & ~n7165 ) | ( n7166 & n7167 ) | ( ~n7165 & n7167 ) ;
  assign n7170 = ( x26 & n7056 ) | ( x26 & n7168 ) | ( n7056 & n7168 ) ;
  assign n7169 = ( n7056 & ~x26 ) | ( n7056 & n7168 ) | ( ~x26 & n7168 ) ;
  assign n7171 = ( x26 & ~n7170 ) | ( x26 & n7169 ) | ( ~n7170 & n7169 ) ;
  assign n7199 = ~n2178 & n5135 ;
  assign n7196 = n2392 | n5010 ;
  assign n7197 = n2296 | n5067 ;
  assign n7198 = n7196 &  n7197 ;
  assign n7200 = ( n2178 & n7199 ) | ( n2178 & n7198 ) | ( n7199 & n7198 ) ;
  assign n7201 = n5012 | n5269 ;
  assign n7202 = n7200 &  n7201 ;
  assign n7203 = x23 &  n7202 ;
  assign n7204 = x23 | n7202 ;
  assign n7205 = ~n7203 & n7204 ;
  assign n7206 = ( n7195 & ~n7171 ) | ( n7195 & n7205 ) | ( ~n7171 & n7205 ) ;
  assign n7207 = ( n7159 & ~n7162 ) | ( n7159 & n7206 ) | ( ~n7162 & n7206 ) ;
  assign n7144 = ( n6945 & n7020 ) | ( n6945 & n7061 ) | ( n7020 & n7061 ) ;
  assign n7145 = ( n7020 & ~n6945 ) | ( n7020 & n7061 ) | ( ~n6945 & n7061 ) ;
  assign n7146 = ( n6945 & ~n7144 ) | ( n6945 & n7145 ) | ( ~n7144 & n7145 ) ;
  assign n7148 = ( x23 & n7068 ) | ( x23 & n7146 ) | ( n7068 & n7146 ) ;
  assign n7147 = ( n7068 & ~x23 ) | ( n7068 & n7146 ) | ( ~x23 & n7146 ) ;
  assign n7149 = ( x23 & ~n7148 ) | ( x23 & n7147 ) | ( ~n7148 & n7147 ) ;
  assign n7208 = ~n1940 & n5339 ;
  assign n7209 = n1875 | n5761 ;
  assign n7210 = ~n7208 & n7209 ;
  assign n7211 = ~n1748 & n5837 ;
  assign n7212 = ( n1748 & n7210 ) | ( n1748 & n7211 ) | ( n7210 & n7211 ) ;
  assign n7213 = n4743 | n5341 ;
  assign n7214 = n7212 &  n7213 ;
  assign n7215 = x20 &  n7214 ;
  assign n7216 = x20 | n7214 ;
  assign n7217 = ~n7215 & n7216 ;
  assign n7218 = ( n7207 & ~n7149 ) | ( n7207 & n7217 ) | ( ~n7149 & n7217 ) ;
  assign n7141 = ( n7017 & n7072 ) | ( n7017 & n7082 ) | ( n7072 & n7082 ) ;
  assign n7142 = ( n7017 & ~n7072 ) | ( n7017 & n7082 ) | ( ~n7072 & n7082 ) ;
  assign n7143 = ( n7072 & ~n7141 ) | ( n7072 & n7142 ) | ( ~n7141 & n7142 ) ;
  assign n7219 = n1378 | n6395 ;
  assign n7220 = n1566 | n5970 ;
  assign n7221 = n7219 &  n7220 ;
  assign n7222 = n1483 &  n6170 ;
  assign n7223 = ( n7221 & ~n1483 ) | ( n7221 & n7222 ) | ( ~n1483 & n7222 ) ;
  assign n7224 = ( n5038 & ~n5972 ) | ( n5038 & 1'b0 ) | ( ~n5972 & 1'b0 ) ;
  assign n7225 = ( n7223 & ~n7224 ) | ( n7223 & 1'b0 ) | ( ~n7224 & 1'b0 ) ;
  assign n7226 = x17 &  n7225 ;
  assign n7227 = x17 | n7225 ;
  assign n7228 = ~n7226 & n7227 ;
  assign n7229 = ( n7218 & ~n7143 ) | ( n7218 & n7228 ) | ( ~n7143 & n7228 ) ;
  assign n7230 = ( n7138 & n7140 ) | ( n7138 & n7229 ) | ( n7140 & n7229 ) ;
  assign n7231 = ( n7128 & ~n7230 ) | ( n7128 & 1'b0 ) | ( ~n7230 & 1'b0 ) ;
  assign n7240 = ~n7128 & n7230 ;
  assign n7241 = ( n7238 & ~x14 ) | ( n7238 & n7240 ) | ( ~x14 & n7240 ) ;
  assign n7242 = ( n7239 & ~n7231 ) | ( n7239 & n7241 ) | ( ~n7231 & n7241 ) ;
  assign n7261 = n7096 | n7106 ;
  assign n7262 = ( x14 & ~n7261 ) | ( x14 & n7104 ) | ( ~n7261 & n7104 ) ;
  assign n7263 = ( n7104 & ~x14 ) | ( n7104 & n7261 ) | ( ~x14 & n7261 ) ;
  assign n7264 = ( n7262 & ~n7104 ) | ( n7262 & n7263 ) | ( ~n7104 & n7263 ) ;
  assign n7243 = ~x9 & x10 ;
  assign n7244 = ( x9 & ~x10 ) | ( x9 & 1'b0 ) | ( ~x10 & 1'b0 ) ;
  assign n7245 = n7243 | n7244 ;
  assign n7249 = ( x8 & ~x9 ) | ( x8 & 1'b0 ) | ( ~x9 & 1'b0 ) ;
  assign n7250 = ~x8 & x9 ;
  assign n7251 = n7249 | n7250 ;
  assign n7246 = ( x10 & ~x11 ) | ( x10 & 1'b0 ) | ( ~x11 & 1'b0 ) ;
  assign n7247 = ~x10 & x11 ;
  assign n7248 = n7246 | n7247 ;
  assign n7252 = ( n7245 & ~n7251 ) | ( n7245 & n7248 ) | ( ~n7251 & n7248 ) ;
  assign n7253 = ~n7245 & n7252 ;
  assign n7254 = ~n599 & n7253 ;
  assign n7255 = ~n7248 | ~n7251 ;
  assign n7256 = ( n7254 & ~n3637 ) | ( n7254 & n7255 ) | ( ~n3637 & n7255 ) ;
  assign n7257 = n3637 | n7256 ;
  assign n7258 = ( x11 & ~n7254 ) | ( x11 & n7257 ) | ( ~n7254 & n7257 ) ;
  assign n7259 = ( n7254 & ~x11 ) | ( n7254 & n7257 ) | ( ~x11 & n7257 ) ;
  assign n7260 = ( n7258 & ~n7257 ) | ( n7258 & n7259 ) | ( ~n7257 & n7259 ) ;
  assign n7265 = ( n7242 & ~n7264 ) | ( n7242 & n7260 ) | ( ~n7264 & n7260 ) ;
  assign n7266 = ( n7108 & ~n7118 ) | ( n7108 & n7121 ) | ( ~n7118 & n7121 ) ;
  assign n7267 = ( n7118 & ~n7122 ) | ( n7118 & n7266 ) | ( ~n7122 & n7266 ) ;
  assign n7271 = ( n7138 & ~n7229 ) | ( n7138 & n7140 ) | ( ~n7229 & n7140 ) ;
  assign n7272 = ( n7140 & ~n7138 ) | ( n7140 & n7229 ) | ( ~n7138 & n7229 ) ;
  assign n7273 = ( n7271 & ~n7140 ) | ( n7271 & n7272 ) | ( ~n7140 & n7272 ) ;
  assign n7277 = ~n946 & n7097 ;
  assign n7274 = n1151 | n6530 ;
  assign n7275 = n1043 | n6983 ;
  assign n7276 = n7274 &  n7275 ;
  assign n7278 = ( n946 & n7277 ) | ( n946 & n7276 ) | ( n7277 & n7276 ) ;
  assign n7279 = ( n6532 & ~n4038 ) | ( n6532 & n7278 ) | ( ~n4038 & n7278 ) ;
  assign n7280 = ~n6532 & n7279 ;
  assign n7281 = ( x14 & ~n7278 ) | ( x14 & n7280 ) | ( ~n7278 & n7280 ) ;
  assign n7282 = ( n7278 & ~x14 ) | ( n7278 & n7280 ) | ( ~x14 & n7280 ) ;
  assign n7283 = ( n7281 & ~n7280 ) | ( n7281 & n7282 ) | ( ~n7280 & n7282 ) ;
  assign n7299 = ~n1875 & n5837 ;
  assign n7296 = ~n2022 & n5339 ;
  assign n7297 = n1940 | n5761 ;
  assign n7298 = ~n7296 & n7297 ;
  assign n7300 = ( n1875 & n7299 ) | ( n1875 & n7298 ) | ( n7299 & n7298 ) ;
  assign n7301 = ( n5341 & ~n5381 ) | ( n5341 & n7300 ) | ( ~n5381 & n7300 ) ;
  assign n7302 = ~n5341 & n7301 ;
  assign n7303 = ( x20 & ~n7300 ) | ( x20 & n7302 ) | ( ~n7300 & n7302 ) ;
  assign n7304 = ( n7300 & ~x20 ) | ( n7300 & n7302 ) | ( ~x20 & n7302 ) ;
  assign n7305 = ( n7303 & ~n7302 ) | ( n7303 & n7304 ) | ( ~n7302 & n7304 ) ;
  assign n7293 = ( n7162 & ~n7159 ) | ( n7162 & n7206 ) | ( ~n7159 & n7206 ) ;
  assign n7294 = ( n7159 & ~n7206 ) | ( n7159 & n7162 ) | ( ~n7206 & n7162 ) ;
  assign n7295 = ( n7293 & ~n7162 ) | ( n7293 & n7294 ) | ( ~n7162 & n7294 ) ;
  assign n7315 = ( n6660 & ~n6649 ) | ( n6660 & n6906 ) | ( ~n6649 & n6906 ) ;
  assign n7316 = ( n6649 & ~n6906 ) | ( n6649 & n6660 ) | ( ~n6906 & n6660 ) ;
  assign n7317 = ( n7315 & ~n6660 ) | ( n7315 & n7316 ) | ( ~n6660 & n7316 ) ;
  assign n7321 = ~n2839 & n4430 ;
  assign n7318 = n523 | n3030 ;
  assign n7319 = n2995 | n3939 ;
  assign n7320 = n7318 &  n7319 ;
  assign n7322 = ( n2839 & n7321 ) | ( n2839 & n7320 ) | ( n7321 & n7320 ) ;
  assign n7323 = ~n3610 & n6591 ;
  assign n7324 = n6592 | n7323 ;
  assign n7325 = ( n7322 & ~n601 ) | ( n7322 & n7324 ) | ( ~n601 & n7324 ) ;
  assign n7326 = ~n7324 & n7325 ;
  assign n7327 = ( x29 & ~n7322 ) | ( x29 & n7326 ) | ( ~n7322 & n7326 ) ;
  assign n7328 = ( n7322 & ~x29 ) | ( n7322 & n7326 ) | ( ~x29 & n7326 ) ;
  assign n7329 = ( n7327 & ~n7326 ) | ( n7327 & n7328 ) | ( ~n7326 & n7328 ) ;
  assign n7330 = ( n6711 & ~n6700 ) | ( n6711 & n6905 ) | ( ~n6700 & n6905 ) ;
  assign n7331 = ( n6700 & ~n6905 ) | ( n6700 & n6711 ) | ( ~n6905 & n6711 ) ;
  assign n7332 = ( n7330 & ~n6711 ) | ( n7330 & n7331 ) | ( ~n6711 & n7331 ) ;
  assign n7333 = n523 | n3106 ;
  assign n7334 = n3030 | n3939 ;
  assign n7335 = n7333 &  n7334 ;
  assign n7336 = ~n2995 & n4430 ;
  assign n7337 = ( n2995 & n7335 ) | ( n2995 & n7336 ) | ( n7335 & n7336 ) ;
  assign n7338 = ~n3609 & n6604 ;
  assign n7339 = n6605 | n7338 ;
  assign n7340 = ( n7337 & ~n601 ) | ( n7337 & n7339 ) | ( ~n601 & n7339 ) ;
  assign n7341 = ~n7339 & n7340 ;
  assign n7342 = ( x29 & ~n7337 ) | ( x29 & n7341 ) | ( ~n7337 & n7341 ) ;
  assign n7343 = ( n7337 & ~x29 ) | ( n7337 & n7341 ) | ( ~x29 & n7341 ) ;
  assign n7344 = ( n7342 & ~n7341 ) | ( n7342 & n7343 ) | ( ~n7341 & n7343 ) ;
  assign n7348 = ~n3030 & n4430 ;
  assign n7345 = n523 | n3197 ;
  assign n7346 = n3106 | n3939 ;
  assign n7347 = n7345 &  n7346 ;
  assign n7349 = ( n3030 & n7348 ) | ( n3030 & n7347 ) | ( n7348 & n7347 ) ;
  assign n7350 = ( n6314 & ~n601 ) | ( n6314 & n7349 ) | ( ~n601 & n7349 ) ;
  assign n7351 = ~n6314 & n7350 ;
  assign n7352 = ( x29 & ~n7349 ) | ( x29 & n7351 ) | ( ~n7349 & n7351 ) ;
  assign n7353 = ( n7349 & ~x29 ) | ( n7349 & n7351 ) | ( ~x29 & n7351 ) ;
  assign n7354 = ( n7352 & ~n7351 ) | ( n7352 & n7353 ) | ( ~n7351 & n7353 ) ;
  assign n7355 = ( n6748 & n6759 ) | ( n6748 & n6904 ) | ( n6759 & n6904 ) ;
  assign n7356 = ( n6759 & ~n7355 ) | ( n6759 & n6905 ) | ( ~n7355 & n6905 ) ;
  assign n7360 = n3266 | n523 ;
  assign n7357 = n3106 | n4430 ;
  assign n7358 = n3197 | n3939 ;
  assign n7359 = n7357 &  n7358 ;
  assign n7361 = ( n523 & ~n7360 ) | ( n523 & n7359 ) | ( ~n7360 & n7359 ) ;
  assign n7362 = ~n3607 & n6654 ;
  assign n7363 = n6655 | n7362 ;
  assign n7364 = ( n7361 & ~n601 ) | ( n7361 & n7363 ) | ( ~n601 & n7363 ) ;
  assign n7365 = ~n7363 & n7364 ;
  assign n7366 = ( x29 & ~n7361 ) | ( x29 & n7365 ) | ( ~n7361 & n7365 ) ;
  assign n7367 = ( n7361 & ~x29 ) | ( n7361 & n7365 ) | ( ~x29 & n7365 ) ;
  assign n7368 = ( n7366 & ~n7365 ) | ( n7366 & n7367 ) | ( ~n7365 & n7367 ) ;
  assign n7369 = ( n6795 & ~n6806 ) | ( n6795 & n6903 ) | ( ~n6806 & n6903 ) ;
  assign n7370 = ( n6806 & ~n6904 ) | ( n6806 & n7369 ) | ( ~n6904 & n7369 ) ;
  assign n7371 = n3197 | n4430 ;
  assign n7372 = n523 | n3325 ;
  assign n7373 = n7371 &  n7372 ;
  assign n7374 = n3266 &  n3939 ;
  assign n7375 = ( n7373 & ~n3266 ) | ( n7373 & n7374 ) | ( ~n3266 & n7374 ) ;
  assign n7376 = n3606 | n6705 ;
  assign n7377 = ~n6706 & n7376 ;
  assign n7378 = ( n601 & ~n7375 ) | ( n601 & n7377 ) | ( ~n7375 & n7377 ) ;
  assign n7379 = ( n7377 & ~n7378 ) | ( n7377 & 1'b0 ) | ( ~n7378 & 1'b0 ) ;
  assign n7380 = ( x29 & ~n7375 ) | ( x29 & n7379 ) | ( ~n7375 & n7379 ) ;
  assign n7381 = ( n7375 & ~x29 ) | ( n7375 & n7379 ) | ( ~x29 & n7379 ) ;
  assign n7382 = ( n7380 & ~n7379 ) | ( n7380 & n7381 ) | ( ~n7379 & n7381 ) ;
  assign n7383 = ( n6893 & ~n6852 ) | ( n6893 & n6902 ) | ( ~n6852 & n6902 ) ;
  assign n7384 = ( n6852 & ~n6903 ) | ( n6852 & n7383 ) | ( ~n6903 & n7383 ) ;
  assign n7385 = n523 | n3361 ;
  assign n7386 = n3325 | n3939 ;
  assign n7387 = n7385 &  n7386 ;
  assign n7388 = n3266 &  n4430 ;
  assign n7389 = ( n7387 & ~n3266 ) | ( n7387 & n7388 ) | ( ~n3266 & n7388 ) ;
  assign n7390 = n3605 | n6753 ;
  assign n7391 = ~n6754 & n7390 ;
  assign n7392 = ( n601 & ~n7389 ) | ( n601 & n7391 ) | ( ~n7389 & n7391 ) ;
  assign n7393 = ( n7391 & ~n7392 ) | ( n7391 & 1'b0 ) | ( ~n7392 & 1'b0 ) ;
  assign n7394 = ( x29 & ~n7389 ) | ( x29 & n7393 ) | ( ~n7389 & n7393 ) ;
  assign n7395 = ( n7389 & ~x29 ) | ( n7389 & n7393 ) | ( ~x29 & n7393 ) ;
  assign n7396 = ( n7394 & ~n7393 ) | ( n7394 & n7395 ) | ( ~n7393 & n7395 ) ;
  assign n7397 = ( n6881 & ~n6892 ) | ( n6881 & 1'b0 ) | ( ~n6892 & 1'b0 ) ;
  assign n7398 = ( n6893 & ~n6881 ) | ( n6893 & n7397 ) | ( ~n6881 & n7397 ) ;
  assign n7402 = ~n523 & n3460 ;
  assign n7399 = n3325 | n4430 ;
  assign n7400 = n3361 | n3939 ;
  assign n7401 = n7399 &  n7400 ;
  assign n7403 = ( n523 & n7402 ) | ( n523 & n7401 ) | ( n7402 & n7401 ) ;
  assign n7404 = ~n3604 & n6800 ;
  assign n7405 = n6801 | n7404 ;
  assign n7406 = ( n7403 & ~n601 ) | ( n7403 & n7405 ) | ( ~n601 & n7405 ) ;
  assign n7407 = ~n7405 & n7406 ;
  assign n7408 = ( x29 & ~n7403 ) | ( x29 & n7407 ) | ( ~n7403 & n7407 ) ;
  assign n7409 = ( n7403 & ~x29 ) | ( n7403 & n7407 ) | ( ~x29 & n7407 ) ;
  assign n7410 = ( n7408 & ~n7407 ) | ( n7408 & n7409 ) | ( ~n7407 & n7409 ) ;
  assign n7418 = ~n3547 & n3643 ;
  assign n7439 = ~n3460 & n3939 ;
  assign n7436 = n3361 | n4430 ;
  assign n7437 = n523 | n3601 ;
  assign n7438 = n7436 &  n7437 ;
  assign n7440 = ( n3460 & n7439 ) | ( n3460 & n7438 ) | ( n7439 & n7438 ) ;
  assign n7441 = ( n6895 & ~n601 ) | ( n6895 & n7440 ) | ( ~n601 & n7440 ) ;
  assign n7442 = ~n6895 & n7441 ;
  assign n7443 = ( x29 & ~n7440 ) | ( x29 & n7442 ) | ( ~n7440 & n7442 ) ;
  assign n7444 = ( n7440 & ~x29 ) | ( n7440 & n7442 ) | ( ~x29 & n7442 ) ;
  assign n7445 = ( n7443 & ~n7442 ) | ( n7443 & n7444 ) | ( ~n7442 & n7444 ) ;
  assign n7432 = ~n601 & n6886 ;
  assign n7430 = ~n3460 & n4430 ;
  assign n7427 = n523 | n3547 ;
  assign n7428 = n3601 | n3939 ;
  assign n7429 = n7427 &  n7428 ;
  assign n7431 = ( n3460 & n7430 ) | ( n3460 & n7429 ) | ( n7430 & n7429 ) ;
  assign n7433 = ( n601 & n7432 ) | ( n601 & n7431 ) | ( n7432 & n7431 ) ;
  assign n7411 = ~n3547 & n3601 ;
  assign n7412 = n6883 | n7411 ;
  assign n7422 = n7412 | n601 ;
  assign n7419 = n3547 | n3939 ;
  assign n7420 = n3601 | n4430 ;
  assign n7421 = n7419 &  n7420 ;
  assign n7423 = ( n601 & ~n7422 ) | ( n601 & n7421 ) | ( ~n7422 & n7421 ) ;
  assign n7424 = ( n521 & ~n3547 ) | ( n521 & 1'b0 ) | ( ~n3547 & 1'b0 ) ;
  assign n7425 = ( x29 & ~n7423 ) | ( x29 & n7424 ) | ( ~n7423 & n7424 ) ;
  assign n7434 = ( x29 & ~n7433 ) | ( x29 & n7425 ) | ( ~n7433 & n7425 ) ;
  assign n7435 = ( x29 & ~n7434 ) | ( x29 & 1'b0 ) | ( ~n7434 & 1'b0 ) ;
  assign n7446 = ( n7418 & ~n7445 ) | ( n7418 & n7435 ) | ( ~n7445 & n7435 ) ;
  assign n7416 = n7412 | n3644 ;
  assign n7413 = ~n3547 & n3657 ;
  assign n7414 = n3601 | n3653 ;
  assign n7415 = ~n7413 & n7414 ;
  assign n7417 = ( n3644 & ~n7416 ) | ( n3644 & n7415 ) | ( ~n7416 & n7415 ) ;
  assign n7447 = ( n7410 & ~n7446 ) | ( n7410 & n7417 ) | ( ~n7446 & n7417 ) ;
  assign n7448 = ( n7396 & ~n7398 ) | ( n7396 & n7447 ) | ( ~n7398 & n7447 ) ;
  assign n7449 = ( n7382 & n7384 ) | ( n7382 & n7448 ) | ( n7384 & n7448 ) ;
  assign n7450 = ( n7368 & n7370 ) | ( n7368 & n7449 ) | ( n7370 & n7449 ) ;
  assign n7451 = ( n7354 & ~n7356 ) | ( n7354 & n7450 ) | ( ~n7356 & n7450 ) ;
  assign n7452 = ( n7332 & n7344 ) | ( n7332 & n7451 ) | ( n7344 & n7451 ) ;
  assign n7453 = ( n7317 & n7329 ) | ( n7317 & n7452 ) | ( n7329 & n7452 ) ;
  assign n7454 = n6613 | n6907 ;
  assign n7455 = n6613 &  n6907 ;
  assign n7456 = ( n7454 & ~n7455 ) | ( n7454 & 1'b0 ) | ( ~n7455 & 1'b0 ) ;
  assign n7457 = ~n6917 & n7456 ;
  assign n7458 = n6917 | n7456 ;
  assign n7459 = ( n7457 & ~n7456 ) | ( n7457 & n7458 ) | ( ~n7456 & n7458 ) ;
  assign n7463 = ~n2751 & n4495 ;
  assign n7460 = n2665 | n4962 ;
  assign n7461 = n2783 | n4482 ;
  assign n7462 = n7460 &  n7461 ;
  assign n7464 = ( n2751 & n7463 ) | ( n2751 & n7462 ) | ( n7463 & n7462 ) ;
  assign n7465 = n4478 | n6119 ;
  assign n7466 = n7464 &  n7465 ;
  assign n7467 = x26 &  n7466 ;
  assign n7468 = x26 | n7466 ;
  assign n7469 = ~n7467 & n7468 ;
  assign n7470 = ( n7453 & ~n7459 ) | ( n7453 & n7469 ) | ( ~n7459 & n7469 ) ;
  assign n7312 = ( n7174 & n7184 ) | ( n7174 & n7194 ) | ( n7184 & n7194 ) ;
  assign n7313 = ( n7174 & ~n7184 ) | ( n7174 & n7194 ) | ( ~n7184 & n7194 ) ;
  assign n7314 = ( n7184 & ~n7312 ) | ( n7184 & n7313 ) | ( ~n7312 & n7313 ) ;
  assign n7474 = ~n2296 & n5135 ;
  assign n7471 = n2483 | n5010 ;
  assign n7472 = n2392 | n5067 ;
  assign n7473 = n7471 &  n7472 ;
  assign n7475 = ( n2296 & n7474 ) | ( n2296 & n7473 ) | ( n7474 & n7473 ) ;
  assign n7476 = ( n5500 & ~n5012 ) | ( n5500 & n7475 ) | ( ~n5012 & n7475 ) ;
  assign n7477 = ~n5500 & n7476 ;
  assign n7478 = ( x23 & ~n7475 ) | ( x23 & n7477 ) | ( ~n7475 & n7477 ) ;
  assign n7479 = ( n7475 & ~x23 ) | ( n7475 & n7477 ) | ( ~x23 & n7477 ) ;
  assign n7480 = ( n7478 & ~n7477 ) | ( n7478 & n7479 ) | ( ~n7477 & n7479 ) ;
  assign n7481 = ( n7470 & ~n7314 ) | ( n7470 & n7480 ) | ( ~n7314 & n7480 ) ;
  assign n7306 = ( n7059 & n7168 ) | ( n7059 & n7195 ) | ( n7168 & n7195 ) ;
  assign n7307 = ( n7168 & ~n7059 ) | ( n7168 & n7195 ) | ( ~n7059 & n7195 ) ;
  assign n7308 = ( n7059 & ~n7306 ) | ( n7059 & n7307 ) | ( ~n7306 & n7307 ) ;
  assign n7310 = ( x23 & n7202 ) | ( x23 & n7308 ) | ( n7202 & n7308 ) ;
  assign n7309 = ( n7202 & ~x23 ) | ( n7202 & n7308 ) | ( ~x23 & n7308 ) ;
  assign n7311 = ( x23 & ~n7310 ) | ( x23 & n7309 ) | ( ~n7310 & n7309 ) ;
  assign n7482 = ~n2127 & n5339 ;
  assign n7483 = n2022 | n5761 ;
  assign n7484 = ~n7482 & n7483 ;
  assign n7485 = ~n1940 & n5837 ;
  assign n7486 = ( n1940 & n7484 ) | ( n1940 & n7485 ) | ( n7484 & n7485 ) ;
  assign n7487 = n5341 | n5799 ;
  assign n7488 = n7486 &  n7487 ;
  assign n7489 = x20 &  n7488 ;
  assign n7490 = x20 | n7488 ;
  assign n7491 = ~n7489 & n7490 ;
  assign n7492 = ( n7481 & ~n7311 ) | ( n7481 & n7491 ) | ( ~n7311 & n7491 ) ;
  assign n7493 = ( n7305 & ~n7295 ) | ( n7305 & n7492 ) | ( ~n7295 & n7492 ) ;
  assign n7287 = ( n7071 & n7146 ) | ( n7071 & n7207 ) | ( n7146 & n7207 ) ;
  assign n7288 = ( n7146 & ~n7071 ) | ( n7146 & n7207 ) | ( ~n7071 & n7207 ) ;
  assign n7289 = ( n7071 & ~n7287 ) | ( n7071 & n7288 ) | ( ~n7287 & n7288 ) ;
  assign n7291 = ( x20 & n7214 ) | ( x20 & n7289 ) | ( n7214 & n7289 ) ;
  assign n7290 = ( n7214 & ~x20 ) | ( n7214 & n7289 ) | ( ~x20 & n7289 ) ;
  assign n7292 = ( x20 & ~n7291 ) | ( x20 & n7290 ) | ( ~n7291 & n7290 ) ;
  assign n7494 = n1671 | n5970 ;
  assign n7495 = n1566 | n6170 ;
  assign n7496 = n7494 &  n7495 ;
  assign n7497 = n1483 &  n6395 ;
  assign n7498 = ( n7496 & ~n1483 ) | ( n7496 & n7497 ) | ( ~n1483 & n7497 ) ;
  assign n7499 = ( n4274 & ~n5972 ) | ( n4274 & 1'b0 ) | ( ~n5972 & 1'b0 ) ;
  assign n7500 = ( n7498 & ~n7499 ) | ( n7498 & 1'b0 ) | ( ~n7499 & 1'b0 ) ;
  assign n7501 = x17 &  n7500 ;
  assign n7502 = x17 | n7500 ;
  assign n7503 = ~n7501 & n7502 ;
  assign n7504 = ( n7493 & ~n7292 ) | ( n7493 & n7503 ) | ( ~n7292 & n7503 ) ;
  assign n7284 = ( n7143 & n7218 ) | ( n7143 & n7228 ) | ( n7218 & n7228 ) ;
  assign n7285 = ( n7143 & ~n7218 ) | ( n7143 & n7228 ) | ( ~n7218 & n7228 ) ;
  assign n7286 = ( n7218 & ~n7284 ) | ( n7218 & n7285 ) | ( ~n7284 & n7285 ) ;
  assign n7505 = n1043 | n7097 ;
  assign n7506 = n1151 | n6983 ;
  assign n7507 = n7505 &  n7506 ;
  assign n7508 = n1267 &  n6530 ;
  assign n7509 = ( n7507 & ~n1267 ) | ( n7507 & n7508 ) | ( ~n1267 & n7508 ) ;
  assign n7510 = n3952 | n6532 ;
  assign n7511 = n7509 &  n7510 ;
  assign n7512 = x14 &  n7511 ;
  assign n7513 = x14 | n7511 ;
  assign n7514 = ~n7512 & n7513 ;
  assign n7515 = ( n7504 & ~n7286 ) | ( n7504 & n7514 ) | ( ~n7286 & n7514 ) ;
  assign n7516 = ( n7273 & n7283 ) | ( n7273 & n7515 ) | ( n7283 & n7515 ) ;
  assign n7526 = n7231 | n7240 ;
  assign n7527 = ( x14 & ~n7526 ) | ( x14 & n7238 ) | ( ~n7526 & n7238 ) ;
  assign n7528 = ( n7238 & ~x14 ) | ( n7238 & n7526 ) | ( ~x14 & n7526 ) ;
  assign n7529 = ( n7527 & ~n7238 ) | ( n7527 & n7528 ) | ( ~n7238 & n7528 ) ;
  assign n7517 = ~n702 & n7253 ;
  assign n7518 = ~n7245 |  n7251 ;
  assign n7519 = n599 | n7518 ;
  assign n7520 = ~n7517 & n7519 ;
  assign n7521 = ( n3937 & n7255 ) | ( n3937 & n7520 ) | ( n7255 & n7520 ) ;
  assign n7522 = ~n7255 & n7521 ;
  assign n7523 = ( x11 & ~n7520 ) | ( x11 & n7522 ) | ( ~n7520 & n7522 ) ;
  assign n7524 = ( n7520 & ~x11 ) | ( n7520 & n7522 ) | ( ~x11 & n7522 ) ;
  assign n7525 = ( n7523 & ~n7522 ) | ( n7523 & n7524 ) | ( ~n7522 & n7524 ) ;
  assign n7530 = ( n7516 & ~n7529 ) | ( n7516 & n7525 ) | ( ~n7529 & n7525 ) ;
  assign n7269 = ( n7242 & n7260 ) | ( n7242 & n7264 ) | ( n7260 & n7264 ) ;
  assign n7268 = ( n7242 & ~n7260 ) | ( n7242 & n7264 ) | ( ~n7260 & n7264 ) ;
  assign n7270 = ( n7260 & ~n7269 ) | ( n7260 & n7268 ) | ( ~n7269 & n7268 ) ;
  assign n7782 = n946 &  n7253 ;
  assign n7783 = ~n7251 |  n7248 ;
  assign n7784 = n702 | n7783 ;
  assign n7785 = n863 | n7518 ;
  assign n7786 = n7784 &  n7785 ;
  assign n7787 = ( n7782 & ~n7253 ) | ( n7782 & n7786 ) | ( ~n7253 & n7786 ) ;
  assign n7788 = n3650 | n7255 ;
  assign n7789 = n7787 &  n7788 ;
  assign n7790 = ( x11 & ~n7789 ) | ( x11 & 1'b0 ) | ( ~n7789 & 1'b0 ) ;
  assign n7531 = ( n7286 & n7504 ) | ( n7286 & n7514 ) | ( n7504 & n7514 ) ;
  assign n7532 = ( n7286 & ~n7504 ) | ( n7286 & n7514 ) | ( ~n7504 & n7514 ) ;
  assign n7533 = ( n7504 & ~n7531 ) | ( n7504 & n7532 ) | ( ~n7531 & n7532 ) ;
  assign n7543 = ~n1566 & n6395 ;
  assign n7540 = n1748 | n5970 ;
  assign n7541 = n1671 | n6170 ;
  assign n7542 = n7540 &  n7541 ;
  assign n7544 = ( n1566 & n7543 ) | ( n1566 & n7542 ) | ( n7543 & n7542 ) ;
  assign n7545 = n4597 | n5972 ;
  assign n7546 = n7544 &  n7545 ;
  assign n7547 = x17 &  n7546 ;
  assign n7548 = x17 | n7546 ;
  assign n7549 = ~n7547 & n7548 ;
  assign n7550 = ( n7295 & ~n7492 ) | ( n7295 & n7305 ) | ( ~n7492 & n7305 ) ;
  assign n7551 = ( n7493 & ~n7305 ) | ( n7493 & n7550 ) | ( ~n7305 & n7550 ) ;
  assign n7561 = ( n7329 & ~n7317 ) | ( n7329 & n7452 ) | ( ~n7317 & n7452 ) ;
  assign n7562 = ( n7317 & ~n7452 ) | ( n7317 & n7329 ) | ( ~n7452 & n7329 ) ;
  assign n7563 = ( n7561 & ~n7329 ) | ( n7561 & n7562 ) | ( ~n7329 & n7562 ) ;
  assign n7564 = n2751 | n4962 ;
  assign n7565 = n2783 | n4495 ;
  assign n7566 = n7564 &  n7565 ;
  assign n7567 = n2910 &  n4482 ;
  assign n7568 = ( n7566 & ~n2910 ) | ( n7566 & n7567 ) | ( ~n2910 & n7567 ) ;
  assign n7569 = ( n6226 & ~n4478 ) | ( n6226 & n7568 ) | ( ~n4478 & n7568 ) ;
  assign n7570 = ~n6226 & n7569 ;
  assign n7571 = ( x26 & ~n7568 ) | ( x26 & n7570 ) | ( ~n7568 & n7570 ) ;
  assign n7572 = ( n7568 & ~x26 ) | ( n7568 & n7570 ) | ( ~x26 & n7570 ) ;
  assign n7573 = ( n7571 & ~n7570 ) | ( n7571 & n7572 ) | ( ~n7570 & n7572 ) ;
  assign n7574 = ( n7344 & ~n7332 ) | ( n7344 & n7451 ) | ( ~n7332 & n7451 ) ;
  assign n7575 = ( n7332 & ~n7451 ) | ( n7332 & n7344 ) | ( ~n7451 & n7344 ) ;
  assign n7576 = ( n7574 & ~n7344 ) | ( n7574 & n7575 ) | ( ~n7344 & n7575 ) ;
  assign n7577 = n2783 | n4962 ;
  assign n7578 = n2839 | n4482 ;
  assign n7579 = n7577 &  n7578 ;
  assign n7580 = n2910 &  n4495 ;
  assign n7581 = ( n7579 & ~n2910 ) | ( n7579 & n7580 ) | ( ~n2910 & n7580 ) ;
  assign n7582 = ( n4478 & ~n7581 ) | ( n4478 & n6104 ) | ( ~n7581 & n6104 ) ;
  assign n7583 = ( n6104 & ~n7582 ) | ( n6104 & 1'b0 ) | ( ~n7582 & 1'b0 ) ;
  assign n7584 = ( x26 & ~n7581 ) | ( x26 & n7583 ) | ( ~n7581 & n7583 ) ;
  assign n7585 = ( n7581 & ~x26 ) | ( n7581 & n7583 ) | ( ~x26 & n7583 ) ;
  assign n7586 = ( n7584 & ~n7583 ) | ( n7584 & n7585 ) | ( ~n7583 & n7585 ) ;
  assign n7590 = n2995 | n4482 ;
  assign n7591 = n2839 | n4495 ;
  assign n7592 = n7590 &  n7591 ;
  assign n7593 = n2910 &  n4962 ;
  assign n7594 = ( n7592 & ~n2910 ) | ( n7592 & n7593 ) | ( ~n2910 & n7593 ) ;
  assign n7595 = ( n4478 & ~n7594 ) | ( n4478 & n6330 ) | ( ~n7594 & n6330 ) ;
  assign n7596 = ( n6330 & ~n7595 ) | ( n6330 & 1'b0 ) | ( ~n7595 & 1'b0 ) ;
  assign n7597 = ( x26 & ~n7594 ) | ( x26 & n7596 ) | ( ~n7594 & n7596 ) ;
  assign n7598 = ( n7594 & ~x26 ) | ( n7594 & n7596 ) | ( ~x26 & n7596 ) ;
  assign n7599 = ( n7597 & ~n7596 ) | ( n7597 & n7598 ) | ( ~n7596 & n7598 ) ;
  assign n7587 = ( n7354 & ~n7450 ) | ( n7354 & n7356 ) | ( ~n7450 & n7356 ) ;
  assign n7588 = ( n7356 & ~n7354 ) | ( n7356 & n7450 ) | ( ~n7354 & n7450 ) ;
  assign n7589 = ( n7587 & ~n7356 ) | ( n7587 & n7588 ) | ( ~n7356 & n7588 ) ;
  assign n7600 = ( n7370 & ~n7368 ) | ( n7370 & n7449 ) | ( ~n7368 & n7449 ) ;
  assign n7601 = ( n7368 & ~n7449 ) | ( n7368 & n7370 ) | ( ~n7449 & n7370 ) ;
  assign n7602 = ( n7600 & ~n7370 ) | ( n7600 & n7601 ) | ( ~n7370 & n7601 ) ;
  assign n7606 = ~n2839 & n4962 ;
  assign n7603 = n3030 | n4482 ;
  assign n7604 = n2995 | n4495 ;
  assign n7605 = n7603 &  n7604 ;
  assign n7607 = ( n2839 & n7606 ) | ( n2839 & n7605 ) | ( n7606 & n7605 ) ;
  assign n7608 = ( n7324 & ~n4478 ) | ( n7324 & n7607 ) | ( ~n4478 & n7607 ) ;
  assign n7609 = ~n7324 & n7608 ;
  assign n7610 = ( x26 & ~n7607 ) | ( x26 & n7609 ) | ( ~n7607 & n7609 ) ;
  assign n7611 = ( n7607 & ~x26 ) | ( n7607 & n7609 ) | ( ~x26 & n7609 ) ;
  assign n7612 = ( n7610 & ~n7609 ) | ( n7610 & n7611 ) | ( ~n7609 & n7611 ) ;
  assign n7613 = ( n7384 & ~n7382 ) | ( n7384 & n7448 ) | ( ~n7382 & n7448 ) ;
  assign n7614 = ( n7382 & ~n7448 ) | ( n7382 & n7384 ) | ( ~n7448 & n7384 ) ;
  assign n7615 = ( n7613 & ~n7384 ) | ( n7613 & n7614 ) | ( ~n7384 & n7614 ) ;
  assign n7616 = n3106 | n4482 ;
  assign n7617 = n3030 | n4495 ;
  assign n7618 = n7616 &  n7617 ;
  assign n7619 = ~n2995 & n4962 ;
  assign n7620 = ( n2995 & n7618 ) | ( n2995 & n7619 ) | ( n7618 & n7619 ) ;
  assign n7621 = ( n7339 & ~n4478 ) | ( n7339 & n7620 ) | ( ~n4478 & n7620 ) ;
  assign n7622 = ~n7339 & n7621 ;
  assign n7623 = ( x26 & ~n7620 ) | ( x26 & n7622 ) | ( ~n7620 & n7622 ) ;
  assign n7624 = ( n7620 & ~x26 ) | ( n7620 & n7622 ) | ( ~x26 & n7622 ) ;
  assign n7625 = ( n7623 & ~n7622 ) | ( n7623 & n7624 ) | ( ~n7622 & n7624 ) ;
  assign n7632 = ~n3030 & n4962 ;
  assign n7629 = n3197 | n4482 ;
  assign n7630 = n3106 | n4495 ;
  assign n7631 = n7629 &  n7630 ;
  assign n7633 = ( n3030 & n7632 ) | ( n3030 & n7631 ) | ( n7632 & n7631 ) ;
  assign n7634 = ( n6314 & ~n4478 ) | ( n6314 & n7633 ) | ( ~n4478 & n7633 ) ;
  assign n7635 = ~n6314 & n7634 ;
  assign n7636 = ( x26 & ~n7633 ) | ( x26 & n7635 ) | ( ~n7633 & n7635 ) ;
  assign n7637 = ( n7633 & ~x26 ) | ( n7633 & n7635 ) | ( ~x26 & n7635 ) ;
  assign n7638 = ( n7636 & ~n7635 ) | ( n7636 & n7637 ) | ( ~n7635 & n7637 ) ;
  assign n7626 = ( n7396 & ~n7447 ) | ( n7396 & n7398 ) | ( ~n7447 & n7398 ) ;
  assign n7627 = ( n7398 & ~n7396 ) | ( n7398 & n7447 ) | ( ~n7396 & n7447 ) ;
  assign n7628 = ( n7626 & ~n7398 ) | ( n7626 & n7627 ) | ( ~n7398 & n7627 ) ;
  assign n7642 = n3106 | n4962 ;
  assign n7643 = n3197 | n4495 ;
  assign n7644 = n7642 &  n7643 ;
  assign n7645 = n3266 &  n4482 ;
  assign n7646 = ( n7644 & ~n3266 ) | ( n7644 & n7645 ) | ( ~n3266 & n7645 ) ;
  assign n7647 = ( n7363 & ~n4478 ) | ( n7363 & n7646 ) | ( ~n4478 & n7646 ) ;
  assign n7648 = ~n7363 & n7647 ;
  assign n7649 = ( x26 & ~n7646 ) | ( x26 & n7648 ) | ( ~n7646 & n7648 ) ;
  assign n7650 = ( n7646 & ~x26 ) | ( n7646 & n7648 ) | ( ~x26 & n7648 ) ;
  assign n7651 = ( n7649 & ~n7648 ) | ( n7649 & n7650 ) | ( ~n7648 & n7650 ) ;
  assign n7640 = ( n7410 & n7417 ) | ( n7410 & n7446 ) | ( n7417 & n7446 ) ;
  assign n7639 = ( n7410 & ~n7417 ) | ( n7410 & n7446 ) | ( ~n7417 & n7446 ) ;
  assign n7641 = ( n7417 & ~n7640 ) | ( n7417 & n7639 ) | ( ~n7640 & n7639 ) ;
  assign n7652 = n3197 | n4962 ;
  assign n7653 = n3325 | n4482 ;
  assign n7654 = n7652 &  n7653 ;
  assign n7655 = n3266 &  n4495 ;
  assign n7656 = ( n7654 & ~n3266 ) | ( n7654 & n7655 ) | ( ~n3266 & n7655 ) ;
  assign n7657 = ( n4478 & ~n7656 ) | ( n4478 & n7377 ) | ( ~n7656 & n7377 ) ;
  assign n7658 = ( n7377 & ~n7657 ) | ( n7377 & 1'b0 ) | ( ~n7657 & 1'b0 ) ;
  assign n7659 = ( x26 & ~n7656 ) | ( x26 & n7658 ) | ( ~n7656 & n7658 ) ;
  assign n7660 = ( n7656 & ~x26 ) | ( n7656 & n7658 ) | ( ~x26 & n7658 ) ;
  assign n7661 = ( n7659 & ~n7658 ) | ( n7659 & n7660 ) | ( ~n7658 & n7660 ) ;
  assign n7663 = ( n7418 & n7435 ) | ( n7418 & n7445 ) | ( n7435 & n7445 ) ;
  assign n7662 = ( n7418 & ~n7435 ) | ( n7418 & n7445 ) | ( ~n7435 & n7445 ) ;
  assign n7664 = ( n7435 & ~n7663 ) | ( n7435 & n7662 ) | ( ~n7663 & n7662 ) ;
  assign n7665 = n3361 | n4482 ;
  assign n7666 = n3325 | n4495 ;
  assign n7667 = n7665 &  n7666 ;
  assign n7668 = n3266 &  n4962 ;
  assign n7669 = ( n7667 & ~n3266 ) | ( n7667 & n7668 ) | ( ~n3266 & n7668 ) ;
  assign n7670 = ( n4478 & ~n7669 ) | ( n4478 & n7391 ) | ( ~n7669 & n7391 ) ;
  assign n7671 = ( n7391 & ~n7670 ) | ( n7391 & 1'b0 ) | ( ~n7670 & 1'b0 ) ;
  assign n7672 = ( x26 & ~n7669 ) | ( x26 & n7671 ) | ( ~n7669 & n7671 ) ;
  assign n7673 = ( n7669 & ~x26 ) | ( n7669 & n7671 ) | ( ~x26 & n7671 ) ;
  assign n7674 = ( n7672 & ~n7671 ) | ( n7672 & n7673 ) | ( ~n7671 & n7673 ) ;
  assign n7426 = ( x29 & ~n7425 ) | ( x29 & 1'b0 ) | ( ~n7425 & 1'b0 ) ;
  assign n7676 = ( x29 & n7426 ) | ( x29 & n7433 ) | ( n7426 & n7433 ) ;
  assign n7675 = ( x29 & ~n7426 ) | ( x29 & n7433 ) | ( ~n7426 & n7433 ) ;
  assign n7677 = ( n7426 & ~n7676 ) | ( n7426 & n7675 ) | ( ~n7676 & n7675 ) ;
  assign n7678 = x29 &  n7424 ;
  assign n7679 = n7423 &  n7678 ;
  assign n7680 = n7423 | n7678 ;
  assign n7681 = ~n7679 & n7680 ;
  assign n7712 = ~n3460 & n4495 ;
  assign n7709 = n3361 | n4962 ;
  assign n7710 = n3601 | n4482 ;
  assign n7711 = n7709 &  n7710 ;
  assign n7713 = ( n3460 & n7712 ) | ( n3460 & n7711 ) | ( n7712 & n7711 ) ;
  assign n7714 = ( n6895 & ~n4478 ) | ( n6895 & n7713 ) | ( ~n4478 & n7713 ) ;
  assign n7715 = ~n6895 & n7714 ;
  assign n7716 = ( x26 & ~n7713 ) | ( x26 & n7715 ) | ( ~n7713 & n7715 ) ;
  assign n7717 = ( n7713 & ~x26 ) | ( n7713 & n7715 ) | ( ~x26 & n7715 ) ;
  assign n7718 = ( n7716 & ~n7715 ) | ( n7716 & n7717 ) | ( ~n7715 & n7717 ) ;
  assign n7705 = ~n4478 & n6886 ;
  assign n7703 = ~n3460 & n4962 ;
  assign n7700 = n3547 | n4482 ;
  assign n7701 = n3601 | n4495 ;
  assign n7702 = n7700 &  n7701 ;
  assign n7704 = ( n3460 & n7703 ) | ( n3460 & n7702 ) | ( n7703 & n7702 ) ;
  assign n7706 = ( n4478 & n7705 ) | ( n4478 & n7704 ) | ( n7705 & n7704 ) ;
  assign n7695 = n7412 | n4478 ;
  assign n7692 = n3547 | n4495 ;
  assign n7693 = n3601 | n4962 ;
  assign n7694 = n7692 &  n7693 ;
  assign n7696 = ( n4478 & ~n7695 ) | ( n4478 & n7694 ) | ( ~n7695 & n7694 ) ;
  assign n7697 = ~n3547 & n4474 ;
  assign n7698 = ( x26 & ~n7696 ) | ( x26 & n7697 ) | ( ~n7696 & n7697 ) ;
  assign n7707 = ( x26 & ~n7706 ) | ( x26 & n7698 ) | ( ~n7706 & n7698 ) ;
  assign n7708 = ( x26 & ~n7707 ) | ( x26 & 1'b0 ) | ( ~n7707 & 1'b0 ) ;
  assign n7719 = ( n7424 & ~n7718 ) | ( n7424 & n7708 ) | ( ~n7718 & n7708 ) ;
  assign n7685 = ~n3460 & n4482 ;
  assign n7682 = n3325 | n4962 ;
  assign n7683 = n3361 | n4495 ;
  assign n7684 = n7682 &  n7683 ;
  assign n7686 = ( n3460 & n7685 ) | ( n3460 & n7684 ) | ( n7685 & n7684 ) ;
  assign n7687 = ( n7405 & ~n4478 ) | ( n7405 & n7686 ) | ( ~n4478 & n7686 ) ;
  assign n7688 = ~n7405 & n7687 ;
  assign n7689 = ( x26 & ~n7686 ) | ( x26 & n7688 ) | ( ~n7686 & n7688 ) ;
  assign n7690 = ( n7686 & ~x26 ) | ( n7686 & n7688 ) | ( ~x26 & n7688 ) ;
  assign n7691 = ( n7689 & ~n7688 ) | ( n7689 & n7690 ) | ( ~n7688 & n7690 ) ;
  assign n7720 = ( n7681 & ~n7719 ) | ( n7681 & n7691 ) | ( ~n7719 & n7691 ) ;
  assign n7721 = ( n7674 & n7677 ) | ( n7674 & n7720 ) | ( n7677 & n7720 ) ;
  assign n7722 = ( n7661 & n7664 ) | ( n7661 & n7721 ) | ( n7664 & n7721 ) ;
  assign n7723 = ( n7651 & ~n7641 ) | ( n7651 & n7722 ) | ( ~n7641 & n7722 ) ;
  assign n7724 = ( n7638 & ~n7628 ) | ( n7638 & n7723 ) | ( ~n7628 & n7723 ) ;
  assign n7725 = ( n7615 & n7625 ) | ( n7615 & n7724 ) | ( n7625 & n7724 ) ;
  assign n7726 = ( n7602 & n7612 ) | ( n7602 & n7725 ) | ( n7612 & n7725 ) ;
  assign n7727 = ( n7599 & ~n7589 ) | ( n7599 & n7726 ) | ( ~n7589 & n7726 ) ;
  assign n7728 = ( n7576 & n7586 ) | ( n7576 & n7727 ) | ( n7586 & n7727 ) ;
  assign n7729 = ( n7563 & n7573 ) | ( n7563 & n7728 ) | ( n7573 & n7728 ) ;
  assign n7730 = ( n6917 & n7453 ) | ( n6917 & n7456 ) | ( n7453 & n7456 ) ;
  assign n7731 = ( n7453 & ~n6917 ) | ( n7453 & n7456 ) | ( ~n6917 & n7456 ) ;
  assign n7732 = ( n6917 & ~n7730 ) | ( n6917 & n7731 ) | ( ~n7730 & n7731 ) ;
  assign n7733 = ( x26 & ~n7466 ) | ( x26 & n7732 ) | ( ~n7466 & n7732 ) ;
  assign n7734 = ( n7466 & ~x26 ) | ( n7466 & n7732 ) | ( ~x26 & n7732 ) ;
  assign n7735 = ( n7733 & ~n7732 ) | ( n7733 & n7734 ) | ( ~n7732 & n7734 ) ;
  assign n7739 = ~n2392 & n5135 ;
  assign n7736 = n2569 | n5010 ;
  assign n7737 = n2483 | n5067 ;
  assign n7738 = n7736 &  n7737 ;
  assign n7740 = ( n2392 & n7739 ) | ( n2392 & n7738 ) | ( n7739 & n7738 ) ;
  assign n7741 = n5012 | n6212 ;
  assign n7742 = n7740 &  n7741 ;
  assign n7743 = x23 &  n7742 ;
  assign n7744 = x23 | n7742 ;
  assign n7745 = ~n7743 & n7744 ;
  assign n7746 = ( n7729 & ~n7735 ) | ( n7729 & n7745 ) | ( ~n7735 & n7745 ) ;
  assign n7558 = ( n7314 & n7470 ) | ( n7314 & n7480 ) | ( n7470 & n7480 ) ;
  assign n7559 = ( n7314 & ~n7470 ) | ( n7314 & n7480 ) | ( ~n7470 & n7480 ) ;
  assign n7560 = ( n7470 & ~n7558 ) | ( n7470 & n7559 ) | ( ~n7558 & n7559 ) ;
  assign n7747 = ~n2178 & n5339 ;
  assign n7748 = n2127 | n5761 ;
  assign n7749 = ~n7747 & n7748 ;
  assign n7750 = ~n2022 & n5837 ;
  assign n7751 = ( n2022 & n7749 ) | ( n2022 & n7750 ) | ( n7749 & n7750 ) ;
  assign n7752 = ( n5341 & ~n4934 ) | ( n5341 & n7751 ) | ( ~n4934 & n7751 ) ;
  assign n7753 = ~n5341 & n7752 ;
  assign n7754 = ( x20 & ~n7751 ) | ( x20 & n7753 ) | ( ~n7751 & n7753 ) ;
  assign n7755 = ( n7751 & ~x20 ) | ( n7751 & n7753 ) | ( ~x20 & n7753 ) ;
  assign n7756 = ( n7754 & ~n7753 ) | ( n7754 & n7755 ) | ( ~n7753 & n7755 ) ;
  assign n7757 = ( n7746 & ~n7560 ) | ( n7746 & n7756 ) | ( ~n7560 & n7756 ) ;
  assign n7552 = ( n7205 & n7308 ) | ( n7205 & n7481 ) | ( n7308 & n7481 ) ;
  assign n7553 = ( n7308 & ~n7205 ) | ( n7308 & n7481 ) | ( ~n7205 & n7481 ) ;
  assign n7554 = ( n7205 & ~n7552 ) | ( n7205 & n7553 ) | ( ~n7552 & n7553 ) ;
  assign n7556 = ( x20 & n7488 ) | ( x20 & n7554 ) | ( n7488 & n7554 ) ;
  assign n7555 = ( n7488 & ~x20 ) | ( n7488 & n7554 ) | ( ~x20 & n7554 ) ;
  assign n7557 = ( x20 & ~n7556 ) | ( x20 & n7555 ) | ( ~n7556 & n7555 ) ;
  assign n7761 = ~n1875 & n5970 ;
  assign n7758 = n1671 | n6395 ;
  assign n7759 = n1748 | n6170 ;
  assign n7760 = n7758 &  n7759 ;
  assign n7762 = ( n1875 & n7761 ) | ( n1875 & n7760 ) | ( n7761 & n7760 ) ;
  assign n7763 = n4580 | n5972 ;
  assign n7764 = n7762 &  n7763 ;
  assign n7765 = x17 &  n7764 ;
  assign n7766 = x17 | n7764 ;
  assign n7767 = ~n7765 & n7766 ;
  assign n7768 = ( n7757 & ~n7557 ) | ( n7757 & n7767 ) | ( ~n7557 & n7767 ) ;
  assign n7769 = ( n7549 & ~n7551 ) | ( n7549 & n7768 ) | ( ~n7551 & n7768 ) ;
  assign n7534 = ( n7217 & n7289 ) | ( n7217 & n7493 ) | ( n7289 & n7493 ) ;
  assign n7535 = ( n7289 & ~n7217 ) | ( n7289 & n7493 ) | ( ~n7217 & n7493 ) ;
  assign n7536 = ( n7217 & ~n7534 ) | ( n7217 & n7535 ) | ( ~n7534 & n7535 ) ;
  assign n7538 = ( x17 & n7500 ) | ( x17 & n7536 ) | ( n7500 & n7536 ) ;
  assign n7537 = ( n7500 & ~x17 ) | ( n7500 & n7536 ) | ( ~x17 & n7536 ) ;
  assign n7539 = ( x17 & ~n7538 ) | ( x17 & n7537 ) | ( ~n7538 & n7537 ) ;
  assign n7770 = n1151 | n7097 ;
  assign n7771 = n1378 | n6530 ;
  assign n7772 = n7770 &  n7771 ;
  assign n7773 = n1267 &  n6983 ;
  assign n7774 = ( n7772 & ~n1267 ) | ( n7772 & n7773 ) | ( ~n1267 & n7773 ) ;
  assign n7775 = ( n4061 & ~n6532 ) | ( n4061 & 1'b0 ) | ( ~n6532 & 1'b0 ) ;
  assign n7776 = ( n7774 & ~n7775 ) | ( n7774 & 1'b0 ) | ( ~n7775 & 1'b0 ) ;
  assign n7777 = x14 &  n7776 ;
  assign n7778 = x14 | n7776 ;
  assign n7779 = ~n7777 & n7778 ;
  assign n7780 = ( n7769 & ~n7539 ) | ( n7769 & n7779 ) | ( ~n7539 & n7779 ) ;
  assign n7781 = ( n7533 & ~n7780 ) | ( n7533 & 1'b0 ) | ( ~n7780 & 1'b0 ) ;
  assign n7791 = ~n7533 & n7780 ;
  assign n7792 = ( n7789 & ~x11 ) | ( n7789 & n7791 ) | ( ~x11 & n7791 ) ;
  assign n7793 = ( n7790 & ~n7781 ) | ( n7790 & n7792 ) | ( ~n7781 & n7792 ) ;
  assign n7794 = n863 &  n7253 ;
  assign n7795 = n599 | n7783 ;
  assign n7796 = n702 | n7518 ;
  assign n7797 = n7795 &  n7796 ;
  assign n7798 = ( n7794 & ~n7253 ) | ( n7794 & n7797 ) | ( ~n7253 & n7797 ) ;
  assign n7799 = ( n7255 & ~n4452 ) | ( n7255 & n7798 ) | ( ~n4452 & n7798 ) ;
  assign n7800 = ~n7255 & n7799 ;
  assign n7801 = ( x11 & ~n7798 ) | ( x11 & n7800 ) | ( ~n7798 & n7800 ) ;
  assign n7802 = ( n7798 & ~x11 ) | ( n7798 & n7800 ) | ( ~x11 & n7800 ) ;
  assign n7803 = ( n7801 & ~n7800 ) | ( n7801 & n7802 ) | ( ~n7800 & n7802 ) ;
  assign n7804 = ( n7273 & ~n7283 ) | ( n7273 & n7515 ) | ( ~n7283 & n7515 ) ;
  assign n7805 = ( n7283 & ~n7516 ) | ( n7283 & n7804 ) | ( ~n7516 & n7804 ) ;
  assign n7806 = ( n7793 & n7803 ) | ( n7793 & n7805 ) | ( n7803 & n7805 ) ;
  assign n7808 = ( n7516 & n7525 ) | ( n7516 & n7529 ) | ( n7525 & n7529 ) ;
  assign n7807 = ( n7516 & ~n7525 ) | ( n7516 & n7529 ) | ( ~n7525 & n7529 ) ;
  assign n7809 = ( n7525 & ~n7808 ) | ( n7525 & n7807 ) | ( ~n7808 & n7807 ) ;
  assign n7810 = ( n7803 & ~n7793 ) | ( n7803 & n7805 ) | ( ~n7793 & n7805 ) ;
  assign n7811 = ( n7793 & ~n7805 ) | ( n7793 & n7803 ) | ( ~n7805 & n7803 ) ;
  assign n7812 = ( n7810 & ~n7803 ) | ( n7810 & n7811 ) | ( ~n7803 & n7811 ) ;
  assign n7819 = ( n1483 & ~n6530 ) | ( n1483 & 1'b0 ) | ( ~n6530 & 1'b0 ) ;
  assign n7820 = n1378 | n6983 ;
  assign n7821 = ~n7819 & n7820 ;
  assign n7822 = n1267 &  n7097 ;
  assign n7823 = ( n7821 & ~n1267 ) | ( n7821 & n7822 ) | ( ~n1267 & n7822 ) ;
  assign n7824 = ( n4422 & n6532 ) | ( n4422 & n7823 ) | ( n6532 & n7823 ) ;
  assign n7825 = ~n6532 & n7824 ;
  assign n7826 = ( x14 & ~n7823 ) | ( x14 & n7825 ) | ( ~n7823 & n7825 ) ;
  assign n7827 = ( n7823 & ~x14 ) | ( n7823 & n7825 ) | ( ~x14 & n7825 ) ;
  assign n7828 = ( n7826 & ~n7825 ) | ( n7826 & n7827 ) | ( ~n7825 & n7827 ) ;
  assign n7816 = ( n7551 & ~n7549 ) | ( n7551 & n7768 ) | ( ~n7549 & n7768 ) ;
  assign n7817 = ( n7549 & ~n7768 ) | ( n7549 & n7551 ) | ( ~n7768 & n7551 ) ;
  assign n7818 = ( n7816 & ~n7551 ) | ( n7816 & n7817 ) | ( ~n7551 & n7817 ) ;
  assign n7838 = ( n7469 & ~n7729 ) | ( n7469 & n7732 ) | ( ~n7729 & n7732 ) ;
  assign n7839 = ( n7729 & ~n7469 ) | ( n7729 & n7732 ) | ( ~n7469 & n7732 ) ;
  assign n7840 = ( n7838 & ~n7732 ) | ( n7838 & n7839 ) | ( ~n7732 & n7839 ) ;
  assign n8046 = n7745 &  n7840 ;
  assign n7844 = ~n2665 & n5010 ;
  assign n7841 = n2483 | n5135 ;
  assign n7842 = n2569 | n5067 ;
  assign n7843 = n7841 &  n7842 ;
  assign n7845 = ( n2665 & n7844 ) | ( n2665 & n7843 ) | ( n7844 & n7843 ) ;
  assign n7846 = ( n6465 & ~n5012 ) | ( n6465 & n7845 ) | ( ~n5012 & n7845 ) ;
  assign n7847 = ~n6465 & n7846 ;
  assign n7848 = ( x23 & ~n7845 ) | ( x23 & n7847 ) | ( ~n7845 & n7847 ) ;
  assign n7849 = ( n7845 & ~x23 ) | ( n7845 & n7847 ) | ( ~x23 & n7847 ) ;
  assign n7850 = ( n7848 & ~n7847 ) | ( n7848 & n7849 ) | ( ~n7847 & n7849 ) ;
  assign n7851 = ( n7563 & ~n7573 ) | ( n7563 & n7728 ) | ( ~n7573 & n7728 ) ;
  assign n7852 = ( n7573 & ~n7729 ) | ( n7573 & n7851 ) | ( ~n7729 & n7851 ) ;
  assign n7856 = ~n2751 & n5010 ;
  assign n7853 = n2569 | n5135 ;
  assign n7854 = n2665 | n5067 ;
  assign n7855 = n7853 &  n7854 ;
  assign n7857 = ( n2751 & n7856 ) | ( n2751 & n7855 ) | ( n7856 & n7855 ) ;
  assign n7858 = ( n5705 & ~n5012 ) | ( n5705 & n7857 ) | ( ~n5012 & n7857 ) ;
  assign n7859 = ~n5705 & n7858 ;
  assign n7860 = ( x23 & ~n7857 ) | ( x23 & n7859 ) | ( ~n7857 & n7859 ) ;
  assign n7861 = ( n7857 & ~x23 ) | ( n7857 & n7859 ) | ( ~x23 & n7859 ) ;
  assign n7862 = ( n7860 & ~n7859 ) | ( n7860 & n7861 ) | ( ~n7859 & n7861 ) ;
  assign n7863 = ( n7576 & ~n7586 ) | ( n7576 & n7727 ) | ( ~n7586 & n7727 ) ;
  assign n7864 = ( n7586 & ~n7728 ) | ( n7586 & n7863 ) | ( ~n7728 & n7863 ) ;
  assign n7868 = ~n2751 & n5067 ;
  assign n7865 = n2665 | n5135 ;
  assign n7866 = n2783 | n5010 ;
  assign n7867 = n7865 &  n7866 ;
  assign n7869 = ( n2751 & n7868 ) | ( n2751 & n7867 ) | ( n7868 & n7867 ) ;
  assign n7870 = ( n6119 & ~n5012 ) | ( n6119 & n7869 ) | ( ~n5012 & n7869 ) ;
  assign n7871 = ~n6119 & n7870 ;
  assign n7872 = ( x23 & ~n7869 ) | ( x23 & n7871 ) | ( ~n7869 & n7871 ) ;
  assign n7873 = ( n7869 & ~x23 ) | ( n7869 & n7871 ) | ( ~x23 & n7871 ) ;
  assign n7874 = ( n7872 & ~n7871 ) | ( n7872 & n7873 ) | ( ~n7871 & n7873 ) ;
  assign n7875 = ( n7589 & ~n7726 ) | ( n7589 & n7599 ) | ( ~n7726 & n7599 ) ;
  assign n7876 = ( n7727 & ~n7599 ) | ( n7727 & n7875 ) | ( ~n7599 & n7875 ) ;
  assign n7877 = n2751 | n5135 ;
  assign n7878 = n2783 | n5067 ;
  assign n7879 = n7877 &  n7878 ;
  assign n7880 = n2910 &  n5010 ;
  assign n7881 = ( n7879 & ~n2910 ) | ( n7879 & n7880 ) | ( ~n2910 & n7880 ) ;
  assign n7882 = ( n6226 & ~n5012 ) | ( n6226 & n7881 ) | ( ~n5012 & n7881 ) ;
  assign n7883 = ~n6226 & n7882 ;
  assign n7884 = ( x23 & ~n7881 ) | ( x23 & n7883 ) | ( ~n7881 & n7883 ) ;
  assign n7885 = ( n7881 & ~x23 ) | ( n7881 & n7883 ) | ( ~x23 & n7883 ) ;
  assign n7886 = ( n7884 & ~n7883 ) | ( n7884 & n7885 ) | ( ~n7883 & n7885 ) ;
  assign n7887 = ( n7602 & ~n7612 ) | ( n7602 & n7725 ) | ( ~n7612 & n7725 ) ;
  assign n7888 = ( n7612 & ~n7726 ) | ( n7612 & n7887 ) | ( ~n7726 & n7887 ) ;
  assign n7889 = n2783 | n5135 ;
  assign n7890 = n2839 | n5010 ;
  assign n7891 = n7889 &  n7890 ;
  assign n7892 = n2910 &  n5067 ;
  assign n7893 = ( n7891 & ~n2910 ) | ( n7891 & n7892 ) | ( ~n2910 & n7892 ) ;
  assign n7894 = ~n5012 & n6104 ;
  assign n7895 = ( n7893 & ~n7894 ) | ( n7893 & 1'b0 ) | ( ~n7894 & 1'b0 ) ;
  assign n7896 = x23 &  n7895 ;
  assign n7897 = x23 | n7895 ;
  assign n7898 = ~n7896 & n7897 ;
  assign n7899 = ( n7615 & ~n7625 ) | ( n7615 & n7724 ) | ( ~n7625 & n7724 ) ;
  assign n7900 = ( n7625 & ~n7725 ) | ( n7625 & n7899 ) | ( ~n7725 & n7899 ) ;
  assign n7901 = n2995 | n5010 ;
  assign n7902 = n2839 | n5067 ;
  assign n7903 = n7901 &  n7902 ;
  assign n7904 = n2910 &  n5135 ;
  assign n7905 = ( n7903 & ~n2910 ) | ( n7903 & n7904 ) | ( ~n2910 & n7904 ) ;
  assign n7906 = ( n5012 & ~n7905 ) | ( n5012 & n6330 ) | ( ~n7905 & n6330 ) ;
  assign n7907 = ( n6330 & ~n7906 ) | ( n6330 & 1'b0 ) | ( ~n7906 & 1'b0 ) ;
  assign n7908 = ( x23 & ~n7905 ) | ( x23 & n7907 ) | ( ~n7905 & n7907 ) ;
  assign n7909 = ( n7905 & ~x23 ) | ( n7905 & n7907 ) | ( ~x23 & n7907 ) ;
  assign n7910 = ( n7908 & ~n7907 ) | ( n7908 & n7909 ) | ( ~n7907 & n7909 ) ;
  assign n7911 = ( n7628 & ~n7723 ) | ( n7628 & n7638 ) | ( ~n7723 & n7638 ) ;
  assign n7912 = ( n7724 & ~n7638 ) | ( n7724 & n7911 ) | ( ~n7638 & n7911 ) ;
  assign n7916 = ~n2839 & n5135 ;
  assign n7913 = n3030 | n5010 ;
  assign n7914 = n2995 | n5067 ;
  assign n7915 = n7913 &  n7914 ;
  assign n7917 = ( n2839 & n7916 ) | ( n2839 & n7915 ) | ( n7916 & n7915 ) ;
  assign n7918 = ( n7324 & ~n5012 ) | ( n7324 & n7917 ) | ( ~n5012 & n7917 ) ;
  assign n7919 = ~n7324 & n7918 ;
  assign n7920 = ( x23 & ~n7917 ) | ( x23 & n7919 ) | ( ~n7917 & n7919 ) ;
  assign n7921 = ( n7917 & ~x23 ) | ( n7917 & n7919 ) | ( ~x23 & n7919 ) ;
  assign n7922 = ( n7920 & ~n7919 ) | ( n7920 & n7921 ) | ( ~n7919 & n7921 ) ;
  assign n7923 = ( n7641 & n7651 ) | ( n7641 & n7722 ) | ( n7651 & n7722 ) ;
  assign n7924 = ( n7641 & ~n7651 ) | ( n7641 & n7722 ) | ( ~n7651 & n7722 ) ;
  assign n7925 = ( n7651 & ~n7923 ) | ( n7651 & n7924 ) | ( ~n7923 & n7924 ) ;
  assign n7926 = ( n7661 & ~n7721 ) | ( n7661 & n7664 ) | ( ~n7721 & n7664 ) ;
  assign n7927 = ( n7664 & ~n7661 ) | ( n7664 & n7721 ) | ( ~n7661 & n7721 ) ;
  assign n7928 = ( n7926 & ~n7664 ) | ( n7926 & n7927 ) | ( ~n7664 & n7927 ) ;
  assign n7929 = n3106 | n5010 ;
  assign n7930 = n3030 | n5067 ;
  assign n7931 = n7929 &  n7930 ;
  assign n7932 = ~n2995 & n5135 ;
  assign n7933 = ( n2995 & n7931 ) | ( n2995 & n7932 ) | ( n7931 & n7932 ) ;
  assign n7934 = ( n7339 & ~n5012 ) | ( n7339 & n7933 ) | ( ~n5012 & n7933 ) ;
  assign n7935 = ~n7339 & n7934 ;
  assign n7936 = ( x23 & ~n7933 ) | ( x23 & n7935 ) | ( ~n7933 & n7935 ) ;
  assign n7937 = ( n7933 & ~x23 ) | ( n7933 & n7935 ) | ( ~x23 & n7935 ) ;
  assign n7938 = ( n7936 & ~n7935 ) | ( n7936 & n7937 ) | ( ~n7935 & n7937 ) ;
  assign n7939 = ( n7674 & ~n7720 ) | ( n7674 & n7677 ) | ( ~n7720 & n7677 ) ;
  assign n7940 = ( n7677 & ~n7674 ) | ( n7677 & n7720 ) | ( ~n7674 & n7720 ) ;
  assign n7941 = ( n7939 & ~n7677 ) | ( n7939 & n7940 ) | ( ~n7677 & n7940 ) ;
  assign n7945 = ~n3030 & n5135 ;
  assign n7942 = n3197 | n5010 ;
  assign n7943 = n3106 | n5067 ;
  assign n7944 = n7942 &  n7943 ;
  assign n7946 = ( n3030 & n7945 ) | ( n3030 & n7944 ) | ( n7945 & n7944 ) ;
  assign n7947 = ( n6314 & ~n5012 ) | ( n6314 & n7946 ) | ( ~n5012 & n7946 ) ;
  assign n7948 = ~n6314 & n7947 ;
  assign n7949 = ( x23 & ~n7946 ) | ( x23 & n7948 ) | ( ~n7946 & n7948 ) ;
  assign n7950 = ( n7946 & ~x23 ) | ( n7946 & n7948 ) | ( ~x23 & n7948 ) ;
  assign n7951 = ( n7949 & ~n7948 ) | ( n7949 & n7950 ) | ( ~n7948 & n7950 ) ;
  assign n7952 = n3106 | n5135 ;
  assign n7953 = n3197 | n5067 ;
  assign n7954 = n7952 &  n7953 ;
  assign n7955 = n3266 &  n5010 ;
  assign n7956 = ( n7954 & ~n3266 ) | ( n7954 & n7955 ) | ( ~n3266 & n7955 ) ;
  assign n7957 = ( n7363 & ~n5012 ) | ( n7363 & n7956 ) | ( ~n5012 & n7956 ) ;
  assign n7958 = ~n7363 & n7957 ;
  assign n7959 = ( x23 & ~n7956 ) | ( x23 & n7958 ) | ( ~n7956 & n7958 ) ;
  assign n7960 = ( n7956 & ~x23 ) | ( n7956 & n7958 ) | ( ~x23 & n7958 ) ;
  assign n7961 = ( n7959 & ~n7958 ) | ( n7959 & n7960 ) | ( ~n7958 & n7960 ) ;
  assign n7962 = ( n7691 & ~n7681 ) | ( n7691 & n7719 ) | ( ~n7681 & n7719 ) ;
  assign n7963 = ( n7720 & ~n7691 ) | ( n7720 & n7962 ) | ( ~n7691 & n7962 ) ;
  assign n7965 = ( n7424 & n7708 ) | ( n7424 & n7718 ) | ( n7708 & n7718 ) ;
  assign n7964 = ( n7424 & ~n7708 ) | ( n7424 & n7718 ) | ( ~n7708 & n7718 ) ;
  assign n7966 = ( n7708 & ~n7965 ) | ( n7708 & n7964 ) | ( ~n7965 & n7964 ) ;
  assign n7967 = n3197 | n5135 ;
  assign n7968 = n3325 | n5010 ;
  assign n7969 = n7967 &  n7968 ;
  assign n7970 = n3266 &  n5067 ;
  assign n7971 = ( n7969 & ~n3266 ) | ( n7969 & n7970 ) | ( ~n3266 & n7970 ) ;
  assign n7972 = ( n5012 & ~n7971 ) | ( n5012 & n7377 ) | ( ~n7971 & n7377 ) ;
  assign n7973 = ( n7377 & ~n7972 ) | ( n7377 & 1'b0 ) | ( ~n7972 & 1'b0 ) ;
  assign n7974 = ( x23 & ~n7971 ) | ( x23 & n7973 ) | ( ~n7971 & n7973 ) ;
  assign n7975 = ( n7971 & ~x23 ) | ( n7971 & n7973 ) | ( ~x23 & n7973 ) ;
  assign n7976 = ( n7974 & ~n7973 ) | ( n7974 & n7975 ) | ( ~n7973 & n7975 ) ;
  assign n7977 = n3361 | n5010 ;
  assign n7978 = n3325 | n5067 ;
  assign n7979 = n7977 &  n7978 ;
  assign n7980 = n3266 &  n5135 ;
  assign n7981 = ( n7979 & ~n3266 ) | ( n7979 & n7980 ) | ( ~n3266 & n7980 ) ;
  assign n7982 = ( n5012 & ~n7981 ) | ( n5012 & n7391 ) | ( ~n7981 & n7391 ) ;
  assign n7983 = ( n7391 & ~n7982 ) | ( n7391 & 1'b0 ) | ( ~n7982 & 1'b0 ) ;
  assign n7984 = ( x23 & ~n7981 ) | ( x23 & n7983 ) | ( ~n7981 & n7983 ) ;
  assign n7985 = ( n7981 & ~x23 ) | ( n7981 & n7983 ) | ( ~x23 & n7983 ) ;
  assign n7986 = ( n7984 & ~n7983 ) | ( n7984 & n7985 ) | ( ~n7983 & n7985 ) ;
  assign n7699 = ( x26 & ~n7698 ) | ( x26 & 1'b0 ) | ( ~n7698 & 1'b0 ) ;
  assign n7988 = ( x26 & n7699 ) | ( x26 & n7706 ) | ( n7699 & n7706 ) ;
  assign n7987 = ( x26 & ~n7699 ) | ( x26 & n7706 ) | ( ~n7699 & n7706 ) ;
  assign n7989 = ( n7699 & ~n7988 ) | ( n7699 & n7987 ) | ( ~n7988 & n7987 ) ;
  assign n7990 = x26 &  n7697 ;
  assign n7991 = n7696 &  n7990 ;
  assign n7992 = n7696 | n7990 ;
  assign n7993 = ~n7991 & n7992 ;
  assign n8024 = ~n3460 & n5067 ;
  assign n8021 = n3361 | n5135 ;
  assign n8022 = n3601 | n5010 ;
  assign n8023 = n8021 &  n8022 ;
  assign n8025 = ( n3460 & n8024 ) | ( n3460 & n8023 ) | ( n8024 & n8023 ) ;
  assign n8026 = ( n6895 & ~n5012 ) | ( n6895 & n8025 ) | ( ~n5012 & n8025 ) ;
  assign n8027 = ~n6895 & n8026 ;
  assign n8028 = ( x23 & ~n8025 ) | ( x23 & n8027 ) | ( ~n8025 & n8027 ) ;
  assign n8029 = ( n8025 & ~x23 ) | ( n8025 & n8027 ) | ( ~x23 & n8027 ) ;
  assign n8030 = ( n8028 & ~n8027 ) | ( n8028 & n8029 ) | ( ~n8027 & n8029 ) ;
  assign n8017 = ~n5012 & n6886 ;
  assign n8015 = ~n3460 & n5135 ;
  assign n8012 = n3547 | n5010 ;
  assign n8013 = n3601 | n5067 ;
  assign n8014 = n8012 &  n8013 ;
  assign n8016 = ( n3460 & n8015 ) | ( n3460 & n8014 ) | ( n8015 & n8014 ) ;
  assign n8018 = ( n5012 & n8017 ) | ( n5012 & n8016 ) | ( n8017 & n8016 ) ;
  assign n8007 = n7412 | n5012 ;
  assign n8004 = n3547 | n5067 ;
  assign n8005 = n3601 | n5135 ;
  assign n8006 = n8004 &  n8005 ;
  assign n8008 = ( n5012 & ~n8007 ) | ( n5012 & n8006 ) | ( ~n8007 & n8006 ) ;
  assign n8009 = ~n3547 & n5005 ;
  assign n8010 = ( x23 & ~n8008 ) | ( x23 & n8009 ) | ( ~n8008 & n8009 ) ;
  assign n8019 = ( x23 & ~n8018 ) | ( x23 & n8010 ) | ( ~n8018 & n8010 ) ;
  assign n8020 = ( x23 & ~n8019 ) | ( x23 & 1'b0 ) | ( ~n8019 & 1'b0 ) ;
  assign n8031 = ( n7697 & ~n8030 ) | ( n7697 & n8020 ) | ( ~n8030 & n8020 ) ;
  assign n7997 = ~n3460 & n5010 ;
  assign n7994 = n3325 | n5135 ;
  assign n7995 = n3361 | n5067 ;
  assign n7996 = n7994 &  n7995 ;
  assign n7998 = ( n3460 & n7997 ) | ( n3460 & n7996 ) | ( n7997 & n7996 ) ;
  assign n7999 = ( n7405 & ~n5012 ) | ( n7405 & n7998 ) | ( ~n5012 & n7998 ) ;
  assign n8000 = ~n7405 & n7999 ;
  assign n8001 = ( x23 & ~n7998 ) | ( x23 & n8000 ) | ( ~n7998 & n8000 ) ;
  assign n8002 = ( n7998 & ~x23 ) | ( n7998 & n8000 ) | ( ~x23 & n8000 ) ;
  assign n8003 = ( n8001 & ~n8000 ) | ( n8001 & n8002 ) | ( ~n8000 & n8002 ) ;
  assign n8032 = ( n7993 & ~n8031 ) | ( n7993 & n8003 ) | ( ~n8031 & n8003 ) ;
  assign n8033 = ( n7986 & n7989 ) | ( n7986 & n8032 ) | ( n7989 & n8032 ) ;
  assign n8034 = ( n7966 & n7976 ) | ( n7966 & n8033 ) | ( n7976 & n8033 ) ;
  assign n8035 = ( n7961 & ~n7963 ) | ( n7961 & n8034 ) | ( ~n7963 & n8034 ) ;
  assign n8036 = ( n7941 & n7951 ) | ( n7941 & n8035 ) | ( n7951 & n8035 ) ;
  assign n8037 = ( n7928 & n7938 ) | ( n7928 & n8036 ) | ( n7938 & n8036 ) ;
  assign n8038 = ( n7922 & ~n7925 ) | ( n7922 & n8037 ) | ( ~n7925 & n8037 ) ;
  assign n8039 = ( n7910 & ~n7912 ) | ( n7910 & n8038 ) | ( ~n7912 & n8038 ) ;
  assign n8040 = ( n7898 & n7900 ) | ( n7898 & n8039 ) | ( n7900 & n8039 ) ;
  assign n8041 = ( n7886 & n7888 ) | ( n7886 & n8040 ) | ( n7888 & n8040 ) ;
  assign n8042 = ( n7874 & ~n7876 ) | ( n7874 & n8041 ) | ( ~n7876 & n8041 ) ;
  assign n8043 = ( n7862 & n7864 ) | ( n7862 & n8042 ) | ( n7864 & n8042 ) ;
  assign n8044 = ( n7850 & n7852 ) | ( n7850 & n8043 ) | ( n7852 & n8043 ) ;
  assign n8045 = ( n7745 & ~n8044 ) | ( n7745 & n7840 ) | ( ~n8044 & n7840 ) ;
  assign n8047 = n2296 &  n5339 ;
  assign n8048 = n2127 | n5837 ;
  assign n8049 = n2178 | n5761 ;
  assign n8050 = n8048 &  n8049 ;
  assign n8051 = ( n8047 & ~n5339 ) | ( n8047 & n8050 ) | ( ~n5339 & n8050 ) ;
  assign n8052 = n5283 | n5341 ;
  assign n8053 = n8051 &  n8052 ;
  assign n8054 = x20 &  n8053 ;
  assign n8055 = x20 | n8053 ;
  assign n8056 = ~n8054 & n8055 ;
  assign n8057 = ( n7840 & ~n7745 ) | ( n7840 & n8044 ) | ( ~n7745 & n8044 ) ;
  assign n8058 = ( n8045 & ~n7840 ) | ( n8045 & n8057 ) | ( ~n7840 & n8057 ) ;
  assign n8059 = n8056 | n8058 ;
  assign n8060 = ( n8046 & ~n8045 ) | ( n8046 & n8059 ) | ( ~n8045 & n8059 ) ;
  assign n7835 = ( n7560 & n7746 ) | ( n7560 & n7756 ) | ( n7746 & n7756 ) ;
  assign n7836 = ( n7560 & ~n7746 ) | ( n7560 & n7756 ) | ( ~n7746 & n7756 ) ;
  assign n7837 = ( n7746 & ~n7835 ) | ( n7746 & n7836 ) | ( ~n7835 & n7836 ) ;
  assign n8061 = n1940 | n5970 ;
  assign n8062 = n1875 | n6170 ;
  assign n8063 = n8061 &  n8062 ;
  assign n8064 = ~n1748 & n6395 ;
  assign n8065 = ( n1748 & n8063 ) | ( n1748 & n8064 ) | ( n8063 & n8064 ) ;
  assign n8066 = ( n5972 & ~n4743 ) | ( n5972 & n8065 ) | ( ~n4743 & n8065 ) ;
  assign n8067 = ~n5972 & n8066 ;
  assign n8068 = ( x17 & ~n8065 ) | ( x17 & n8067 ) | ( ~n8065 & n8067 ) ;
  assign n8069 = ( n8065 & ~x17 ) | ( n8065 & n8067 ) | ( ~x17 & n8067 ) ;
  assign n8070 = ( n8068 & ~n8067 ) | ( n8068 & n8069 ) | ( ~n8067 & n8069 ) ;
  assign n8071 = ( n8060 & ~n7837 ) | ( n8060 & n8070 ) | ( ~n7837 & n8070 ) ;
  assign n7829 = ( n7491 & n7554 ) | ( n7491 & n7757 ) | ( n7554 & n7757 ) ;
  assign n7830 = ( n7554 & ~n7491 ) | ( n7554 & n7757 ) | ( ~n7491 & n7757 ) ;
  assign n7831 = ( n7491 & ~n7829 ) | ( n7491 & n7830 ) | ( ~n7829 & n7830 ) ;
  assign n7833 = ( x17 & n7764 ) | ( x17 & n7831 ) | ( n7764 & n7831 ) ;
  assign n7832 = ( n7764 & ~x17 ) | ( n7764 & n7831 ) | ( ~x17 & n7831 ) ;
  assign n7834 = ( x17 & ~n7833 ) | ( x17 & n7832 ) | ( ~n7833 & n7832 ) ;
  assign n8072 = n1378 | n7097 ;
  assign n8073 = n1566 | n6530 ;
  assign n8074 = n8072 &  n8073 ;
  assign n8075 = n1483 &  n6983 ;
  assign n8076 = ( n8074 & ~n1483 ) | ( n8074 & n8075 ) | ( ~n1483 & n8075 ) ;
  assign n8077 = ( n5038 & ~n6532 ) | ( n5038 & 1'b0 ) | ( ~n6532 & 1'b0 ) ;
  assign n8078 = ( n8076 & ~n8077 ) | ( n8076 & 1'b0 ) | ( ~n8077 & 1'b0 ) ;
  assign n8079 = x14 &  n8078 ;
  assign n8080 = x14 | n8078 ;
  assign n8081 = ~n8079 & n8080 ;
  assign n8082 = ( n8071 & ~n7834 ) | ( n8071 & n8081 ) | ( ~n7834 & n8081 ) ;
  assign n8083 = ( n7828 & ~n7818 ) | ( n7828 & n8082 ) | ( ~n7818 & n8082 ) ;
  assign n7813 = ( n7539 & n7769 ) | ( n7539 & n7779 ) | ( n7769 & n7779 ) ;
  assign n7814 = ( n7539 & ~n7769 ) | ( n7539 & n7779 ) | ( ~n7769 & n7779 ) ;
  assign n7815 = ( n7769 & ~n7813 ) | ( n7769 & n7814 ) | ( ~n7813 & n7814 ) ;
  assign n8087 = ~n946 & n7518 ;
  assign n8084 = n863 | n7783 ;
  assign n8085 = ~n1043 & n7253 ;
  assign n8086 = ( n8084 & ~n8085 ) | ( n8084 & 1'b0 ) | ( ~n8085 & 1'b0 ) ;
  assign n8088 = ( n946 & n8087 ) | ( n946 & n8086 ) | ( n8087 & n8086 ) ;
  assign n8089 = n3914 | n7255 ;
  assign n8090 = n8088 &  n8089 ;
  assign n8091 = x11 &  n8090 ;
  assign n8092 = x11 | n8090 ;
  assign n8093 = ~n8091 & n8092 ;
  assign n8094 = ( n8083 & ~n7815 ) | ( n8083 & n8093 ) | ( ~n7815 & n8093 ) ;
  assign n8113 = n7781 | n7791 ;
  assign n8114 = ( x11 & ~n8113 ) | ( x11 & n7789 ) | ( ~n8113 & n7789 ) ;
  assign n8115 = ( n7789 & ~x11 ) | ( n7789 & n8113 ) | ( ~x11 & n8113 ) ;
  assign n8116 = ( n8114 & ~n7789 ) | ( n8114 & n8115 ) | ( ~n7789 & n8115 ) ;
  assign n8095 = ~x6 & x7 ;
  assign n8096 = ( x6 & ~x7 ) | ( x6 & 1'b0 ) | ( ~x7 & 1'b0 ) ;
  assign n8097 = n8095 | n8096 ;
  assign n8101 = ( x5 & ~x6 ) | ( x5 & 1'b0 ) | ( ~x6 & 1'b0 ) ;
  assign n8102 = ~x5 & x6 ;
  assign n8103 = n8101 | n8102 ;
  assign n8098 = ( x7 & ~x8 ) | ( x7 & 1'b0 ) | ( ~x8 & 1'b0 ) ;
  assign n8099 = ~x7 & x8 ;
  assign n8100 = n8098 | n8099 ;
  assign n8104 = ( n8097 & ~n8103 ) | ( n8097 & n8100 ) | ( ~n8103 & n8100 ) ;
  assign n8105 = ~n8097 & n8104 ;
  assign n8106 = ~n599 & n8105 ;
  assign n8107 = ~n8100 | ~n8103 ;
  assign n8108 = ( n8106 & ~n3637 ) | ( n8106 & n8107 ) | ( ~n3637 & n8107 ) ;
  assign n8109 = n3637 | n8108 ;
  assign n8110 = ( x8 & ~n8106 ) | ( x8 & n8109 ) | ( ~n8106 & n8109 ) ;
  assign n8111 = ( n8106 & ~x8 ) | ( n8106 & n8109 ) | ( ~x8 & n8109 ) ;
  assign n8112 = ( n8110 & ~n8109 ) | ( n8110 & n8111 ) | ( ~n8109 & n8111 ) ;
  assign n8117 = ( n8094 & ~n8116 ) | ( n8094 & n8112 ) | ( ~n8116 & n8112 ) ;
  assign n8132 = ( n7852 & ~n7850 ) | ( n7852 & n8043 ) | ( ~n7850 & n8043 ) ;
  assign n8133 = ( n7850 & ~n8043 ) | ( n7850 & n7852 ) | ( ~n8043 & n7852 ) ;
  assign n8134 = ( n8132 & ~n7852 ) | ( n8132 & n8133 ) | ( ~n7852 & n8133 ) ;
  assign n8138 = ~n2178 & n5837 ;
  assign n8135 = ~n2392 & n5339 ;
  assign n8136 = n2296 | n5761 ;
  assign n8137 = ~n8135 & n8136 ;
  assign n8139 = ( n2178 & n8138 ) | ( n2178 & n8137 ) | ( n8138 & n8137 ) ;
  assign n8140 = ( n5341 & ~n5269 ) | ( n5341 & n8139 ) | ( ~n5269 & n8139 ) ;
  assign n8141 = ~n5341 & n8140 ;
  assign n8142 = ( x20 & ~n8139 ) | ( x20 & n8141 ) | ( ~n8139 & n8141 ) ;
  assign n8143 = ( n8139 & ~x20 ) | ( n8139 & n8141 ) | ( ~x20 & n8141 ) ;
  assign n8144 = ( n8142 & ~n8141 ) | ( n8142 & n8143 ) | ( ~n8141 & n8143 ) ;
  assign n8145 = ( n7864 & ~n7862 ) | ( n7864 & n8042 ) | ( ~n7862 & n8042 ) ;
  assign n8146 = ( n7862 & ~n8042 ) | ( n7862 & n7864 ) | ( ~n8042 & n7864 ) ;
  assign n8147 = ( n8145 & ~n7864 ) | ( n8145 & n8146 ) | ( ~n7864 & n8146 ) ;
  assign n8151 = ~n2296 & n5837 ;
  assign n8148 = ~n2483 & n5339 ;
  assign n8149 = n2392 | n5761 ;
  assign n8150 = ~n8148 & n8149 ;
  assign n8152 = ( n2296 & n8151 ) | ( n2296 & n8150 ) | ( n8151 & n8150 ) ;
  assign n8153 = ( n5500 & ~n5341 ) | ( n5500 & n8152 ) | ( ~n5341 & n8152 ) ;
  assign n8154 = ~n5500 & n8153 ;
  assign n8155 = ( x20 & ~n8152 ) | ( x20 & n8154 ) | ( ~n8152 & n8154 ) ;
  assign n8156 = ( n8152 & ~x20 ) | ( n8152 & n8154 ) | ( ~x20 & n8154 ) ;
  assign n8157 = ( n8155 & ~n8154 ) | ( n8155 & n8156 ) | ( ~n8154 & n8156 ) ;
  assign n8164 = ~n2392 & n5837 ;
  assign n8161 = ~n2569 & n5339 ;
  assign n8162 = n2483 | n5761 ;
  assign n8163 = ~n8161 & n8162 ;
  assign n8165 = ( n2392 & n8164 ) | ( n2392 & n8163 ) | ( n8164 & n8163 ) ;
  assign n8166 = ( n6212 & ~n5341 ) | ( n6212 & n8165 ) | ( ~n5341 & n8165 ) ;
  assign n8167 = ~n6212 & n8166 ;
  assign n8168 = ( x20 & ~n8165 ) | ( x20 & n8167 ) | ( ~n8165 & n8167 ) ;
  assign n8169 = ( n8165 & ~x20 ) | ( n8165 & n8167 ) | ( ~x20 & n8167 ) ;
  assign n8170 = ( n8168 & ~n8167 ) | ( n8168 & n8169 ) | ( ~n8167 & n8169 ) ;
  assign n8158 = ( n7874 & ~n8041 ) | ( n7874 & n7876 ) | ( ~n8041 & n7876 ) ;
  assign n8159 = ( n7876 & ~n7874 ) | ( n7876 & n8041 ) | ( ~n7874 & n8041 ) ;
  assign n8160 = ( n8158 & ~n7876 ) | ( n8158 & n8159 ) | ( ~n7876 & n8159 ) ;
  assign n8171 = ( n7888 & ~n7886 ) | ( n7888 & n8040 ) | ( ~n7886 & n8040 ) ;
  assign n8172 = ( n7886 & ~n8040 ) | ( n7886 & n7888 ) | ( ~n8040 & n7888 ) ;
  assign n8173 = ( n8171 & ~n7888 ) | ( n8171 & n8172 ) | ( ~n7888 & n8172 ) ;
  assign n8174 = n2665 &  n5339 ;
  assign n8175 = n2483 | n5837 ;
  assign n8176 = n2569 | n5761 ;
  assign n8177 = n8175 &  n8176 ;
  assign n8178 = ( n8174 & ~n5339 ) | ( n8174 & n8177 ) | ( ~n5339 & n8177 ) ;
  assign n8179 = ( n6465 & ~n5341 ) | ( n6465 & n8178 ) | ( ~n5341 & n8178 ) ;
  assign n8180 = ~n6465 & n8179 ;
  assign n8181 = ( x20 & ~n8178 ) | ( x20 & n8180 ) | ( ~n8178 & n8180 ) ;
  assign n8182 = ( n8178 & ~x20 ) | ( n8178 & n8180 ) | ( ~x20 & n8180 ) ;
  assign n8183 = ( n8181 & ~n8180 ) | ( n8181 & n8182 ) | ( ~n8180 & n8182 ) ;
  assign n8184 = ( n7900 & ~n7898 ) | ( n7900 & n8039 ) | ( ~n7898 & n8039 ) ;
  assign n8185 = ( n7898 & ~n8039 ) | ( n7898 & n7900 ) | ( ~n8039 & n7900 ) ;
  assign n8186 = ( n8184 & ~n7900 ) | ( n8184 & n8185 ) | ( ~n7900 & n8185 ) ;
  assign n8187 = n2751 &  n5339 ;
  assign n8188 = n2569 | n5837 ;
  assign n8189 = n2665 | n5761 ;
  assign n8190 = n8188 &  n8189 ;
  assign n8191 = ( n8187 & ~n5339 ) | ( n8187 & n8190 ) | ( ~n5339 & n8190 ) ;
  assign n8192 = ( n5705 & ~n5341 ) | ( n5705 & n8191 ) | ( ~n5341 & n8191 ) ;
  assign n8193 = ~n5705 & n8192 ;
  assign n8194 = ( x20 & ~n8191 ) | ( x20 & n8193 ) | ( ~n8191 & n8193 ) ;
  assign n8195 = ( n8191 & ~x20 ) | ( n8191 & n8193 ) | ( ~x20 & n8193 ) ;
  assign n8196 = ( n8194 & ~n8193 ) | ( n8194 & n8195 ) | ( ~n8193 & n8195 ) ;
  assign n8203 = ~n2751 & n5761 ;
  assign n8200 = n2665 | n5837 ;
  assign n8201 = ~n2783 & n5339 ;
  assign n8202 = ( n8200 & ~n8201 ) | ( n8200 & 1'b0 ) | ( ~n8201 & 1'b0 ) ;
  assign n8204 = ( n2751 & n8203 ) | ( n2751 & n8202 ) | ( n8203 & n8202 ) ;
  assign n8205 = ( n6119 & ~n5341 ) | ( n6119 & n8204 ) | ( ~n5341 & n8204 ) ;
  assign n8206 = ~n6119 & n8205 ;
  assign n8207 = ( x20 & ~n8204 ) | ( x20 & n8206 ) | ( ~n8204 & n8206 ) ;
  assign n8208 = ( n8204 & ~x20 ) | ( n8204 & n8206 ) | ( ~x20 & n8206 ) ;
  assign n8209 = ( n8207 & ~n8206 ) | ( n8207 & n8208 ) | ( ~n8206 & n8208 ) ;
  assign n8197 = ( n7910 & ~n8038 ) | ( n7910 & n7912 ) | ( ~n8038 & n7912 ) ;
  assign n8198 = ( n7912 & ~n7910 ) | ( n7912 & n8038 ) | ( ~n7910 & n8038 ) ;
  assign n8199 = ( n8197 & ~n7912 ) | ( n8197 & n8198 ) | ( ~n7912 & n8198 ) ;
  assign n8216 = ~n5339 & n2910 ;
  assign n8213 = n2751 | n5837 ;
  assign n8214 = n2783 | n5761 ;
  assign n8215 = n8213 &  n8214 ;
  assign n8217 = ( n8216 & ~n2910 ) | ( n8216 & n8215 ) | ( ~n2910 & n8215 ) ;
  assign n8218 = ( n6226 & ~n5341 ) | ( n6226 & n8217 ) | ( ~n5341 & n8217 ) ;
  assign n8219 = ~n6226 & n8218 ;
  assign n8220 = ( x20 & ~n8217 ) | ( x20 & n8219 ) | ( ~n8217 & n8219 ) ;
  assign n8221 = ( n8217 & ~x20 ) | ( n8217 & n8219 ) | ( ~x20 & n8219 ) ;
  assign n8222 = ( n8220 & ~n8219 ) | ( n8220 & n8221 ) | ( ~n8219 & n8221 ) ;
  assign n8210 = ( n7922 & ~n8037 ) | ( n7922 & n7925 ) | ( ~n8037 & n7925 ) ;
  assign n8211 = ( n7925 & ~n7922 ) | ( n7925 & n8037 ) | ( ~n7922 & n8037 ) ;
  assign n8212 = ( n8210 & ~n7925 ) | ( n8210 & n8211 ) | ( ~n7925 & n8211 ) ;
  assign n8223 = n2783 | n5837 ;
  assign n8224 = ~n2839 & n5339 ;
  assign n8225 = ( n8223 & ~n8224 ) | ( n8223 & 1'b0 ) | ( ~n8224 & 1'b0 ) ;
  assign n8226 = n2910 &  n5761 ;
  assign n8227 = ( n8225 & ~n2910 ) | ( n8225 & n8226 ) | ( ~n2910 & n8226 ) ;
  assign n8228 = ~n5341 & n6104 ;
  assign n8229 = ( n8227 & ~n8228 ) | ( n8227 & 1'b0 ) | ( ~n8228 & 1'b0 ) ;
  assign n8230 = x20 &  n8229 ;
  assign n8231 = x20 | n8229 ;
  assign n8232 = ~n8230 & n8231 ;
  assign n8233 = ( n7928 & ~n7938 ) | ( n7928 & n8036 ) | ( ~n7938 & n8036 ) ;
  assign n8234 = ( n7938 & ~n8037 ) | ( n7938 & n8233 ) | ( ~n8037 & n8233 ) ;
  assign n8235 = ~n2995 & n5339 ;
  assign n8236 = n2839 | n5761 ;
  assign n8237 = ~n8235 & n8236 ;
  assign n8238 = n2910 &  n5837 ;
  assign n8239 = ( n8237 & ~n2910 ) | ( n8237 & n8238 ) | ( ~n2910 & n8238 ) ;
  assign n8240 = ( n5341 & ~n8239 ) | ( n5341 & n6330 ) | ( ~n8239 & n6330 ) ;
  assign n8241 = ( n6330 & ~n8240 ) | ( n6330 & 1'b0 ) | ( ~n8240 & 1'b0 ) ;
  assign n8242 = ( x20 & ~n8239 ) | ( x20 & n8241 ) | ( ~n8239 & n8241 ) ;
  assign n8243 = ( n8239 & ~x20 ) | ( n8239 & n8241 ) | ( ~x20 & n8241 ) ;
  assign n8244 = ( n8242 & ~n8241 ) | ( n8242 & n8243 ) | ( ~n8241 & n8243 ) ;
  assign n8245 = ( n7941 & ~n7951 ) | ( n7941 & n8035 ) | ( ~n7951 & n8035 ) ;
  assign n8246 = ( n7951 & ~n8036 ) | ( n7951 & n8245 ) | ( ~n8036 & n8245 ) ;
  assign n8253 = ~n2839 & n5837 ;
  assign n8250 = ~n3030 & n5339 ;
  assign n8251 = n2995 | n5761 ;
  assign n8252 = ~n8250 & n8251 ;
  assign n8254 = ( n2839 & n8253 ) | ( n2839 & n8252 ) | ( n8253 & n8252 ) ;
  assign n8255 = ( n7324 & ~n5341 ) | ( n7324 & n8254 ) | ( ~n5341 & n8254 ) ;
  assign n8256 = ~n7324 & n8255 ;
  assign n8257 = ( x20 & ~n8254 ) | ( x20 & n8256 ) | ( ~n8254 & n8256 ) ;
  assign n8258 = ( n8254 & ~x20 ) | ( n8254 & n8256 ) | ( ~x20 & n8256 ) ;
  assign n8259 = ( n8257 & ~n8256 ) | ( n8257 & n8258 ) | ( ~n8256 & n8258 ) ;
  assign n8247 = ( n7963 & ~n7961 ) | ( n7963 & n8034 ) | ( ~n7961 & n8034 ) ;
  assign n8248 = ( n7961 & ~n8034 ) | ( n7961 & n7963 ) | ( ~n8034 & n7963 ) ;
  assign n8249 = ( n8247 & ~n7963 ) | ( n8247 & n8248 ) | ( ~n7963 & n8248 ) ;
  assign n8260 = ( n7976 & ~n7966 ) | ( n7976 & n8033 ) | ( ~n7966 & n8033 ) ;
  assign n8261 = ( n7966 & ~n8033 ) | ( n7966 & n7976 ) | ( ~n8033 & n7976 ) ;
  assign n8262 = ( n8260 & ~n7976 ) | ( n8260 & n8261 ) | ( ~n7976 & n8261 ) ;
  assign n8263 = ~n3106 & n5339 ;
  assign n8264 = n3030 | n5761 ;
  assign n8265 = ~n8263 & n8264 ;
  assign n8266 = ~n2995 & n5837 ;
  assign n8267 = ( n2995 & n8265 ) | ( n2995 & n8266 ) | ( n8265 & n8266 ) ;
  assign n8268 = ( n7339 & ~n5341 ) | ( n7339 & n8267 ) | ( ~n5341 & n8267 ) ;
  assign n8269 = ~n7339 & n8268 ;
  assign n8270 = ( x20 & ~n8267 ) | ( x20 & n8269 ) | ( ~n8267 & n8269 ) ;
  assign n8271 = ( n8267 & ~x20 ) | ( n8267 & n8269 ) | ( ~x20 & n8269 ) ;
  assign n8272 = ( n8270 & ~n8269 ) | ( n8270 & n8271 ) | ( ~n8269 & n8271 ) ;
  assign n8273 = ( n7986 & ~n8032 ) | ( n7986 & n7989 ) | ( ~n8032 & n7989 ) ;
  assign n8274 = ( n7989 & ~n7986 ) | ( n7989 & n8032 ) | ( ~n7986 & n8032 ) ;
  assign n8275 = ( n8273 & ~n7989 ) | ( n8273 & n8274 ) | ( ~n7989 & n8274 ) ;
  assign n8279 = ~n3030 & n5837 ;
  assign n8276 = ~n3197 & n5339 ;
  assign n8277 = n3106 | n5761 ;
  assign n8278 = ~n8276 & n8277 ;
  assign n8280 = ( n3030 & n8279 ) | ( n3030 & n8278 ) | ( n8279 & n8278 ) ;
  assign n8281 = ( n6314 & ~n5341 ) | ( n6314 & n8280 ) | ( ~n5341 & n8280 ) ;
  assign n8282 = ~n6314 & n8281 ;
  assign n8283 = ( x20 & ~n8280 ) | ( x20 & n8282 ) | ( ~n8280 & n8282 ) ;
  assign n8284 = ( n8280 & ~x20 ) | ( n8280 & n8282 ) | ( ~x20 & n8282 ) ;
  assign n8285 = ( n8283 & ~n8282 ) | ( n8283 & n8284 ) | ( ~n8282 & n8284 ) ;
  assign n8289 = ~n5339 & n3266 ;
  assign n8286 = n3106 | n5837 ;
  assign n8287 = n3197 | n5761 ;
  assign n8288 = n8286 &  n8287 ;
  assign n8290 = ( n8289 & ~n3266 ) | ( n8289 & n8288 ) | ( ~n3266 & n8288 ) ;
  assign n8291 = ( n7363 & ~n5341 ) | ( n7363 & n8290 ) | ( ~n5341 & n8290 ) ;
  assign n8292 = ~n7363 & n8291 ;
  assign n8293 = ( x20 & ~n8290 ) | ( x20 & n8292 ) | ( ~n8290 & n8292 ) ;
  assign n8294 = ( n8290 & ~x20 ) | ( n8290 & n8292 ) | ( ~x20 & n8292 ) ;
  assign n8295 = ( n8293 & ~n8292 ) | ( n8293 & n8294 ) | ( ~n8292 & n8294 ) ;
  assign n8296 = ( n8003 & ~n7993 ) | ( n8003 & n8031 ) | ( ~n7993 & n8031 ) ;
  assign n8297 = ( n8032 & ~n8003 ) | ( n8032 & n8296 ) | ( ~n8003 & n8296 ) ;
  assign n8299 = ( n7697 & n8020 ) | ( n7697 & n8030 ) | ( n8020 & n8030 ) ;
  assign n8298 = ( n7697 & ~n8020 ) | ( n7697 & n8030 ) | ( ~n8020 & n8030 ) ;
  assign n8300 = ( n8020 & ~n8299 ) | ( n8020 & n8298 ) | ( ~n8299 & n8298 ) ;
  assign n8301 = n3197 | n5837 ;
  assign n8302 = ~n3325 & n5339 ;
  assign n8303 = ( n8301 & ~n8302 ) | ( n8301 & 1'b0 ) | ( ~n8302 & 1'b0 ) ;
  assign n8304 = n3266 &  n5761 ;
  assign n8305 = ( n8303 & ~n3266 ) | ( n8303 & n8304 ) | ( ~n3266 & n8304 ) ;
  assign n8306 = ( n5341 & ~n8305 ) | ( n5341 & n7377 ) | ( ~n8305 & n7377 ) ;
  assign n8307 = ( n7377 & ~n8306 ) | ( n7377 & 1'b0 ) | ( ~n8306 & 1'b0 ) ;
  assign n8308 = ( x20 & ~n8305 ) | ( x20 & n8307 ) | ( ~n8305 & n8307 ) ;
  assign n8309 = ( n8305 & ~x20 ) | ( n8305 & n8307 ) | ( ~x20 & n8307 ) ;
  assign n8310 = ( n8308 & ~n8307 ) | ( n8308 & n8309 ) | ( ~n8307 & n8309 ) ;
  assign n8311 = ~n3361 & n5339 ;
  assign n8312 = n3325 | n5761 ;
  assign n8313 = ~n8311 & n8312 ;
  assign n8314 = n3266 &  n5837 ;
  assign n8315 = ( n8313 & ~n3266 ) | ( n8313 & n8314 ) | ( ~n3266 & n8314 ) ;
  assign n8316 = ( n5341 & ~n8315 ) | ( n5341 & n7391 ) | ( ~n8315 & n7391 ) ;
  assign n8317 = ( n7391 & ~n8316 ) | ( n7391 & 1'b0 ) | ( ~n8316 & 1'b0 ) ;
  assign n8318 = ( x20 & ~n8315 ) | ( x20 & n8317 ) | ( ~n8315 & n8317 ) ;
  assign n8319 = ( n8315 & ~x20 ) | ( n8315 & n8317 ) | ( ~x20 & n8317 ) ;
  assign n8320 = ( n8318 & ~n8317 ) | ( n8318 & n8319 ) | ( ~n8317 & n8319 ) ;
  assign n8011 = ( x23 & ~n8010 ) | ( x23 & 1'b0 ) | ( ~n8010 & 1'b0 ) ;
  assign n8322 = ( x23 & n8011 ) | ( x23 & n8018 ) | ( n8011 & n8018 ) ;
  assign n8321 = ( x23 & ~n8011 ) | ( x23 & n8018 ) | ( ~n8011 & n8018 ) ;
  assign n8323 = ( n8011 & ~n8322 ) | ( n8011 & n8321 ) | ( ~n8322 & n8321 ) ;
  assign n8324 = x23 &  n8009 ;
  assign n8325 = n8008 &  n8324 ;
  assign n8326 = n8008 | n8324 ;
  assign n8327 = ~n8325 & n8326 ;
  assign n8358 = ~n3460 & n5761 ;
  assign n8355 = n3361 | n5837 ;
  assign n8356 = ~n3601 & n5339 ;
  assign n8357 = ( n8355 & ~n8356 ) | ( n8355 & 1'b0 ) | ( ~n8356 & 1'b0 ) ;
  assign n8359 = ( n3460 & n8358 ) | ( n3460 & n8357 ) | ( n8358 & n8357 ) ;
  assign n8360 = ( n6895 & ~n5341 ) | ( n6895 & n8359 ) | ( ~n5341 & n8359 ) ;
  assign n8361 = ~n6895 & n8360 ;
  assign n8362 = ( x20 & ~n8359 ) | ( x20 & n8361 ) | ( ~n8359 & n8361 ) ;
  assign n8363 = ( n8359 & ~x20 ) | ( n8359 & n8361 ) | ( ~x20 & n8361 ) ;
  assign n8364 = ( n8362 & ~n8361 ) | ( n8362 & n8363 ) | ( ~n8361 & n8363 ) ;
  assign n8351 = ~n5341 & n6886 ;
  assign n8349 = ~n3460 & n5837 ;
  assign n8346 = ~n3547 & n5339 ;
  assign n8347 = n3601 | n5761 ;
  assign n8348 = ~n8346 & n8347 ;
  assign n8350 = ( n3460 & n8349 ) | ( n3460 & n8348 ) | ( n8349 & n8348 ) ;
  assign n8352 = ( n5341 & n8351 ) | ( n5341 & n8350 ) | ( n8351 & n8350 ) ;
  assign n8341 = n7412 | n5341 ;
  assign n8338 = n3547 | n5761 ;
  assign n8339 = n3601 | n5837 ;
  assign n8340 = n8338 &  n8339 ;
  assign n8342 = ( n5341 & ~n8341 ) | ( n5341 & n8340 ) | ( ~n8341 & n8340 ) ;
  assign n8343 = ~n3547 & n5337 ;
  assign n8344 = ( x20 & ~n8342 ) | ( x20 & n8343 ) | ( ~n8342 & n8343 ) ;
  assign n8353 = ( x20 & ~n8352 ) | ( x20 & n8344 ) | ( ~n8352 & n8344 ) ;
  assign n8354 = ( x20 & ~n8353 ) | ( x20 & 1'b0 ) | ( ~n8353 & 1'b0 ) ;
  assign n8365 = ( n8009 & ~n8364 ) | ( n8009 & n8354 ) | ( ~n8364 & n8354 ) ;
  assign n8328 = n3460 &  n5339 ;
  assign n8329 = n3325 | n5837 ;
  assign n8330 = n3361 | n5761 ;
  assign n8331 = n8329 &  n8330 ;
  assign n8332 = ( n8328 & ~n5339 ) | ( n8328 & n8331 ) | ( ~n5339 & n8331 ) ;
  assign n8333 = ( n7405 & ~n5341 ) | ( n7405 & n8332 ) | ( ~n5341 & n8332 ) ;
  assign n8334 = ~n7405 & n8333 ;
  assign n8335 = ( x20 & ~n8332 ) | ( x20 & n8334 ) | ( ~n8332 & n8334 ) ;
  assign n8336 = ( n8332 & ~x20 ) | ( n8332 & n8334 ) | ( ~x20 & n8334 ) ;
  assign n8337 = ( n8335 & ~n8334 ) | ( n8335 & n8336 ) | ( ~n8334 & n8336 ) ;
  assign n8366 = ( n8327 & ~n8365 ) | ( n8327 & n8337 ) | ( ~n8365 & n8337 ) ;
  assign n8367 = ( n8320 & n8323 ) | ( n8320 & n8366 ) | ( n8323 & n8366 ) ;
  assign n8368 = ( n8300 & n8310 ) | ( n8300 & n8367 ) | ( n8310 & n8367 ) ;
  assign n8369 = ( n8295 & ~n8297 ) | ( n8295 & n8368 ) | ( ~n8297 & n8368 ) ;
  assign n8370 = ( n8275 & n8285 ) | ( n8275 & n8369 ) | ( n8285 & n8369 ) ;
  assign n8371 = ( n8262 & n8272 ) | ( n8262 & n8370 ) | ( n8272 & n8370 ) ;
  assign n8372 = ( n8259 & ~n8249 ) | ( n8259 & n8371 ) | ( ~n8249 & n8371 ) ;
  assign n8373 = ( n8244 & n8246 ) | ( n8244 & n8372 ) | ( n8246 & n8372 ) ;
  assign n8374 = ( n8232 & n8234 ) | ( n8232 & n8373 ) | ( n8234 & n8373 ) ;
  assign n8375 = ( n8222 & ~n8212 ) | ( n8222 & n8374 ) | ( ~n8212 & n8374 ) ;
  assign n8376 = ( n8209 & ~n8199 ) | ( n8209 & n8375 ) | ( ~n8199 & n8375 ) ;
  assign n8377 = ( n8186 & n8196 ) | ( n8186 & n8376 ) | ( n8196 & n8376 ) ;
  assign n8378 = ( n8173 & n8183 ) | ( n8173 & n8377 ) | ( n8183 & n8377 ) ;
  assign n8379 = ( n8170 & ~n8160 ) | ( n8170 & n8378 ) | ( ~n8160 & n8378 ) ;
  assign n8380 = ( n8147 & n8157 ) | ( n8147 & n8379 ) | ( n8157 & n8379 ) ;
  assign n8381 = ( n8134 & n8144 ) | ( n8134 & n8380 ) | ( n8144 & n8380 ) ;
  assign n8130 = n8056 &  n8058 ;
  assign n8131 = ( n8059 & ~n8130 ) | ( n8059 & 1'b0 ) | ( ~n8130 & 1'b0 ) ;
  assign n8385 = ~n1875 & n6395 ;
  assign n8382 = n2022 | n5970 ;
  assign n8383 = n1940 | n6170 ;
  assign n8384 = n8382 &  n8383 ;
  assign n8386 = ( n1875 & n8385 ) | ( n1875 & n8384 ) | ( n8385 & n8384 ) ;
  assign n8387 = n5381 | n5972 ;
  assign n8388 = n8386 &  n8387 ;
  assign n8389 = x17 &  n8388 ;
  assign n8390 = x17 | n8388 ;
  assign n8391 = ~n8389 & n8390 ;
  assign n8392 = ( n8381 & ~n8131 ) | ( n8381 & n8391 ) | ( ~n8131 & n8391 ) ;
  assign n8127 = ( n7837 & n8060 ) | ( n7837 & n8070 ) | ( n8060 & n8070 ) ;
  assign n8128 = ( n7837 & ~n8060 ) | ( n7837 & n8070 ) | ( ~n8060 & n8070 ) ;
  assign n8129 = ( n8060 & ~n8127 ) | ( n8060 & n8128 ) | ( ~n8127 & n8128 ) ;
  assign n8393 = n1671 | n6530 ;
  assign n8394 = n1566 | n6983 ;
  assign n8395 = n8393 &  n8394 ;
  assign n8396 = n1483 &  n7097 ;
  assign n8397 = ( n8395 & ~n1483 ) | ( n8395 & n8396 ) | ( ~n1483 & n8396 ) ;
  assign n8398 = ( n4274 & n6532 ) | ( n4274 & n8397 ) | ( n6532 & n8397 ) ;
  assign n8399 = ~n6532 & n8398 ;
  assign n8400 = ( x14 & ~n8397 ) | ( x14 & n8399 ) | ( ~n8397 & n8399 ) ;
  assign n8401 = ( n8397 & ~x14 ) | ( n8397 & n8399 ) | ( ~x14 & n8399 ) ;
  assign n8402 = ( n8400 & ~n8399 ) | ( n8400 & n8401 ) | ( ~n8399 & n8401 ) ;
  assign n8403 = ( n8392 & ~n8129 ) | ( n8392 & n8402 ) | ( ~n8129 & n8402 ) ;
  assign n8121 = ( n7767 & n7831 ) | ( n7767 & n8071 ) | ( n7831 & n8071 ) ;
  assign n8122 = ( n7831 & ~n7767 ) | ( n7831 & n8071 ) | ( ~n7767 & n8071 ) ;
  assign n8123 = ( n7767 & ~n8121 ) | ( n7767 & n8122 ) | ( ~n8121 & n8122 ) ;
  assign n8125 = ( x14 & n8078 ) | ( x14 & n8123 ) | ( n8078 & n8123 ) ;
  assign n8124 = ( n8078 & ~x14 ) | ( n8078 & n8123 ) | ( ~x14 & n8123 ) ;
  assign n8126 = ( x14 & ~n8125 ) | ( x14 & n8124 ) | ( ~n8125 & n8124 ) ;
  assign n8407 = ~n7253 & n1267 ;
  assign n8404 = n1043 | n7783 ;
  assign n8405 = n1151 | n7518 ;
  assign n8406 = n8404 &  n8405 ;
  assign n8408 = ( n8407 & ~n1267 ) | ( n8407 & n8406 ) | ( ~n1267 & n8406 ) ;
  assign n8409 = n3952 | n7255 ;
  assign n8410 = n8408 &  n8409 ;
  assign n8411 = x11 &  n8410 ;
  assign n8412 = x11 | n8410 ;
  assign n8413 = ~n8411 & n8412 ;
  assign n8414 = ( n8403 & ~n8126 ) | ( n8403 & n8413 ) | ( ~n8126 & n8413 ) ;
  assign n8425 = ( n7818 & ~n8082 ) | ( n7818 & n7828 ) | ( ~n8082 & n7828 ) ;
  assign n8426 = ( n8083 & ~n7828 ) | ( n8083 & n8425 ) | ( ~n7828 & n8425 ) ;
  assign n8418 = ~n946 & n7783 ;
  assign n8415 = ~n1151 & n7253 ;
  assign n8416 = n1043 | n7518 ;
  assign n8417 = ~n8415 & n8416 ;
  assign n8419 = ( n946 & n8418 ) | ( n946 & n8417 ) | ( n8418 & n8417 ) ;
  assign n8420 = ( n7255 & ~n4038 ) | ( n7255 & n8419 ) | ( ~n4038 & n8419 ) ;
  assign n8421 = ~n7255 & n8420 ;
  assign n8422 = ( x11 & ~n8419 ) | ( x11 & n8421 ) | ( ~n8419 & n8421 ) ;
  assign n8423 = ( n8419 & ~x11 ) | ( n8419 & n8421 ) | ( ~x11 & n8421 ) ;
  assign n8424 = ( n8422 & ~n8421 ) | ( n8422 & n8423 ) | ( ~n8421 & n8423 ) ;
  assign n8427 = ( n8414 & ~n8426 ) | ( n8414 & n8424 ) | ( ~n8426 & n8424 ) ;
  assign n8437 = ( n7815 & n8083 ) | ( n7815 & n8093 ) | ( n8083 & n8093 ) ;
  assign n8438 = ( n7815 & ~n8083 ) | ( n7815 & n8093 ) | ( ~n8083 & n8093 ) ;
  assign n8439 = ( n8083 & ~n8437 ) | ( n8083 & n8438 ) | ( ~n8437 & n8438 ) ;
  assign n8428 = ~n702 & n8105 ;
  assign n8429 = ~n8097 |  n8103 ;
  assign n8430 = n599 | n8429 ;
  assign n8431 = ~n8428 & n8430 ;
  assign n8432 = ( n3937 & n8107 ) | ( n3937 & n8431 ) | ( n8107 & n8431 ) ;
  assign n8433 = ~n8107 & n8432 ;
  assign n8434 = ( x8 & ~n8431 ) | ( x8 & n8433 ) | ( ~n8431 & n8433 ) ;
  assign n8435 = ( n8431 & ~x8 ) | ( n8431 & n8433 ) | ( ~x8 & n8433 ) ;
  assign n8436 = ( n8434 & ~n8433 ) | ( n8434 & n8435 ) | ( ~n8433 & n8435 ) ;
  assign n8440 = ( n8427 & ~n8439 ) | ( n8427 & n8436 ) | ( ~n8439 & n8436 ) ;
  assign n8119 = ( n8094 & n8112 ) | ( n8094 & n8116 ) | ( n8112 & n8116 ) ;
  assign n8118 = ( n8094 & ~n8112 ) | ( n8094 & n8116 ) | ( ~n8112 & n8116 ) ;
  assign n8120 = ( n8112 & ~n8119 ) | ( n8112 & n8118 ) | ( ~n8119 & n8118 ) ;
  assign n8449 = ( n8056 & ~n8381 ) | ( n8056 & n8058 ) | ( ~n8381 & n8058 ) ;
  assign n8450 = ( n8058 & ~n8056 ) | ( n8058 & n8381 ) | ( ~n8056 & n8381 ) ;
  assign n8451 = ( n8449 & ~n8058 ) | ( n8449 & n8450 ) | ( ~n8058 & n8450 ) ;
  assign n8737 = n8391 &  n8451 ;
  assign n8452 = n2127 | n5970 ;
  assign n8453 = n2022 | n6170 ;
  assign n8454 = n8452 &  n8453 ;
  assign n8455 = ~n1940 & n6395 ;
  assign n8456 = ( n1940 & n8454 ) | ( n1940 & n8455 ) | ( n8454 & n8455 ) ;
  assign n8457 = ( n5972 & ~n5799 ) | ( n5972 & n8456 ) | ( ~n5799 & n8456 ) ;
  assign n8458 = ~n5972 & n8457 ;
  assign n8459 = ( x17 & ~n8456 ) | ( x17 & n8458 ) | ( ~n8456 & n8458 ) ;
  assign n8460 = ( n8456 & ~x17 ) | ( n8456 & n8458 ) | ( ~x17 & n8458 ) ;
  assign n8461 = ( n8459 & ~n8458 ) | ( n8459 & n8460 ) | ( ~n8458 & n8460 ) ;
  assign n8462 = ( n8134 & ~n8144 ) | ( n8134 & n8380 ) | ( ~n8144 & n8380 ) ;
  assign n8463 = ( n8144 & ~n8381 ) | ( n8144 & n8462 ) | ( ~n8381 & n8462 ) ;
  assign n8464 = n2178 | n5970 ;
  assign n8465 = n2127 | n6170 ;
  assign n8466 = n8464 &  n8465 ;
  assign n8467 = ~n2022 & n6395 ;
  assign n8468 = ( n2022 & n8466 ) | ( n2022 & n8467 ) | ( n8466 & n8467 ) ;
  assign n8469 = ( n5972 & ~n4934 ) | ( n5972 & n8468 ) | ( ~n4934 & n8468 ) ;
  assign n8470 = ~n5972 & n8469 ;
  assign n8471 = ( x17 & ~n8468 ) | ( x17 & n8470 ) | ( ~n8468 & n8470 ) ;
  assign n8472 = ( n8468 & ~x17 ) | ( n8468 & n8470 ) | ( ~x17 & n8470 ) ;
  assign n8473 = ( n8471 & ~n8470 ) | ( n8471 & n8472 ) | ( ~n8470 & n8472 ) ;
  assign n8474 = ( n8147 & ~n8157 ) | ( n8147 & n8379 ) | ( ~n8157 & n8379 ) ;
  assign n8475 = ( n8157 & ~n8380 ) | ( n8157 & n8474 ) | ( ~n8380 & n8474 ) ;
  assign n8479 = ~n2296 & n5970 ;
  assign n8476 = n2127 | n6395 ;
  assign n8477 = n2178 | n6170 ;
  assign n8478 = n8476 &  n8477 ;
  assign n8480 = ( n2296 & n8479 ) | ( n2296 & n8478 ) | ( n8479 & n8478 ) ;
  assign n8481 = ( n5972 & ~n5283 ) | ( n5972 & n8480 ) | ( ~n5283 & n8480 ) ;
  assign n8482 = ~n5972 & n8481 ;
  assign n8483 = ( x17 & ~n8480 ) | ( x17 & n8482 ) | ( ~n8480 & n8482 ) ;
  assign n8484 = ( n8480 & ~x17 ) | ( n8480 & n8482 ) | ( ~x17 & n8482 ) ;
  assign n8485 = ( n8483 & ~n8482 ) | ( n8483 & n8484 ) | ( ~n8482 & n8484 ) ;
  assign n8486 = ( n8160 & ~n8378 ) | ( n8160 & n8170 ) | ( ~n8378 & n8170 ) ;
  assign n8487 = ( n8379 & ~n8170 ) | ( n8379 & n8486 ) | ( ~n8170 & n8486 ) ;
  assign n8491 = ~n2178 & n6395 ;
  assign n8488 = n2392 | n5970 ;
  assign n8489 = n2296 | n6170 ;
  assign n8490 = n8488 &  n8489 ;
  assign n8492 = ( n2178 & n8491 ) | ( n2178 & n8490 ) | ( n8491 & n8490 ) ;
  assign n8493 = ( n5972 & ~n5269 ) | ( n5972 & n8492 ) | ( ~n5269 & n8492 ) ;
  assign n8494 = ~n5972 & n8493 ;
  assign n8495 = ( x17 & ~n8492 ) | ( x17 & n8494 ) | ( ~n8492 & n8494 ) ;
  assign n8496 = ( n8492 & ~x17 ) | ( n8492 & n8494 ) | ( ~x17 & n8494 ) ;
  assign n8497 = ( n8495 & ~n8494 ) | ( n8495 & n8496 ) | ( ~n8494 & n8496 ) ;
  assign n8498 = ( n8173 & ~n8183 ) | ( n8173 & n8377 ) | ( ~n8183 & n8377 ) ;
  assign n8499 = ( n8183 & ~n8378 ) | ( n8183 & n8498 ) | ( ~n8378 & n8498 ) ;
  assign n8503 = ~n2296 & n6395 ;
  assign n8500 = n2483 | n5970 ;
  assign n8501 = n2392 | n6170 ;
  assign n8502 = n8500 &  n8501 ;
  assign n8504 = ( n2296 & n8503 ) | ( n2296 & n8502 ) | ( n8503 & n8502 ) ;
  assign n8505 = ( n5972 & ~n5500 ) | ( n5972 & n8504 ) | ( ~n5500 & n8504 ) ;
  assign n8506 = ~n5972 & n8505 ;
  assign n8507 = ( x17 & ~n8504 ) | ( x17 & n8506 ) | ( ~n8504 & n8506 ) ;
  assign n8508 = ( n8504 & ~x17 ) | ( n8504 & n8506 ) | ( ~x17 & n8506 ) ;
  assign n8509 = ( n8507 & ~n8506 ) | ( n8507 & n8508 ) | ( ~n8506 & n8508 ) ;
  assign n8510 = ( n8186 & ~n8196 ) | ( n8186 & n8376 ) | ( ~n8196 & n8376 ) ;
  assign n8511 = ( n8196 & ~n8377 ) | ( n8196 & n8510 ) | ( ~n8377 & n8510 ) ;
  assign n8515 = ~n2392 & n6395 ;
  assign n8512 = n2569 | n5970 ;
  assign n8513 = n2483 | n6170 ;
  assign n8514 = n8512 &  n8513 ;
  assign n8516 = ( n2392 & n8515 ) | ( n2392 & n8514 ) | ( n8515 & n8514 ) ;
  assign n8517 = ( n5972 & ~n6212 ) | ( n5972 & n8516 ) | ( ~n6212 & n8516 ) ;
  assign n8518 = ~n5972 & n8517 ;
  assign n8519 = ( x17 & ~n8516 ) | ( x17 & n8518 ) | ( ~n8516 & n8518 ) ;
  assign n8520 = ( n8516 & ~x17 ) | ( n8516 & n8518 ) | ( ~x17 & n8518 ) ;
  assign n8521 = ( n8519 & ~n8518 ) | ( n8519 & n8520 ) | ( ~n8518 & n8520 ) ;
  assign n8522 = ( n8199 & ~n8375 ) | ( n8199 & n8209 ) | ( ~n8375 & n8209 ) ;
  assign n8523 = ( n8376 & ~n8209 ) | ( n8376 & n8522 ) | ( ~n8209 & n8522 ) ;
  assign n8527 = ~n2665 & n5970 ;
  assign n8524 = n2483 | n6395 ;
  assign n8525 = n2569 | n6170 ;
  assign n8526 = n8524 &  n8525 ;
  assign n8528 = ( n2665 & n8527 ) | ( n2665 & n8526 ) | ( n8527 & n8526 ) ;
  assign n8529 = ( n5972 & ~n6465 ) | ( n5972 & n8528 ) | ( ~n6465 & n8528 ) ;
  assign n8530 = ~n5972 & n8529 ;
  assign n8531 = ( x17 & ~n8528 ) | ( x17 & n8530 ) | ( ~n8528 & n8530 ) ;
  assign n8532 = ( n8528 & ~x17 ) | ( n8528 & n8530 ) | ( ~x17 & n8530 ) ;
  assign n8533 = ( n8531 & ~n8530 ) | ( n8531 & n8532 ) | ( ~n8530 & n8532 ) ;
  assign n8534 = ( n8212 & ~n8374 ) | ( n8212 & n8222 ) | ( ~n8374 & n8222 ) ;
  assign n8535 = ( n8375 & ~n8222 ) | ( n8375 & n8534 ) | ( ~n8222 & n8534 ) ;
  assign n8536 = ( n8232 & ~n8373 ) | ( n8232 & n8234 ) | ( ~n8373 & n8234 ) ;
  assign n8537 = ( n8234 & ~n8232 ) | ( n8234 & n8373 ) | ( ~n8232 & n8373 ) ;
  assign n8538 = ( n8536 & ~n8234 ) | ( n8536 & n8537 ) | ( ~n8234 & n8537 ) ;
  assign n8542 = ~n2751 & n5970 ;
  assign n8539 = n2569 | n6395 ;
  assign n8540 = n2665 | n6170 ;
  assign n8541 = n8539 &  n8540 ;
  assign n8543 = ( n2751 & n8542 ) | ( n2751 & n8541 ) | ( n8542 & n8541 ) ;
  assign n8544 = ( n5972 & ~n5705 ) | ( n5972 & n8543 ) | ( ~n5705 & n8543 ) ;
  assign n8545 = ~n5972 & n8544 ;
  assign n8546 = ( x17 & ~n8543 ) | ( x17 & n8545 ) | ( ~n8543 & n8545 ) ;
  assign n8547 = ( n8543 & ~x17 ) | ( n8543 & n8545 ) | ( ~x17 & n8545 ) ;
  assign n8548 = ( n8546 & ~n8545 ) | ( n8546 & n8547 ) | ( ~n8545 & n8547 ) ;
  assign n8549 = ( n8246 & ~n8244 ) | ( n8246 & n8372 ) | ( ~n8244 & n8372 ) ;
  assign n8550 = ( n8244 & ~n8372 ) | ( n8244 & n8246 ) | ( ~n8372 & n8246 ) ;
  assign n8551 = ( n8549 & ~n8246 ) | ( n8549 & n8550 ) | ( ~n8246 & n8550 ) ;
  assign n8555 = ~n2751 & n6170 ;
  assign n8552 = n2665 | n6395 ;
  assign n8553 = n2783 | n5970 ;
  assign n8554 = n8552 &  n8553 ;
  assign n8556 = ( n2751 & n8555 ) | ( n2751 & n8554 ) | ( n8555 & n8554 ) ;
  assign n8557 = ( n6119 & ~n5972 ) | ( n6119 & n8556 ) | ( ~n5972 & n8556 ) ;
  assign n8558 = ~n6119 & n8557 ;
  assign n8559 = ( x17 & ~n8556 ) | ( x17 & n8558 ) | ( ~n8556 & n8558 ) ;
  assign n8560 = ( n8556 & ~x17 ) | ( n8556 & n8558 ) | ( ~x17 & n8558 ) ;
  assign n8561 = ( n8559 & ~n8558 ) | ( n8559 & n8560 ) | ( ~n8558 & n8560 ) ;
  assign n8562 = n2751 | n6395 ;
  assign n8563 = n2783 | n6170 ;
  assign n8564 = n8562 &  n8563 ;
  assign n8565 = n2910 &  n5970 ;
  assign n8566 = ( n8564 & ~n2910 ) | ( n8564 & n8565 ) | ( ~n2910 & n8565 ) ;
  assign n8567 = ( n6226 & ~n5972 ) | ( n6226 & n8566 ) | ( ~n5972 & n8566 ) ;
  assign n8568 = ~n6226 & n8567 ;
  assign n8569 = ( x17 & ~n8566 ) | ( x17 & n8568 ) | ( ~n8566 & n8568 ) ;
  assign n8570 = ( n8566 & ~x17 ) | ( n8566 & n8568 ) | ( ~x17 & n8568 ) ;
  assign n8571 = ( n8569 & ~n8568 ) | ( n8569 & n8570 ) | ( ~n8568 & n8570 ) ;
  assign n8572 = ( n8249 & ~n8371 ) | ( n8249 & n8259 ) | ( ~n8371 & n8259 ) ;
  assign n8573 = ( n8372 & ~n8259 ) | ( n8372 & n8572 ) | ( ~n8259 & n8572 ) ;
  assign n8574 = n2783 | n6395 ;
  assign n8575 = n2839 | n5970 ;
  assign n8576 = n8574 &  n8575 ;
  assign n8577 = n2910 &  n6170 ;
  assign n8578 = ( n8576 & ~n2910 ) | ( n8576 & n8577 ) | ( ~n2910 & n8577 ) ;
  assign n8579 = ~n5972 & n6104 ;
  assign n8580 = ( n8578 & ~n8579 ) | ( n8578 & 1'b0 ) | ( ~n8579 & 1'b0 ) ;
  assign n8581 = x17 &  n8580 ;
  assign n8582 = x17 | n8580 ;
  assign n8583 = ~n8581 & n8582 ;
  assign n8584 = ( n8262 & ~n8272 ) | ( n8262 & n8370 ) | ( ~n8272 & n8370 ) ;
  assign n8585 = ( n8272 & ~n8371 ) | ( n8272 & n8584 ) | ( ~n8371 & n8584 ) ;
  assign n8586 = n2995 | n5970 ;
  assign n8587 = n2839 | n6170 ;
  assign n8588 = n8586 &  n8587 ;
  assign n8589 = n2910 &  n6395 ;
  assign n8590 = ( n8588 & ~n2910 ) | ( n8588 & n8589 ) | ( ~n2910 & n8589 ) ;
  assign n8591 = ( n5972 & ~n8590 ) | ( n5972 & n6330 ) | ( ~n8590 & n6330 ) ;
  assign n8592 = ( n6330 & ~n8591 ) | ( n6330 & 1'b0 ) | ( ~n8591 & 1'b0 ) ;
  assign n8593 = ( x17 & ~n8590 ) | ( x17 & n8592 ) | ( ~n8590 & n8592 ) ;
  assign n8594 = ( n8590 & ~x17 ) | ( n8590 & n8592 ) | ( ~x17 & n8592 ) ;
  assign n8595 = ( n8593 & ~n8592 ) | ( n8593 & n8594 ) | ( ~n8592 & n8594 ) ;
  assign n8596 = ( n8275 & ~n8285 ) | ( n8275 & n8369 ) | ( ~n8285 & n8369 ) ;
  assign n8597 = ( n8285 & ~n8370 ) | ( n8285 & n8596 ) | ( ~n8370 & n8596 ) ;
  assign n8604 = ~n2839 & n6395 ;
  assign n8601 = n3030 | n5970 ;
  assign n8602 = n2995 | n6170 ;
  assign n8603 = n8601 &  n8602 ;
  assign n8605 = ( n2839 & n8604 ) | ( n2839 & n8603 ) | ( n8604 & n8603 ) ;
  assign n8606 = ( n7324 & ~n5972 ) | ( n7324 & n8605 ) | ( ~n5972 & n8605 ) ;
  assign n8607 = ~n7324 & n8606 ;
  assign n8608 = ( x17 & ~n8605 ) | ( x17 & n8607 ) | ( ~n8605 & n8607 ) ;
  assign n8609 = ( n8605 & ~x17 ) | ( n8605 & n8607 ) | ( ~x17 & n8607 ) ;
  assign n8610 = ( n8608 & ~n8607 ) | ( n8608 & n8609 ) | ( ~n8607 & n8609 ) ;
  assign n8598 = ( n8297 & ~n8295 ) | ( n8297 & n8368 ) | ( ~n8295 & n8368 ) ;
  assign n8599 = ( n8295 & ~n8368 ) | ( n8295 & n8297 ) | ( ~n8368 & n8297 ) ;
  assign n8600 = ( n8598 & ~n8297 ) | ( n8598 & n8599 ) | ( ~n8297 & n8599 ) ;
  assign n8611 = ( n8310 & ~n8300 ) | ( n8310 & n8367 ) | ( ~n8300 & n8367 ) ;
  assign n8612 = ( n8300 & ~n8367 ) | ( n8300 & n8310 ) | ( ~n8367 & n8310 ) ;
  assign n8613 = ( n8611 & ~n8310 ) | ( n8611 & n8612 ) | ( ~n8310 & n8612 ) ;
  assign n8614 = n3106 | n5970 ;
  assign n8615 = n3030 | n6170 ;
  assign n8616 = n8614 &  n8615 ;
  assign n8617 = ~n2995 & n6395 ;
  assign n8618 = ( n2995 & n8616 ) | ( n2995 & n8617 ) | ( n8616 & n8617 ) ;
  assign n8619 = ( n7339 & ~n5972 ) | ( n7339 & n8618 ) | ( ~n5972 & n8618 ) ;
  assign n8620 = ~n7339 & n8619 ;
  assign n8621 = ( x17 & ~n8618 ) | ( x17 & n8620 ) | ( ~n8618 & n8620 ) ;
  assign n8622 = ( n8618 & ~x17 ) | ( n8618 & n8620 ) | ( ~x17 & n8620 ) ;
  assign n8623 = ( n8621 & ~n8620 ) | ( n8621 & n8622 ) | ( ~n8620 & n8622 ) ;
  assign n8624 = ( n8320 & ~n8366 ) | ( n8320 & n8323 ) | ( ~n8366 & n8323 ) ;
  assign n8625 = ( n8323 & ~n8320 ) | ( n8323 & n8366 ) | ( ~n8320 & n8366 ) ;
  assign n8626 = ( n8624 & ~n8323 ) | ( n8624 & n8625 ) | ( ~n8323 & n8625 ) ;
  assign n8630 = ~n3030 & n6395 ;
  assign n8627 = n3197 | n5970 ;
  assign n8628 = n3106 | n6170 ;
  assign n8629 = n8627 &  n8628 ;
  assign n8631 = ( n3030 & n8630 ) | ( n3030 & n8629 ) | ( n8630 & n8629 ) ;
  assign n8632 = ( n6314 & ~n5972 ) | ( n6314 & n8631 ) | ( ~n5972 & n8631 ) ;
  assign n8633 = ~n6314 & n8632 ;
  assign n8634 = ( x17 & ~n8631 ) | ( x17 & n8633 ) | ( ~n8631 & n8633 ) ;
  assign n8635 = ( n8631 & ~x17 ) | ( n8631 & n8633 ) | ( ~x17 & n8633 ) ;
  assign n8636 = ( n8634 & ~n8633 ) | ( n8634 & n8635 ) | ( ~n8633 & n8635 ) ;
  assign n8637 = n3106 | n6395 ;
  assign n8638 = n3197 | n6170 ;
  assign n8639 = n8637 &  n8638 ;
  assign n8640 = n3266 &  n5970 ;
  assign n8641 = ( n8639 & ~n3266 ) | ( n8639 & n8640 ) | ( ~n3266 & n8640 ) ;
  assign n8642 = ( n7363 & ~n5972 ) | ( n7363 & n8641 ) | ( ~n5972 & n8641 ) ;
  assign n8643 = ~n7363 & n8642 ;
  assign n8644 = ( x17 & ~n8641 ) | ( x17 & n8643 ) | ( ~n8641 & n8643 ) ;
  assign n8645 = ( n8641 & ~x17 ) | ( n8641 & n8643 ) | ( ~x17 & n8643 ) ;
  assign n8646 = ( n8644 & ~n8643 ) | ( n8644 & n8645 ) | ( ~n8643 & n8645 ) ;
  assign n8647 = ( n8337 & ~n8327 ) | ( n8337 & n8365 ) | ( ~n8327 & n8365 ) ;
  assign n8648 = ( n8366 & ~n8337 ) | ( n8366 & n8647 ) | ( ~n8337 & n8647 ) ;
  assign n8650 = ( n8009 & n8354 ) | ( n8009 & n8364 ) | ( n8354 & n8364 ) ;
  assign n8649 = ( n8009 & ~n8354 ) | ( n8009 & n8364 ) | ( ~n8354 & n8364 ) ;
  assign n8651 = ( n8354 & ~n8650 ) | ( n8354 & n8649 ) | ( ~n8650 & n8649 ) ;
  assign n8652 = n3197 | n6395 ;
  assign n8653 = n3325 | n5970 ;
  assign n8654 = n8652 &  n8653 ;
  assign n8655 = n3266 &  n6170 ;
  assign n8656 = ( n8654 & ~n3266 ) | ( n8654 & n8655 ) | ( ~n3266 & n8655 ) ;
  assign n8657 = ( n5972 & ~n8656 ) | ( n5972 & n7377 ) | ( ~n8656 & n7377 ) ;
  assign n8658 = ( n7377 & ~n8657 ) | ( n7377 & 1'b0 ) | ( ~n8657 & 1'b0 ) ;
  assign n8659 = ( x17 & ~n8656 ) | ( x17 & n8658 ) | ( ~n8656 & n8658 ) ;
  assign n8660 = ( n8656 & ~x17 ) | ( n8656 & n8658 ) | ( ~x17 & n8658 ) ;
  assign n8661 = ( n8659 & ~n8658 ) | ( n8659 & n8660 ) | ( ~n8658 & n8660 ) ;
  assign n8662 = n3361 | n5970 ;
  assign n8663 = n3325 | n6170 ;
  assign n8664 = n8662 &  n8663 ;
  assign n8665 = n3266 &  n6395 ;
  assign n8666 = ( n8664 & ~n3266 ) | ( n8664 & n8665 ) | ( ~n3266 & n8665 ) ;
  assign n8667 = ( n5972 & ~n8666 ) | ( n5972 & n7391 ) | ( ~n8666 & n7391 ) ;
  assign n8668 = ( n7391 & ~n8667 ) | ( n7391 & 1'b0 ) | ( ~n8667 & 1'b0 ) ;
  assign n8669 = ( x17 & ~n8666 ) | ( x17 & n8668 ) | ( ~n8666 & n8668 ) ;
  assign n8670 = ( n8666 & ~x17 ) | ( n8666 & n8668 ) | ( ~x17 & n8668 ) ;
  assign n8671 = ( n8669 & ~n8668 ) | ( n8669 & n8670 ) | ( ~n8668 & n8670 ) ;
  assign n8345 = ( x20 & ~n8344 ) | ( x20 & 1'b0 ) | ( ~n8344 & 1'b0 ) ;
  assign n8673 = ( x20 & n8345 ) | ( x20 & n8352 ) | ( n8345 & n8352 ) ;
  assign n8672 = ( x20 & ~n8345 ) | ( x20 & n8352 ) | ( ~n8345 & n8352 ) ;
  assign n8674 = ( n8345 & ~n8673 ) | ( n8345 & n8672 ) | ( ~n8673 & n8672 ) ;
  assign n8675 = x20 &  n8343 ;
  assign n8676 = n8342 &  n8675 ;
  assign n8677 = n8342 | n8675 ;
  assign n8678 = ~n8676 & n8677 ;
  assign n8709 = ~n3460 & n6170 ;
  assign n8706 = n3361 | n6395 ;
  assign n8707 = n3601 | n5970 ;
  assign n8708 = n8706 &  n8707 ;
  assign n8710 = ( n3460 & n8709 ) | ( n3460 & n8708 ) | ( n8709 & n8708 ) ;
  assign n8711 = ( n6895 & ~n5972 ) | ( n6895 & n8710 ) | ( ~n5972 & n8710 ) ;
  assign n8712 = ~n6895 & n8711 ;
  assign n8713 = ( x17 & ~n8710 ) | ( x17 & n8712 ) | ( ~n8710 & n8712 ) ;
  assign n8714 = ( n8710 & ~x17 ) | ( n8710 & n8712 ) | ( ~x17 & n8712 ) ;
  assign n8715 = ( n8713 & ~n8712 ) | ( n8713 & n8714 ) | ( ~n8712 & n8714 ) ;
  assign n8702 = ~n5972 & n6886 ;
  assign n8700 = ~n3460 & n6395 ;
  assign n8697 = n3547 | n5970 ;
  assign n8698 = n3601 | n6170 ;
  assign n8699 = n8697 &  n8698 ;
  assign n8701 = ( n3460 & n8700 ) | ( n3460 & n8699 ) | ( n8700 & n8699 ) ;
  assign n8703 = ( n5972 & n8702 ) | ( n5972 & n8701 ) | ( n8702 & n8701 ) ;
  assign n8692 = n7412 | n5972 ;
  assign n8689 = n3547 | n6170 ;
  assign n8690 = n3601 | n6395 ;
  assign n8691 = n8689 &  n8690 ;
  assign n8693 = ( n5972 & ~n8692 ) | ( n5972 & n8691 ) | ( ~n8692 & n8691 ) ;
  assign n8694 = ~n3547 & n5965 ;
  assign n8695 = ( x17 & ~n8693 ) | ( x17 & n8694 ) | ( ~n8693 & n8694 ) ;
  assign n8704 = ( x17 & ~n8703 ) | ( x17 & n8695 ) | ( ~n8703 & n8695 ) ;
  assign n8705 = ( x17 & ~n8704 ) | ( x17 & 1'b0 ) | ( ~n8704 & 1'b0 ) ;
  assign n8716 = ( n8343 & ~n8715 ) | ( n8343 & n8705 ) | ( ~n8715 & n8705 ) ;
  assign n8682 = ~n3460 & n5970 ;
  assign n8679 = n3325 | n6395 ;
  assign n8680 = n3361 | n6170 ;
  assign n8681 = n8679 &  n8680 ;
  assign n8683 = ( n3460 & n8682 ) | ( n3460 & n8681 ) | ( n8682 & n8681 ) ;
  assign n8684 = ( n7405 & ~n5972 ) | ( n7405 & n8683 ) | ( ~n5972 & n8683 ) ;
  assign n8685 = ~n7405 & n8684 ;
  assign n8686 = ( x17 & ~n8683 ) | ( x17 & n8685 ) | ( ~n8683 & n8685 ) ;
  assign n8687 = ( n8683 & ~x17 ) | ( n8683 & n8685 ) | ( ~x17 & n8685 ) ;
  assign n8688 = ( n8686 & ~n8685 ) | ( n8686 & n8687 ) | ( ~n8685 & n8687 ) ;
  assign n8717 = ( n8678 & ~n8716 ) | ( n8678 & n8688 ) | ( ~n8716 & n8688 ) ;
  assign n8718 = ( n8671 & n8674 ) | ( n8671 & n8717 ) | ( n8674 & n8717 ) ;
  assign n8719 = ( n8651 & n8661 ) | ( n8651 & n8718 ) | ( n8661 & n8718 ) ;
  assign n8720 = ( n8646 & ~n8648 ) | ( n8646 & n8719 ) | ( ~n8648 & n8719 ) ;
  assign n8721 = ( n8626 & n8636 ) | ( n8626 & n8720 ) | ( n8636 & n8720 ) ;
  assign n8722 = ( n8613 & n8623 ) | ( n8613 & n8721 ) | ( n8623 & n8721 ) ;
  assign n8723 = ( n8610 & ~n8600 ) | ( n8610 & n8722 ) | ( ~n8600 & n8722 ) ;
  assign n8724 = ( n8595 & n8597 ) | ( n8595 & n8723 ) | ( n8597 & n8723 ) ;
  assign n8725 = ( n8583 & n8585 ) | ( n8583 & n8724 ) | ( n8585 & n8724 ) ;
  assign n8726 = ( n8571 & ~n8573 ) | ( n8571 & n8725 ) | ( ~n8573 & n8725 ) ;
  assign n8727 = ( n8551 & n8561 ) | ( n8551 & n8726 ) | ( n8561 & n8726 ) ;
  assign n8728 = ( n8538 & n8548 ) | ( n8538 & n8727 ) | ( n8548 & n8727 ) ;
  assign n8729 = ( n8533 & ~n8535 ) | ( n8533 & n8728 ) | ( ~n8535 & n8728 ) ;
  assign n8730 = ( n8521 & ~n8523 ) | ( n8521 & n8729 ) | ( ~n8523 & n8729 ) ;
  assign n8731 = ( n8509 & n8511 ) | ( n8509 & n8730 ) | ( n8511 & n8730 ) ;
  assign n8732 = ( n8497 & n8499 ) | ( n8497 & n8731 ) | ( n8499 & n8731 ) ;
  assign n8733 = ( n8485 & ~n8487 ) | ( n8485 & n8732 ) | ( ~n8487 & n8732 ) ;
  assign n8734 = ( n8473 & n8475 ) | ( n8473 & n8733 ) | ( n8475 & n8733 ) ;
  assign n8735 = ( n8461 & n8463 ) | ( n8461 & n8734 ) | ( n8463 & n8734 ) ;
  assign n8736 = ( n8391 & ~n8735 ) | ( n8391 & n8451 ) | ( ~n8735 & n8451 ) ;
  assign n8741 = ~n1566 & n7097 ;
  assign n8738 = n1748 | n6530 ;
  assign n8739 = n1671 | n6983 ;
  assign n8740 = n8738 &  n8739 ;
  assign n8742 = ( n1566 & n8741 ) | ( n1566 & n8740 ) | ( n8741 & n8740 ) ;
  assign n8743 = n4597 | n6532 ;
  assign n8744 = n8742 &  n8743 ;
  assign n8745 = x14 &  n8744 ;
  assign n8746 = x14 | n8744 ;
  assign n8747 = ~n8745 & n8746 ;
  assign n8748 = ( n8451 & ~n8391 ) | ( n8451 & n8735 ) | ( ~n8391 & n8735 ) ;
  assign n8749 = ( n8736 & ~n8451 ) | ( n8736 & n8748 ) | ( ~n8451 & n8748 ) ;
  assign n8750 = n8747 | n8749 ;
  assign n8751 = ( n8737 & ~n8736 ) | ( n8737 & n8750 ) | ( ~n8736 & n8750 ) ;
  assign n8446 = ( n8129 & n8392 ) | ( n8129 & n8402 ) | ( n8392 & n8402 ) ;
  assign n8447 = ( n8129 & ~n8392 ) | ( n8129 & n8402 ) | ( ~n8392 & n8402 ) ;
  assign n8448 = ( n8392 & ~n8446 ) | ( n8392 & n8447 ) | ( ~n8446 & n8447 ) ;
  assign n8752 = n1151 | n7783 ;
  assign n8753 = ~n1378 & n7253 ;
  assign n8754 = ( n8752 & ~n8753 ) | ( n8752 & 1'b0 ) | ( ~n8753 & 1'b0 ) ;
  assign n8755 = n1267 &  n7518 ;
  assign n8756 = ( n8754 & ~n1267 ) | ( n8754 & n8755 ) | ( ~n1267 & n8755 ) ;
  assign n8757 = ( n4061 & n7255 ) | ( n4061 & n8756 ) | ( n7255 & n8756 ) ;
  assign n8758 = ~n7255 & n8757 ;
  assign n8759 = ( x11 & ~n8756 ) | ( x11 & n8758 ) | ( ~n8756 & n8758 ) ;
  assign n8760 = ( n8756 & ~x11 ) | ( n8756 & n8758 ) | ( ~x11 & n8758 ) ;
  assign n8761 = ( n8759 & ~n8758 ) | ( n8759 & n8760 ) | ( ~n8758 & n8760 ) ;
  assign n8762 = ( n8751 & ~n8448 ) | ( n8751 & n8761 ) | ( ~n8448 & n8761 ) ;
  assign n8441 = ( x14 & ~n8123 ) | ( x14 & n8078 ) | ( ~n8123 & n8078 ) ;
  assign n8442 = ( n8124 & ~n8078 ) | ( n8124 & n8441 ) | ( ~n8078 & n8441 ) ;
  assign n8443 = ( n8413 & ~n8403 ) | ( n8413 & n8442 ) | ( ~n8403 & n8442 ) ;
  assign n8444 = ( n8403 & ~n8413 ) | ( n8403 & n8442 ) | ( ~n8413 & n8442 ) ;
  assign n8445 = ( n8443 & ~n8442 ) | ( n8443 & n8444 ) | ( ~n8442 & n8444 ) ;
  assign n8763 = n946 &  n8105 ;
  assign n8764 = ~n8103 |  n8100 ;
  assign n8765 = n702 | n8764 ;
  assign n8766 = n863 | n8429 ;
  assign n8767 = n8765 &  n8766 ;
  assign n8768 = ( n8763 & ~n8105 ) | ( n8763 & n8767 ) | ( ~n8105 & n8767 ) ;
  assign n8769 = ( n8107 & ~n3650 ) | ( n8107 & n8768 ) | ( ~n3650 & n8768 ) ;
  assign n8770 = ~n8107 & n8769 ;
  assign n8771 = ( x8 & ~n8768 ) | ( x8 & n8770 ) | ( ~n8768 & n8770 ) ;
  assign n8772 = ( n8768 & ~x8 ) | ( n8768 & n8770 ) | ( ~x8 & n8770 ) ;
  assign n8773 = ( n8771 & ~n8770 ) | ( n8771 & n8772 ) | ( ~n8770 & n8772 ) ;
  assign n8774 = ( n8762 & ~n8445 ) | ( n8762 & n8773 ) | ( ~n8445 & n8773 ) ;
  assign n8785 = ( n8424 & ~n8414 ) | ( n8424 & n8426 ) | ( ~n8414 & n8426 ) ;
  assign n8786 = ( n8427 & ~n8424 ) | ( n8427 & n8785 ) | ( ~n8424 & n8785 ) ;
  assign n8775 = n863 &  n8105 ;
  assign n8776 = n599 | n8764 ;
  assign n8777 = n702 | n8429 ;
  assign n8778 = n8776 &  n8777 ;
  assign n8779 = ( n8775 & ~n8105 ) | ( n8775 & n8778 ) | ( ~n8105 & n8778 ) ;
  assign n8780 = ( n8107 & ~n4452 ) | ( n8107 & n8779 ) | ( ~n4452 & n8779 ) ;
  assign n8781 = ~n8107 & n8780 ;
  assign n8782 = ( x8 & ~n8779 ) | ( x8 & n8781 ) | ( ~n8779 & n8781 ) ;
  assign n8783 = ( n8779 & ~x8 ) | ( n8779 & n8781 ) | ( ~x8 & n8781 ) ;
  assign n8784 = ( n8782 & ~n8781 ) | ( n8782 & n8783 ) | ( ~n8781 & n8783 ) ;
  assign n8787 = ( n8774 & ~n8786 ) | ( n8774 & n8784 ) | ( ~n8786 & n8784 ) ;
  assign n8789 = ( n8427 & n8436 ) | ( n8427 & n8439 ) | ( n8436 & n8439 ) ;
  assign n8788 = ( n8427 & ~n8436 ) | ( n8427 & n8439 ) | ( ~n8436 & n8439 ) ;
  assign n8790 = ( n8436 & ~n8789 ) | ( n8436 & n8788 ) | ( ~n8789 & n8788 ) ;
  assign n8794 = ( n8463 & ~n8461 ) | ( n8463 & n8734 ) | ( ~n8461 & n8734 ) ;
  assign n8795 = ( n8461 & ~n8734 ) | ( n8461 & n8463 ) | ( ~n8734 & n8463 ) ;
  assign n8796 = ( n8794 & ~n8463 ) | ( n8794 & n8795 ) | ( ~n8463 & n8795 ) ;
  assign n8800 = ~n1875 & n6530 ;
  assign n8797 = n1671 | n7097 ;
  assign n8798 = n1748 | n6983 ;
  assign n8799 = n8797 &  n8798 ;
  assign n8801 = ( n1875 & n8800 ) | ( n1875 & n8799 ) | ( n8800 & n8799 ) ;
  assign n8802 = ( n6532 & ~n4580 ) | ( n6532 & n8801 ) | ( ~n4580 & n8801 ) ;
  assign n8803 = ~n6532 & n8802 ;
  assign n8804 = ( x14 & ~n8801 ) | ( x14 & n8803 ) | ( ~n8801 & n8803 ) ;
  assign n8805 = ( n8801 & ~x14 ) | ( n8801 & n8803 ) | ( ~x14 & n8803 ) ;
  assign n8806 = ( n8804 & ~n8803 ) | ( n8804 & n8805 ) | ( ~n8803 & n8805 ) ;
  assign n8807 = ( n8475 & ~n8473 ) | ( n8475 & n8733 ) | ( ~n8473 & n8733 ) ;
  assign n8808 = ( n8473 & ~n8733 ) | ( n8473 & n8475 ) | ( ~n8733 & n8475 ) ;
  assign n8809 = ( n8807 & ~n8475 ) | ( n8807 & n8808 ) | ( ~n8475 & n8808 ) ;
  assign n8810 = n1940 | n6530 ;
  assign n8811 = n1875 | n6983 ;
  assign n8812 = n8810 &  n8811 ;
  assign n8813 = ~n1748 & n7097 ;
  assign n8814 = ( n1748 & n8812 ) | ( n1748 & n8813 ) | ( n8812 & n8813 ) ;
  assign n8815 = ( n6532 & ~n4743 ) | ( n6532 & n8814 ) | ( ~n4743 & n8814 ) ;
  assign n8816 = ~n6532 & n8815 ;
  assign n8817 = ( x14 & ~n8814 ) | ( x14 & n8816 ) | ( ~n8814 & n8816 ) ;
  assign n8818 = ( n8814 & ~x14 ) | ( n8814 & n8816 ) | ( ~x14 & n8816 ) ;
  assign n8819 = ( n8817 & ~n8816 ) | ( n8817 & n8818 ) | ( ~n8816 & n8818 ) ;
  assign n8826 = ~n1875 & n7097 ;
  assign n8823 = n2022 | n6530 ;
  assign n8824 = n1940 | n6983 ;
  assign n8825 = n8823 &  n8824 ;
  assign n8827 = ( n1875 & n8826 ) | ( n1875 & n8825 ) | ( n8826 & n8825 ) ;
  assign n8828 = ( n6532 & ~n5381 ) | ( n6532 & n8827 ) | ( ~n5381 & n8827 ) ;
  assign n8829 = ~n6532 & n8828 ;
  assign n8830 = ( x14 & ~n8827 ) | ( x14 & n8829 ) | ( ~n8827 & n8829 ) ;
  assign n8831 = ( n8827 & ~x14 ) | ( n8827 & n8829 ) | ( ~x14 & n8829 ) ;
  assign n8832 = ( n8830 & ~n8829 ) | ( n8830 & n8831 ) | ( ~n8829 & n8831 ) ;
  assign n8820 = ( n8485 & ~n8732 ) | ( n8485 & n8487 ) | ( ~n8732 & n8487 ) ;
  assign n8821 = ( n8487 & ~n8485 ) | ( n8487 & n8732 ) | ( ~n8485 & n8732 ) ;
  assign n8822 = ( n8820 & ~n8487 ) | ( n8820 & n8821 ) | ( ~n8487 & n8821 ) ;
  assign n8833 = ( n8499 & ~n8497 ) | ( n8499 & n8731 ) | ( ~n8497 & n8731 ) ;
  assign n8834 = ( n8497 & ~n8731 ) | ( n8497 & n8499 ) | ( ~n8731 & n8499 ) ;
  assign n8835 = ( n8833 & ~n8499 ) | ( n8833 & n8834 ) | ( ~n8499 & n8834 ) ;
  assign n8836 = n2127 | n6530 ;
  assign n8837 = n2022 | n6983 ;
  assign n8838 = n8836 &  n8837 ;
  assign n8839 = ~n1940 & n7097 ;
  assign n8840 = ( n1940 & n8838 ) | ( n1940 & n8839 ) | ( n8838 & n8839 ) ;
  assign n8841 = ( n6532 & ~n5799 ) | ( n6532 & n8840 ) | ( ~n5799 & n8840 ) ;
  assign n8842 = ~n6532 & n8841 ;
  assign n8843 = ( x14 & ~n8840 ) | ( x14 & n8842 ) | ( ~n8840 & n8842 ) ;
  assign n8844 = ( n8840 & ~x14 ) | ( n8840 & n8842 ) | ( ~x14 & n8842 ) ;
  assign n8845 = ( n8843 & ~n8842 ) | ( n8843 & n8844 ) | ( ~n8842 & n8844 ) ;
  assign n8846 = ( n8511 & ~n8509 ) | ( n8511 & n8730 ) | ( ~n8509 & n8730 ) ;
  assign n8847 = ( n8509 & ~n8730 ) | ( n8509 & n8511 ) | ( ~n8730 & n8511 ) ;
  assign n8848 = ( n8846 & ~n8511 ) | ( n8846 & n8847 ) | ( ~n8511 & n8847 ) ;
  assign n8849 = n2178 | n6530 ;
  assign n8850 = n2127 | n6983 ;
  assign n8851 = n8849 &  n8850 ;
  assign n8852 = ~n2022 & n7097 ;
  assign n8853 = ( n2022 & n8851 ) | ( n2022 & n8852 ) | ( n8851 & n8852 ) ;
  assign n8854 = ( n6532 & ~n4934 ) | ( n6532 & n8853 ) | ( ~n4934 & n8853 ) ;
  assign n8855 = ~n6532 & n8854 ;
  assign n8856 = ( x14 & ~n8853 ) | ( x14 & n8855 ) | ( ~n8853 & n8855 ) ;
  assign n8857 = ( n8853 & ~x14 ) | ( n8853 & n8855 ) | ( ~x14 & n8855 ) ;
  assign n8858 = ( n8856 & ~n8855 ) | ( n8856 & n8857 ) | ( ~n8855 & n8857 ) ;
  assign n8865 = ~n2296 & n6530 ;
  assign n8862 = n2127 | n7097 ;
  assign n8863 = n2178 | n6983 ;
  assign n8864 = n8862 &  n8863 ;
  assign n8866 = ( n2296 & n8865 ) | ( n2296 & n8864 ) | ( n8865 & n8864 ) ;
  assign n8867 = ( n6532 & ~n5283 ) | ( n6532 & n8866 ) | ( ~n5283 & n8866 ) ;
  assign n8868 = ~n6532 & n8867 ;
  assign n8869 = ( x14 & ~n8866 ) | ( x14 & n8868 ) | ( ~n8866 & n8868 ) ;
  assign n8870 = ( n8866 & ~x14 ) | ( n8866 & n8868 ) | ( ~x14 & n8868 ) ;
  assign n8871 = ( n8869 & ~n8868 ) | ( n8869 & n8870 ) | ( ~n8868 & n8870 ) ;
  assign n8859 = ( n8521 & ~n8729 ) | ( n8521 & n8523 ) | ( ~n8729 & n8523 ) ;
  assign n8860 = ( n8523 & ~n8521 ) | ( n8523 & n8729 ) | ( ~n8521 & n8729 ) ;
  assign n8861 = ( n8859 & ~n8523 ) | ( n8859 & n8860 ) | ( ~n8523 & n8860 ) ;
  assign n8878 = ~n2178 & n7097 ;
  assign n8875 = n2392 | n6530 ;
  assign n8876 = n2296 | n6983 ;
  assign n8877 = n8875 &  n8876 ;
  assign n8879 = ( n2178 & n8878 ) | ( n2178 & n8877 ) | ( n8878 & n8877 ) ;
  assign n8880 = ( n6532 & ~n5269 ) | ( n6532 & n8879 ) | ( ~n5269 & n8879 ) ;
  assign n8881 = ~n6532 & n8880 ;
  assign n8882 = ( x14 & ~n8879 ) | ( x14 & n8881 ) | ( ~n8879 & n8881 ) ;
  assign n8883 = ( n8879 & ~x14 ) | ( n8879 & n8881 ) | ( ~x14 & n8881 ) ;
  assign n8884 = ( n8882 & ~n8881 ) | ( n8882 & n8883 ) | ( ~n8881 & n8883 ) ;
  assign n8872 = ( n8533 & ~n8728 ) | ( n8533 & n8535 ) | ( ~n8728 & n8535 ) ;
  assign n8873 = ( n8535 & ~n8533 ) | ( n8535 & n8728 ) | ( ~n8533 & n8728 ) ;
  assign n8874 = ( n8872 & ~n8535 ) | ( n8872 & n8873 ) | ( ~n8535 & n8873 ) ;
  assign n8888 = ~n2296 & n7097 ;
  assign n8885 = n2483 | n6530 ;
  assign n8886 = n2392 | n6983 ;
  assign n8887 = n8885 &  n8886 ;
  assign n8889 = ( n2296 & n8888 ) | ( n2296 & n8887 ) | ( n8888 & n8887 ) ;
  assign n8890 = ( n6532 & ~n5500 ) | ( n6532 & n8889 ) | ( ~n5500 & n8889 ) ;
  assign n8891 = ~n6532 & n8890 ;
  assign n8892 = ( x14 & ~n8889 ) | ( x14 & n8891 ) | ( ~n8889 & n8891 ) ;
  assign n8893 = ( n8889 & ~x14 ) | ( n8889 & n8891 ) | ( ~x14 & n8891 ) ;
  assign n8894 = ( n8892 & ~n8891 ) | ( n8892 & n8893 ) | ( ~n8891 & n8893 ) ;
  assign n8895 = ( n8538 & ~n8548 ) | ( n8538 & n8727 ) | ( ~n8548 & n8727 ) ;
  assign n8896 = ( n8548 & ~n8728 ) | ( n8548 & n8895 ) | ( ~n8728 & n8895 ) ;
  assign n8900 = ~n2392 & n7097 ;
  assign n8897 = n2569 | n6530 ;
  assign n8898 = n2483 | n6983 ;
  assign n8899 = n8897 &  n8898 ;
  assign n8901 = ( n2392 & n8900 ) | ( n2392 & n8899 ) | ( n8900 & n8899 ) ;
  assign n8902 = ( n6532 & ~n6212 ) | ( n6532 & n8901 ) | ( ~n6212 & n8901 ) ;
  assign n8903 = ~n6532 & n8902 ;
  assign n8904 = ( x14 & ~n8901 ) | ( x14 & n8903 ) | ( ~n8901 & n8903 ) ;
  assign n8905 = ( n8901 & ~x14 ) | ( n8901 & n8903 ) | ( ~x14 & n8903 ) ;
  assign n8906 = ( n8904 & ~n8903 ) | ( n8904 & n8905 ) | ( ~n8903 & n8905 ) ;
  assign n8907 = ( n8551 & ~n8561 ) | ( n8551 & n8726 ) | ( ~n8561 & n8726 ) ;
  assign n8908 = ( n8561 & ~n8727 ) | ( n8561 & n8907 ) | ( ~n8727 & n8907 ) ;
  assign n8915 = ~n2665 & n6530 ;
  assign n8912 = n2483 | n7097 ;
  assign n8913 = n2569 | n6983 ;
  assign n8914 = n8912 &  n8913 ;
  assign n8916 = ( n2665 & n8915 ) | ( n2665 & n8914 ) | ( n8915 & n8914 ) ;
  assign n8917 = ( n6532 & ~n6465 ) | ( n6532 & n8916 ) | ( ~n6465 & n8916 ) ;
  assign n8918 = ~n6532 & n8917 ;
  assign n8919 = ( x14 & ~n8916 ) | ( x14 & n8918 ) | ( ~n8916 & n8918 ) ;
  assign n8920 = ( n8916 & ~x14 ) | ( n8916 & n8918 ) | ( ~x14 & n8918 ) ;
  assign n8921 = ( n8919 & ~n8918 ) | ( n8919 & n8920 ) | ( ~n8918 & n8920 ) ;
  assign n8909 = ( n8573 & ~n8571 ) | ( n8573 & n8725 ) | ( ~n8571 & n8725 ) ;
  assign n8910 = ( n8571 & ~n8725 ) | ( n8571 & n8573 ) | ( ~n8725 & n8573 ) ;
  assign n8911 = ( n8909 & ~n8573 ) | ( n8909 & n8910 ) | ( ~n8573 & n8910 ) ;
  assign n8922 = ( n8585 & ~n8583 ) | ( n8585 & n8724 ) | ( ~n8583 & n8724 ) ;
  assign n8923 = ( n8583 & ~n8724 ) | ( n8583 & n8585 ) | ( ~n8724 & n8585 ) ;
  assign n8924 = ( n8922 & ~n8585 ) | ( n8922 & n8923 ) | ( ~n8585 & n8923 ) ;
  assign n8928 = ~n2751 & n6530 ;
  assign n8925 = n2569 | n7097 ;
  assign n8926 = n2665 | n6983 ;
  assign n8927 = n8925 &  n8926 ;
  assign n8929 = ( n2751 & n8928 ) | ( n2751 & n8927 ) | ( n8928 & n8927 ) ;
  assign n8930 = ( n6532 & ~n5705 ) | ( n6532 & n8929 ) | ( ~n5705 & n8929 ) ;
  assign n8931 = ~n6532 & n8930 ;
  assign n8932 = ( x14 & ~n8929 ) | ( x14 & n8931 ) | ( ~n8929 & n8931 ) ;
  assign n8933 = ( n8929 & ~x14 ) | ( n8929 & n8931 ) | ( ~x14 & n8931 ) ;
  assign n8934 = ( n8932 & ~n8931 ) | ( n8932 & n8933 ) | ( ~n8931 & n8933 ) ;
  assign n8935 = ( n8597 & ~n8595 ) | ( n8597 & n8723 ) | ( ~n8595 & n8723 ) ;
  assign n8936 = ( n8595 & ~n8723 ) | ( n8595 & n8597 ) | ( ~n8723 & n8597 ) ;
  assign n8937 = ( n8935 & ~n8597 ) | ( n8935 & n8936 ) | ( ~n8597 & n8936 ) ;
  assign n8941 = ~n2751 & n6983 ;
  assign n8938 = n2665 | n7097 ;
  assign n8939 = n2783 | n6530 ;
  assign n8940 = n8938 &  n8939 ;
  assign n8942 = ( n2751 & n8941 ) | ( n2751 & n8940 ) | ( n8941 & n8940 ) ;
  assign n8943 = ( n6532 & ~n6119 ) | ( n6532 & n8942 ) | ( ~n6119 & n8942 ) ;
  assign n8944 = ~n6532 & n8943 ;
  assign n8945 = ( x14 & ~n8942 ) | ( x14 & n8944 ) | ( ~n8942 & n8944 ) ;
  assign n8946 = ( n8942 & ~x14 ) | ( n8942 & n8944 ) | ( ~x14 & n8944 ) ;
  assign n8947 = ( n8945 & ~n8944 ) | ( n8945 & n8946 ) | ( ~n8944 & n8946 ) ;
  assign n8948 = n2751 | n7097 ;
  assign n8949 = n2783 | n6983 ;
  assign n8950 = n8948 &  n8949 ;
  assign n8951 = n2910 &  n6530 ;
  assign n8952 = ( n8950 & ~n2910 ) | ( n8950 & n8951 ) | ( ~n2910 & n8951 ) ;
  assign n8953 = ( n6532 & ~n6226 ) | ( n6532 & n8952 ) | ( ~n6226 & n8952 ) ;
  assign n8954 = ~n6532 & n8953 ;
  assign n8955 = ( x14 & ~n8952 ) | ( x14 & n8954 ) | ( ~n8952 & n8954 ) ;
  assign n8956 = ( n8952 & ~x14 ) | ( n8952 & n8954 ) | ( ~x14 & n8954 ) ;
  assign n8957 = ( n8955 & ~n8954 ) | ( n8955 & n8956 ) | ( ~n8954 & n8956 ) ;
  assign n8958 = ( n8600 & ~n8722 ) | ( n8600 & n8610 ) | ( ~n8722 & n8610 ) ;
  assign n8959 = ( n8723 & ~n8610 ) | ( n8723 & n8958 ) | ( ~n8610 & n8958 ) ;
  assign n8960 = n2783 | n7097 ;
  assign n8961 = n2839 | n6530 ;
  assign n8962 = n8960 &  n8961 ;
  assign n8963 = n2910 &  n6983 ;
  assign n8964 = ( n8962 & ~n2910 ) | ( n8962 & n8963 ) | ( ~n2910 & n8963 ) ;
  assign n8965 = ( n6104 & ~n6532 ) | ( n6104 & 1'b0 ) | ( ~n6532 & 1'b0 ) ;
  assign n8966 = ( n8964 & ~n8965 ) | ( n8964 & 1'b0 ) | ( ~n8965 & 1'b0 ) ;
  assign n8967 = x14 &  n8966 ;
  assign n8968 = x14 | n8966 ;
  assign n8969 = ~n8967 & n8968 ;
  assign n8970 = ( n8613 & ~n8623 ) | ( n8613 & n8721 ) | ( ~n8623 & n8721 ) ;
  assign n8971 = ( n8623 & ~n8722 ) | ( n8623 & n8970 ) | ( ~n8722 & n8970 ) ;
  assign n8972 = n2995 | n6530 ;
  assign n8973 = n2839 | n6983 ;
  assign n8974 = n8972 &  n8973 ;
  assign n8975 = n2910 &  n7097 ;
  assign n8976 = ( n8974 & ~n2910 ) | ( n8974 & n8975 ) | ( ~n2910 & n8975 ) ;
  assign n8977 = ( n6330 & n6532 ) | ( n6330 & n8976 ) | ( n6532 & n8976 ) ;
  assign n8978 = ~n6532 & n8977 ;
  assign n8979 = ( x14 & ~n8976 ) | ( x14 & n8978 ) | ( ~n8976 & n8978 ) ;
  assign n8980 = ( n8976 & ~x14 ) | ( n8976 & n8978 ) | ( ~x14 & n8978 ) ;
  assign n8981 = ( n8979 & ~n8978 ) | ( n8979 & n8980 ) | ( ~n8978 & n8980 ) ;
  assign n8982 = ( n8626 & ~n8636 ) | ( n8626 & n8720 ) | ( ~n8636 & n8720 ) ;
  assign n8983 = ( n8636 & ~n8721 ) | ( n8636 & n8982 ) | ( ~n8721 & n8982 ) ;
  assign n8990 = ~n2839 & n7097 ;
  assign n8987 = n3030 | n6530 ;
  assign n8988 = n2995 | n6983 ;
  assign n8989 = n8987 &  n8988 ;
  assign n8991 = ( n2839 & n8990 ) | ( n2839 & n8989 ) | ( n8990 & n8989 ) ;
  assign n8992 = ( n7324 & ~n6532 ) | ( n7324 & n8991 ) | ( ~n6532 & n8991 ) ;
  assign n8993 = ~n7324 & n8992 ;
  assign n8994 = ( x14 & ~n8991 ) | ( x14 & n8993 ) | ( ~n8991 & n8993 ) ;
  assign n8995 = ( n8991 & ~x14 ) | ( n8991 & n8993 ) | ( ~x14 & n8993 ) ;
  assign n8996 = ( n8994 & ~n8993 ) | ( n8994 & n8995 ) | ( ~n8993 & n8995 ) ;
  assign n8984 = ( n8648 & ~n8646 ) | ( n8648 & n8719 ) | ( ~n8646 & n8719 ) ;
  assign n8985 = ( n8646 & ~n8719 ) | ( n8646 & n8648 ) | ( ~n8719 & n8648 ) ;
  assign n8986 = ( n8984 & ~n8648 ) | ( n8984 & n8985 ) | ( ~n8648 & n8985 ) ;
  assign n8997 = ( n8661 & ~n8651 ) | ( n8661 & n8718 ) | ( ~n8651 & n8718 ) ;
  assign n8998 = ( n8651 & ~n8718 ) | ( n8651 & n8661 ) | ( ~n8718 & n8661 ) ;
  assign n8999 = ( n8997 & ~n8661 ) | ( n8997 & n8998 ) | ( ~n8661 & n8998 ) ;
  assign n9000 = n3106 | n6530 ;
  assign n9001 = n3030 | n6983 ;
  assign n9002 = n9000 &  n9001 ;
  assign n9003 = ~n2995 & n7097 ;
  assign n9004 = ( n2995 & n9002 ) | ( n2995 & n9003 ) | ( n9002 & n9003 ) ;
  assign n9005 = ( n7339 & ~n6532 ) | ( n7339 & n9004 ) | ( ~n6532 & n9004 ) ;
  assign n9006 = ~n7339 & n9005 ;
  assign n9007 = ( x14 & ~n9004 ) | ( x14 & n9006 ) | ( ~n9004 & n9006 ) ;
  assign n9008 = ( n9004 & ~x14 ) | ( n9004 & n9006 ) | ( ~x14 & n9006 ) ;
  assign n9009 = ( n9007 & ~n9006 ) | ( n9007 & n9008 ) | ( ~n9006 & n9008 ) ;
  assign n9010 = ( n8671 & ~n8717 ) | ( n8671 & n8674 ) | ( ~n8717 & n8674 ) ;
  assign n9011 = ( n8674 & ~n8671 ) | ( n8674 & n8717 ) | ( ~n8671 & n8717 ) ;
  assign n9012 = ( n9010 & ~n8674 ) | ( n9010 & n9011 ) | ( ~n8674 & n9011 ) ;
  assign n9016 = ~n3030 & n7097 ;
  assign n9013 = n3197 | n6530 ;
  assign n9014 = n3106 | n6983 ;
  assign n9015 = n9013 &  n9014 ;
  assign n9017 = ( n3030 & n9016 ) | ( n3030 & n9015 ) | ( n9016 & n9015 ) ;
  assign n9018 = ( n6532 & ~n6314 ) | ( n6532 & n9017 ) | ( ~n6314 & n9017 ) ;
  assign n9019 = ~n6532 & n9018 ;
  assign n9020 = ( x14 & ~n9017 ) | ( x14 & n9019 ) | ( ~n9017 & n9019 ) ;
  assign n9021 = ( n9017 & ~x14 ) | ( n9017 & n9019 ) | ( ~x14 & n9019 ) ;
  assign n9022 = ( n9020 & ~n9019 ) | ( n9020 & n9021 ) | ( ~n9019 & n9021 ) ;
  assign n9023 = n3106 | n7097 ;
  assign n9024 = n3197 | n6983 ;
  assign n9025 = n9023 &  n9024 ;
  assign n9026 = n3266 &  n6530 ;
  assign n9027 = ( n9025 & ~n3266 ) | ( n9025 & n9026 ) | ( ~n3266 & n9026 ) ;
  assign n9028 = ( n7363 & ~n6532 ) | ( n7363 & n9027 ) | ( ~n6532 & n9027 ) ;
  assign n9029 = ~n7363 & n9028 ;
  assign n9030 = ( x14 & ~n9027 ) | ( x14 & n9029 ) | ( ~n9027 & n9029 ) ;
  assign n9031 = ( n9027 & ~x14 ) | ( n9027 & n9029 ) | ( ~x14 & n9029 ) ;
  assign n9032 = ( n9030 & ~n9029 ) | ( n9030 & n9031 ) | ( ~n9029 & n9031 ) ;
  assign n9033 = ( n8688 & ~n8678 ) | ( n8688 & n8716 ) | ( ~n8678 & n8716 ) ;
  assign n9034 = ( n8717 & ~n8688 ) | ( n8717 & n9033 ) | ( ~n8688 & n9033 ) ;
  assign n9036 = ( n8343 & n8705 ) | ( n8343 & n8715 ) | ( n8705 & n8715 ) ;
  assign n9035 = ( n8343 & ~n8705 ) | ( n8343 & n8715 ) | ( ~n8705 & n8715 ) ;
  assign n9037 = ( n8705 & ~n9036 ) | ( n8705 & n9035 ) | ( ~n9036 & n9035 ) ;
  assign n9038 = n3197 | n7097 ;
  assign n9039 = n3325 | n6530 ;
  assign n9040 = n9038 &  n9039 ;
  assign n9041 = n3266 &  n6983 ;
  assign n9042 = ( n9040 & ~n3266 ) | ( n9040 & n9041 ) | ( ~n3266 & n9041 ) ;
  assign n9043 = ( n6532 & ~n9042 ) | ( n6532 & n7377 ) | ( ~n9042 & n7377 ) ;
  assign n9044 = ( n7377 & ~n9043 ) | ( n7377 & 1'b0 ) | ( ~n9043 & 1'b0 ) ;
  assign n9045 = ( x14 & ~n9042 ) | ( x14 & n9044 ) | ( ~n9042 & n9044 ) ;
  assign n9046 = ( n9042 & ~x14 ) | ( n9042 & n9044 ) | ( ~x14 & n9044 ) ;
  assign n9047 = ( n9045 & ~n9044 ) | ( n9045 & n9046 ) | ( ~n9044 & n9046 ) ;
  assign n9048 = n3361 | n6530 ;
  assign n9049 = n3325 | n6983 ;
  assign n9050 = n9048 &  n9049 ;
  assign n9051 = n3266 &  n7097 ;
  assign n9052 = ( n9050 & ~n3266 ) | ( n9050 & n9051 ) | ( ~n3266 & n9051 ) ;
  assign n9053 = ( n6532 & ~n9052 ) | ( n6532 & n7391 ) | ( ~n9052 & n7391 ) ;
  assign n9054 = ( n7391 & ~n9053 ) | ( n7391 & 1'b0 ) | ( ~n9053 & 1'b0 ) ;
  assign n9055 = ( x14 & ~n9052 ) | ( x14 & n9054 ) | ( ~n9052 & n9054 ) ;
  assign n9056 = ( n9052 & ~x14 ) | ( n9052 & n9054 ) | ( ~x14 & n9054 ) ;
  assign n9057 = ( n9055 & ~n9054 ) | ( n9055 & n9056 ) | ( ~n9054 & n9056 ) ;
  assign n8696 = ( x17 & ~n8695 ) | ( x17 & 1'b0 ) | ( ~n8695 & 1'b0 ) ;
  assign n9059 = ( x17 & n8696 ) | ( x17 & n8703 ) | ( n8696 & n8703 ) ;
  assign n9058 = ( x17 & ~n8696 ) | ( x17 & n8703 ) | ( ~n8696 & n8703 ) ;
  assign n9060 = ( n8696 & ~n9059 ) | ( n8696 & n9058 ) | ( ~n9059 & n9058 ) ;
  assign n9061 = x17 &  n8694 ;
  assign n9062 = n8693 &  n9061 ;
  assign n9063 = n8693 | n9061 ;
  assign n9064 = ~n9062 & n9063 ;
  assign n9095 = ~n3460 & n6983 ;
  assign n9092 = n3361 | n7097 ;
  assign n9093 = n3601 | n6530 ;
  assign n9094 = n9092 &  n9093 ;
  assign n9096 = ( n3460 & n9095 ) | ( n3460 & n9094 ) | ( n9095 & n9094 ) ;
  assign n9097 = ( n6895 & ~n6532 ) | ( n6895 & n9096 ) | ( ~n6532 & n9096 ) ;
  assign n9098 = ~n6895 & n9097 ;
  assign n9099 = ( x14 & ~n9096 ) | ( x14 & n9098 ) | ( ~n9096 & n9098 ) ;
  assign n9100 = ( n9096 & ~x14 ) | ( n9096 & n9098 ) | ( ~x14 & n9098 ) ;
  assign n9101 = ( n9099 & ~n9098 ) | ( n9099 & n9100 ) | ( ~n9098 & n9100 ) ;
  assign n9088 = ~n6532 & n6886 ;
  assign n9086 = ~n3460 & n7097 ;
  assign n9083 = n3547 | n6530 ;
  assign n9084 = n3601 | n6983 ;
  assign n9085 = n9083 &  n9084 ;
  assign n9087 = ( n3460 & n9086 ) | ( n3460 & n9085 ) | ( n9086 & n9085 ) ;
  assign n9089 = ( n6532 & n9088 ) | ( n6532 & n9087 ) | ( n9088 & n9087 ) ;
  assign n9078 = n7412 | n6532 ;
  assign n9075 = n3547 | n6983 ;
  assign n9076 = n3601 | n7097 ;
  assign n9077 = n9075 &  n9076 ;
  assign n9079 = ( n6532 & ~n9078 ) | ( n6532 & n9077 ) | ( ~n9078 & n9077 ) ;
  assign n9080 = ~n3547 & n6525 ;
  assign n9081 = ( x14 & ~n9079 ) | ( x14 & n9080 ) | ( ~n9079 & n9080 ) ;
  assign n9090 = ( x14 & ~n9089 ) | ( x14 & n9081 ) | ( ~n9089 & n9081 ) ;
  assign n9091 = ( x14 & ~n9090 ) | ( x14 & 1'b0 ) | ( ~n9090 & 1'b0 ) ;
  assign n9102 = ( n8694 & ~n9101 ) | ( n8694 & n9091 ) | ( ~n9101 & n9091 ) ;
  assign n9068 = ~n3460 & n6530 ;
  assign n9065 = n3325 | n7097 ;
  assign n9066 = n3361 | n6983 ;
  assign n9067 = n9065 &  n9066 ;
  assign n9069 = ( n3460 & n9068 ) | ( n3460 & n9067 ) | ( n9068 & n9067 ) ;
  assign n9070 = ( n7405 & ~n6532 ) | ( n7405 & n9069 ) | ( ~n6532 & n9069 ) ;
  assign n9071 = ~n7405 & n9070 ;
  assign n9072 = ( x14 & ~n9069 ) | ( x14 & n9071 ) | ( ~n9069 & n9071 ) ;
  assign n9073 = ( n9069 & ~x14 ) | ( n9069 & n9071 ) | ( ~x14 & n9071 ) ;
  assign n9074 = ( n9072 & ~n9071 ) | ( n9072 & n9073 ) | ( ~n9071 & n9073 ) ;
  assign n9103 = ( n9064 & ~n9102 ) | ( n9064 & n9074 ) | ( ~n9102 & n9074 ) ;
  assign n9104 = ( n9057 & n9060 ) | ( n9057 & n9103 ) | ( n9060 & n9103 ) ;
  assign n9105 = ( n9037 & n9047 ) | ( n9037 & n9104 ) | ( n9047 & n9104 ) ;
  assign n9106 = ( n9032 & ~n9034 ) | ( n9032 & n9105 ) | ( ~n9034 & n9105 ) ;
  assign n9107 = ( n9012 & n9022 ) | ( n9012 & n9106 ) | ( n9022 & n9106 ) ;
  assign n9108 = ( n8999 & n9009 ) | ( n8999 & n9107 ) | ( n9009 & n9107 ) ;
  assign n9109 = ( n8996 & ~n8986 ) | ( n8996 & n9108 ) | ( ~n8986 & n9108 ) ;
  assign n9110 = ( n8981 & n8983 ) | ( n8981 & n9109 ) | ( n8983 & n9109 ) ;
  assign n9111 = ( n8969 & n8971 ) | ( n8969 & n9110 ) | ( n8971 & n9110 ) ;
  assign n9112 = ( n8957 & ~n8959 ) | ( n8957 & n9111 ) | ( ~n8959 & n9111 ) ;
  assign n9113 = ( n8937 & n8947 ) | ( n8937 & n9112 ) | ( n8947 & n9112 ) ;
  assign n9114 = ( n8924 & n8934 ) | ( n8924 & n9113 ) | ( n8934 & n9113 ) ;
  assign n9115 = ( n8921 & ~n8911 ) | ( n8921 & n9114 ) | ( ~n8911 & n9114 ) ;
  assign n9116 = ( n8906 & n8908 ) | ( n8906 & n9115 ) | ( n8908 & n9115 ) ;
  assign n9117 = ( n8894 & n8896 ) | ( n8894 & n9116 ) | ( n8896 & n9116 ) ;
  assign n9118 = ( n8884 & ~n8874 ) | ( n8884 & n9117 ) | ( ~n8874 & n9117 ) ;
  assign n9119 = ( n8871 & ~n8861 ) | ( n8871 & n9118 ) | ( ~n8861 & n9118 ) ;
  assign n9120 = ( n8848 & n8858 ) | ( n8848 & n9119 ) | ( n8858 & n9119 ) ;
  assign n9121 = ( n8835 & n8845 ) | ( n8835 & n9120 ) | ( n8845 & n9120 ) ;
  assign n9122 = ( n8832 & ~n8822 ) | ( n8832 & n9121 ) | ( ~n8822 & n9121 ) ;
  assign n9123 = ( n8809 & n8819 ) | ( n8809 & n9122 ) | ( n8819 & n9122 ) ;
  assign n9124 = ( n8796 & n8806 ) | ( n8796 & n9123 ) | ( n8806 & n9123 ) ;
  assign n9125 = n8747 &  n8749 ;
  assign n9126 = ( n8750 & ~n9125 ) | ( n8750 & 1'b0 ) | ( ~n9125 & 1'b0 ) ;
  assign n9127 = n1483 &  n7253 ;
  assign n9128 = n1378 | n7518 ;
  assign n9129 = ~n9127 & n9128 ;
  assign n9130 = n1267 &  n7783 ;
  assign n9131 = ( n9129 & ~n1267 ) | ( n9129 & n9130 ) | ( ~n1267 & n9130 ) ;
  assign n9132 = ( n4422 & n7255 ) | ( n4422 & n9131 ) | ( n7255 & n9131 ) ;
  assign n9133 = ~n7255 & n9132 ;
  assign n9134 = ( x11 & ~n9131 ) | ( x11 & n9133 ) | ( ~n9131 & n9133 ) ;
  assign n9135 = ( n9131 & ~x11 ) | ( n9131 & n9133 ) | ( ~x11 & n9133 ) ;
  assign n9136 = ( n9134 & ~n9133 ) | ( n9134 & n9135 ) | ( ~n9133 & n9135 ) ;
  assign n9137 = ( n9124 & ~n9126 ) | ( n9124 & n9136 ) | ( ~n9126 & n9136 ) ;
  assign n8791 = ( n8448 & n8751 ) | ( n8448 & n8761 ) | ( n8751 & n8761 ) ;
  assign n8792 = ( n8448 & ~n8751 ) | ( n8448 & n8761 ) | ( ~n8751 & n8761 ) ;
  assign n8793 = ( n8751 & ~n8791 ) | ( n8751 & n8792 ) | ( ~n8791 & n8792 ) ;
  assign n9141 = ~n946 & n8429 ;
  assign n9138 = n863 | n8764 ;
  assign n9139 = ~n1043 & n8105 ;
  assign n9140 = ( n9138 & ~n9139 ) | ( n9138 & 1'b0 ) | ( ~n9139 & 1'b0 ) ;
  assign n9142 = ( n946 & n9141 ) | ( n946 & n9140 ) | ( n9141 & n9140 ) ;
  assign n9143 = ( n8107 & ~n3914 ) | ( n8107 & n9142 ) | ( ~n3914 & n9142 ) ;
  assign n9144 = ~n8107 & n9143 ;
  assign n9145 = ( x8 & ~n9142 ) | ( x8 & n9144 ) | ( ~n9142 & n9144 ) ;
  assign n9146 = ( n9142 & ~x8 ) | ( n9142 & n9144 ) | ( ~x8 & n9144 ) ;
  assign n9147 = ( n9145 & ~n9144 ) | ( n9145 & n9146 ) | ( ~n9144 & n9146 ) ;
  assign n9148 = ( n9137 & ~n8793 ) | ( n9137 & n9147 ) | ( ~n8793 & n9147 ) ;
  assign n9167 = ( n8445 & n8762 ) | ( n8445 & n8773 ) | ( n8762 & n8773 ) ;
  assign n9168 = ( n8445 & ~n8762 ) | ( n8445 & n8773 ) | ( ~n8762 & n8773 ) ;
  assign n9169 = ( n8762 & ~n9167 ) | ( n8762 & n9168 ) | ( ~n9167 & n9168 ) ;
  assign n9149 = ( x4 & ~x5 ) | ( x4 & 1'b0 ) | ( ~x5 & 1'b0 ) ;
  assign n9150 = ~x4 & x5 ;
  assign n9151 = n9149 | n9150 ;
  assign n9152 = ( x2 & ~x3 ) | ( x2 & 1'b0 ) | ( ~x3 & 1'b0 ) ;
  assign n9153 = ~x2 & x3 ;
  assign n9154 = n9152 | n9153 ;
  assign n9159 = ( n9151 & ~n9154 ) | ( n9151 & 1'b0 ) | ( ~n9154 & 1'b0 ) ;
  assign n9156 = ~x3 & x4 ;
  assign n9157 = ( x3 & ~x4 ) | ( x3 & 1'b0 ) | ( ~x4 & 1'b0 ) ;
  assign n9158 = n9156 | n9157 ;
  assign n9160 = ~n9159 |  n9158 ;
  assign n9161 = n599 | n9160 ;
  assign n9155 = ~n9151 | ~n9154 ;
  assign n9162 = ~n3637 & n9155 ;
  assign n9163 = ( n3637 & n9161 ) | ( n3637 & n9162 ) | ( n9161 & n9162 ) ;
  assign n9164 = x5 &  n9163 ;
  assign n9165 = x5 | n9163 ;
  assign n9166 = ~n9164 & n9165 ;
  assign n9170 = ( n9148 & ~n9169 ) | ( n9148 & n9166 ) | ( ~n9169 & n9166 ) ;
  assign n9171 = ( n8784 & ~n8774 ) | ( n8784 & n8786 ) | ( ~n8774 & n8786 ) ;
  assign n9172 = ( n8787 & ~n8784 ) | ( n8787 & n9171 ) | ( ~n8784 & n9171 ) ;
  assign n9175 = n1378 | n7783 ;
  assign n9176 = ~n1566 & n7253 ;
  assign n9177 = ( n9175 & ~n9176 ) | ( n9175 & 1'b0 ) | ( ~n9176 & 1'b0 ) ;
  assign n9178 = n1483 &  n7518 ;
  assign n9179 = ( n9177 & ~n1483 ) | ( n9177 & n9178 ) | ( ~n1483 & n9178 ) ;
  assign n9180 = ( n5038 & n7255 ) | ( n5038 & n9179 ) | ( n7255 & n9179 ) ;
  assign n9181 = ~n7255 & n9180 ;
  assign n9182 = ( x11 & ~n9179 ) | ( x11 & n9181 ) | ( ~n9179 & n9181 ) ;
  assign n9183 = ( n9179 & ~x11 ) | ( n9179 & n9181 ) | ( ~x11 & n9181 ) ;
  assign n9184 = ( n9182 & ~n9181 ) | ( n9182 & n9183 ) | ( ~n9181 & n9183 ) ;
  assign n9185 = ( n8796 & ~n8806 ) | ( n8796 & n9123 ) | ( ~n8806 & n9123 ) ;
  assign n9186 = ( n8806 & ~n9124 ) | ( n8806 & n9185 ) | ( ~n9124 & n9185 ) ;
  assign n9187 = ~n1671 & n7253 ;
  assign n9188 = n1566 | n7518 ;
  assign n9189 = ~n9187 & n9188 ;
  assign n9190 = n1483 &  n7783 ;
  assign n9191 = ( n9189 & ~n1483 ) | ( n9189 & n9190 ) | ( ~n1483 & n9190 ) ;
  assign n9192 = ( n4274 & n7255 ) | ( n4274 & n9191 ) | ( n7255 & n9191 ) ;
  assign n9193 = ~n7255 & n9192 ;
  assign n9194 = ( x11 & ~n9191 ) | ( x11 & n9193 ) | ( ~n9191 & n9193 ) ;
  assign n9195 = ( n9191 & ~x11 ) | ( n9191 & n9193 ) | ( ~x11 & n9193 ) ;
  assign n9196 = ( n9194 & ~n9193 ) | ( n9194 & n9195 ) | ( ~n9193 & n9195 ) ;
  assign n9197 = ( n8809 & ~n8819 ) | ( n8809 & n9122 ) | ( ~n8819 & n9122 ) ;
  assign n9198 = ( n8819 & ~n9123 ) | ( n8819 & n9197 ) | ( ~n9123 & n9197 ) ;
  assign n9202 = ~n1566 & n7783 ;
  assign n9199 = ~n1748 & n7253 ;
  assign n9200 = n1671 | n7518 ;
  assign n9201 = ~n9199 & n9200 ;
  assign n9203 = ( n1566 & n9202 ) | ( n1566 & n9201 ) | ( n9202 & n9201 ) ;
  assign n9204 = ( n7255 & ~n4597 ) | ( n7255 & n9203 ) | ( ~n4597 & n9203 ) ;
  assign n9205 = ~n7255 & n9204 ;
  assign n9206 = ( x11 & ~n9203 ) | ( x11 & n9205 ) | ( ~n9203 & n9205 ) ;
  assign n9207 = ( n9203 & ~x11 ) | ( n9203 & n9205 ) | ( ~x11 & n9205 ) ;
  assign n9208 = ( n9206 & ~n9205 ) | ( n9206 & n9207 ) | ( ~n9205 & n9207 ) ;
  assign n9209 = ( n8822 & ~n9121 ) | ( n8822 & n8832 ) | ( ~n9121 & n8832 ) ;
  assign n9210 = ( n9122 & ~n8832 ) | ( n9122 & n9209 ) | ( ~n8832 & n9209 ) ;
  assign n9211 = n1875 &  n7253 ;
  assign n9212 = n1671 | n7783 ;
  assign n9213 = n1748 | n7518 ;
  assign n9214 = n9212 &  n9213 ;
  assign n9215 = ( n9211 & ~n7253 ) | ( n9211 & n9214 ) | ( ~n7253 & n9214 ) ;
  assign n9216 = ( n7255 & ~n4580 ) | ( n7255 & n9215 ) | ( ~n4580 & n9215 ) ;
  assign n9217 = ~n7255 & n9216 ;
  assign n9218 = ( x11 & ~n9215 ) | ( x11 & n9217 ) | ( ~n9215 & n9217 ) ;
  assign n9219 = ( n9215 & ~x11 ) | ( n9215 & n9217 ) | ( ~x11 & n9217 ) ;
  assign n9220 = ( n9218 & ~n9217 ) | ( n9218 & n9219 ) | ( ~n9217 & n9219 ) ;
  assign n9221 = ( n8835 & ~n8845 ) | ( n8835 & n9120 ) | ( ~n8845 & n9120 ) ;
  assign n9222 = ( n8845 & ~n9121 ) | ( n8845 & n9221 ) | ( ~n9121 & n9221 ) ;
  assign n9223 = ~n1940 & n7253 ;
  assign n9224 = n1875 | n7518 ;
  assign n9225 = ~n9223 & n9224 ;
  assign n9226 = ~n1748 & n7783 ;
  assign n9227 = ( n1748 & n9225 ) | ( n1748 & n9226 ) | ( n9225 & n9226 ) ;
  assign n9228 = ( n7255 & ~n4743 ) | ( n7255 & n9227 ) | ( ~n4743 & n9227 ) ;
  assign n9229 = ~n7255 & n9228 ;
  assign n9230 = ( x11 & ~n9227 ) | ( x11 & n9229 ) | ( ~n9227 & n9229 ) ;
  assign n9231 = ( n9227 & ~x11 ) | ( n9227 & n9229 ) | ( ~x11 & n9229 ) ;
  assign n9232 = ( n9230 & ~n9229 ) | ( n9230 & n9231 ) | ( ~n9229 & n9231 ) ;
  assign n9233 = ( n8848 & ~n8858 ) | ( n8848 & n9119 ) | ( ~n8858 & n9119 ) ;
  assign n9234 = ( n8858 & ~n9120 ) | ( n8858 & n9233 ) | ( ~n9120 & n9233 ) ;
  assign n9238 = ~n1875 & n7783 ;
  assign n9235 = ~n2022 & n7253 ;
  assign n9236 = n1940 | n7518 ;
  assign n9237 = ~n9235 & n9236 ;
  assign n9239 = ( n1875 & n9238 ) | ( n1875 & n9237 ) | ( n9238 & n9237 ) ;
  assign n9240 = ( n7255 & ~n5381 ) | ( n7255 & n9239 ) | ( ~n5381 & n9239 ) ;
  assign n9241 = ~n7255 & n9240 ;
  assign n9242 = ( x11 & ~n9239 ) | ( x11 & n9241 ) | ( ~n9239 & n9241 ) ;
  assign n9243 = ( n9239 & ~x11 ) | ( n9239 & n9241 ) | ( ~x11 & n9241 ) ;
  assign n9244 = ( n9242 & ~n9241 ) | ( n9242 & n9243 ) | ( ~n9241 & n9243 ) ;
  assign n9245 = ( n8861 & ~n9118 ) | ( n8861 & n8871 ) | ( ~n9118 & n8871 ) ;
  assign n9246 = ( n9119 & ~n8871 ) | ( n9119 & n9245 ) | ( ~n8871 & n9245 ) ;
  assign n9247 = ~n2127 & n7253 ;
  assign n9248 = n2022 | n7518 ;
  assign n9249 = ~n9247 & n9248 ;
  assign n9250 = ~n1940 & n7783 ;
  assign n9251 = ( n1940 & n9249 ) | ( n1940 & n9250 ) | ( n9249 & n9250 ) ;
  assign n9252 = n5799 | n7255 ;
  assign n9253 = n9251 &  n9252 ;
  assign n9254 = x11 | n9253 ;
  assign n9255 = x11 &  n9253 ;
  assign n9256 = ( n9254 & ~n9255 ) | ( n9254 & 1'b0 ) | ( ~n9255 & 1'b0 ) ;
  assign n9257 = ( n8874 & ~n9117 ) | ( n8874 & n8884 ) | ( ~n9117 & n8884 ) ;
  assign n9258 = ( n9118 & ~n8884 ) | ( n9118 & n9257 ) | ( ~n8884 & n9257 ) ;
  assign n9259 = ( n8894 & ~n9116 ) | ( n8894 & n8896 ) | ( ~n9116 & n8896 ) ;
  assign n9260 = ( n8896 & ~n8894 ) | ( n8896 & n9116 ) | ( ~n8894 & n9116 ) ;
  assign n9261 = ( n9259 & ~n8896 ) | ( n9259 & n9260 ) | ( ~n8896 & n9260 ) ;
  assign n9262 = ~n2178 & n7253 ;
  assign n9263 = n2127 | n7518 ;
  assign n9264 = ~n9262 & n9263 ;
  assign n9265 = ~n2022 & n7783 ;
  assign n9266 = ( n2022 & n9264 ) | ( n2022 & n9265 ) | ( n9264 & n9265 ) ;
  assign n9267 = ( n4931 & ~n3621 ) | ( n4931 & n7255 ) | ( ~n3621 & n7255 ) ;
  assign n9268 = ( n4933 & n9266 ) | ( n4933 & n9267 ) | ( n9266 & n9267 ) ;
  assign n9269 = x11 &  n9268 ;
  assign n9270 = x11 | n9268 ;
  assign n9271 = ~n9269 & n9270 ;
  assign n9272 = ( n8908 & ~n8906 ) | ( n8908 & n9115 ) | ( ~n8906 & n9115 ) ;
  assign n9273 = ( n8906 & ~n9115 ) | ( n8906 & n8908 ) | ( ~n9115 & n8908 ) ;
  assign n9274 = ( n9272 & ~n8908 ) | ( n9272 & n9273 ) | ( ~n8908 & n9273 ) ;
  assign n9275 = n2296 &  n7253 ;
  assign n9276 = n2127 | n7783 ;
  assign n9277 = n2178 | n7518 ;
  assign n9278 = n9276 &  n9277 ;
  assign n9279 = ( n9275 & ~n7253 ) | ( n9275 & n9278 ) | ( ~n7253 & n9278 ) ;
  assign n9280 = ( n5280 & ~n3620 ) | ( n5280 & n7255 ) | ( ~n3620 & n7255 ) ;
  assign n9281 = ( n5282 & n9279 ) | ( n5282 & n9280 ) | ( n9279 & n9280 ) ;
  assign n9282 = x11 &  n9281 ;
  assign n9283 = x11 | n9281 ;
  assign n9284 = ~n9282 & n9283 ;
  assign n9288 = ~n2178 & n7783 ;
  assign n9285 = ~n2392 & n7253 ;
  assign n9286 = n2296 | n7518 ;
  assign n9287 = ~n9285 & n9286 ;
  assign n9289 = ( n2178 & n9288 ) | ( n2178 & n9287 ) | ( n9288 & n9287 ) ;
  assign n9290 = n5269 | n7255 ;
  assign n9291 = n9289 &  n9290 ;
  assign n9292 = x11 | n9291 ;
  assign n9293 = x11 &  n9291 ;
  assign n9294 = ( n9292 & ~n9293 ) | ( n9292 & 1'b0 ) | ( ~n9293 & 1'b0 ) ;
  assign n9295 = ( n8911 & ~n9114 ) | ( n8911 & n8921 ) | ( ~n9114 & n8921 ) ;
  assign n9296 = ( n9115 & ~n8921 ) | ( n9115 & n9295 ) | ( ~n8921 & n9295 ) ;
  assign n9300 = ~n2296 & n7783 ;
  assign n9297 = ~n2483 & n7253 ;
  assign n9298 = n2392 | n7518 ;
  assign n9299 = ~n9297 & n9298 ;
  assign n9301 = ( n2296 & n9300 ) | ( n2296 & n9299 ) | ( n9300 & n9299 ) ;
  assign n9302 = n5500 | n7255 ;
  assign n9303 = n9301 &  n9302 ;
  assign n9304 = x11 | n9303 ;
  assign n9305 = x11 &  n9303 ;
  assign n9306 = ( n9304 & ~n9305 ) | ( n9304 & 1'b0 ) | ( ~n9305 & 1'b0 ) ;
  assign n9307 = ( n8924 & ~n8934 ) | ( n8924 & n9113 ) | ( ~n8934 & n9113 ) ;
  assign n9308 = ( n8934 & ~n9114 ) | ( n8934 & n9307 ) | ( ~n9114 & n9307 ) ;
  assign n9312 = ~n2392 & n7783 ;
  assign n9309 = ~n2569 & n7253 ;
  assign n9310 = n2483 | n7518 ;
  assign n9311 = ~n9309 & n9310 ;
  assign n9313 = ( n2392 & n9312 ) | ( n2392 & n9311 ) | ( n9312 & n9311 ) ;
  assign n9314 = n6212 | n7255 ;
  assign n9315 = n9313 &  n9314 ;
  assign n9316 = x11 | n9315 ;
  assign n9317 = x11 &  n9315 ;
  assign n9318 = ( n9316 & ~n9317 ) | ( n9316 & 1'b0 ) | ( ~n9317 & 1'b0 ) ;
  assign n9319 = ( n8937 & ~n8947 ) | ( n8937 & n9112 ) | ( ~n8947 & n9112 ) ;
  assign n9320 = ( n8947 & ~n9113 ) | ( n8947 & n9319 ) | ( ~n9113 & n9319 ) ;
  assign n9324 = n2665 &  n7253 ;
  assign n9325 = n2483 | n7783 ;
  assign n9326 = n2569 | n7518 ;
  assign n9327 = n9325 &  n9326 ;
  assign n9328 = ( n9324 & ~n7253 ) | ( n9324 & n9327 ) | ( ~n7253 & n9327 ) ;
  assign n9329 = ( n5886 & ~n3616 ) | ( n5886 & n7255 ) | ( ~n3616 & n7255 ) ;
  assign n9330 = ( n5887 & n9328 ) | ( n5887 & n9329 ) | ( n9328 & n9329 ) ;
  assign n9331 = x11 &  n9330 ;
  assign n9332 = x11 | n9330 ;
  assign n9333 = ~n9331 & n9332 ;
  assign n9321 = ( n8959 & ~n8957 ) | ( n8959 & n9111 ) | ( ~n8957 & n9111 ) ;
  assign n9322 = ( n8957 & ~n9111 ) | ( n8957 & n8959 ) | ( ~n9111 & n8959 ) ;
  assign n9323 = ( n9321 & ~n8959 ) | ( n9321 & n9322 ) | ( ~n8959 & n9322 ) ;
  assign n9334 = ( n8971 & ~n8969 ) | ( n8971 & n9110 ) | ( ~n8969 & n9110 ) ;
  assign n9335 = ( n8969 & ~n9110 ) | ( n8969 & n8971 ) | ( ~n9110 & n8971 ) ;
  assign n9336 = ( n9334 & ~n8971 ) | ( n9334 & n9335 ) | ( ~n8971 & n9335 ) ;
  assign n9337 = n2751 &  n7253 ;
  assign n9338 = n2569 | n7783 ;
  assign n9339 = n2665 | n7518 ;
  assign n9340 = n9338 &  n9339 ;
  assign n9341 = ( n9337 & ~n7253 ) | ( n9337 & n9340 ) | ( ~n7253 & n9340 ) ;
  assign n9342 = ( n5702 & ~n3615 ) | ( n5702 & n7255 ) | ( ~n3615 & n7255 ) ;
  assign n9343 = ( n5704 & n9341 ) | ( n5704 & n9342 ) | ( n9341 & n9342 ) ;
  assign n9344 = x11 &  n9343 ;
  assign n9345 = x11 | n9343 ;
  assign n9346 = ~n9344 & n9345 ;
  assign n9347 = ( n8983 & ~n8981 ) | ( n8983 & n9109 ) | ( ~n8981 & n9109 ) ;
  assign n9348 = ( n8981 & ~n9109 ) | ( n8981 & n8983 ) | ( ~n9109 & n8983 ) ;
  assign n9349 = ( n9347 & ~n8983 ) | ( n9347 & n9348 ) | ( ~n8983 & n9348 ) ;
  assign n9353 = ~n2751 & n7518 ;
  assign n9350 = n2665 | n7783 ;
  assign n9351 = ~n2783 & n7253 ;
  assign n9352 = ( n9350 & ~n9351 ) | ( n9350 & 1'b0 ) | ( ~n9351 & 1'b0 ) ;
  assign n9354 = ( n2751 & n9353 ) | ( n2751 & n9352 ) | ( n9353 & n9352 ) ;
  assign n9355 = ( n6116 & ~n3614 ) | ( n6116 & n7255 ) | ( ~n3614 & n7255 ) ;
  assign n9356 = ( n6118 & n9354 ) | ( n6118 & n9355 ) | ( n9354 & n9355 ) ;
  assign n9357 = x11 &  n9356 ;
  assign n9358 = x11 | n9356 ;
  assign n9359 = ~n9357 & n9358 ;
  assign n9363 = ~n7253 & n2910 ;
  assign n9360 = n2751 | n7783 ;
  assign n9361 = n2783 | n7518 ;
  assign n9362 = n9360 &  n9361 ;
  assign n9364 = ( n9363 & ~n2910 ) | ( n9363 & n9362 ) | ( ~n2910 & n9362 ) ;
  assign n9365 = n6226 | n7255 ;
  assign n9366 = n9364 &  n9365 ;
  assign n9367 = x11 | n9366 ;
  assign n9368 = x11 &  n9366 ;
  assign n9369 = ( n9367 & ~n9368 ) | ( n9367 & 1'b0 ) | ( ~n9368 & 1'b0 ) ;
  assign n9370 = ( n8986 & ~n9108 ) | ( n8986 & n8996 ) | ( ~n9108 & n8996 ) ;
  assign n9371 = ( n9109 & ~n8996 ) | ( n9109 & n9370 ) | ( ~n8996 & n9370 ) ;
  assign n9372 = n2783 | n7783 ;
  assign n9373 = ~n2839 & n7253 ;
  assign n9374 = ( n9372 & ~n9373 ) | ( n9372 & 1'b0 ) | ( ~n9373 & 1'b0 ) ;
  assign n9375 = n2910 &  n7518 ;
  assign n9376 = ( n9374 & ~n2910 ) | ( n9374 & n9375 ) | ( ~n2910 & n9375 ) ;
  assign n9377 = ( n6104 & ~n7255 ) | ( n6104 & 1'b0 ) | ( ~n7255 & 1'b0 ) ;
  assign n9378 = ( n9376 & ~n9377 ) | ( n9376 & 1'b0 ) | ( ~n9377 & 1'b0 ) ;
  assign n9379 = x11 | n9378 ;
  assign n9380 = x11 &  n9378 ;
  assign n9381 = ( n9379 & ~n9380 ) | ( n9379 & 1'b0 ) | ( ~n9380 & 1'b0 ) ;
  assign n9382 = ( n8999 & ~n9009 ) | ( n8999 & n9107 ) | ( ~n9009 & n9107 ) ;
  assign n9383 = ( n9009 & ~n9108 ) | ( n9009 & n9382 ) | ( ~n9108 & n9382 ) ;
  assign n9384 = ~n2995 & n7253 ;
  assign n9385 = n2839 | n7518 ;
  assign n9386 = ~n9384 & n9385 ;
  assign n9387 = n2910 &  n7783 ;
  assign n9388 = ( n9386 & ~n2910 ) | ( n9386 & n9387 ) | ( ~n2910 & n9387 ) ;
  assign n9389 = ( n6330 & ~n7255 ) | ( n6330 & 1'b0 ) | ( ~n7255 & 1'b0 ) ;
  assign n9390 = ( n9388 & ~n9389 ) | ( n9388 & 1'b0 ) | ( ~n9389 & 1'b0 ) ;
  assign n9391 = x11 | n9390 ;
  assign n9392 = x11 &  n9390 ;
  assign n9393 = ( n9391 & ~n9392 ) | ( n9391 & 1'b0 ) | ( ~n9392 & 1'b0 ) ;
  assign n9394 = ( n9012 & ~n9022 ) | ( n9012 & n9106 ) | ( ~n9022 & n9106 ) ;
  assign n9395 = ( n9022 & ~n9107 ) | ( n9022 & n9394 ) | ( ~n9107 & n9394 ) ;
  assign n9402 = ~n2839 & n7783 ;
  assign n9399 = ~n3030 & n7253 ;
  assign n9400 = n2995 | n7518 ;
  assign n9401 = ~n9399 & n9400 ;
  assign n9403 = ( n2839 & n9402 ) | ( n2839 & n9401 ) | ( n9402 & n9401 ) ;
  assign n9404 = ( n6591 & ~n3610 ) | ( n6591 & n7255 ) | ( ~n3610 & n7255 ) ;
  assign n9405 = ( n6592 & n9403 ) | ( n6592 & n9404 ) | ( n9403 & n9404 ) ;
  assign n9406 = x11 &  n9405 ;
  assign n9407 = x11 | n9405 ;
  assign n9408 = ~n9406 & n9407 ;
  assign n9396 = ( n9034 & ~n9032 ) | ( n9034 & n9105 ) | ( ~n9032 & n9105 ) ;
  assign n9397 = ( n9032 & ~n9105 ) | ( n9032 & n9034 ) | ( ~n9105 & n9034 ) ;
  assign n9398 = ( n9396 & ~n9034 ) | ( n9396 & n9397 ) | ( ~n9034 & n9397 ) ;
  assign n9409 = ( n9047 & ~n9037 ) | ( n9047 & n9104 ) | ( ~n9037 & n9104 ) ;
  assign n9410 = ( n9037 & ~n9104 ) | ( n9037 & n9047 ) | ( ~n9104 & n9047 ) ;
  assign n9411 = ( n9409 & ~n9047 ) | ( n9409 & n9410 ) | ( ~n9047 & n9410 ) ;
  assign n9412 = ~n3106 & n7253 ;
  assign n9413 = n3030 | n7518 ;
  assign n9414 = ~n9412 & n9413 ;
  assign n9415 = ~n2995 & n7783 ;
  assign n9416 = ( n2995 & n9414 ) | ( n2995 & n9415 ) | ( n9414 & n9415 ) ;
  assign n9417 = ( n6604 & ~n3609 ) | ( n6604 & n7255 ) | ( ~n3609 & n7255 ) ;
  assign n9418 = ( n6605 & n9416 ) | ( n6605 & n9417 ) | ( n9416 & n9417 ) ;
  assign n9419 = x11 &  n9418 ;
  assign n9420 = x11 | n9418 ;
  assign n9421 = ~n9419 & n9420 ;
  assign n9422 = ( n9057 & ~n9103 ) | ( n9057 & n9060 ) | ( ~n9103 & n9060 ) ;
  assign n9423 = ( n9060 & ~n9057 ) | ( n9060 & n9103 ) | ( ~n9057 & n9103 ) ;
  assign n9424 = ( n9422 & ~n9060 ) | ( n9422 & n9423 ) | ( ~n9060 & n9423 ) ;
  assign n9428 = ~n3030 & n7783 ;
  assign n9425 = ~n3197 & n7253 ;
  assign n9426 = n3106 | n7518 ;
  assign n9427 = ~n9425 & n9426 ;
  assign n9429 = ( n3030 & n9428 ) | ( n3030 & n9427 ) | ( n9428 & n9427 ) ;
  assign n9430 = ( n6311 & ~n3608 ) | ( n6311 & n7255 ) | ( ~n3608 & n7255 ) ;
  assign n9431 = ( n6313 & n9429 ) | ( n6313 & n9430 ) | ( n9429 & n9430 ) ;
  assign n9432 = x11 &  n9431 ;
  assign n9433 = x11 | n9431 ;
  assign n9434 = ~n9432 & n9433 ;
  assign n9438 = ~n7253 & n3266 ;
  assign n9435 = n3106 | n7783 ;
  assign n9436 = n3197 | n7518 ;
  assign n9437 = n9435 &  n9436 ;
  assign n9439 = ( n9438 & ~n3266 ) | ( n9438 & n9437 ) | ( ~n3266 & n9437 ) ;
  assign n9440 = n7255 | n7363 ;
  assign n9441 = n9439 &  n9440 ;
  assign n9442 = x11 | n9441 ;
  assign n9443 = x11 &  n9441 ;
  assign n9444 = ( n9442 & ~n9443 ) | ( n9442 & 1'b0 ) | ( ~n9443 & 1'b0 ) ;
  assign n9445 = ( n9074 & ~n9064 ) | ( n9074 & n9102 ) | ( ~n9064 & n9102 ) ;
  assign n9446 = ( n9103 & ~n9074 ) | ( n9103 & n9445 ) | ( ~n9074 & n9445 ) ;
  assign n9448 = ( n8694 & n9091 ) | ( n8694 & n9101 ) | ( n9091 & n9101 ) ;
  assign n9447 = ( n8694 & ~n9091 ) | ( n8694 & n9101 ) | ( ~n9091 & n9101 ) ;
  assign n9449 = ( n9091 & ~n9448 ) | ( n9091 & n9447 ) | ( ~n9448 & n9447 ) ;
  assign n9455 = n7255 | n7377 ;
  assign n9450 = n3197 | n7783 ;
  assign n9451 = ~n3325 & n7253 ;
  assign n9452 = ( n9450 & ~n9451 ) | ( n9450 & 1'b0 ) | ( ~n9451 & 1'b0 ) ;
  assign n9453 = n3266 &  n7518 ;
  assign n9454 = ( n9452 & ~n3266 ) | ( n9452 & n9453 ) | ( ~n3266 & n9453 ) ;
  assign n9456 = ( n7255 & ~n9455 ) | ( n7255 & n9454 ) | ( ~n9455 & n9454 ) ;
  assign n9457 = x11 &  n9456 ;
  assign n9458 = x11 | n9456 ;
  assign n9459 = ~n9457 & n9458 ;
  assign n9465 = ( n3605 & ~n7255 ) | ( n3605 & n6753 ) | ( ~n7255 & n6753 ) ;
  assign n9460 = ~n3361 & n7253 ;
  assign n9461 = n3325 | n7518 ;
  assign n9462 = ~n9460 & n9461 ;
  assign n9463 = n3266 &  n7783 ;
  assign n9464 = ( n9462 & ~n3266 ) | ( n9462 & n9463 ) | ( ~n3266 & n9463 ) ;
  assign n9466 = ( n6754 & ~n9465 ) | ( n6754 & n9464 ) | ( ~n9465 & n9464 ) ;
  assign n9467 = x11 | n9466 ;
  assign n9468 = ( x11 & ~n9466 ) | ( x11 & 1'b0 ) | ( ~n9466 & 1'b0 ) ;
  assign n9469 = ( n9467 & ~x11 ) | ( n9467 & n9468 ) | ( ~x11 & n9468 ) ;
  assign n9082 = ( x14 & ~n9081 ) | ( x14 & 1'b0 ) | ( ~n9081 & 1'b0 ) ;
  assign n9471 = ( x14 & n9082 ) | ( x14 & n9089 ) | ( n9082 & n9089 ) ;
  assign n9470 = ( x14 & ~n9082 ) | ( x14 & n9089 ) | ( ~n9082 & n9089 ) ;
  assign n9472 = ( n9082 & ~n9471 ) | ( n9082 & n9470 ) | ( ~n9471 & n9470 ) ;
  assign n9473 = x14 &  n9080 ;
  assign n9474 = n9079 &  n9473 ;
  assign n9475 = n9079 | n9473 ;
  assign n9476 = ~n9474 & n9475 ;
  assign n9506 = ~n3460 & n7518 ;
  assign n9503 = n3361 | n7783 ;
  assign n9504 = ~n3601 & n7253 ;
  assign n9505 = ( n9503 & ~n9504 ) | ( n9503 & 1'b0 ) | ( ~n9504 & 1'b0 ) ;
  assign n9507 = ( n3460 & n9506 ) | ( n3460 & n9505 ) | ( n9506 & n9505 ) ;
  assign n9508 = n3361 | n3460 ;
  assign n9509 = n3361 &  n3460 ;
  assign n9510 = ( n9508 & ~n9509 ) | ( n9508 & 1'b0 ) | ( ~n9509 & 1'b0 ) ;
  assign n9511 = ( n3603 & ~n9510 ) | ( n3603 & 1'b0 ) | ( ~n9510 & 1'b0 ) ;
  assign n9512 = ( n7255 & ~n3603 ) | ( n7255 & n9510 ) | ( ~n3603 & n9510 ) ;
  assign n9513 = ( n9507 & n9511 ) | ( n9507 & n9512 ) | ( n9511 & n9512 ) ;
  assign n9514 = x11 | n9513 ;
  assign n9515 = ( x11 & ~n9513 ) | ( x11 & 1'b0 ) | ( ~n9513 & 1'b0 ) ;
  assign n9516 = ( n9514 & ~x11 ) | ( n9514 & n9515 ) | ( ~x11 & n9515 ) ;
  assign n9497 = n7412 | n7255 ;
  assign n9494 = n3547 | n7518 ;
  assign n9495 = n3601 | n7783 ;
  assign n9496 = n9494 &  n9495 ;
  assign n9498 = ( n7255 & ~n9497 ) | ( n7255 & n9496 ) | ( ~n9497 & n9496 ) ;
  assign n9492 = ~n6886 & n7255 ;
  assign n9490 = ~n3460 & n7783 ;
  assign n9487 = ~n3547 & n7253 ;
  assign n9488 = n3601 | n7518 ;
  assign n9489 = ~n9487 & n9488 ;
  assign n9491 = ( n3460 & n9490 ) | ( n3460 & n9489 ) | ( n9490 & n9489 ) ;
  assign n9493 = ( n6886 & n9492 ) | ( n6886 & n9491 ) | ( n9492 & n9491 ) ;
  assign n9499 = ~n3547 & n7251 ;
  assign n9500 = ( n9498 & ~n9493 ) | ( n9498 & n9499 ) | ( ~n9493 & n9499 ) ;
  assign n9501 = ( x11 & ~n9498 ) | ( x11 & n9500 ) | ( ~n9498 & n9500 ) ;
  assign n9502 = ( x11 & ~n9501 ) | ( x11 & 1'b0 ) | ( ~n9501 & 1'b0 ) ;
  assign n9517 = ( n9080 & ~n9516 ) | ( n9080 & n9502 ) | ( ~n9516 & n9502 ) ;
  assign n9477 = n3460 &  n7253 ;
  assign n9478 = n3325 | n7783 ;
  assign n9479 = n3361 | n7518 ;
  assign n9480 = n9478 &  n9479 ;
  assign n9481 = ( n9477 & ~n7253 ) | ( n9477 & n9480 ) | ( ~n7253 & n9480 ) ;
  assign n9482 = ( n6800 & ~n3604 ) | ( n6800 & n7255 ) | ( ~n3604 & n7255 ) ;
  assign n9483 = ( n6801 & n9481 ) | ( n6801 & n9482 ) | ( n9481 & n9482 ) ;
  assign n9485 = x11 &  n9483 ;
  assign n9484 = ~x11 & n9483 ;
  assign n9486 = ( x11 & ~n9485 ) | ( x11 & n9484 ) | ( ~n9485 & n9484 ) ;
  assign n9518 = ( n9476 & ~n9517 ) | ( n9476 & n9486 ) | ( ~n9517 & n9486 ) ;
  assign n9519 = ( n9469 & n9472 ) | ( n9469 & n9518 ) | ( n9472 & n9518 ) ;
  assign n9520 = ( n9449 & n9459 ) | ( n9449 & n9519 ) | ( n9459 & n9519 ) ;
  assign n9521 = ( n9444 & ~n9446 ) | ( n9444 & n9520 ) | ( ~n9446 & n9520 ) ;
  assign n9522 = ( n9424 & n9434 ) | ( n9424 & n9521 ) | ( n9434 & n9521 ) ;
  assign n9523 = ( n9411 & n9421 ) | ( n9411 & n9522 ) | ( n9421 & n9522 ) ;
  assign n9524 = ( n9408 & ~n9398 ) | ( n9408 & n9523 ) | ( ~n9398 & n9523 ) ;
  assign n9525 = ( n9393 & n9395 ) | ( n9393 & n9524 ) | ( n9395 & n9524 ) ;
  assign n9526 = ( n9381 & n9383 ) | ( n9381 & n9525 ) | ( n9383 & n9525 ) ;
  assign n9527 = ( n9369 & ~n9371 ) | ( n9369 & n9526 ) | ( ~n9371 & n9526 ) ;
  assign n9528 = ( n9349 & n9359 ) | ( n9349 & n9527 ) | ( n9359 & n9527 ) ;
  assign n9529 = ( n9336 & n9346 ) | ( n9336 & n9528 ) | ( n9346 & n9528 ) ;
  assign n9530 = ( n9333 & ~n9323 ) | ( n9333 & n9529 ) | ( ~n9323 & n9529 ) ;
  assign n9531 = ( n9318 & n9320 ) | ( n9318 & n9530 ) | ( n9320 & n9530 ) ;
  assign n9532 = ( n9306 & n9308 ) | ( n9306 & n9531 ) | ( n9308 & n9531 ) ;
  assign n9533 = ( n9294 & ~n9296 ) | ( n9294 & n9532 ) | ( ~n9296 & n9532 ) ;
  assign n9534 = ( n9274 & n9284 ) | ( n9274 & n9533 ) | ( n9284 & n9533 ) ;
  assign n9535 = ( n9261 & n9271 ) | ( n9261 & n9534 ) | ( n9271 & n9534 ) ;
  assign n9536 = ( n9256 & ~n9258 ) | ( n9256 & n9535 ) | ( ~n9258 & n9535 ) ;
  assign n9537 = ( n9244 & ~n9246 ) | ( n9244 & n9536 ) | ( ~n9246 & n9536 ) ;
  assign n9538 = ( n9232 & n9234 ) | ( n9232 & n9537 ) | ( n9234 & n9537 ) ;
  assign n9539 = ( n9220 & n9222 ) | ( n9220 & n9538 ) | ( n9222 & n9538 ) ;
  assign n9540 = ( n9208 & ~n9210 ) | ( n9208 & n9539 ) | ( ~n9210 & n9539 ) ;
  assign n9541 = ( n9196 & n9198 ) | ( n9196 & n9540 ) | ( n9198 & n9540 ) ;
  assign n9542 = ( n9184 & n9186 ) | ( n9184 & n9541 ) | ( n9186 & n9541 ) ;
  assign n9543 = ( n9124 & n9126 ) | ( n9124 & n9136 ) | ( n9126 & n9136 ) ;
  assign n9544 = ( n9124 & ~n9136 ) | ( n9124 & n9126 ) | ( ~n9136 & n9126 ) ;
  assign n9545 = ( n9136 & ~n9543 ) | ( n9136 & n9544 ) | ( ~n9543 & n9544 ) ;
  assign n9549 = ~n946 & n8764 ;
  assign n9546 = ~n1151 & n8105 ;
  assign n9547 = n1043 | n8429 ;
  assign n9548 = ~n9546 & n9547 ;
  assign n9550 = ( n946 & n9549 ) | ( n946 & n9548 ) | ( n9549 & n9548 ) ;
  assign n9551 = ( n8107 & ~n4038 ) | ( n8107 & n9550 ) | ( ~n4038 & n9550 ) ;
  assign n9552 = ~n8107 & n9551 ;
  assign n9553 = ( x8 & ~n9550 ) | ( x8 & n9552 ) | ( ~n9550 & n9552 ) ;
  assign n9554 = ( n9550 & ~x8 ) | ( n9550 & n9552 ) | ( ~x8 & n9552 ) ;
  assign n9555 = ( n9553 & ~n9552 ) | ( n9553 & n9554 ) | ( ~n9552 & n9554 ) ;
  assign n9556 = ( n9542 & ~n9545 ) | ( n9542 & n9555 ) | ( ~n9545 & n9555 ) ;
  assign n9566 = ( n8793 & n9137 ) | ( n8793 & n9147 ) | ( n9137 & n9147 ) ;
  assign n9567 = ( n8793 & ~n9137 ) | ( n8793 & n9147 ) | ( ~n9137 & n9147 ) ;
  assign n9568 = ( n9137 & ~n9566 ) | ( n9137 & n9567 ) | ( ~n9566 & n9567 ) ;
  assign n9557 = n702 | n9160 ;
  assign n9558 = ~n9158 |  n9154 ;
  assign n9559 = n599 | n9558 ;
  assign n9560 = n9557 &  n9559 ;
  assign n9561 = n3937 &  n9155 ;
  assign n9562 = ( n9560 & ~n3937 ) | ( n9560 & n9561 ) | ( ~n3937 & n9561 ) ;
  assign n9563 = x5 &  n9562 ;
  assign n9564 = x5 | n9562 ;
  assign n9565 = ~n9563 & n9564 ;
  assign n9569 = ( n9556 & ~n9568 ) | ( n9556 & n9565 ) | ( ~n9568 & n9565 ) ;
  assign n9173 = ( n9148 & n9166 ) | ( n9148 & n9169 ) | ( n9166 & n9169 ) ;
  assign n9174 = ( n9169 & ~n9173 ) | ( n9169 & n9170 ) | ( ~n9173 & n9170 ) ;
  assign n9570 = ( n9186 & ~n9184 ) | ( n9186 & n9541 ) | ( ~n9184 & n9541 ) ;
  assign n9571 = ( n9184 & ~n9541 ) | ( n9184 & n9186 ) | ( ~n9541 & n9186 ) ;
  assign n9572 = ( n9570 & ~n9186 ) | ( n9570 & n9571 ) | ( ~n9186 & n9571 ) ;
  assign n9576 = ~n8105 & n1267 ;
  assign n9573 = n1043 | n8764 ;
  assign n9574 = n1151 | n8429 ;
  assign n9575 = n9573 &  n9574 ;
  assign n9577 = ( n9576 & ~n1267 ) | ( n9576 & n9575 ) | ( ~n1267 & n9575 ) ;
  assign n9578 = ( n8107 & ~n3952 ) | ( n8107 & n9577 ) | ( ~n3952 & n9577 ) ;
  assign n9579 = ~n8107 & n9578 ;
  assign n9580 = ( x8 & ~n9577 ) | ( x8 & n9579 ) | ( ~n9577 & n9579 ) ;
  assign n9581 = ( n9577 & ~x8 ) | ( n9577 & n9579 ) | ( ~x8 & n9579 ) ;
  assign n9582 = ( n9580 & ~n9579 ) | ( n9580 & n9581 ) | ( ~n9579 & n9581 ) ;
  assign n9583 = ( n9198 & ~n9196 ) | ( n9198 & n9540 ) | ( ~n9196 & n9540 ) ;
  assign n9584 = ( n9196 & ~n9540 ) | ( n9196 & n9198 ) | ( ~n9540 & n9198 ) ;
  assign n9585 = ( n9583 & ~n9198 ) | ( n9583 & n9584 ) | ( ~n9198 & n9584 ) ;
  assign n9586 = n1151 | n8764 ;
  assign n9587 = ~n1378 & n8105 ;
  assign n9588 = ( n9586 & ~n9587 ) | ( n9586 & 1'b0 ) | ( ~n9587 & 1'b0 ) ;
  assign n9589 = n1267 &  n8429 ;
  assign n9590 = ( n9588 & ~n1267 ) | ( n9588 & n9589 ) | ( ~n1267 & n9589 ) ;
  assign n9591 = ( n4061 & n8107 ) | ( n4061 & n9590 ) | ( n8107 & n9590 ) ;
  assign n9592 = ~n8107 & n9591 ;
  assign n9593 = ( x8 & ~n9590 ) | ( x8 & n9592 ) | ( ~n9590 & n9592 ) ;
  assign n9594 = ( n9590 & ~x8 ) | ( n9590 & n9592 ) | ( ~x8 & n9592 ) ;
  assign n9595 = ( n9593 & ~n9592 ) | ( n9593 & n9594 ) | ( ~n9592 & n9594 ) ;
  assign n9599 = n1483 &  n8105 ;
  assign n9600 = n1378 | n8429 ;
  assign n9601 = ~n9599 & n9600 ;
  assign n9602 = n1267 &  n8764 ;
  assign n9603 = ( n9601 & ~n1267 ) | ( n9601 & n9602 ) | ( ~n1267 & n9602 ) ;
  assign n9604 = ( n4422 & n8107 ) | ( n4422 & n9603 ) | ( n8107 & n9603 ) ;
  assign n9605 = ~n8107 & n9604 ;
  assign n9606 = ( x8 & ~n9603 ) | ( x8 & n9605 ) | ( ~n9603 & n9605 ) ;
  assign n9607 = ( n9603 & ~x8 ) | ( n9603 & n9605 ) | ( ~x8 & n9605 ) ;
  assign n9608 = ( n9606 & ~n9605 ) | ( n9606 & n9607 ) | ( ~n9605 & n9607 ) ;
  assign n9596 = ( n9208 & ~n9539 ) | ( n9208 & n9210 ) | ( ~n9539 & n9210 ) ;
  assign n9597 = ( n9210 & ~n9208 ) | ( n9210 & n9539 ) | ( ~n9208 & n9539 ) ;
  assign n9598 = ( n9596 & ~n9210 ) | ( n9596 & n9597 ) | ( ~n9210 & n9597 ) ;
  assign n9609 = ( n9222 & ~n9220 ) | ( n9222 & n9538 ) | ( ~n9220 & n9538 ) ;
  assign n9610 = ( n9220 & ~n9538 ) | ( n9220 & n9222 ) | ( ~n9538 & n9222 ) ;
  assign n9611 = ( n9609 & ~n9222 ) | ( n9609 & n9610 ) | ( ~n9222 & n9610 ) ;
  assign n9612 = n1378 | n8764 ;
  assign n9613 = ~n1566 & n8105 ;
  assign n9614 = ( n9612 & ~n9613 ) | ( n9612 & 1'b0 ) | ( ~n9613 & 1'b0 ) ;
  assign n9615 = n1483 &  n8429 ;
  assign n9616 = ( n9614 & ~n1483 ) | ( n9614 & n9615 ) | ( ~n1483 & n9615 ) ;
  assign n9617 = ( n5038 & n8107 ) | ( n5038 & n9616 ) | ( n8107 & n9616 ) ;
  assign n9618 = ~n8107 & n9617 ;
  assign n9619 = ( x8 & ~n9616 ) | ( x8 & n9618 ) | ( ~n9616 & n9618 ) ;
  assign n9620 = ( n9616 & ~x8 ) | ( n9616 & n9618 ) | ( ~x8 & n9618 ) ;
  assign n9621 = ( n9619 & ~n9618 ) | ( n9619 & n9620 ) | ( ~n9618 & n9620 ) ;
  assign n9622 = ( n9234 & ~n9232 ) | ( n9234 & n9537 ) | ( ~n9232 & n9537 ) ;
  assign n9623 = ( n9232 & ~n9537 ) | ( n9232 & n9234 ) | ( ~n9537 & n9234 ) ;
  assign n9624 = ( n9622 & ~n9234 ) | ( n9622 & n9623 ) | ( ~n9234 & n9623 ) ;
  assign n9625 = ~n1671 & n8105 ;
  assign n9626 = n1566 | n8429 ;
  assign n9627 = ~n9625 & n9626 ;
  assign n9628 = n1483 &  n8764 ;
  assign n9629 = ( n9627 & ~n1483 ) | ( n9627 & n9628 ) | ( ~n1483 & n9628 ) ;
  assign n9630 = ( n4274 & n8107 ) | ( n4274 & n9629 ) | ( n8107 & n9629 ) ;
  assign n9631 = ~n8107 & n9630 ;
  assign n9632 = ( x8 & ~n9629 ) | ( x8 & n9631 ) | ( ~n9629 & n9631 ) ;
  assign n9633 = ( n9629 & ~x8 ) | ( n9629 & n9631 ) | ( ~x8 & n9631 ) ;
  assign n9634 = ( n9632 & ~n9631 ) | ( n9632 & n9633 ) | ( ~n9631 & n9633 ) ;
  assign n9641 = ~n1566 & n8764 ;
  assign n9638 = ~n1748 & n8105 ;
  assign n9639 = n1671 | n8429 ;
  assign n9640 = ~n9638 & n9639 ;
  assign n9642 = ( n1566 & n9641 ) | ( n1566 & n9640 ) | ( n9641 & n9640 ) ;
  assign n9643 = ( n8107 & ~n4597 ) | ( n8107 & n9642 ) | ( ~n4597 & n9642 ) ;
  assign n9644 = ~n8107 & n9643 ;
  assign n9645 = ( x8 & ~n9642 ) | ( x8 & n9644 ) | ( ~n9642 & n9644 ) ;
  assign n9646 = ( n9642 & ~x8 ) | ( n9642 & n9644 ) | ( ~x8 & n9644 ) ;
  assign n9647 = ( n9645 & ~n9644 ) | ( n9645 & n9646 ) | ( ~n9644 & n9646 ) ;
  assign n9635 = ( n9244 & ~n9536 ) | ( n9244 & n9246 ) | ( ~n9536 & n9246 ) ;
  assign n9636 = ( n9246 & ~n9244 ) | ( n9246 & n9536 ) | ( ~n9244 & n9536 ) ;
  assign n9637 = ( n9635 & ~n9246 ) | ( n9635 & n9636 ) | ( ~n9246 & n9636 ) ;
  assign n9650 = n1875 &  n8105 ;
  assign n9651 = n1671 | n8764 ;
  assign n9652 = n1748 | n8429 ;
  assign n9653 = n9651 &  n9652 ;
  assign n9654 = ( n9650 & ~n8105 ) | ( n9650 & n9653 ) | ( ~n8105 & n9653 ) ;
  assign n9655 = ( n4577 & ~n3625 ) | ( n4577 & n8107 ) | ( ~n3625 & n8107 ) ;
  assign n9656 = ( n4579 & n9654 ) | ( n4579 & n9655 ) | ( n9654 & n9655 ) ;
  assign n9657 = x8 &  n9656 ;
  assign n9658 = x8 | n9656 ;
  assign n9659 = ~n9657 & n9658 ;
  assign n9648 = ( n9256 & n9258 ) | ( n9256 & n9535 ) | ( n9258 & n9535 ) ;
  assign n9649 = ( n9258 & ~n9648 ) | ( n9258 & n9536 ) | ( ~n9648 & n9536 ) ;
  assign n9660 = ~n1940 & n8105 ;
  assign n9661 = n1875 | n8429 ;
  assign n9662 = ~n9660 & n9661 ;
  assign n9663 = ~n1748 & n8764 ;
  assign n9664 = ( n1748 & n9662 ) | ( n1748 & n9663 ) | ( n9662 & n9663 ) ;
  assign n9665 = ( n4740 & ~n3624 ) | ( n4740 & n8107 ) | ( ~n3624 & n8107 ) ;
  assign n9666 = ( n4742 & n9664 ) | ( n4742 & n9665 ) | ( n9664 & n9665 ) ;
  assign n9667 = x8 | n9666 ;
  assign n9668 = ( x8 & ~n9666 ) | ( x8 & 1'b0 ) | ( ~n9666 & 1'b0 ) ;
  assign n9669 = ( n9667 & ~x8 ) | ( n9667 & n9668 ) | ( ~x8 & n9668 ) ;
  assign n9670 = ( n9271 & ~n9261 ) | ( n9271 & n9534 ) | ( ~n9261 & n9534 ) ;
  assign n9671 = ( n9261 & ~n9271 ) | ( n9261 & n9534 ) | ( ~n9271 & n9534 ) ;
  assign n9672 = ( n9670 & ~n9534 ) | ( n9670 & n9671 ) | ( ~n9534 & n9671 ) ;
  assign n9676 = ~n1875 & n8764 ;
  assign n9673 = ~n2022 & n8105 ;
  assign n9674 = n1940 | n8429 ;
  assign n9675 = ~n9673 & n9674 ;
  assign n9677 = ( n1875 & n9676 ) | ( n1875 & n9675 ) | ( n9676 & n9675 ) ;
  assign n9678 = ( n4761 & ~n3623 ) | ( n4761 & n8107 ) | ( ~n3623 & n8107 ) ;
  assign n9679 = ( n4762 & n9677 ) | ( n4762 & n9678 ) | ( n9677 & n9678 ) ;
  assign n9680 = x8 | n9679 ;
  assign n9681 = ( x8 & ~n9679 ) | ( x8 & 1'b0 ) | ( ~n9679 & 1'b0 ) ;
  assign n9682 = ( n9680 & ~x8 ) | ( n9680 & n9681 ) | ( ~x8 & n9681 ) ;
  assign n9683 = ( n9284 & ~n9274 ) | ( n9284 & n9533 ) | ( ~n9274 & n9533 ) ;
  assign n9684 = ( n9274 & ~n9284 ) | ( n9274 & n9533 ) | ( ~n9284 & n9533 ) ;
  assign n9685 = ( n9683 & ~n9533 ) | ( n9683 & n9684 ) | ( ~n9533 & n9684 ) ;
  assign n9688 = ~n2127 & n8105 ;
  assign n9689 = n2022 | n8429 ;
  assign n9690 = ~n9688 & n9689 ;
  assign n9691 = ~n1940 & n8764 ;
  assign n9692 = ( n1940 & n9690 ) | ( n1940 & n9691 ) | ( n9690 & n9691 ) ;
  assign n9693 = ( n5085 & ~n3622 ) | ( n5085 & n8107 ) | ( ~n3622 & n8107 ) ;
  assign n9694 = ( n5086 & n9692 ) | ( n5086 & n9693 ) | ( n9692 & n9693 ) ;
  assign n9695 = x8 &  n9694 ;
  assign n9696 = x8 | n9694 ;
  assign n9697 = ~n9695 & n9696 ;
  assign n9686 = ( n9294 & n9296 ) | ( n9294 & n9532 ) | ( n9296 & n9532 ) ;
  assign n9687 = ( n9296 & ~n9686 ) | ( n9296 & n9533 ) | ( ~n9686 & n9533 ) ;
  assign n9698 = ( n9306 & ~n9308 ) | ( n9306 & n9531 ) | ( ~n9308 & n9531 ) ;
  assign n9699 = ( n9308 & ~n9532 ) | ( n9308 & n9698 ) | ( ~n9532 & n9698 ) ;
  assign n9700 = ~n2178 & n8105 ;
  assign n9701 = n2127 | n8429 ;
  assign n9702 = ~n9700 & n9701 ;
  assign n9703 = ~n2022 & n8764 ;
  assign n9704 = ( n2022 & n9702 ) | ( n2022 & n9703 ) | ( n9702 & n9703 ) ;
  assign n9705 = ( n4931 & ~n3621 ) | ( n4931 & n8107 ) | ( ~n3621 & n8107 ) ;
  assign n9706 = ( n4933 & n9704 ) | ( n4933 & n9705 ) | ( n9704 & n9705 ) ;
  assign n9707 = x8 &  n9706 ;
  assign n9708 = x8 | n9706 ;
  assign n9709 = ~n9707 & n9708 ;
  assign n9710 = ( n9318 & ~n9320 ) | ( n9318 & n9530 ) | ( ~n9320 & n9530 ) ;
  assign n9711 = ( n9320 & ~n9531 ) | ( n9320 & n9710 ) | ( ~n9531 & n9710 ) ;
  assign n9712 = n2296 &  n8105 ;
  assign n9713 = n2127 | n8764 ;
  assign n9714 = n2178 | n8429 ;
  assign n9715 = n9713 &  n9714 ;
  assign n9716 = ( n9712 & ~n8105 ) | ( n9712 & n9715 ) | ( ~n8105 & n9715 ) ;
  assign n9717 = ( n5280 & ~n3620 ) | ( n5280 & n8107 ) | ( ~n3620 & n8107 ) ;
  assign n9718 = ( n5282 & n9716 ) | ( n5282 & n9717 ) | ( n9716 & n9717 ) ;
  assign n9719 = x8 &  n9718 ;
  assign n9720 = x8 | n9718 ;
  assign n9721 = ~n9719 & n9720 ;
  assign n9725 = ~n2178 & n8764 ;
  assign n9722 = ~n2392 & n8105 ;
  assign n9723 = n2296 | n8429 ;
  assign n9724 = ~n9722 & n9723 ;
  assign n9726 = ( n2178 & n9725 ) | ( n2178 & n9724 ) | ( n9725 & n9724 ) ;
  assign n9727 = ( n5266 & ~n3619 ) | ( n5266 & n8107 ) | ( ~n3619 & n8107 ) ;
  assign n9728 = ( n5268 & n9726 ) | ( n5268 & n9727 ) | ( n9726 & n9727 ) ;
  assign n9729 = x8 | n9728 ;
  assign n9730 = ( x8 & ~n9728 ) | ( x8 & 1'b0 ) | ( ~n9728 & 1'b0 ) ;
  assign n9731 = ( n9729 & ~x8 ) | ( n9729 & n9730 ) | ( ~x8 & n9730 ) ;
  assign n9732 = ( n9323 & n9333 ) | ( n9323 & n9529 ) | ( n9333 & n9529 ) ;
  assign n9733 = ( n9323 & ~n9529 ) | ( n9323 & n9333 ) | ( ~n9529 & n9333 ) ;
  assign n9734 = ( n9529 & ~n9732 ) | ( n9529 & n9733 ) | ( ~n9732 & n9733 ) ;
  assign n9738 = ~n2296 & n8764 ;
  assign n9735 = ~n2483 & n8105 ;
  assign n9736 = n2392 | n8429 ;
  assign n9737 = ~n9735 & n9736 ;
  assign n9739 = ( n2296 & n9738 ) | ( n2296 & n9737 ) | ( n9738 & n9737 ) ;
  assign n9740 = ( n5497 & ~n3618 ) | ( n5497 & n8107 ) | ( ~n3618 & n8107 ) ;
  assign n9741 = ( n5499 & n9739 ) | ( n5499 & n9740 ) | ( n9739 & n9740 ) ;
  assign n9742 = x8 | n9741 ;
  assign n9743 = ( x8 & ~n9741 ) | ( x8 & 1'b0 ) | ( ~n9741 & 1'b0 ) ;
  assign n9744 = ( n9742 & ~x8 ) | ( n9742 & n9743 ) | ( ~x8 & n9743 ) ;
  assign n9745 = ( n9346 & ~n9336 ) | ( n9346 & n9528 ) | ( ~n9336 & n9528 ) ;
  assign n9746 = ( n9336 & ~n9346 ) | ( n9336 & n9528 ) | ( ~n9346 & n9528 ) ;
  assign n9747 = ( n9745 & ~n9528 ) | ( n9745 & n9746 ) | ( ~n9528 & n9746 ) ;
  assign n9751 = ~n2392 & n8764 ;
  assign n9748 = ~n2569 & n8105 ;
  assign n9749 = n2483 | n8429 ;
  assign n9750 = ~n9748 & n9749 ;
  assign n9752 = ( n2392 & n9751 ) | ( n2392 & n9750 ) | ( n9751 & n9750 ) ;
  assign n9753 = ( n5519 & ~n3617 ) | ( n5519 & n8107 ) | ( ~n3617 & n8107 ) ;
  assign n9754 = ( n5520 & n9752 ) | ( n5520 & n9753 ) | ( n9752 & n9753 ) ;
  assign n9755 = x8 | n9754 ;
  assign n9756 = ( x8 & ~n9754 ) | ( x8 & 1'b0 ) | ( ~n9754 & 1'b0 ) ;
  assign n9757 = ( n9755 & ~x8 ) | ( n9755 & n9756 ) | ( ~x8 & n9756 ) ;
  assign n9758 = ( n9359 & ~n9349 ) | ( n9359 & n9527 ) | ( ~n9349 & n9527 ) ;
  assign n9759 = ( n9349 & ~n9359 ) | ( n9349 & n9527 ) | ( ~n9359 & n9527 ) ;
  assign n9760 = ( n9758 & ~n9527 ) | ( n9758 & n9759 ) | ( ~n9527 & n9759 ) ;
  assign n9763 = n2665 &  n8105 ;
  assign n9764 = n2483 | n8764 ;
  assign n9765 = n2569 | n8429 ;
  assign n9766 = n9764 &  n9765 ;
  assign n9767 = ( n9763 & ~n8105 ) | ( n9763 & n9766 ) | ( ~n8105 & n9766 ) ;
  assign n9768 = ( n5886 & ~n3616 ) | ( n5886 & n8107 ) | ( ~n3616 & n8107 ) ;
  assign n9769 = ( n5887 & n9767 ) | ( n5887 & n9768 ) | ( n9767 & n9768 ) ;
  assign n9770 = x8 &  n9769 ;
  assign n9771 = x8 | n9769 ;
  assign n9772 = ~n9770 & n9771 ;
  assign n9761 = ( n9369 & n9371 ) | ( n9369 & n9526 ) | ( n9371 & n9526 ) ;
  assign n9762 = ( n9371 & ~n9761 ) | ( n9371 & n9527 ) | ( ~n9761 & n9527 ) ;
  assign n9773 = ( n9381 & ~n9383 ) | ( n9381 & n9525 ) | ( ~n9383 & n9525 ) ;
  assign n9774 = ( n9383 & ~n9526 ) | ( n9383 & n9773 ) | ( ~n9526 & n9773 ) ;
  assign n9775 = n2751 &  n8105 ;
  assign n9776 = n2569 | n8764 ;
  assign n9777 = n2665 | n8429 ;
  assign n9778 = n9776 &  n9777 ;
  assign n9779 = ( n9775 & ~n8105 ) | ( n9775 & n9778 ) | ( ~n8105 & n9778 ) ;
  assign n9780 = ( n5702 & ~n3615 ) | ( n5702 & n8107 ) | ( ~n3615 & n8107 ) ;
  assign n9781 = ( n5704 & n9779 ) | ( n5704 & n9780 ) | ( n9779 & n9780 ) ;
  assign n9782 = x8 &  n9781 ;
  assign n9783 = x8 | n9781 ;
  assign n9784 = ~n9782 & n9783 ;
  assign n9785 = ( n9393 & ~n9395 ) | ( n9393 & n9524 ) | ( ~n9395 & n9524 ) ;
  assign n9786 = ( n9395 & ~n9525 ) | ( n9395 & n9785 ) | ( ~n9525 & n9785 ) ;
  assign n9790 = ~n2751 & n8429 ;
  assign n9787 = n2665 | n8764 ;
  assign n9788 = ~n2783 & n8105 ;
  assign n9789 = ( n9787 & ~n9788 ) | ( n9787 & 1'b0 ) | ( ~n9788 & 1'b0 ) ;
  assign n9791 = ( n2751 & n9790 ) | ( n2751 & n9789 ) | ( n9790 & n9789 ) ;
  assign n9792 = ( n6116 & ~n3614 ) | ( n6116 & n8107 ) | ( ~n3614 & n8107 ) ;
  assign n9793 = ( n6118 & n9791 ) | ( n6118 & n9792 ) | ( n9791 & n9792 ) ;
  assign n9794 = x8 &  n9793 ;
  assign n9795 = x8 | n9793 ;
  assign n9796 = ~n9794 & n9795 ;
  assign n9800 = ~n8105 & n2910 ;
  assign n9797 = n2751 | n8764 ;
  assign n9798 = n2783 | n8429 ;
  assign n9799 = n9797 &  n9798 ;
  assign n9801 = ( n9800 & ~n2910 ) | ( n9800 & n9799 ) | ( ~n2910 & n9799 ) ;
  assign n9802 = n2751 | n2783 ;
  assign n9803 = ( n2751 & ~n2783 ) | ( n2751 & 1'b0 ) | ( ~n2783 & 1'b0 ) ;
  assign n9804 = ( n9802 & ~n2751 ) | ( n9802 & n9803 ) | ( ~n2751 & n9803 ) ;
  assign n9805 = ( n3613 & ~n9804 ) | ( n3613 & 1'b0 ) | ( ~n9804 & 1'b0 ) ;
  assign n9806 = ( n8107 & ~n3613 ) | ( n8107 & n9804 ) | ( ~n3613 & n9804 ) ;
  assign n9807 = ( n9801 & n9805 ) | ( n9801 & n9806 ) | ( n9805 & n9806 ) ;
  assign n9808 = x8 | n9807 ;
  assign n9809 = ( x8 & ~n9807 ) | ( x8 & 1'b0 ) | ( ~n9807 & 1'b0 ) ;
  assign n9810 = ( n9808 & ~x8 ) | ( n9808 & n9809 ) | ( ~x8 & n9809 ) ;
  assign n9811 = ( n9398 & n9408 ) | ( n9398 & n9523 ) | ( n9408 & n9523 ) ;
  assign n9812 = ( n9398 & ~n9523 ) | ( n9398 & n9408 ) | ( ~n9523 & n9408 ) ;
  assign n9813 = ( n9523 & ~n9811 ) | ( n9523 & n9812 ) | ( ~n9811 & n9812 ) ;
  assign n9814 = n2783 | n8764 ;
  assign n9815 = ~n2839 & n8105 ;
  assign n9816 = ( n9814 & ~n9815 ) | ( n9814 & 1'b0 ) | ( ~n9815 & 1'b0 ) ;
  assign n9817 = n2910 &  n8429 ;
  assign n9818 = ( n9816 & ~n2910 ) | ( n9816 & n9817 ) | ( ~n2910 & n9817 ) ;
  assign n9819 = ( n6104 & ~n8107 ) | ( n6104 & 1'b0 ) | ( ~n8107 & 1'b0 ) ;
  assign n9820 = ( n9818 & ~n9819 ) | ( n9818 & 1'b0 ) | ( ~n9819 & 1'b0 ) ;
  assign n9821 = x8 | n9820 ;
  assign n9822 = x8 &  n9820 ;
  assign n9823 = ( n9821 & ~n9822 ) | ( n9821 & 1'b0 ) | ( ~n9822 & 1'b0 ) ;
  assign n9824 = ( n9421 & ~n9411 ) | ( n9421 & n9522 ) | ( ~n9411 & n9522 ) ;
  assign n9825 = ( n9411 & ~n9421 ) | ( n9411 & n9522 ) | ( ~n9421 & n9522 ) ;
  assign n9826 = ( n9824 & ~n9522 ) | ( n9824 & n9825 ) | ( ~n9522 & n9825 ) ;
  assign n9827 = ~n2995 & n8105 ;
  assign n9828 = n2839 | n8429 ;
  assign n9829 = ~n9827 & n9828 ;
  assign n9830 = n2910 &  n8764 ;
  assign n9831 = ( n9829 & ~n2910 ) | ( n9829 & n9830 ) | ( ~n2910 & n9830 ) ;
  assign n9832 = ~n2839 & n2910 ;
  assign n9833 = ( n2839 & ~n2910 ) | ( n2839 & 1'b0 ) | ( ~n2910 & 1'b0 ) ;
  assign n9834 = n9832 | n9833 ;
  assign n9836 = ( n3611 & ~n8107 ) | ( n3611 & n9834 ) | ( ~n8107 & n9834 ) ;
  assign n9835 = n3611 &  n9834 ;
  assign n9837 = ( n9831 & ~n9836 ) | ( n9831 & n9835 ) | ( ~n9836 & n9835 ) ;
  assign n9838 = x8 | n9837 ;
  assign n9839 = x8 &  n9837 ;
  assign n9840 = ( n9838 & ~n9839 ) | ( n9838 & 1'b0 ) | ( ~n9839 & 1'b0 ) ;
  assign n9841 = ( n9434 & ~n9424 ) | ( n9434 & n9521 ) | ( ~n9424 & n9521 ) ;
  assign n9842 = ( n9424 & ~n9434 ) | ( n9424 & n9521 ) | ( ~n9434 & n9521 ) ;
  assign n9843 = ( n9841 & ~n9521 ) | ( n9841 & n9842 ) | ( ~n9521 & n9842 ) ;
  assign n9849 = ~n2839 & n8764 ;
  assign n9846 = ~n3030 & n8105 ;
  assign n9847 = n2995 | n8429 ;
  assign n9848 = ~n9846 & n9847 ;
  assign n9850 = ( n2839 & n9849 ) | ( n2839 & n9848 ) | ( n9849 & n9848 ) ;
  assign n9851 = ( n6591 & ~n3610 ) | ( n6591 & n8107 ) | ( ~n3610 & n8107 ) ;
  assign n9852 = ( n6592 & n9850 ) | ( n6592 & n9851 ) | ( n9850 & n9851 ) ;
  assign n9853 = x8 &  n9852 ;
  assign n9854 = x8 | n9852 ;
  assign n9855 = ~n9853 & n9854 ;
  assign n9844 = ( n9444 & n9446 ) | ( n9444 & n9520 ) | ( n9446 & n9520 ) ;
  assign n9845 = ( n9446 & ~n9844 ) | ( n9446 & n9521 ) | ( ~n9844 & n9521 ) ;
  assign n9856 = ( n9449 & ~n9519 ) | ( n9449 & n9459 ) | ( ~n9519 & n9459 ) ;
  assign n9857 = ( n9519 & ~n9520 ) | ( n9519 & n9856 ) | ( ~n9520 & n9856 ) ;
  assign n9858 = ~n3106 & n8105 ;
  assign n9859 = n3030 | n8429 ;
  assign n9860 = ~n9858 & n9859 ;
  assign n9861 = ~n2995 & n8764 ;
  assign n9862 = ( n2995 & n9860 ) | ( n2995 & n9861 ) | ( n9860 & n9861 ) ;
  assign n9863 = ( n6604 & ~n3609 ) | ( n6604 & n8107 ) | ( ~n3609 & n8107 ) ;
  assign n9864 = ( n6605 & n9862 ) | ( n6605 & n9863 ) | ( n9862 & n9863 ) ;
  assign n9865 = x8 &  n9864 ;
  assign n9866 = x8 | n9864 ;
  assign n9867 = ~n9865 & n9866 ;
  assign n9868 = ( n9469 & ~n9518 ) | ( n9469 & n9472 ) | ( ~n9518 & n9472 ) ;
  assign n9869 = ( n9472 & ~n9469 ) | ( n9472 & n9518 ) | ( ~n9469 & n9518 ) ;
  assign n9870 = ( n9868 & ~n9472 ) | ( n9868 & n9869 ) | ( ~n9472 & n9869 ) ;
  assign n9874 = ~n3030 & n8764 ;
  assign n9871 = ~n3197 & n8105 ;
  assign n9872 = n3106 | n8429 ;
  assign n9873 = ~n9871 & n9872 ;
  assign n9875 = ( n3030 & n9874 ) | ( n3030 & n9873 ) | ( n9874 & n9873 ) ;
  assign n9876 = ( n6311 & ~n3608 ) | ( n6311 & n8107 ) | ( ~n3608 & n8107 ) ;
  assign n9877 = ( n6313 & n9875 ) | ( n6313 & n9876 ) | ( n9875 & n9876 ) ;
  assign n9878 = x8 &  n9877 ;
  assign n9879 = x8 | n9877 ;
  assign n9880 = ~n9878 & n9879 ;
  assign n9884 = ~n8105 & n3266 ;
  assign n9881 = n3106 | n8764 ;
  assign n9882 = n3197 | n8429 ;
  assign n9883 = n9881 &  n9882 ;
  assign n9885 = ( n9884 & ~n3266 ) | ( n9884 & n9883 ) | ( ~n3266 & n9883 ) ;
  assign n9886 = ( n6654 & ~n3607 ) | ( n6654 & n8107 ) | ( ~n3607 & n8107 ) ;
  assign n9887 = ( n6655 & n9885 ) | ( n6655 & n9886 ) | ( n9885 & n9886 ) ;
  assign n9888 = x8 | n9887 ;
  assign n9889 = ( x8 & ~n9887 ) | ( x8 & 1'b0 ) | ( ~n9887 & 1'b0 ) ;
  assign n9890 = ( n9888 & ~x8 ) | ( n9888 & n9889 ) | ( ~x8 & n9889 ) ;
  assign n9891 = ( n9486 & ~n9476 ) | ( n9486 & n9517 ) | ( ~n9476 & n9517 ) ;
  assign n9892 = ( n9518 & ~n9486 ) | ( n9518 & n9891 ) | ( ~n9486 & n9891 ) ;
  assign n9894 = ( n9080 & n9502 ) | ( n9080 & n9516 ) | ( n9502 & n9516 ) ;
  assign n9893 = ( n9080 & ~n9502 ) | ( n9080 & n9516 ) | ( ~n9502 & n9516 ) ;
  assign n9895 = ( n9502 & ~n9894 ) | ( n9502 & n9893 ) | ( ~n9894 & n9893 ) ;
  assign n9901 = ( n3606 & ~n8107 ) | ( n3606 & n6705 ) | ( ~n8107 & n6705 ) ;
  assign n9896 = n3197 | n8764 ;
  assign n9897 = ~n3325 & n8105 ;
  assign n9898 = ( n9896 & ~n9897 ) | ( n9896 & 1'b0 ) | ( ~n9897 & 1'b0 ) ;
  assign n9899 = n3266 &  n8429 ;
  assign n9900 = ( n9898 & ~n3266 ) | ( n9898 & n9899 ) | ( ~n3266 & n9899 ) ;
  assign n9902 = ( n6706 & ~n9901 ) | ( n6706 & n9900 ) | ( ~n9901 & n9900 ) ;
  assign n9904 = x8 &  n9902 ;
  assign n9903 = ~x8 & n9902 ;
  assign n9905 = ( x8 & ~n9904 ) | ( x8 & n9903 ) | ( ~n9904 & n9903 ) ;
  assign n9911 = ( n3605 & ~n8107 ) | ( n3605 & n6753 ) | ( ~n8107 & n6753 ) ;
  assign n9906 = ~n3361 & n8105 ;
  assign n9907 = n3325 | n8429 ;
  assign n9908 = ~n9906 & n9907 ;
  assign n9909 = n3266 &  n8764 ;
  assign n9910 = ( n9908 & ~n3266 ) | ( n9908 & n9909 ) | ( ~n3266 & n9909 ) ;
  assign n9912 = ( n6754 & ~n9911 ) | ( n6754 & n9910 ) | ( ~n9911 & n9910 ) ;
  assign n9913 = x8 | n9912 ;
  assign n9914 = x8 &  n9912 ;
  assign n9915 = ( n9913 & ~n9914 ) | ( n9913 & 1'b0 ) | ( ~n9914 & 1'b0 ) ;
  assign n9916 = ( x11 & ~n9498 ) | ( x11 & n9499 ) | ( ~n9498 & n9499 ) ;
  assign n9917 = ( x11 & ~n9916 ) | ( x11 & 1'b0 ) | ( ~n9916 & 1'b0 ) ;
  assign n9918 = ( x11 & ~n9917 ) | ( x11 & n9493 ) | ( ~n9917 & n9493 ) ;
  assign n9919 = ( n9493 & ~x11 ) | ( n9493 & n9917 ) | ( ~x11 & n9917 ) ;
  assign n9920 = ( n9918 & ~n9493 ) | ( n9918 & n9919 ) | ( ~n9493 & n9919 ) ;
  assign n9921 = x11 &  n9499 ;
  assign n9922 = ~n9498 & n9921 ;
  assign n9923 = ( n9498 & ~n9921 ) | ( n9498 & 1'b0 ) | ( ~n9921 & 1'b0 ) ;
  assign n9924 = n9922 | n9923 ;
  assign n9958 = ~n3460 & n8429 ;
  assign n9955 = n3361 | n8764 ;
  assign n9956 = ~n3601 & n8105 ;
  assign n9957 = ( n9955 & ~n9956 ) | ( n9955 & 1'b0 ) | ( ~n9956 & 1'b0 ) ;
  assign n9959 = ( n3460 & n9958 ) | ( n3460 & n9957 ) | ( n9958 & n9957 ) ;
  assign n9960 = ( n8107 & ~n3603 ) | ( n8107 & n9510 ) | ( ~n3603 & n9510 ) ;
  assign n9961 = ( n9511 & n9959 ) | ( n9511 & n9960 ) | ( n9959 & n9960 ) ;
  assign n9962 = x8 | n9961 ;
  assign n9963 = ( x8 & ~n9961 ) | ( x8 & 1'b0 ) | ( ~n9961 & 1'b0 ) ;
  assign n9964 = ( n9962 & ~x8 ) | ( n9962 & n9963 ) | ( ~x8 & n9963 ) ;
  assign n9940 = ~n6886 & n8107 ;
  assign n9938 = ~n3460 & n8764 ;
  assign n9935 = ~n3547 & n8105 ;
  assign n9936 = n3601 | n8429 ;
  assign n9937 = ~n9935 & n9936 ;
  assign n9939 = ( n3460 & n9938 ) | ( n3460 & n9937 ) | ( n9938 & n9937 ) ;
  assign n9941 = ( n6886 & n9940 ) | ( n6886 & n9939 ) | ( n9940 & n9939 ) ;
  assign n9945 = n8107 &  n7412 ;
  assign n9942 = n3547 | n8429 ;
  assign n9943 = n3601 | n8764 ;
  assign n9944 = n9942 &  n9943 ;
  assign n9946 = ( n9945 & ~n7412 ) | ( n9945 & n9944 ) | ( ~n7412 & n9944 ) ;
  assign n9947 = x8 &  n9946 ;
  assign n9948 = x8 | n9946 ;
  assign n9949 = ~n9947 & n9948 ;
  assign n9950 = ( x8 & ~n9941 ) | ( x8 & n9949 ) | ( ~n9941 & n9949 ) ;
  assign n9951 = ~n3547 & n8103 ;
  assign n9952 = ( x8 & ~n9951 ) | ( x8 & 1'b0 ) | ( ~n9951 & 1'b0 ) ;
  assign n9953 = ( x8 & ~n9941 ) | ( x8 & n9952 ) | ( ~n9941 & n9952 ) ;
  assign n9954 = ~n9950 & n9953 ;
  assign n9965 = ( n9499 & ~n9964 ) | ( n9499 & n9954 ) | ( ~n9964 & n9954 ) ;
  assign n9925 = n3460 &  n8105 ;
  assign n9926 = n3325 | n8764 ;
  assign n9927 = n3361 | n8429 ;
  assign n9928 = n9926 &  n9927 ;
  assign n9929 = ( n9925 & ~n8105 ) | ( n9925 & n9928 ) | ( ~n8105 & n9928 ) ;
  assign n9930 = ( n6800 & ~n3604 ) | ( n6800 & n8107 ) | ( ~n3604 & n8107 ) ;
  assign n9931 = ( n6801 & n9929 ) | ( n6801 & n9930 ) | ( n9929 & n9930 ) ;
  assign n9932 = x8 &  n9931 ;
  assign n9933 = x8 | n9931 ;
  assign n9934 = ~n9932 & n9933 ;
  assign n9966 = ( n9924 & ~n9965 ) | ( n9924 & n9934 ) | ( ~n9965 & n9934 ) ;
  assign n9967 = ( n9915 & n9920 ) | ( n9915 & n9966 ) | ( n9920 & n9966 ) ;
  assign n9968 = ( n9895 & n9905 ) | ( n9895 & n9967 ) | ( n9905 & n9967 ) ;
  assign n9969 = ( n9890 & ~n9892 ) | ( n9890 & n9968 ) | ( ~n9892 & n9968 ) ;
  assign n9970 = ( n9870 & n9880 ) | ( n9870 & n9969 ) | ( n9880 & n9969 ) ;
  assign n9971 = ( n9857 & n9867 ) | ( n9857 & n9970 ) | ( n9867 & n9970 ) ;
  assign n9972 = ( n9855 & ~n9845 ) | ( n9855 & n9971 ) | ( ~n9845 & n9971 ) ;
  assign n9973 = ( n9840 & n9843 ) | ( n9840 & n9972 ) | ( n9843 & n9972 ) ;
  assign n9974 = ( n9823 & n9826 ) | ( n9823 & n9973 ) | ( n9826 & n9973 ) ;
  assign n9975 = ( n9810 & ~n9813 ) | ( n9810 & n9974 ) | ( ~n9813 & n9974 ) ;
  assign n9976 = ( n9786 & n9796 ) | ( n9786 & n9975 ) | ( n9796 & n9975 ) ;
  assign n9977 = ( n9774 & n9784 ) | ( n9774 & n9976 ) | ( n9784 & n9976 ) ;
  assign n9978 = ( n9772 & ~n9762 ) | ( n9772 & n9977 ) | ( ~n9762 & n9977 ) ;
  assign n9979 = ( n9757 & n9760 ) | ( n9757 & n9978 ) | ( n9760 & n9978 ) ;
  assign n9980 = ( n9744 & n9747 ) | ( n9744 & n9979 ) | ( n9747 & n9979 ) ;
  assign n9981 = ( n9731 & ~n9734 ) | ( n9731 & n9980 ) | ( ~n9734 & n9980 ) ;
  assign n9982 = ( n9711 & n9721 ) | ( n9711 & n9981 ) | ( n9721 & n9981 ) ;
  assign n9983 = ( n9699 & n9709 ) | ( n9699 & n9982 ) | ( n9709 & n9982 ) ;
  assign n9984 = ( n9697 & ~n9687 ) | ( n9697 & n9983 ) | ( ~n9687 & n9983 ) ;
  assign n9985 = ( n9682 & n9685 ) | ( n9682 & n9984 ) | ( n9685 & n9984 ) ;
  assign n9986 = ( n9669 & n9672 ) | ( n9669 & n9985 ) | ( n9672 & n9985 ) ;
  assign n9987 = ( n9659 & ~n9649 ) | ( n9659 & n9986 ) | ( ~n9649 & n9986 ) ;
  assign n9988 = ( n9647 & ~n9637 ) | ( n9647 & n9987 ) | ( ~n9637 & n9987 ) ;
  assign n9989 = ( n9624 & n9634 ) | ( n9624 & n9988 ) | ( n9634 & n9988 ) ;
  assign n9990 = ( n9611 & n9621 ) | ( n9611 & n9989 ) | ( n9621 & n9989 ) ;
  assign n9991 = ( n9608 & ~n9598 ) | ( n9608 & n9990 ) | ( ~n9598 & n9990 ) ;
  assign n9992 = ( n9585 & n9595 ) | ( n9585 & n9991 ) | ( n9595 & n9991 ) ;
  assign n9993 = ( n9572 & n9582 ) | ( n9572 & n9992 ) | ( n9582 & n9992 ) ;
  assign n9994 = ( n9545 & ~n9542 ) | ( n9545 & n9555 ) | ( ~n9542 & n9555 ) ;
  assign n9995 = ( n9542 & ~n9555 ) | ( n9542 & n9545 ) | ( ~n9555 & n9545 ) ;
  assign n9996 = ( n9994 & ~n9545 ) | ( n9994 & n9995 ) | ( ~n9545 & n9995 ) ;
  assign n10001 = ~n863 & n9160 ;
  assign n9997 = ~n9154 |  n9151 ;
  assign n9998 = n599 | n9997 ;
  assign n9999 = n702 | n9558 ;
  assign n10000 = n9998 &  n9999 ;
  assign n10002 = ( n863 & n10001 ) | ( n863 & n10000 ) | ( n10001 & n10000 ) ;
  assign n10003 = n4452 | n9155 ;
  assign n10004 = n10002 &  n10003 ;
  assign n10005 = x5 | n10004 ;
  assign n10006 = x5 &  n10004 ;
  assign n10007 = ( n10005 & ~n10006 ) | ( n10005 & 1'b0 ) | ( ~n10006 & 1'b0 ) ;
  assign n10008 = ( n9993 & ~n9996 ) | ( n9993 & n10007 ) | ( ~n9996 & n10007 ) ;
  assign n10009 = ( n9556 & n9565 ) | ( n9556 & n9568 ) | ( n9565 & n9568 ) ;
  assign n10010 = ( n9568 & ~n10009 ) | ( n9568 & n9569 ) | ( ~n10009 & n9569 ) ;
  assign n10014 = ( x0 & ~x1 ) | ( x0 & x2 ) | ( ~x1 & x2 ) ;
  assign n10015 = ~n10014 |  x0 ;
  assign n10016 = n599 | n10015 ;
  assign n10019 = ~n3635 & n702 ;
  assign n10011 = ( x1 & ~x2 ) | ( x1 & 1'b0 ) | ( ~x2 & 1'b0 ) ;
  assign n10012 = ~x1 & x2 ;
  assign n10013 = n10011 | n10012 ;
  assign n10017 = ~x0 | ~n10013 ;
  assign n10018 = n599 | n10017 ;
  assign n10020 = ( n702 & ~n10019 ) | ( n702 & n10018 ) | ( ~n10019 & n10018 ) ;
  assign n10021 = n10016 &  n10020 ;
  assign n10022 = x2 | n10021 ;
  assign n10023 = x2 &  n10021 ;
  assign n10024 = ( n10022 & ~n10023 ) | ( n10022 & 1'b0 ) | ( ~n10023 & 1'b0 ) ;
  assign n10028 = ~n946 & n9160 ;
  assign n10025 = n702 | n9997 ;
  assign n10026 = n863 | n9558 ;
  assign n10027 = n10025 &  n10026 ;
  assign n10029 = ( n946 & n10028 ) | ( n946 & n10027 ) | ( n10028 & n10027 ) ;
  assign n10030 = ( n9155 & ~n3650 ) | ( n9155 & n10029 ) | ( ~n3650 & n10029 ) ;
  assign n10031 = ~n9155 & n10030 ;
  assign n10032 = ( x5 & ~n10029 ) | ( x5 & n10031 ) | ( ~n10029 & n10031 ) ;
  assign n10033 = ( n10029 & ~x5 ) | ( n10029 & n10031 ) | ( ~x5 & n10031 ) ;
  assign n10034 = ( n10032 & ~n10031 ) | ( n10032 & n10033 ) | ( ~n10031 & n10033 ) ;
  assign n10035 = ( n9572 & ~n9582 ) | ( n9572 & n9992 ) | ( ~n9582 & n9992 ) ;
  assign n10036 = ( n9582 & ~n9993 ) | ( n9582 & n10035 ) | ( ~n9993 & n10035 ) ;
  assign n10037 = ( n10024 & n10034 ) | ( n10024 & n10036 ) | ( n10034 & n10036 ) ;
  assign n10038 = ( n9993 & n9996 ) | ( n9993 & n10007 ) | ( n9996 & n10007 ) ;
  assign n10039 = ( n9996 & ~n9993 ) | ( n9996 & n10007 ) | ( ~n9993 & n10007 ) ;
  assign n10040 = ( n9993 & ~n10038 ) | ( n9993 & n10039 ) | ( ~n10038 & n10039 ) ;
  assign n10041 = ( n10024 & ~n10034 ) | ( n10024 & n10036 ) | ( ~n10034 & n10036 ) ;
  assign n10042 = ( n10034 & ~n10037 ) | ( n10034 & n10041 ) | ( ~n10037 & n10041 ) ;
  assign n10046 = ~n946 & n9558 ;
  assign n10043 = n863 | n9997 ;
  assign n10044 = n1043 | n9160 ;
  assign n10045 = n10043 &  n10044 ;
  assign n10047 = ( n946 & n10046 ) | ( n946 & n10045 ) | ( n10046 & n10045 ) ;
  assign n10048 = ( n3911 & ~n3633 ) | ( n3911 & n9155 ) | ( ~n3633 & n9155 ) ;
  assign n10049 = ( n3913 & n10047 ) | ( n3913 & n10048 ) | ( n10047 & n10048 ) ;
  assign n10050 = x5 | n10049 ;
  assign n10051 = x5 &  n10049 ;
  assign n10052 = ( n10050 & ~n10051 ) | ( n10050 & 1'b0 ) | ( ~n10051 & 1'b0 ) ;
  assign n10053 = ( n9585 & ~n9595 ) | ( n9585 & n9991 ) | ( ~n9595 & n9991 ) ;
  assign n10054 = ( n9595 & ~n9992 ) | ( n9595 & n10053 ) | ( ~n9992 & n10053 ) ;
  assign n10058 = ~n946 & n9997 ;
  assign n10055 = n1151 | n9160 ;
  assign n10056 = n1043 | n9558 ;
  assign n10057 = n10055 &  n10056 ;
  assign n10059 = ( n946 & n10058 ) | ( n946 & n10057 ) | ( n10058 & n10057 ) ;
  assign n10060 = ( n4035 & ~n3632 ) | ( n4035 & n9155 ) | ( ~n3632 & n9155 ) ;
  assign n10061 = ( n4037 & n10059 ) | ( n4037 & n10060 ) | ( n10059 & n10060 ) ;
  assign n10062 = x5 | n10061 ;
  assign n10063 = x5 &  n10061 ;
  assign n10064 = ( n10062 & ~n10063 ) | ( n10062 & 1'b0 ) | ( ~n10063 & 1'b0 ) ;
  assign n10065 = ( n9598 & ~n9990 ) | ( n9598 & n9608 ) | ( ~n9990 & n9608 ) ;
  assign n10066 = ( n9991 & ~n9608 ) | ( n9991 & n10065 ) | ( ~n9608 & n10065 ) ;
  assign n10067 = n1043 | n9997 ;
  assign n10068 = n1151 | n9558 ;
  assign n10069 = n10067 &  n10068 ;
  assign n10070 = n1267 &  n9160 ;
  assign n10071 = ( n10069 & ~n1267 ) | ( n10069 & n10070 ) | ( ~n1267 & n10070 ) ;
  assign n10072 = ( n3949 & ~n3631 ) | ( n3949 & n9155 ) | ( ~n3631 & n9155 ) ;
  assign n10073 = ( n3951 & n10071 ) | ( n3951 & n10072 ) | ( n10071 & n10072 ) ;
  assign n10074 = x5 | n10073 ;
  assign n10075 = x5 &  n10073 ;
  assign n10076 = ( n10074 & ~n10075 ) | ( n10074 & 1'b0 ) | ( ~n10075 & 1'b0 ) ;
  assign n10077 = ( n9611 & ~n9621 ) | ( n9611 & n9989 ) | ( ~n9621 & n9989 ) ;
  assign n10078 = ( n9621 & ~n9990 ) | ( n9621 & n10077 ) | ( ~n9990 & n10077 ) ;
  assign n10084 = ( n3630 & ~n9155 ) | ( n3630 & n4058 ) | ( ~n9155 & n4058 ) ;
  assign n10079 = n1151 | n9997 ;
  assign n10080 = n1378 | n9160 ;
  assign n10081 = n10079 &  n10080 ;
  assign n10082 = n1267 &  n9558 ;
  assign n10083 = ( n10081 & ~n1267 ) | ( n10081 & n10082 ) | ( ~n1267 & n10082 ) ;
  assign n10085 = ( n4060 & ~n10084 ) | ( n4060 & n10083 ) | ( ~n10084 & n10083 ) ;
  assign n10086 = x5 | n10085 ;
  assign n10087 = x5 &  n10085 ;
  assign n10088 = ( n10086 & ~n10087 ) | ( n10086 & 1'b0 ) | ( ~n10087 & 1'b0 ) ;
  assign n10089 = ( n9624 & ~n9634 ) | ( n9624 & n9988 ) | ( ~n9634 & n9988 ) ;
  assign n10090 = ( n9634 & ~n9989 ) | ( n9634 & n10089 ) | ( ~n9989 & n10089 ) ;
  assign n10096 = ( n3629 & ~n9155 ) | ( n3629 & n4419 ) | ( ~n9155 & n4419 ) ;
  assign n10091 = ( n1483 & ~n9160 ) | ( n1483 & 1'b0 ) | ( ~n9160 & 1'b0 ) ;
  assign n10092 = n1378 | n9558 ;
  assign n10093 = ~n10091 & n10092 ;
  assign n10094 = n1267 &  n9997 ;
  assign n10095 = ( n10093 & ~n1267 ) | ( n10093 & n10094 ) | ( ~n1267 & n10094 ) ;
  assign n10097 = ( n4421 & ~n10096 ) | ( n4421 & n10095 ) | ( ~n10096 & n10095 ) ;
  assign n10098 = x5 | n10097 ;
  assign n10099 = x5 &  n10097 ;
  assign n10100 = ( n10098 & ~n10099 ) | ( n10098 & 1'b0 ) | ( ~n10099 & 1'b0 ) ;
  assign n10101 = ( n9637 & ~n9987 ) | ( n9637 & n9647 ) | ( ~n9987 & n9647 ) ;
  assign n10102 = ( n9988 & ~n9647 ) | ( n9988 & n10101 ) | ( ~n9647 & n10101 ) ;
  assign n10103 = n1378 | n9997 ;
  assign n10104 = n1566 | n9160 ;
  assign n10105 = n10103 &  n10104 ;
  assign n10106 = n1483 &  n9558 ;
  assign n10107 = ( n10105 & ~n1483 ) | ( n10105 & n10106 ) | ( ~n1483 & n10106 ) ;
  assign n10108 = ( n5038 & n9155 ) | ( n5038 & n10107 ) | ( n9155 & n10107 ) ;
  assign n10109 = ~n9155 & n10108 ;
  assign n10110 = ( x5 & ~n10107 ) | ( x5 & n10109 ) | ( ~n10107 & n10109 ) ;
  assign n10111 = ( n10107 & ~x5 ) | ( n10107 & n10109 ) | ( ~x5 & n10109 ) ;
  assign n10112 = ( n10110 & ~n10109 ) | ( n10110 & n10111 ) | ( ~n10109 & n10111 ) ;
  assign n10113 = ( n9649 & n9659 ) | ( n9649 & n9986 ) | ( n9659 & n9986 ) ;
  assign n10114 = ( n9649 & ~n9986 ) | ( n9649 & n9659 ) | ( ~n9986 & n9659 ) ;
  assign n10115 = ( n9986 & ~n10113 ) | ( n9986 & n10114 ) | ( ~n10113 & n10114 ) ;
  assign n10116 = ( n9669 & ~n9985 ) | ( n9669 & n9672 ) | ( ~n9985 & n9672 ) ;
  assign n10117 = ( n9672 & ~n9669 ) | ( n9672 & n9985 ) | ( ~n9669 & n9985 ) ;
  assign n10118 = ( n10116 & ~n9672 ) | ( n10116 & n10117 ) | ( ~n9672 & n10117 ) ;
  assign n10124 = ( n3627 & ~n9155 ) | ( n3627 & n4271 ) | ( ~n9155 & n4271 ) ;
  assign n10119 = n1671 | n9160 ;
  assign n10120 = n1566 | n9558 ;
  assign n10121 = n10119 &  n10120 ;
  assign n10122 = n1483 &  n9997 ;
  assign n10123 = ( n10121 & ~n1483 ) | ( n10121 & n10122 ) | ( ~n1483 & n10122 ) ;
  assign n10125 = ( n4273 & ~n10124 ) | ( n4273 & n10123 ) | ( ~n10124 & n10123 ) ;
  assign n10126 = x5 &  n10125 ;
  assign n10127 = x5 | n10125 ;
  assign n10128 = ~n10126 & n10127 ;
  assign n10129 = ( n9685 & ~n9682 ) | ( n9685 & n9984 ) | ( ~n9682 & n9984 ) ;
  assign n10130 = ( n9682 & ~n9984 ) | ( n9682 & n9685 ) | ( ~n9984 & n9685 ) ;
  assign n10131 = ( n10129 & ~n9685 ) | ( n10129 & n10130 ) | ( ~n9685 & n10130 ) ;
  assign n10135 = ~n1566 & n9997 ;
  assign n10132 = n1748 | n9160 ;
  assign n10133 = n1671 | n9558 ;
  assign n10134 = n10132 &  n10133 ;
  assign n10136 = ( n1566 & n10135 ) | ( n1566 & n10134 ) | ( n10135 & n10134 ) ;
  assign n10137 = ( n4594 & ~n3626 ) | ( n4594 & n9155 ) | ( ~n3626 & n9155 ) ;
  assign n10138 = ( n4596 & n10136 ) | ( n4596 & n10137 ) | ( n10136 & n10137 ) ;
  assign n10139 = x5 &  n10138 ;
  assign n10140 = x5 | n10138 ;
  assign n10141 = ~n10139 & n10140 ;
  assign n10145 = ~n1875 & n9160 ;
  assign n10142 = n1671 | n9997 ;
  assign n10143 = n1748 | n9558 ;
  assign n10144 = n10142 &  n10143 ;
  assign n10146 = ( n1875 & n10145 ) | ( n1875 & n10144 ) | ( n10145 & n10144 ) ;
  assign n10147 = ( n9155 & ~n4580 ) | ( n9155 & n10146 ) | ( ~n4580 & n10146 ) ;
  assign n10148 = ~n9155 & n10147 ;
  assign n10149 = ( x5 & ~n10146 ) | ( x5 & n10148 ) | ( ~n10146 & n10148 ) ;
  assign n10150 = ( n10146 & ~x5 ) | ( n10146 & n10148 ) | ( ~x5 & n10148 ) ;
  assign n10151 = ( n10149 & ~n10148 ) | ( n10149 & n10150 ) | ( ~n10148 & n10150 ) ;
  assign n10152 = ( n9687 & n9697 ) | ( n9687 & n9983 ) | ( n9697 & n9983 ) ;
  assign n10153 = ( n9687 & ~n9983 ) | ( n9687 & n9697 ) | ( ~n9983 & n9697 ) ;
  assign n10154 = ( n9983 & ~n10152 ) | ( n9983 & n10153 ) | ( ~n10152 & n10153 ) ;
  assign n10155 = ~n1748 & n9997 ;
  assign n10156 = n1940 | n9160 ;
  assign n10157 = n1875 | n9558 ;
  assign n10158 = n10156 &  n10157 ;
  assign n10159 = ( n1748 & n10155 ) | ( n1748 & n10158 ) | ( n10155 & n10158 ) ;
  assign n10160 = ( n9155 & ~n4743 ) | ( n9155 & n10159 ) | ( ~n4743 & n10159 ) ;
  assign n10161 = ~n9155 & n10160 ;
  assign n10162 = ( x5 & ~n10159 ) | ( x5 & n10161 ) | ( ~n10159 & n10161 ) ;
  assign n10163 = ( n10159 & ~x5 ) | ( n10159 & n10161 ) | ( ~x5 & n10161 ) ;
  assign n10164 = ( n10162 & ~n10161 ) | ( n10162 & n10163 ) | ( ~n10161 & n10163 ) ;
  assign n10165 = ( n9709 & ~n9699 ) | ( n9709 & n9982 ) | ( ~n9699 & n9982 ) ;
  assign n10166 = ( n9699 & ~n9709 ) | ( n9699 & n9982 ) | ( ~n9709 & n9982 ) ;
  assign n10167 = ( n10165 & ~n9982 ) | ( n10165 & n10166 ) | ( ~n9982 & n10166 ) ;
  assign n10171 = ~n1875 & n9997 ;
  assign n10168 = n2022 | n9160 ;
  assign n10169 = n1940 | n9558 ;
  assign n10170 = n10168 &  n10169 ;
  assign n10172 = ( n1875 & n10171 ) | ( n1875 & n10170 ) | ( n10171 & n10170 ) ;
  assign n10173 = ( n9155 & ~n5381 ) | ( n9155 & n10172 ) | ( ~n5381 & n10172 ) ;
  assign n10174 = ~n9155 & n10173 ;
  assign n10175 = ( x5 & ~n10172 ) | ( x5 & n10174 ) | ( ~n10172 & n10174 ) ;
  assign n10176 = ( n10172 & ~x5 ) | ( n10172 & n10174 ) | ( ~x5 & n10174 ) ;
  assign n10177 = ( n10175 & ~n10174 ) | ( n10175 & n10176 ) | ( ~n10174 & n10176 ) ;
  assign n10178 = ( n9721 & ~n9711 ) | ( n9721 & n9981 ) | ( ~n9711 & n9981 ) ;
  assign n10179 = ( n9711 & ~n9721 ) | ( n9711 & n9981 ) | ( ~n9721 & n9981 ) ;
  assign n10180 = ( n10178 & ~n9981 ) | ( n10178 & n10179 ) | ( ~n9981 & n10179 ) ;
  assign n10184 = n2127 | n9160 ;
  assign n10185 = n2022 | n9558 ;
  assign n10186 = n10184 &  n10185 ;
  assign n10187 = ~n1940 & n9997 ;
  assign n10188 = ( n1940 & n10186 ) | ( n1940 & n10187 ) | ( n10186 & n10187 ) ;
  assign n10189 = ( n5085 & ~n3622 ) | ( n5085 & n9155 ) | ( ~n3622 & n9155 ) ;
  assign n10190 = ( n5086 & n10188 ) | ( n5086 & n10189 ) | ( n10188 & n10189 ) ;
  assign n10191 = x5 &  n10190 ;
  assign n10192 = x5 | n10190 ;
  assign n10193 = ~n10191 & n10192 ;
  assign n10181 = ( n9734 & ~n9731 ) | ( n9734 & n9980 ) | ( ~n9731 & n9980 ) ;
  assign n10182 = ( n9731 & ~n9980 ) | ( n9731 & n9734 ) | ( ~n9980 & n9734 ) ;
  assign n10183 = ( n10181 & ~n9734 ) | ( n10181 & n10182 ) | ( ~n9734 & n10182 ) ;
  assign n10194 = ( n9747 & ~n9744 ) | ( n9747 & n9979 ) | ( ~n9744 & n9979 ) ;
  assign n10195 = ( n9744 & ~n9979 ) | ( n9744 & n9747 ) | ( ~n9979 & n9747 ) ;
  assign n10196 = ( n10194 & ~n9747 ) | ( n10194 & n10195 ) | ( ~n9747 & n10195 ) ;
  assign n10197 = n2178 | n9160 ;
  assign n10198 = n2127 | n9558 ;
  assign n10199 = n10197 &  n10198 ;
  assign n10200 = ~n2022 & n9997 ;
  assign n10201 = ( n2022 & n10199 ) | ( n2022 & n10200 ) | ( n10199 & n10200 ) ;
  assign n10202 = ( n4931 & ~n3621 ) | ( n4931 & n9155 ) | ( ~n3621 & n9155 ) ;
  assign n10203 = ( n4933 & n10201 ) | ( n4933 & n10202 ) | ( n10201 & n10202 ) ;
  assign n10204 = x5 &  n10203 ;
  assign n10205 = x5 | n10203 ;
  assign n10206 = ~n10204 & n10205 ;
  assign n10207 = ( n9760 & ~n9757 ) | ( n9760 & n9978 ) | ( ~n9757 & n9978 ) ;
  assign n10208 = ( n9757 & ~n9978 ) | ( n9757 & n9760 ) | ( ~n9978 & n9760 ) ;
  assign n10209 = ( n10207 & ~n9760 ) | ( n10207 & n10208 ) | ( ~n9760 & n10208 ) ;
  assign n10213 = ~n2296 & n9160 ;
  assign n10210 = n2127 | n9997 ;
  assign n10211 = n2178 | n9558 ;
  assign n10212 = n10210 &  n10211 ;
  assign n10214 = ( n2296 & n10213 ) | ( n2296 & n10212 ) | ( n10213 & n10212 ) ;
  assign n10215 = ( n5280 & ~n3620 ) | ( n5280 & n9155 ) | ( ~n3620 & n9155 ) ;
  assign n10216 = ( n5282 & n10214 ) | ( n5282 & n10215 ) | ( n10214 & n10215 ) ;
  assign n10217 = x5 &  n10216 ;
  assign n10218 = x5 | n10216 ;
  assign n10219 = ~n10217 & n10218 ;
  assign n10223 = ~n2178 & n9997 ;
  assign n10220 = n2392 | n9160 ;
  assign n10221 = n2296 | n9558 ;
  assign n10222 = n10220 &  n10221 ;
  assign n10224 = ( n2178 & n10223 ) | ( n2178 & n10222 ) | ( n10223 & n10222 ) ;
  assign n10225 = ( n9155 & ~n5269 ) | ( n9155 & n10224 ) | ( ~n5269 & n10224 ) ;
  assign n10226 = ~n9155 & n10225 ;
  assign n10227 = ( x5 & ~n10224 ) | ( x5 & n10226 ) | ( ~n10224 & n10226 ) ;
  assign n10228 = ( n10224 & ~x5 ) | ( n10224 & n10226 ) | ( ~x5 & n10226 ) ;
  assign n10229 = ( n10227 & ~n10226 ) | ( n10227 & n10228 ) | ( ~n10226 & n10228 ) ;
  assign n10230 = ( n9762 & n9772 ) | ( n9762 & n9977 ) | ( n9772 & n9977 ) ;
  assign n10231 = ( n9762 & ~n9977 ) | ( n9762 & n9772 ) | ( ~n9977 & n9772 ) ;
  assign n10232 = ( n9977 & ~n10230 ) | ( n9977 & n10231 ) | ( ~n10230 & n10231 ) ;
  assign n10236 = ~n2296 & n9997 ;
  assign n10233 = n2483 | n9160 ;
  assign n10234 = n2392 | n9558 ;
  assign n10235 = n10233 &  n10234 ;
  assign n10237 = ( n2296 & n10236 ) | ( n2296 & n10235 ) | ( n10236 & n10235 ) ;
  assign n10238 = ( n9155 & ~n5500 ) | ( n9155 & n10237 ) | ( ~n5500 & n10237 ) ;
  assign n10239 = ~n9155 & n10238 ;
  assign n10240 = ( x5 & ~n10237 ) | ( x5 & n10239 ) | ( ~n10237 & n10239 ) ;
  assign n10241 = ( n10237 & ~x5 ) | ( n10237 & n10239 ) | ( ~x5 & n10239 ) ;
  assign n10242 = ( n10240 & ~n10239 ) | ( n10240 & n10241 ) | ( ~n10239 & n10241 ) ;
  assign n10243 = ( n9784 & ~n9774 ) | ( n9784 & n9976 ) | ( ~n9774 & n9976 ) ;
  assign n10244 = ( n9774 & ~n9784 ) | ( n9774 & n9976 ) | ( ~n9784 & n9976 ) ;
  assign n10245 = ( n10243 & ~n9976 ) | ( n10243 & n10244 ) | ( ~n9976 & n10244 ) ;
  assign n10249 = ~n2392 & n9997 ;
  assign n10246 = n2569 | n9160 ;
  assign n10247 = n2483 | n9558 ;
  assign n10248 = n10246 &  n10247 ;
  assign n10250 = ( n2392 & n10249 ) | ( n2392 & n10248 ) | ( n10249 & n10248 ) ;
  assign n10251 = ( n9155 & ~n6212 ) | ( n9155 & n10250 ) | ( ~n6212 & n10250 ) ;
  assign n10252 = ~n9155 & n10251 ;
  assign n10253 = ( x5 & ~n10250 ) | ( x5 & n10252 ) | ( ~n10250 & n10252 ) ;
  assign n10254 = ( n10250 & ~x5 ) | ( n10250 & n10252 ) | ( ~x5 & n10252 ) ;
  assign n10255 = ( n10253 & ~n10252 ) | ( n10253 & n10254 ) | ( ~n10252 & n10254 ) ;
  assign n10256 = ( n9796 & ~n9786 ) | ( n9796 & n9975 ) | ( ~n9786 & n9975 ) ;
  assign n10257 = ( n9786 & ~n9796 ) | ( n9786 & n9975 ) | ( ~n9796 & n9975 ) ;
  assign n10258 = ( n10256 & ~n9975 ) | ( n10256 & n10257 ) | ( ~n9975 & n10257 ) ;
  assign n10265 = ~n2665 & n9160 ;
  assign n10262 = n2483 | n9997 ;
  assign n10263 = n2569 | n9558 ;
  assign n10264 = n10262 &  n10263 ;
  assign n10266 = ( n2665 & n10265 ) | ( n2665 & n10264 ) | ( n10265 & n10264 ) ;
  assign n10267 = ( n5886 & ~n3616 ) | ( n5886 & n9155 ) | ( ~n3616 & n9155 ) ;
  assign n10268 = ( n5887 & n10266 ) | ( n5887 & n10267 ) | ( n10266 & n10267 ) ;
  assign n10269 = x5 &  n10268 ;
  assign n10270 = x5 | n10268 ;
  assign n10271 = ~n10269 & n10270 ;
  assign n10259 = ( n9813 & ~n9810 ) | ( n9813 & n9974 ) | ( ~n9810 & n9974 ) ;
  assign n10260 = ( n9810 & ~n9974 ) | ( n9810 & n9813 ) | ( ~n9974 & n9813 ) ;
  assign n10261 = ( n10259 & ~n9813 ) | ( n10259 & n10260 ) | ( ~n9813 & n10260 ) ;
  assign n10272 = ( n9823 & ~n9826 ) | ( n9823 & n9973 ) | ( ~n9826 & n9973 ) ;
  assign n10273 = ( n9826 & ~n9974 ) | ( n9826 & n10272 ) | ( ~n9974 & n10272 ) ;
  assign n10277 = ~n2751 & n9160 ;
  assign n10274 = n2569 | n9997 ;
  assign n10275 = n2665 | n9558 ;
  assign n10276 = n10274 &  n10275 ;
  assign n10278 = ( n2751 & n10277 ) | ( n2751 & n10276 ) | ( n10277 & n10276 ) ;
  assign n10279 = ( n5702 & ~n3615 ) | ( n5702 & n9155 ) | ( ~n3615 & n9155 ) ;
  assign n10280 = ( n5704 & n10278 ) | ( n5704 & n10279 ) | ( n10278 & n10279 ) ;
  assign n10281 = x5 &  n10280 ;
  assign n10282 = x5 | n10280 ;
  assign n10283 = ~n10281 & n10282 ;
  assign n10284 = ( n9840 & ~n9843 ) | ( n9840 & n9972 ) | ( ~n9843 & n9972 ) ;
  assign n10285 = ( n9843 & ~n9973 ) | ( n9843 & n10284 ) | ( ~n9973 & n10284 ) ;
  assign n10289 = ~n2751 & n9558 ;
  assign n10286 = n2665 | n9997 ;
  assign n10287 = n2783 | n9160 ;
  assign n10288 = n10286 &  n10287 ;
  assign n10290 = ( n2751 & n10289 ) | ( n2751 & n10288 ) | ( n10289 & n10288 ) ;
  assign n10291 = ( n6116 & ~n3614 ) | ( n6116 & n9155 ) | ( ~n3614 & n9155 ) ;
  assign n10292 = ( n6118 & n10290 ) | ( n6118 & n10291 ) | ( n10290 & n10291 ) ;
  assign n10293 = x5 &  n10292 ;
  assign n10294 = x5 | n10292 ;
  assign n10295 = ~n10293 & n10294 ;
  assign n10296 = n2751 | n9997 ;
  assign n10297 = n2783 | n9558 ;
  assign n10298 = n10296 &  n10297 ;
  assign n10299 = n2910 &  n9160 ;
  assign n10300 = ( n10298 & ~n2910 ) | ( n10298 & n10299 ) | ( ~n2910 & n10299 ) ;
  assign n10301 = ( n9155 & ~n6226 ) | ( n9155 & n10300 ) | ( ~n6226 & n10300 ) ;
  assign n10302 = ~n9155 & n10301 ;
  assign n10303 = ( x5 & ~n10300 ) | ( x5 & n10302 ) | ( ~n10300 & n10302 ) ;
  assign n10304 = ( n10300 & ~x5 ) | ( n10300 & n10302 ) | ( ~x5 & n10302 ) ;
  assign n10305 = ( n10303 & ~n10302 ) | ( n10303 & n10304 ) | ( ~n10302 & n10304 ) ;
  assign n10306 = ( n9845 & n9855 ) | ( n9845 & n9971 ) | ( n9855 & n9971 ) ;
  assign n10307 = ( n9845 & ~n9971 ) | ( n9845 & n9855 ) | ( ~n9971 & n9855 ) ;
  assign n10308 = ( n9971 & ~n10306 ) | ( n9971 & n10307 ) | ( ~n10306 & n10307 ) ;
  assign n10309 = n2783 | n9997 ;
  assign n10310 = n2839 | n9160 ;
  assign n10311 = n10309 &  n10310 ;
  assign n10312 = n2910 &  n9558 ;
  assign n10313 = ( n10311 & ~n2910 ) | ( n10311 & n10312 ) | ( ~n2910 & n10312 ) ;
  assign n10314 = ( n6104 & ~n9155 ) | ( n6104 & 1'b0 ) | ( ~n9155 & 1'b0 ) ;
  assign n10315 = ( n10313 & ~n10314 ) | ( n10313 & 1'b0 ) | ( ~n10314 & 1'b0 ) ;
  assign n10316 = x5 &  n10315 ;
  assign n10317 = x5 | n10315 ;
  assign n10318 = ~n10316 & n10317 ;
  assign n10319 = ( n9867 & ~n9857 ) | ( n9867 & n9970 ) | ( ~n9857 & n9970 ) ;
  assign n10320 = ( n9857 & ~n9867 ) | ( n9857 & n9970 ) | ( ~n9867 & n9970 ) ;
  assign n10321 = ( n10319 & ~n9970 ) | ( n10319 & n10320 ) | ( ~n9970 & n10320 ) ;
  assign n10322 = n2995 | n9160 ;
  assign n10323 = n2839 | n9558 ;
  assign n10324 = n10322 &  n10323 ;
  assign n10325 = n2910 &  n9997 ;
  assign n10326 = ( n10324 & ~n2910 ) | ( n10324 & n10325 ) | ( ~n2910 & n10325 ) ;
  assign n10327 = ( n6330 & n9155 ) | ( n6330 & n10326 ) | ( n9155 & n10326 ) ;
  assign n10328 = ~n9155 & n10327 ;
  assign n10329 = ( x5 & ~n10326 ) | ( x5 & n10328 ) | ( ~n10326 & n10328 ) ;
  assign n10330 = ( n10326 & ~x5 ) | ( n10326 & n10328 ) | ( ~x5 & n10328 ) ;
  assign n10331 = ( n10329 & ~n10328 ) | ( n10329 & n10330 ) | ( ~n10328 & n10330 ) ;
  assign n10332 = ( n9880 & ~n9870 ) | ( n9880 & n9969 ) | ( ~n9870 & n9969 ) ;
  assign n10333 = ( n9870 & ~n9880 ) | ( n9870 & n9969 ) | ( ~n9880 & n9969 ) ;
  assign n10334 = ( n10332 & ~n9969 ) | ( n10332 & n10333 ) | ( ~n9969 & n10333 ) ;
  assign n10341 = ~n2839 & n9997 ;
  assign n10338 = n3030 | n9160 ;
  assign n10339 = n2995 | n9558 ;
  assign n10340 = n10338 &  n10339 ;
  assign n10342 = ( n2839 & n10341 ) | ( n2839 & n10340 ) | ( n10341 & n10340 ) ;
  assign n10343 = ( n6591 & ~n3610 ) | ( n6591 & n9155 ) | ( ~n3610 & n9155 ) ;
  assign n10344 = ( n6592 & n10342 ) | ( n6592 & n10343 ) | ( n10342 & n10343 ) ;
  assign n10345 = x5 &  n10344 ;
  assign n10346 = x5 | n10344 ;
  assign n10347 = ~n10345 & n10346 ;
  assign n10335 = ( n9892 & ~n9890 ) | ( n9892 & n9968 ) | ( ~n9890 & n9968 ) ;
  assign n10336 = ( n9890 & ~n9968 ) | ( n9890 & n9892 ) | ( ~n9968 & n9892 ) ;
  assign n10337 = ( n10335 & ~n9892 ) | ( n10335 & n10336 ) | ( ~n9892 & n10336 ) ;
  assign n10348 = ( n9905 & ~n9895 ) | ( n9905 & n9967 ) | ( ~n9895 & n9967 ) ;
  assign n10349 = ( n9895 & ~n9967 ) | ( n9895 & n9905 ) | ( ~n9967 & n9905 ) ;
  assign n10350 = ( n10348 & ~n9905 ) | ( n10348 & n10349 ) | ( ~n9905 & n10349 ) ;
  assign n10351 = n3106 | n9160 ;
  assign n10352 = n3030 | n9558 ;
  assign n10353 = n10351 &  n10352 ;
  assign n10354 = ~n2995 & n9997 ;
  assign n10355 = ( n2995 & n10353 ) | ( n2995 & n10354 ) | ( n10353 & n10354 ) ;
  assign n10356 = ( n6604 & ~n3609 ) | ( n6604 & n9155 ) | ( ~n3609 & n9155 ) ;
  assign n10357 = ( n6605 & n10355 ) | ( n6605 & n10356 ) | ( n10355 & n10356 ) ;
  assign n10358 = x5 &  n10357 ;
  assign n10359 = x5 | n10357 ;
  assign n10360 = ~n10358 & n10359 ;
  assign n10361 = ( n9915 & ~n9920 ) | ( n9915 & n9966 ) | ( ~n9920 & n9966 ) ;
  assign n10362 = ( n9920 & ~n9967 ) | ( n9920 & n10361 ) | ( ~n9967 & n10361 ) ;
  assign n10366 = ~n3030 & n9997 ;
  assign n10363 = n3197 | n9160 ;
  assign n10364 = n3106 | n9558 ;
  assign n10365 = n10363 &  n10364 ;
  assign n10367 = ( n3030 & n10366 ) | ( n3030 & n10365 ) | ( n10366 & n10365 ) ;
  assign n10368 = ( n6311 & ~n3608 ) | ( n6311 & n9155 ) | ( ~n3608 & n9155 ) ;
  assign n10369 = ( n6313 & n10367 ) | ( n6313 & n10368 ) | ( n10367 & n10368 ) ;
  assign n10370 = x5 &  n10369 ;
  assign n10371 = x5 | n10369 ;
  assign n10372 = ~n10370 & n10371 ;
  assign n10373 = n3106 | n9997 ;
  assign n10374 = n3197 | n9558 ;
  assign n10375 = n10373 &  n10374 ;
  assign n10376 = n3266 &  n9160 ;
  assign n10377 = ( n10375 & ~n3266 ) | ( n10375 & n10376 ) | ( ~n3266 & n10376 ) ;
  assign n10378 = ( n9155 & ~n7363 ) | ( n9155 & n10377 ) | ( ~n7363 & n10377 ) ;
  assign n10379 = ~n9155 & n10378 ;
  assign n10380 = ( x5 & ~n10377 ) | ( x5 & n10379 ) | ( ~n10377 & n10379 ) ;
  assign n10381 = ( n10377 & ~x5 ) | ( n10377 & n10379 ) | ( ~x5 & n10379 ) ;
  assign n10382 = ( n10380 & ~n10379 ) | ( n10380 & n10381 ) | ( ~n10379 & n10381 ) ;
  assign n10383 = ( n9924 & ~n9934 ) | ( n9924 & n9965 ) | ( ~n9934 & n9965 ) ;
  assign n10384 = ( n9934 & ~n9924 ) | ( n9934 & n9965 ) | ( ~n9924 & n9965 ) ;
  assign n10385 = ( n10383 & ~n9965 ) | ( n10383 & n10384 ) | ( ~n9965 & n10384 ) ;
  assign n10387 = ( n9499 & n9954 ) | ( n9499 & n9964 ) | ( n9954 & n9964 ) ;
  assign n10386 = ( n9499 & ~n9954 ) | ( n9499 & n9964 ) | ( ~n9954 & n9964 ) ;
  assign n10388 = ( n9954 & ~n10387 ) | ( n9954 & n10386 ) | ( ~n10387 & n10386 ) ;
  assign n10389 = n3197 | n9997 ;
  assign n10390 = n3325 | n9160 ;
  assign n10391 = n10389 &  n10390 ;
  assign n10392 = n3266 &  n9558 ;
  assign n10393 = ( n10391 & ~n3266 ) | ( n10391 & n10392 ) | ( ~n3266 & n10392 ) ;
  assign n10394 = n7377 &  n9155 ;
  assign n10395 = ( n10393 & ~n7377 ) | ( n10393 & n10394 ) | ( ~n7377 & n10394 ) ;
  assign n10396 = x5 &  n10395 ;
  assign n10397 = x5 | n10395 ;
  assign n10398 = ~n10396 & n10397 ;
  assign n10404 = ( n3605 & ~n9155 ) | ( n3605 & n6753 ) | ( ~n9155 & n6753 ) ;
  assign n10399 = n3361 | n9160 ;
  assign n10400 = n3325 | n9558 ;
  assign n10401 = n10399 &  n10400 ;
  assign n10402 = n3266 &  n9997 ;
  assign n10403 = ( n10401 & ~n3266 ) | ( n10401 & n10402 ) | ( ~n3266 & n10402 ) ;
  assign n10405 = ( n6754 & ~n10404 ) | ( n6754 & n10403 ) | ( ~n10404 & n10403 ) ;
  assign n10406 = x5 | n10405 ;
  assign n10407 = x5 &  n10405 ;
  assign n10408 = ( n10406 & ~n10407 ) | ( n10406 & 1'b0 ) | ( ~n10407 & 1'b0 ) ;
  assign n10409 = ~n9949 & n9952 ;
  assign n10410 = ( x8 & ~n10409 ) | ( x8 & n9941 ) | ( ~n10409 & n9941 ) ;
  assign n10411 = ( n9941 & ~x8 ) | ( n9941 & n10409 ) | ( ~x8 & n10409 ) ;
  assign n10412 = ( n10410 & ~n9941 ) | ( n10410 & n10411 ) | ( ~n9941 & n10411 ) ;
  assign n10413 = ( n9949 & ~n9952 ) | ( n9949 & 1'b0 ) | ( ~n9952 & 1'b0 ) ;
  assign n10414 = n10409 | n10413 ;
  assign n10445 = ~n3460 & n9558 ;
  assign n10442 = n3361 | n9997 ;
  assign n10443 = n3601 | n9160 ;
  assign n10444 = n10442 &  n10443 ;
  assign n10446 = ( n3460 & n10445 ) | ( n3460 & n10444 ) | ( n10445 & n10444 ) ;
  assign n10447 = ( n9155 & ~n6895 ) | ( n9155 & n10446 ) | ( ~n6895 & n10446 ) ;
  assign n10448 = ~n9155 & n10447 ;
  assign n10449 = ( x5 & ~n10446 ) | ( x5 & n10448 ) | ( ~n10446 & n10448 ) ;
  assign n10450 = ( n10446 & ~x5 ) | ( n10446 & n10448 ) | ( ~x5 & n10448 ) ;
  assign n10451 = ( n10449 & ~n10448 ) | ( n10449 & n10450 ) | ( ~n10448 & n10450 ) ;
  assign n10435 = n9155 &  n7412 ;
  assign n10432 = n3547 | n9558 ;
  assign n10433 = n3601 | n9997 ;
  assign n10434 = n10432 &  n10433 ;
  assign n10436 = ( n10435 & ~n7412 ) | ( n10435 & n10434 ) | ( ~n7412 & n10434 ) ;
  assign n10430 = ~n6886 & n9155 ;
  assign n10428 = ~n3460 & n9997 ;
  assign n10425 = n3547 | n9160 ;
  assign n10426 = n3601 | n9558 ;
  assign n10427 = n10425 &  n10426 ;
  assign n10429 = ( n3460 & n10428 ) | ( n3460 & n10427 ) | ( n10428 & n10427 ) ;
  assign n10431 = ( n6886 & n10430 ) | ( n6886 & n10429 ) | ( n10430 & n10429 ) ;
  assign n10437 = ~n3547 & n9154 ;
  assign n10439 = ( n10436 & ~n10431 ) | ( n10436 & n10437 ) | ( ~n10431 & n10437 ) ;
  assign n10440 = ( x5 & ~n10436 ) | ( x5 & n10439 ) | ( ~n10436 & n10439 ) ;
  assign n10441 = ( x5 & ~n10440 ) | ( x5 & 1'b0 ) | ( ~n10440 & 1'b0 ) ;
  assign n10452 = ( n9951 & ~n10451 ) | ( n9951 & n10441 ) | ( ~n10451 & n10441 ) ;
  assign n10418 = ~n3460 & n9160 ;
  assign n10415 = n3325 | n9997 ;
  assign n10416 = n3361 | n9558 ;
  assign n10417 = n10415 &  n10416 ;
  assign n10419 = ( n3460 & n10418 ) | ( n3460 & n10417 ) | ( n10418 & n10417 ) ;
  assign n10420 = ( n9155 & ~n7405 ) | ( n9155 & n10419 ) | ( ~n7405 & n10419 ) ;
  assign n10421 = ~n9155 & n10420 ;
  assign n10422 = ( x5 & ~n10419 ) | ( x5 & n10421 ) | ( ~n10419 & n10421 ) ;
  assign n10423 = ( n10419 & ~x5 ) | ( n10419 & n10421 ) | ( ~x5 & n10421 ) ;
  assign n10424 = ( n10422 & ~n10421 ) | ( n10422 & n10423 ) | ( ~n10421 & n10423 ) ;
  assign n10453 = ( n10414 & ~n10452 ) | ( n10414 & n10424 ) | ( ~n10452 & n10424 ) ;
  assign n10454 = ( n10408 & n10412 ) | ( n10408 & n10453 ) | ( n10412 & n10453 ) ;
  assign n10455 = ( n10388 & n10398 ) | ( n10388 & n10454 ) | ( n10398 & n10454 ) ;
  assign n10456 = ( n10382 & ~n10385 ) | ( n10382 & n10455 ) | ( ~n10385 & n10455 ) ;
  assign n10457 = ( n10362 & n10372 ) | ( n10362 & n10456 ) | ( n10372 & n10456 ) ;
  assign n10458 = ( n10350 & n10360 ) | ( n10350 & n10457 ) | ( n10360 & n10457 ) ;
  assign n10459 = ( n10347 & ~n10337 ) | ( n10347 & n10458 ) | ( ~n10337 & n10458 ) ;
  assign n10460 = ( n10331 & n10334 ) | ( n10331 & n10459 ) | ( n10334 & n10459 ) ;
  assign n10461 = ( n10318 & n10321 ) | ( n10318 & n10460 ) | ( n10321 & n10460 ) ;
  assign n10462 = ( n10305 & ~n10308 ) | ( n10305 & n10461 ) | ( ~n10308 & n10461 ) ;
  assign n10463 = ( n10285 & n10295 ) | ( n10285 & n10462 ) | ( n10295 & n10462 ) ;
  assign n10464 = ( n10273 & n10283 ) | ( n10273 & n10463 ) | ( n10283 & n10463 ) ;
  assign n10465 = ( n10271 & ~n10261 ) | ( n10271 & n10464 ) | ( ~n10261 & n10464 ) ;
  assign n10466 = ( n10255 & n10258 ) | ( n10255 & n10465 ) | ( n10258 & n10465 ) ;
  assign n10467 = ( n10242 & n10245 ) | ( n10242 & n10466 ) | ( n10245 & n10466 ) ;
  assign n10468 = ( n10229 & ~n10232 ) | ( n10229 & n10467 ) | ( ~n10232 & n10467 ) ;
  assign n10469 = ( n10209 & n10219 ) | ( n10209 & n10468 ) | ( n10219 & n10468 ) ;
  assign n10470 = ( n10196 & n10206 ) | ( n10196 & n10469 ) | ( n10206 & n10469 ) ;
  assign n10471 = ( n10193 & ~n10183 ) | ( n10193 & n10470 ) | ( ~n10183 & n10470 ) ;
  assign n10472 = ( n10177 & n10180 ) | ( n10177 & n10471 ) | ( n10180 & n10471 ) ;
  assign n10473 = ( n10164 & n10167 ) | ( n10164 & n10472 ) | ( n10167 & n10472 ) ;
  assign n10474 = ( n10151 & ~n10154 ) | ( n10151 & n10473 ) | ( ~n10154 & n10473 ) ;
  assign n10475 = ( n10131 & n10141 ) | ( n10131 & n10474 ) | ( n10141 & n10474 ) ;
  assign n10476 = ( n10118 & n10128 ) | ( n10118 & n10475 ) | ( n10128 & n10475 ) ;
  assign n10477 = ( n10112 & ~n10115 ) | ( n10112 & n10476 ) | ( ~n10115 & n10476 ) ;
  assign n10478 = ( n10100 & ~n10102 ) | ( n10100 & n10477 ) | ( ~n10102 & n10477 ) ;
  assign n10479 = ( n10088 & n10090 ) | ( n10088 & n10478 ) | ( n10090 & n10478 ) ;
  assign n10480 = ( n10076 & n10078 ) | ( n10076 & n10479 ) | ( n10078 & n10479 ) ;
  assign n10481 = ( n10064 & ~n10066 ) | ( n10064 & n10480 ) | ( ~n10066 & n10480 ) ;
  assign n10482 = ( n10052 & n10054 ) | ( n10052 & n10481 ) | ( n10054 & n10481 ) ;
  assign n10483 = ( n10052 & ~n10054 ) | ( n10052 & n10481 ) | ( ~n10054 & n10481 ) ;
  assign n10484 = ( n10054 & ~n10482 ) | ( n10054 & n10483 ) | ( ~n10482 & n10483 ) ;
  assign n10485 = n702 | n10015 ;
  assign n10486 = ~x1 |  x0 ;
  assign n10487 = n599 | n10486 ;
  assign n10488 = n10485 &  n10487 ;
  assign n10489 = x2 &  n10488 ;
  assign n10490 = n3937 &  n10017 ;
  assign n10491 = ( n10489 & ~n3937 ) | ( n10489 & n10490 ) | ( ~n3937 & n10490 ) ;
  assign n10492 = n10017 &  n10488 ;
  assign n10493 = x2 | n10492 ;
  assign n10494 = n3937 | n10488 ;
  assign n10495 = ( n10493 & ~n3937 ) | ( n10493 & n10494 ) | ( ~n3937 & n10494 ) ;
  assign n10496 = ~n10491 & n10495 ;
  assign n10503 = ~n863 & n10015 ;
  assign n10499 = x0 &  ~n10013 ;
  assign n10500 = ~n599 & n10499 ;
  assign n10501 = n702 | n10486 ;
  assign n10502 = ~n10500 & n10501 ;
  assign n10504 = ( n863 & n10503 ) | ( n863 & n10502 ) | ( n10503 & n10502 ) ;
  assign n10505 = ( n3934 & ~n3635 ) | ( n3934 & n10017 ) | ( ~n3635 & n10017 ) ;
  assign n10506 = ( n4451 & n10504 ) | ( n4451 & n10505 ) | ( n10504 & n10505 ) ;
  assign n10508 = x2 &  n10506 ;
  assign n10507 = ~x2 & n10506 ;
  assign n10509 = ( x2 & ~n10508 ) | ( x2 & n10507 ) | ( ~n10508 & n10507 ) ;
  assign n10497 = ( n10064 & n10066 ) | ( n10064 & n10480 ) | ( n10066 & n10480 ) ;
  assign n10498 = ( n10066 & ~n10497 ) | ( n10066 & n10481 ) | ( ~n10497 & n10481 ) ;
  assign n10510 = ( n10076 & ~n10078 ) | ( n10076 & n10479 ) | ( ~n10078 & n10479 ) ;
  assign n10511 = ( n10078 & ~n10480 ) | ( n10078 & n10510 ) | ( ~n10480 & n10510 ) ;
  assign n10515 = ~n946 & n10015 ;
  assign n10512 = ~n702 & n10499 ;
  assign n10513 = n863 | n10486 ;
  assign n10514 = ~n10512 & n10513 ;
  assign n10516 = ( n946 & n10515 ) | ( n946 & n10514 ) | ( n10515 & n10514 ) ;
  assign n10517 = ( n3647 & ~n3634 ) | ( n3647 & n10017 ) | ( ~n3634 & n10017 ) ;
  assign n10518 = ( n3649 & n10516 ) | ( n3649 & n10517 ) | ( n10516 & n10517 ) ;
  assign n10520 = x2 &  n10518 ;
  assign n10519 = ~x2 & n10518 ;
  assign n10521 = ( x2 & ~n10520 ) | ( x2 & n10519 ) | ( ~n10520 & n10519 ) ;
  assign n10522 = ( n10088 & ~n10090 ) | ( n10088 & n10478 ) | ( ~n10090 & n10478 ) ;
  assign n10523 = ( n10090 & ~n10479 ) | ( n10090 & n10522 ) | ( ~n10479 & n10522 ) ;
  assign n10527 = ~n946 & n10486 ;
  assign n10524 = ~n863 & n10499 ;
  assign n10525 = n1043 | n10015 ;
  assign n10526 = ~n10524 & n10525 ;
  assign n10528 = ( n946 & n10527 ) | ( n946 & n10526 ) | ( n10527 & n10526 ) ;
  assign n10529 = ( n3911 & ~n3633 ) | ( n3911 & n10017 ) | ( ~n3633 & n10017 ) ;
  assign n10530 = ( n3913 & n10528 ) | ( n3913 & n10529 ) | ( n10528 & n10529 ) ;
  assign n10532 = x2 &  n10530 ;
  assign n10531 = ~x2 & n10530 ;
  assign n10533 = ( x2 & ~n10532 ) | ( x2 & n10531 ) | ( ~n10532 & n10531 ) ;
  assign n10536 = n946 &  n10499 ;
  assign n10537 = n1151 | n10015 ;
  assign n10538 = n1043 | n10486 ;
  assign n10539 = n10537 &  n10538 ;
  assign n10540 = ( n10536 & ~n10499 ) | ( n10536 & n10539 ) | ( ~n10499 & n10539 ) ;
  assign n10541 = ( n4035 & ~n3632 ) | ( n4035 & n10017 ) | ( ~n3632 & n10017 ) ;
  assign n10542 = ( n4037 & n10540 ) | ( n4037 & n10541 ) | ( n10540 & n10541 ) ;
  assign n10544 = x2 &  n10542 ;
  assign n10543 = ~x2 & n10542 ;
  assign n10545 = ( x2 & ~n10544 ) | ( x2 & n10543 ) | ( ~n10544 & n10543 ) ;
  assign n10534 = ( n10100 & n10102 ) | ( n10100 & n10477 ) | ( n10102 & n10477 ) ;
  assign n10535 = ( n10102 & ~n10534 ) | ( n10102 & n10478 ) | ( ~n10534 & n10478 ) ;
  assign n10546 = ( n10128 & ~n10118 ) | ( n10128 & n10475 ) | ( ~n10118 & n10475 ) ;
  assign n10547 = ( n10118 & ~n10128 ) | ( n10118 & n10475 ) | ( ~n10128 & n10475 ) ;
  assign n10548 = ( n10546 & ~n10475 ) | ( n10546 & n10547 ) | ( ~n10475 & n10547 ) ;
  assign n10561 = ( x5 & ~n10436 ) | ( x5 & n10437 ) | ( ~n10436 & n10437 ) ;
  assign n10562 = ( x5 & ~n10561 ) | ( x5 & 1'b0 ) | ( ~n10561 & 1'b0 ) ;
  assign n10563 = ( x5 & ~n10562 ) | ( x5 & n10431 ) | ( ~n10562 & n10431 ) ;
  assign n10564 = ( n10431 & ~x5 ) | ( n10431 & n10562 ) | ( ~x5 & n10562 ) ;
  assign n10565 = ( n10563 & ~n10431 ) | ( n10563 & n10564 ) | ( ~n10431 & n10564 ) ;
  assign n10599 = ~n3460 & n10015 ;
  assign n10596 = ~n3325 & n10499 ;
  assign n10597 = n3361 | n10486 ;
  assign n10598 = ~n10596 & n10597 ;
  assign n10600 = ( n3460 & n10599 ) | ( n3460 & n10598 ) | ( n10599 & n10598 ) ;
  assign n10601 = ( n6800 & ~n3604 ) | ( n6800 & n10017 ) | ( ~n3604 & n10017 ) ;
  assign n10602 = ( n6801 & n10600 ) | ( n6801 & n10601 ) | ( n10600 & n10601 ) ;
  assign n10604 = x2 &  n10602 ;
  assign n10603 = ~x2 & n10602 ;
  assign n10605 = ( x2 & ~n10604 ) | ( x2 & n10603 ) | ( ~n10604 & n10603 ) ;
  assign n10588 = ~n3460 & n10486 ;
  assign n10585 = ~n3361 & n10499 ;
  assign n10586 = n3601 | n10015 ;
  assign n10587 = ~n10585 & n10586 ;
  assign n10589 = ( n3460 & n10588 ) | ( n3460 & n10587 ) | ( n10588 & n10587 ) ;
  assign n10590 = ( n9510 & ~n3603 ) | ( n9510 & n10017 ) | ( ~n3603 & n10017 ) ;
  assign n10591 = ( n9511 & n10589 ) | ( n9511 & n10590 ) | ( n10589 & n10590 ) ;
  assign n10592 = x2 | n10591 ;
  assign n10593 = ( x2 & ~n10591 ) | ( x2 & 1'b0 ) | ( ~n10591 & 1'b0 ) ;
  assign n10594 = ( n10592 & ~x2 ) | ( n10592 & n10593 ) | ( ~x2 & n10593 ) ;
  assign n10566 = ( x0 & ~n3547 ) | ( x0 & 1'b0 ) | ( ~n3547 & 1'b0 ) ;
  assign n10567 = ( x2 & ~n10017 ) | ( x2 & 1'b0 ) | ( ~n10017 & 1'b0 ) ;
  assign n10582 = n10567 | n6886 ;
  assign n10568 = n3460 &  n10499 ;
  assign n10569 = n3547 | n10015 ;
  assign n10570 = n3601 | n10486 ;
  assign n10571 = n10569 &  n10570 ;
  assign n10572 = ( n10568 & ~n10499 ) | ( n10568 & n10571 ) | ( ~n10499 & n10571 ) ;
  assign n10573 = ( x2 & ~n10572 ) | ( x2 & 1'b0 ) | ( ~n10572 & 1'b0 ) ;
  assign n10579 = ~n10567 & n7412 ;
  assign n10574 = ( x2 & ~n10486 ) | ( x2 & 1'b0 ) | ( ~n10486 & 1'b0 ) ;
  assign n10575 = ~n3547 & n10574 ;
  assign n10576 = n3601 &  n10499 ;
  assign n10577 = ( x2 & ~n10499 ) | ( x2 & n10576 ) | ( ~n10499 & n10576 ) ;
  assign n10578 = ~n10575 & n10577 ;
  assign n10580 = ( n10579 & ~n7412 ) | ( n10579 & n10578 ) | ( ~n7412 & n10578 ) ;
  assign n10581 = ~n10573 & n10580 ;
  assign n10583 = ( n6886 & ~n10582 ) | ( n6886 & n10581 ) | ( ~n10582 & n10581 ) ;
  assign n10584 = ~n10566 & n10583 ;
  assign n10595 = ( n10437 & ~n10594 ) | ( n10437 & n10584 ) | ( ~n10594 & n10584 ) ;
  assign n10438 = ( x5 & ~n10437 ) | ( x5 & 1'b0 ) | ( ~n10437 & 1'b0 ) ;
  assign n10606 = ( n10436 & ~x5 ) | ( n10436 & n10438 ) | ( ~x5 & n10438 ) ;
  assign n10607 = ( x5 & ~n10438 ) | ( x5 & n10436 ) | ( ~n10438 & n10436 ) ;
  assign n10608 = ( n10606 & ~n10436 ) | ( n10606 & n10607 ) | ( ~n10436 & n10607 ) ;
  assign n10609 = ( n10605 & ~n10595 ) | ( n10605 & n10608 ) | ( ~n10595 & n10608 ) ;
  assign n10615 = ( n3605 & ~n10017 ) | ( n3605 & n6753 ) | ( ~n10017 & n6753 ) ;
  assign n10613 = ~n10499 & n3266 ;
  assign n10610 = n3361 | n10015 ;
  assign n10611 = n3325 | n10486 ;
  assign n10612 = n10610 &  n10611 ;
  assign n10614 = ( n10613 & ~n3266 ) | ( n10613 & n10612 ) | ( ~n3266 & n10612 ) ;
  assign n10616 = ( n6754 & ~n10615 ) | ( n6754 & n10614 ) | ( ~n10615 & n10614 ) ;
  assign n10617 = x2 | n10616 ;
  assign n10618 = ( x2 & ~n10616 ) | ( x2 & 1'b0 ) | ( ~n10616 & 1'b0 ) ;
  assign n10619 = ( n10617 & ~x2 ) | ( n10617 & n10618 ) | ( ~x2 & n10618 ) ;
  assign n10620 = ( n10565 & n10609 ) | ( n10565 & n10619 ) | ( n10609 & n10619 ) ;
  assign n10626 = ( n3606 & ~n10017 ) | ( n3606 & n6705 ) | ( ~n10017 & n6705 ) ;
  assign n10621 = ~n3197 & n10499 ;
  assign n10622 = n3325 | n10015 ;
  assign n10623 = ~n10621 & n10622 ;
  assign n10624 = n3266 &  n10486 ;
  assign n10625 = ( n10623 & ~n3266 ) | ( n10623 & n10624 ) | ( ~n3266 & n10624 ) ;
  assign n10627 = ( n6706 & ~n10626 ) | ( n6706 & n10625 ) | ( ~n10626 & n10625 ) ;
  assign n10629 = x2 &  n10627 ;
  assign n10628 = ~x2 & n10627 ;
  assign n10630 = ( x2 & ~n10629 ) | ( x2 & n10628 ) | ( ~n10629 & n10628 ) ;
  assign n10632 = ( n9951 & n10441 ) | ( n9951 & n10451 ) | ( n10441 & n10451 ) ;
  assign n10631 = ( n9951 & ~n10441 ) | ( n9951 & n10451 ) | ( ~n10441 & n10451 ) ;
  assign n10633 = ( n10441 & ~n10632 ) | ( n10441 & n10631 ) | ( ~n10632 & n10631 ) ;
  assign n10634 = ( n10620 & n10630 ) | ( n10620 & n10633 ) | ( n10630 & n10633 ) ;
  assign n10558 = ( n10414 & n10424 ) | ( n10414 & n10452 ) | ( n10424 & n10452 ) ;
  assign n10559 = ( n10414 & ~n10424 ) | ( n10414 & n10452 ) | ( ~n10424 & n10452 ) ;
  assign n10560 = ( n10424 & ~n10558 ) | ( n10424 & n10559 ) | ( ~n10558 & n10559 ) ;
  assign n10635 = ~n3106 & n10499 ;
  assign n10636 = n3197 | n10486 ;
  assign n10637 = ~n10635 & n10636 ;
  assign n10638 = n3266 &  n10015 ;
  assign n10639 = ( n10637 & ~n3266 ) | ( n10637 & n10638 ) | ( ~n3266 & n10638 ) ;
  assign n10640 = ( n6654 & ~n3607 ) | ( n6654 & n10017 ) | ( ~n3607 & n10017 ) ;
  assign n10641 = ( n6655 & n10639 ) | ( n6655 & n10640 ) | ( n10639 & n10640 ) ;
  assign n10642 = x2 | n10641 ;
  assign n10643 = ( x2 & ~n10641 ) | ( x2 & 1'b0 ) | ( ~n10641 & 1'b0 ) ;
  assign n10644 = ( n10642 & ~x2 ) | ( n10642 & n10643 ) | ( ~x2 & n10643 ) ;
  assign n10645 = ( n10634 & ~n10560 ) | ( n10634 & n10644 ) | ( ~n10560 & n10644 ) ;
  assign n10646 = n3030 &  n10499 ;
  assign n10647 = n3197 | n10015 ;
  assign n10648 = n3106 | n10486 ;
  assign n10649 = n10647 &  n10648 ;
  assign n10650 = ( n10646 & ~n10499 ) | ( n10646 & n10649 ) | ( ~n10499 & n10649 ) ;
  assign n10651 = ( n6311 & ~n3608 ) | ( n6311 & n10017 ) | ( ~n3608 & n10017 ) ;
  assign n10652 = ( n6313 & n10650 ) | ( n6313 & n10651 ) | ( n10650 & n10651 ) ;
  assign n10654 = x2 &  n10652 ;
  assign n10653 = ~x2 & n10652 ;
  assign n10655 = ( x2 & ~n10654 ) | ( x2 & n10653 ) | ( ~n10654 & n10653 ) ;
  assign n10656 = ~x5 & n10405 ;
  assign n10657 = ( n10406 & ~n10405 ) | ( n10406 & n10656 ) | ( ~n10405 & n10656 ) ;
  assign n10659 = ( n10412 & n10453 ) | ( n10412 & n10657 ) | ( n10453 & n10657 ) ;
  assign n10658 = ( n10412 & ~n10657 ) | ( n10412 & n10453 ) | ( ~n10657 & n10453 ) ;
  assign n10660 = ( n10657 & ~n10659 ) | ( n10657 & n10658 ) | ( ~n10659 & n10658 ) ;
  assign n10661 = ( n10645 & n10655 ) | ( n10645 & n10660 ) | ( n10655 & n10660 ) ;
  assign n10665 = n10499 | n2995 ;
  assign n10662 = n3106 | n10015 ;
  assign n10663 = n3030 | n10486 ;
  assign n10664 = n10662 &  n10663 ;
  assign n10666 = ( n2995 & ~n10665 ) | ( n2995 & n10664 ) | ( ~n10665 & n10664 ) ;
  assign n10667 = ( n6604 & ~n3609 ) | ( n6604 & n10017 ) | ( ~n3609 & n10017 ) ;
  assign n10668 = ( n6605 & n10666 ) | ( n6605 & n10667 ) | ( n10666 & n10667 ) ;
  assign n10670 = x2 &  n10668 ;
  assign n10669 = ~x2 & n10668 ;
  assign n10671 = ( x2 & ~n10670 ) | ( x2 & n10669 ) | ( ~n10670 & n10669 ) ;
  assign n10672 = ( n10388 & ~n10454 ) | ( n10388 & n10398 ) | ( ~n10454 & n10398 ) ;
  assign n10673 = ( n10454 & ~n10455 ) | ( n10454 & n10672 ) | ( ~n10455 & n10672 ) ;
  assign n10674 = ( n10661 & n10671 ) | ( n10661 & n10673 ) | ( n10671 & n10673 ) ;
  assign n10685 = n7363 | n9155 ;
  assign n10686 = n10377 &  n10685 ;
  assign n10687 = ( n10385 & ~x5 ) | ( n10385 & n10686 ) | ( ~x5 & n10686 ) ;
  assign n10688 = ( x5 & ~n10686 ) | ( x5 & n10385 ) | ( ~n10686 & n10385 ) ;
  assign n10689 = ( n10687 & ~n10385 ) | ( n10687 & n10688 ) | ( ~n10385 & n10688 ) ;
  assign n10690 = ~n10455 & n10689 ;
  assign n10691 = ( n10455 & ~n10689 ) | ( n10455 & 1'b0 ) | ( ~n10689 & 1'b0 ) ;
  assign n10692 = n10690 | n10691 ;
  assign n10675 = n2839 &  n10499 ;
  assign n10676 = n3030 | n10015 ;
  assign n10677 = n2995 | n10486 ;
  assign n10678 = n10676 &  n10677 ;
  assign n10679 = ( n10675 & ~n10499 ) | ( n10675 & n10678 ) | ( ~n10499 & n10678 ) ;
  assign n10680 = ( n6591 & ~n3610 ) | ( n6591 & n10017 ) | ( ~n3610 & n10017 ) ;
  assign n10681 = ( n6592 & n10679 ) | ( n6592 & n10680 ) | ( n10679 & n10680 ) ;
  assign n10683 = x2 &  n10681 ;
  assign n10682 = ~x2 & n10681 ;
  assign n10684 = ( x2 & ~n10683 ) | ( x2 & n10682 ) | ( ~n10683 & n10682 ) ;
  assign n10693 = ( n10674 & ~n10692 ) | ( n10674 & n10684 ) | ( ~n10692 & n10684 ) ;
  assign n10699 = ( n3611 & ~n10017 ) | ( n3611 & n9834 ) | ( ~n10017 & n9834 ) ;
  assign n10697 = ~n10499 & n2910 ;
  assign n10694 = n2995 | n10015 ;
  assign n10695 = n2839 | n10486 ;
  assign n10696 = n10694 &  n10695 ;
  assign n10698 = ( n10697 & ~n2910 ) | ( n10697 & n10696 ) | ( ~n2910 & n10696 ) ;
  assign n10700 = ( n9835 & ~n10699 ) | ( n9835 & n10698 ) | ( ~n10699 & n10698 ) ;
  assign n10701 = ( x2 & ~n10700 ) | ( x2 & 1'b0 ) | ( ~n10700 & 1'b0 ) ;
  assign n10702 = ~x2 & n10700 ;
  assign n10703 = n10701 | n10702 ;
  assign n10704 = ( n10372 & ~n10362 ) | ( n10372 & n10456 ) | ( ~n10362 & n10456 ) ;
  assign n10705 = ( n10362 & ~n10372 ) | ( n10362 & n10456 ) | ( ~n10372 & n10456 ) ;
  assign n10706 = ( n10704 & ~n10456 ) | ( n10704 & n10705 ) | ( ~n10456 & n10705 ) ;
  assign n10707 = ( n10693 & n10703 ) | ( n10693 & n10706 ) | ( n10703 & n10706 ) ;
  assign n10708 = ( n10360 & ~n10350 ) | ( n10360 & n10457 ) | ( ~n10350 & n10457 ) ;
  assign n10709 = ( n10350 & ~n10360 ) | ( n10350 & n10457 ) | ( ~n10360 & n10457 ) ;
  assign n10710 = ( n10708 & ~n10457 ) | ( n10708 & n10709 ) | ( ~n10457 & n10709 ) ;
  assign n10711 = ~n2783 & n10499 ;
  assign n10712 = n2839 | n10015 ;
  assign n10713 = ~n10711 & n10712 ;
  assign n10714 = n2910 &  n10486 ;
  assign n10715 = ( n10713 & ~n2910 ) | ( n10713 & n10714 ) | ( ~n2910 & n10714 ) ;
  assign n10716 = ( n6104 & n10017 ) | ( n6104 & n10715 ) | ( n10017 & n10715 ) ;
  assign n10717 = ~n10017 & n10716 ;
  assign n10718 = ( x2 & ~n10715 ) | ( x2 & n10717 ) | ( ~n10715 & n10717 ) ;
  assign n10719 = ( n10715 & ~x2 ) | ( n10715 & n10717 ) | ( ~x2 & n10717 ) ;
  assign n10720 = ( n10718 & ~n10717 ) | ( n10718 & n10719 ) | ( ~n10717 & n10719 ) ;
  assign n10721 = ( n10707 & n10710 ) | ( n10707 & n10720 ) | ( n10710 & n10720 ) ;
  assign n10555 = ( n10337 & n10347 ) | ( n10337 & n10458 ) | ( n10347 & n10458 ) ;
  assign n10556 = ( n10337 & ~n10458 ) | ( n10337 & n10347 ) | ( ~n10458 & n10347 ) ;
  assign n10557 = ( n10458 & ~n10555 ) | ( n10458 & n10556 ) | ( ~n10555 & n10556 ) ;
  assign n10722 = ~n2751 & n10499 ;
  assign n10723 = n2783 | n10486 ;
  assign n10724 = ~n10722 & n10723 ;
  assign n10725 = n2910 &  n10015 ;
  assign n10726 = ( n10724 & ~n2910 ) | ( n10724 & n10725 ) | ( ~n2910 & n10725 ) ;
  assign n10727 = ( n9804 & ~n3613 ) | ( n9804 & n10017 ) | ( ~n3613 & n10017 ) ;
  assign n10728 = ( n9805 & n10726 ) | ( n9805 & n10727 ) | ( n10726 & n10727 ) ;
  assign n10729 = x2 | n10728 ;
  assign n10730 = ( x2 & ~n10728 ) | ( x2 & 1'b0 ) | ( ~n10728 & 1'b0 ) ;
  assign n10731 = ( n10729 & ~x2 ) | ( n10729 & n10730 ) | ( ~x2 & n10730 ) ;
  assign n10732 = ( n10721 & ~n10557 ) | ( n10721 & n10731 ) | ( ~n10557 & n10731 ) ;
  assign n10736 = ~n2751 & n10486 ;
  assign n10733 = ~n2665 & n10499 ;
  assign n10734 = n2783 | n10015 ;
  assign n10735 = ~n10733 & n10734 ;
  assign n10737 = ( n2751 & n10736 ) | ( n2751 & n10735 ) | ( n10736 & n10735 ) ;
  assign n10738 = ( n6116 & ~n3614 ) | ( n6116 & n10017 ) | ( ~n3614 & n10017 ) ;
  assign n10739 = ( n6118 & n10737 ) | ( n6118 & n10738 ) | ( n10737 & n10738 ) ;
  assign n10741 = x2 &  n10739 ;
  assign n10740 = ~x2 & n10739 ;
  assign n10742 = ( x2 & ~n10741 ) | ( x2 & n10740 ) | ( ~n10741 & n10740 ) ;
  assign n10743 = ( n6330 & ~n9155 ) | ( n6330 & 1'b0 ) | ( ~n9155 & 1'b0 ) ;
  assign n10744 = ( n10326 & ~n10743 ) | ( n10326 & 1'b0 ) | ( ~n10743 & 1'b0 ) ;
  assign n10745 = ( n10334 & ~x5 ) | ( n10334 & n10744 ) | ( ~x5 & n10744 ) ;
  assign n10746 = ( x5 & ~n10744 ) | ( x5 & n10334 ) | ( ~n10744 & n10334 ) ;
  assign n10747 = ( n10745 & ~n10334 ) | ( n10745 & n10746 ) | ( ~n10334 & n10746 ) ;
  assign n10748 = ~n10459 & n10747 ;
  assign n10749 = ( n10459 & ~n10747 ) | ( n10459 & 1'b0 ) | ( ~n10747 & 1'b0 ) ;
  assign n10750 = n10748 | n10749 ;
  assign n10751 = ( n10732 & n10742 ) | ( n10732 & n10750 ) | ( n10742 & n10750 ) ;
  assign n10755 = ~n2751 & n10015 ;
  assign n10752 = ~n2569 & n10499 ;
  assign n10753 = n2665 | n10486 ;
  assign n10754 = ~n10752 & n10753 ;
  assign n10756 = ( n2751 & n10755 ) | ( n2751 & n10754 ) | ( n10755 & n10754 ) ;
  assign n10757 = ( n5702 & ~n3615 ) | ( n5702 & n10017 ) | ( ~n3615 & n10017 ) ;
  assign n10758 = ( n5704 & n10756 ) | ( n5704 & n10757 ) | ( n10756 & n10757 ) ;
  assign n10760 = x2 &  n10758 ;
  assign n10759 = ~x2 & n10758 ;
  assign n10761 = ( x2 & ~n10760 ) | ( x2 & n10759 ) | ( ~n10760 & n10759 ) ;
  assign n10762 = ( n10315 & ~x5 ) | ( n10315 & n10321 ) | ( ~x5 & n10321 ) ;
  assign n10763 = ( x5 & ~n10315 ) | ( x5 & n10321 ) | ( ~n10315 & n10321 ) ;
  assign n10764 = ( n10762 & ~n10321 ) | ( n10762 & n10763 ) | ( ~n10321 & n10763 ) ;
  assign n10765 = n10460 | n10764 ;
  assign n10766 = n10460 &  n10764 ;
  assign n10767 = ( n10765 & ~n10766 ) | ( n10765 & 1'b0 ) | ( ~n10766 & 1'b0 ) ;
  assign n10768 = ( n10751 & n10761 ) | ( n10751 & n10767 ) | ( n10761 & n10767 ) ;
  assign n10779 = n6226 | n9155 ;
  assign n10780 = n10300 &  n10779 ;
  assign n10781 = ( n10308 & ~x5 ) | ( n10308 & n10780 ) | ( ~x5 & n10780 ) ;
  assign n10782 = ( x5 & ~n10780 ) | ( x5 & n10308 ) | ( ~n10780 & n10308 ) ;
  assign n10783 = ( n10781 & ~n10308 ) | ( n10781 & n10782 ) | ( ~n10308 & n10782 ) ;
  assign n10784 = ~n10461 & n10783 ;
  assign n10785 = ( n10461 & ~n10783 ) | ( n10461 & 1'b0 ) | ( ~n10783 & 1'b0 ) ;
  assign n10786 = n10784 | n10785 ;
  assign n10772 = ~n2665 & n10015 ;
  assign n10769 = ~n2483 & n10499 ;
  assign n10770 = n2569 | n10486 ;
  assign n10771 = ~n10769 & n10770 ;
  assign n10773 = ( n2665 & n10772 ) | ( n2665 & n10771 ) | ( n10772 & n10771 ) ;
  assign n10774 = ( n5886 & ~n3616 ) | ( n5886 & n10017 ) | ( ~n3616 & n10017 ) ;
  assign n10775 = ( n5887 & n10773 ) | ( n5887 & n10774 ) | ( n10773 & n10774 ) ;
  assign n10777 = x2 &  n10775 ;
  assign n10776 = ~x2 & n10775 ;
  assign n10778 = ( x2 & ~n10777 ) | ( x2 & n10776 ) | ( ~n10777 & n10776 ) ;
  assign n10787 = ( n10768 & ~n10786 ) | ( n10768 & n10778 ) | ( ~n10786 & n10778 ) ;
  assign n10788 = ( n10295 & ~n10285 ) | ( n10295 & n10462 ) | ( ~n10285 & n10462 ) ;
  assign n10789 = ( n10285 & ~n10295 ) | ( n10285 & n10462 ) | ( ~n10295 & n10462 ) ;
  assign n10790 = ( n10788 & ~n10462 ) | ( n10788 & n10789 ) | ( ~n10462 & n10789 ) ;
  assign n10791 = n2392 &  n10499 ;
  assign n10792 = n2569 | n10015 ;
  assign n10793 = n2483 | n10486 ;
  assign n10794 = n10792 &  n10793 ;
  assign n10795 = ( n10791 & ~n10499 ) | ( n10791 & n10794 ) | ( ~n10499 & n10794 ) ;
  assign n10796 = ( n5519 & ~n3617 ) | ( n5519 & n10017 ) | ( ~n3617 & n10017 ) ;
  assign n10797 = ( n5520 & n10795 ) | ( n5520 & n10796 ) | ( n10795 & n10796 ) ;
  assign n10798 = x2 | n10797 ;
  assign n10799 = ( x2 & ~n10797 ) | ( x2 & 1'b0 ) | ( ~n10797 & 1'b0 ) ;
  assign n10800 = ( n10798 & ~x2 ) | ( n10798 & n10799 ) | ( ~x2 & n10799 ) ;
  assign n10801 = ( n10787 & n10790 ) | ( n10787 & n10800 ) | ( n10790 & n10800 ) ;
  assign n10802 = ( n10283 & ~n10273 ) | ( n10283 & n10463 ) | ( ~n10273 & n10463 ) ;
  assign n10803 = ( n10273 & ~n10283 ) | ( n10273 & n10463 ) | ( ~n10283 & n10463 ) ;
  assign n10804 = ( n10802 & ~n10463 ) | ( n10802 & n10803 ) | ( ~n10463 & n10803 ) ;
  assign n10805 = n2296 &  n10499 ;
  assign n10806 = n2483 | n10015 ;
  assign n10807 = n2392 | n10486 ;
  assign n10808 = n10806 &  n10807 ;
  assign n10809 = ( n10805 & ~n10499 ) | ( n10805 & n10808 ) | ( ~n10499 & n10808 ) ;
  assign n10810 = ( n5497 & ~n3618 ) | ( n5497 & n10017 ) | ( ~n3618 & n10017 ) ;
  assign n10811 = ( n5499 & n10809 ) | ( n5499 & n10810 ) | ( n10809 & n10810 ) ;
  assign n10812 = x2 | n10811 ;
  assign n10813 = ( x2 & ~n10811 ) | ( x2 & 1'b0 ) | ( ~n10811 & 1'b0 ) ;
  assign n10814 = ( n10812 & ~x2 ) | ( n10812 & n10813 ) | ( ~x2 & n10813 ) ;
  assign n10815 = ( n10801 & n10804 ) | ( n10801 & n10814 ) | ( n10804 & n10814 ) ;
  assign n10552 = ( n10261 & n10271 ) | ( n10261 & n10464 ) | ( n10271 & n10464 ) ;
  assign n10553 = ( n10261 & ~n10464 ) | ( n10261 & n10271 ) | ( ~n10464 & n10271 ) ;
  assign n10554 = ( n10464 & ~n10552 ) | ( n10464 & n10553 ) | ( ~n10552 & n10553 ) ;
  assign n10816 = n2178 &  n10499 ;
  assign n10817 = n2392 | n10015 ;
  assign n10818 = n2296 | n10486 ;
  assign n10819 = n10817 &  n10818 ;
  assign n10820 = ( n10816 & ~n10499 ) | ( n10816 & n10819 ) | ( ~n10499 & n10819 ) ;
  assign n10821 = ( n5266 & ~n3619 ) | ( n5266 & n10017 ) | ( ~n3619 & n10017 ) ;
  assign n10822 = ( n5268 & n10820 ) | ( n5268 & n10821 ) | ( n10820 & n10821 ) ;
  assign n10823 = x2 | n10822 ;
  assign n10824 = ( x2 & ~n10822 ) | ( x2 & 1'b0 ) | ( ~n10822 & 1'b0 ) ;
  assign n10825 = ( n10823 & ~x2 ) | ( n10823 & n10824 ) | ( ~x2 & n10824 ) ;
  assign n10826 = ( n10815 & ~n10554 ) | ( n10815 & n10825 ) | ( ~n10554 & n10825 ) ;
  assign n10830 = ~n2296 & n10015 ;
  assign n10827 = ~n2127 & n10499 ;
  assign n10828 = n2178 | n10486 ;
  assign n10829 = ~n10827 & n10828 ;
  assign n10831 = ( n2296 & n10830 ) | ( n2296 & n10829 ) | ( n10830 & n10829 ) ;
  assign n10832 = ( n5280 & ~n3620 ) | ( n5280 & n10017 ) | ( ~n3620 & n10017 ) ;
  assign n10833 = ( n5282 & n10831 ) | ( n5282 & n10832 ) | ( n10831 & n10832 ) ;
  assign n10835 = x2 &  n10833 ;
  assign n10834 = ~x2 & n10833 ;
  assign n10836 = ( x2 & ~n10835 ) | ( x2 & n10834 ) | ( ~n10835 & n10834 ) ;
  assign n10837 = n6212 | n9155 ;
  assign n10838 = n10250 &  n10837 ;
  assign n10839 = ( n10258 & ~x5 ) | ( n10258 & n10838 ) | ( ~x5 & n10838 ) ;
  assign n10840 = ( x5 & ~n10838 ) | ( x5 & n10258 ) | ( ~n10838 & n10258 ) ;
  assign n10841 = ( n10839 & ~n10258 ) | ( n10839 & n10840 ) | ( ~n10258 & n10840 ) ;
  assign n10842 = ~n10465 & n10841 ;
  assign n10843 = ( n10465 & ~n10841 ) | ( n10465 & 1'b0 ) | ( ~n10841 & 1'b0 ) ;
  assign n10844 = n10842 | n10843 ;
  assign n10845 = ( n10826 & n10836 ) | ( n10826 & n10844 ) | ( n10836 & n10844 ) ;
  assign n10849 = n10499 | n2022 ;
  assign n10846 = n2178 | n10015 ;
  assign n10847 = n2127 | n10486 ;
  assign n10848 = n10846 &  n10847 ;
  assign n10850 = ( n2022 & ~n10849 ) | ( n2022 & n10848 ) | ( ~n10849 & n10848 ) ;
  assign n10851 = ( n4931 & ~n3621 ) | ( n4931 & n10017 ) | ( ~n3621 & n10017 ) ;
  assign n10852 = ( n4933 & n10850 ) | ( n4933 & n10851 ) | ( n10850 & n10851 ) ;
  assign n10854 = x2 &  n10852 ;
  assign n10853 = ~x2 & n10852 ;
  assign n10855 = ( x2 & ~n10854 ) | ( x2 & n10853 ) | ( ~n10854 & n10853 ) ;
  assign n10856 = n5500 | n9155 ;
  assign n10857 = n10237 &  n10856 ;
  assign n10858 = ( n10245 & ~x5 ) | ( n10245 & n10857 ) | ( ~x5 & n10857 ) ;
  assign n10859 = ( x5 & ~n10857 ) | ( x5 & n10245 ) | ( ~n10857 & n10245 ) ;
  assign n10860 = ( n10858 & ~n10245 ) | ( n10858 & n10859 ) | ( ~n10245 & n10859 ) ;
  assign n10861 = n10466 | n10860 ;
  assign n10862 = n10466 &  n10860 ;
  assign n10863 = ( n10861 & ~n10862 ) | ( n10861 & 1'b0 ) | ( ~n10862 & 1'b0 ) ;
  assign n10864 = ( n10845 & n10855 ) | ( n10845 & n10863 ) | ( n10855 & n10863 ) ;
  assign n10875 = n5269 | n9155 ;
  assign n10876 = n10224 &  n10875 ;
  assign n10877 = ( n10232 & ~x5 ) | ( n10232 & n10876 ) | ( ~x5 & n10876 ) ;
  assign n10878 = ( x5 & ~n10876 ) | ( x5 & n10232 ) | ( ~n10876 & n10232 ) ;
  assign n10879 = ( n10877 & ~n10232 ) | ( n10877 & n10878 ) | ( ~n10232 & n10878 ) ;
  assign n10880 = ~n10467 & n10879 ;
  assign n10881 = ( n10467 & ~n10879 ) | ( n10467 & 1'b0 ) | ( ~n10879 & 1'b0 ) ;
  assign n10882 = n10880 | n10881 ;
  assign n10868 = n10499 | n1940 ;
  assign n10865 = n2127 | n10015 ;
  assign n10866 = n2022 | n10486 ;
  assign n10867 = n10865 &  n10866 ;
  assign n10869 = ( n1940 & ~n10868 ) | ( n1940 & n10867 ) | ( ~n10868 & n10867 ) ;
  assign n10870 = ( n5085 & ~n3622 ) | ( n5085 & n10017 ) | ( ~n3622 & n10017 ) ;
  assign n10871 = ( n5086 & n10869 ) | ( n5086 & n10870 ) | ( n10869 & n10870 ) ;
  assign n10873 = x2 &  n10871 ;
  assign n10872 = ~x2 & n10871 ;
  assign n10874 = ( x2 & ~n10873 ) | ( x2 & n10872 ) | ( ~n10873 & n10872 ) ;
  assign n10883 = ( n10864 & ~n10882 ) | ( n10864 & n10874 ) | ( ~n10882 & n10874 ) ;
  assign n10884 = ( n10219 & ~n10209 ) | ( n10219 & n10468 ) | ( ~n10209 & n10468 ) ;
  assign n10885 = ( n10209 & ~n10219 ) | ( n10209 & n10468 ) | ( ~n10219 & n10468 ) ;
  assign n10886 = ( n10884 & ~n10468 ) | ( n10884 & n10885 ) | ( ~n10468 & n10885 ) ;
  assign n10887 = n1875 &  n10499 ;
  assign n10888 = n2022 | n10015 ;
  assign n10889 = n1940 | n10486 ;
  assign n10890 = n10888 &  n10889 ;
  assign n10891 = ( n10887 & ~n10499 ) | ( n10887 & n10890 ) | ( ~n10499 & n10890 ) ;
  assign n10892 = ( n4761 & ~n3623 ) | ( n4761 & n10017 ) | ( ~n3623 & n10017 ) ;
  assign n10893 = ( n4762 & n10891 ) | ( n4762 & n10892 ) | ( n10891 & n10892 ) ;
  assign n10894 = x2 | n10893 ;
  assign n10895 = ( x2 & ~n10893 ) | ( x2 & 1'b0 ) | ( ~n10893 & 1'b0 ) ;
  assign n10896 = ( n10894 & ~x2 ) | ( n10894 & n10895 ) | ( ~x2 & n10895 ) ;
  assign n10897 = ( n10883 & n10886 ) | ( n10883 & n10896 ) | ( n10886 & n10896 ) ;
  assign n10898 = ( n10206 & ~n10196 ) | ( n10206 & n10469 ) | ( ~n10196 & n10469 ) ;
  assign n10899 = ( n10196 & ~n10206 ) | ( n10196 & n10469 ) | ( ~n10206 & n10469 ) ;
  assign n10900 = ( n10898 & ~n10469 ) | ( n10898 & n10899 ) | ( ~n10469 & n10899 ) ;
  assign n10904 = n10499 | n1748 ;
  assign n10901 = n1940 | n10015 ;
  assign n10902 = n1875 | n10486 ;
  assign n10903 = n10901 &  n10902 ;
  assign n10905 = ( n1748 & ~n10904 ) | ( n1748 & n10903 ) | ( ~n10904 & n10903 ) ;
  assign n10906 = ( n4740 & ~n3624 ) | ( n4740 & n10017 ) | ( ~n3624 & n10017 ) ;
  assign n10907 = ( n4742 & n10905 ) | ( n4742 & n10906 ) | ( n10905 & n10906 ) ;
  assign n10908 = x2 | n10907 ;
  assign n10909 = ( x2 & ~n10907 ) | ( x2 & 1'b0 ) | ( ~n10907 & 1'b0 ) ;
  assign n10910 = ( n10908 & ~x2 ) | ( n10908 & n10909 ) | ( ~x2 & n10909 ) ;
  assign n10911 = ( n10897 & n10900 ) | ( n10897 & n10910 ) | ( n10900 & n10910 ) ;
  assign n10549 = ( n10183 & n10193 ) | ( n10183 & n10470 ) | ( n10193 & n10470 ) ;
  assign n10550 = ( n10183 & ~n10470 ) | ( n10183 & n10193 ) | ( ~n10470 & n10193 ) ;
  assign n10551 = ( n10470 & ~n10549 ) | ( n10470 & n10550 ) | ( ~n10549 & n10550 ) ;
  assign n10915 = ~n1875 & n10015 ;
  assign n10912 = ~n1671 & n10499 ;
  assign n10913 = n1748 | n10486 ;
  assign n10914 = ~n10912 & n10913 ;
  assign n10916 = ( n1875 & n10915 ) | ( n1875 & n10914 ) | ( n10915 & n10914 ) ;
  assign n10917 = ( n4577 & ~n3625 ) | ( n4577 & n10017 ) | ( ~n3625 & n10017 ) ;
  assign n10918 = ( n4579 & n10916 ) | ( n4579 & n10917 ) | ( n10916 & n10917 ) ;
  assign n10919 = x2 | n10918 ;
  assign n10920 = ( x2 & ~n10918 ) | ( x2 & 1'b0 ) | ( ~n10918 & 1'b0 ) ;
  assign n10921 = ( n10919 & ~x2 ) | ( n10919 & n10920 ) | ( ~x2 & n10920 ) ;
  assign n10922 = ( n10911 & ~n10551 ) | ( n10911 & n10921 ) | ( ~n10551 & n10921 ) ;
  assign n10923 = n1566 &  n10499 ;
  assign n10924 = n1748 | n10015 ;
  assign n10925 = n1671 | n10486 ;
  assign n10926 = n10924 &  n10925 ;
  assign n10927 = ( n10923 & ~n10499 ) | ( n10923 & n10926 ) | ( ~n10499 & n10926 ) ;
  assign n10928 = ( n4594 & ~n3626 ) | ( n4594 & n10017 ) | ( ~n3626 & n10017 ) ;
  assign n10929 = ( n4596 & n10927 ) | ( n4596 & n10928 ) | ( n10927 & n10928 ) ;
  assign n10931 = x2 &  n10929 ;
  assign n10930 = ~x2 & n10929 ;
  assign n10932 = ( x2 & ~n10931 ) | ( x2 & n10930 ) | ( ~n10931 & n10930 ) ;
  assign n10933 = n5381 | n9155 ;
  assign n10934 = n10172 &  n10933 ;
  assign n10935 = ( n10180 & ~x5 ) | ( n10180 & n10934 ) | ( ~x5 & n10934 ) ;
  assign n10936 = ( x5 & ~n10934 ) | ( x5 & n10180 ) | ( ~n10934 & n10180 ) ;
  assign n10937 = ( n10935 & ~n10180 ) | ( n10935 & n10936 ) | ( ~n10180 & n10936 ) ;
  assign n10938 = ~n10471 & n10937 ;
  assign n10939 = ( n10471 & ~n10937 ) | ( n10471 & 1'b0 ) | ( ~n10937 & 1'b0 ) ;
  assign n10940 = n10938 | n10939 ;
  assign n10941 = ( n10922 & n10932 ) | ( n10922 & n10940 ) | ( n10932 & n10940 ) ;
  assign n10947 = ( n3627 & ~n10017 ) | ( n3627 & n4271 ) | ( ~n10017 & n4271 ) ;
  assign n10945 = ~n10499 & n1483 ;
  assign n10942 = n1671 | n10015 ;
  assign n10943 = n1566 | n10486 ;
  assign n10944 = n10942 &  n10943 ;
  assign n10946 = ( n10945 & ~n1483 ) | ( n10945 & n10944 ) | ( ~n1483 & n10944 ) ;
  assign n10948 = ( n4273 & ~n10947 ) | ( n4273 & n10946 ) | ( ~n10947 & n10946 ) ;
  assign n10950 = x2 &  n10948 ;
  assign n10949 = ~x2 & n10948 ;
  assign n10951 = ( x2 & ~n10950 ) | ( x2 & n10949 ) | ( ~n10950 & n10949 ) ;
  assign n10952 = n4743 | n9155 ;
  assign n10953 = n10159 &  n10952 ;
  assign n10954 = ( n10167 & ~x5 ) | ( n10167 & n10953 ) | ( ~x5 & n10953 ) ;
  assign n10955 = ( x5 & ~n10953 ) | ( x5 & n10167 ) | ( ~n10953 & n10167 ) ;
  assign n10956 = ( n10954 & ~n10167 ) | ( n10954 & n10955 ) | ( ~n10167 & n10955 ) ;
  assign n10957 = n10472 | n10956 ;
  assign n10958 = n10472 &  n10956 ;
  assign n10959 = ( n10957 & ~n10958 ) | ( n10957 & 1'b0 ) | ( ~n10958 & 1'b0 ) ;
  assign n10960 = ( n10941 & n10951 ) | ( n10941 & n10959 ) | ( n10951 & n10959 ) ;
  assign n10971 = n4580 | n9155 ;
  assign n10972 = n10146 &  n10971 ;
  assign n10973 = ( n10154 & ~x5 ) | ( n10154 & n10972 ) | ( ~x5 & n10972 ) ;
  assign n10974 = ( x5 & ~n10972 ) | ( x5 & n10154 ) | ( ~n10972 & n10154 ) ;
  assign n10975 = ( n10973 & ~n10154 ) | ( n10973 & n10974 ) | ( ~n10154 & n10974 ) ;
  assign n10976 = ~n10473 & n10975 ;
  assign n10977 = ( n10473 & ~n10975 ) | ( n10473 & 1'b0 ) | ( ~n10975 & 1'b0 ) ;
  assign n10978 = n10976 | n10977 ;
  assign n10966 = ( n3628 & ~n10017 ) | ( n3628 & n4631 ) | ( ~n10017 & n4631 ) ;
  assign n10961 = ~n1378 & n10499 ;
  assign n10962 = n1566 | n10015 ;
  assign n10963 = ~n10961 & n10962 ;
  assign n10964 = n1483 &  n10486 ;
  assign n10965 = ( n10963 & ~n1483 ) | ( n10963 & n10964 ) | ( ~n1483 & n10964 ) ;
  assign n10967 = ( n4632 & ~n10966 ) | ( n4632 & n10965 ) | ( ~n10966 & n10965 ) ;
  assign n10969 = x2 &  n10967 ;
  assign n10968 = ~x2 & n10967 ;
  assign n10970 = ( x2 & ~n10969 ) | ( x2 & n10968 ) | ( ~n10969 & n10968 ) ;
  assign n10979 = ( n10960 & ~n10978 ) | ( n10960 & n10970 ) | ( ~n10978 & n10970 ) ;
  assign n10980 = ( n10141 & ~n10131 ) | ( n10141 & n10474 ) | ( ~n10131 & n10474 ) ;
  assign n10981 = ( n10131 & ~n10141 ) | ( n10131 & n10474 ) | ( ~n10141 & n10474 ) ;
  assign n10982 = ( n10980 & ~n10474 ) | ( n10980 & n10981 ) | ( ~n10474 & n10981 ) ;
  assign n10988 = ( n3629 & ~n10017 ) | ( n3629 & n4419 ) | ( ~n10017 & n4419 ) ;
  assign n10986 = ~n10499 & n1267 ;
  assign n10983 = ( n1483 & ~n10015 ) | ( n1483 & 1'b0 ) | ( ~n10015 & 1'b0 ) ;
  assign n10984 = n1378 | n10486 ;
  assign n10985 = ~n10983 & n10984 ;
  assign n10987 = ( n10986 & ~n1267 ) | ( n10986 & n10985 ) | ( ~n1267 & n10985 ) ;
  assign n10989 = ( n4421 & ~n10988 ) | ( n4421 & n10987 ) | ( ~n10988 & n10987 ) ;
  assign n10990 = x2 | n10989 ;
  assign n10991 = ( x2 & ~n10989 ) | ( x2 & 1'b0 ) | ( ~n10989 & 1'b0 ) ;
  assign n10992 = ( n10990 & ~x2 ) | ( n10990 & n10991 ) | ( ~x2 & n10991 ) ;
  assign n10993 = ( n10979 & n10982 ) | ( n10979 & n10992 ) | ( n10982 & n10992 ) ;
  assign n10999 = ( n3630 & ~n10017 ) | ( n3630 & n4058 ) | ( ~n10017 & n4058 ) ;
  assign n10994 = ~n1151 & n10499 ;
  assign n10995 = n1378 | n10015 ;
  assign n10996 = ~n10994 & n10995 ;
  assign n10997 = n1267 &  n10486 ;
  assign n10998 = ( n10996 & ~n1267 ) | ( n10996 & n10997 ) | ( ~n1267 & n10997 ) ;
  assign n11000 = ( n4060 & ~n10999 ) | ( n4060 & n10998 ) | ( ~n10999 & n10998 ) ;
  assign n11001 = x2 | n11000 ;
  assign n11002 = ( x2 & ~n11000 ) | ( x2 & 1'b0 ) | ( ~n11000 & 1'b0 ) ;
  assign n11003 = ( n11001 & ~x2 ) | ( n11001 & n11002 ) | ( ~x2 & n11002 ) ;
  assign n11004 = ( n10548 & n10993 ) | ( n10548 & n11003 ) | ( n10993 & n11003 ) ;
  assign n11015 = ( n5038 & ~n9155 ) | ( n5038 & 1'b0 ) | ( ~n9155 & 1'b0 ) ;
  assign n11016 = ( n10107 & ~n11015 ) | ( n10107 & 1'b0 ) | ( ~n11015 & 1'b0 ) ;
  assign n11017 = ( x5 & ~n11016 ) | ( x5 & n10115 ) | ( ~n11016 & n10115 ) ;
  assign n11018 = ( n10115 & ~x5 ) | ( n10115 & n11016 ) | ( ~x5 & n11016 ) ;
  assign n11019 = ( n11017 & ~n10115 ) | ( n11017 & n11018 ) | ( ~n10115 & n11018 ) ;
  assign n11020 = n10476 | n11019 ;
  assign n11021 = n10476 &  n11019 ;
  assign n11022 = ( n11020 & ~n11021 ) | ( n11020 & 1'b0 ) | ( ~n11021 & 1'b0 ) ;
  assign n11005 = ~n1043 & n10499 ;
  assign n11006 = n1151 | n10486 ;
  assign n11007 = ~n11005 & n11006 ;
  assign n11008 = n1267 &  n10015 ;
  assign n11009 = ( n11007 & ~n1267 ) | ( n11007 & n11008 ) | ( ~n1267 & n11008 ) ;
  assign n11010 = ( n3949 & ~n3631 ) | ( n3949 & n10017 ) | ( ~n3631 & n10017 ) ;
  assign n11011 = ( n3951 & n11009 ) | ( n3951 & n11010 ) | ( n11009 & n11010 ) ;
  assign n11013 = x2 &  n11011 ;
  assign n11012 = ~x2 & n11011 ;
  assign n11014 = ( x2 & ~n11013 ) | ( x2 & n11012 ) | ( ~n11013 & n11012 ) ;
  assign n11023 = ( n11004 & ~n11022 ) | ( n11004 & n11014 ) | ( ~n11022 & n11014 ) ;
  assign n11024 = ( n10545 & ~n10535 ) | ( n10545 & n11023 ) | ( ~n10535 & n11023 ) ;
  assign n11025 = ( n10523 & n10533 ) | ( n10523 & n11024 ) | ( n10533 & n11024 ) ;
  assign n11026 = ( n10511 & n10521 ) | ( n10511 & n11025 ) | ( n10521 & n11025 ) ;
  assign n11027 = ( n10509 & ~n10498 ) | ( n10509 & n11026 ) | ( ~n10498 & n11026 ) ;
  assign n11028 = ( n10484 & n10496 ) | ( n10484 & n11027 ) | ( n10496 & n11027 ) ;
  assign n11029 = ( n10042 & n10482 ) | ( n10042 & n11028 ) | ( n10482 & n11028 ) ;
  assign n11030 = ( n10037 & ~n10040 ) | ( n10037 & n11029 ) | ( ~n10040 & n11029 ) ;
  assign n11031 = ( n10008 & ~n10010 ) | ( n10008 & n11030 ) | ( ~n10010 & n11030 ) ;
  assign n11032 = ( n9569 & ~n9174 ) | ( n9569 & n11031 ) | ( ~n9174 & n11031 ) ;
  assign n11033 = ( n9170 & ~n9172 ) | ( n9170 & n11032 ) | ( ~n9172 & n11032 ) ;
  assign n11034 = ( n8787 & ~n8790 ) | ( n8787 & n11033 ) | ( ~n8790 & n11033 ) ;
  assign n11035 = ( n8440 & ~n8120 ) | ( n8440 & n11034 ) | ( ~n8120 & n11034 ) ;
  assign n11036 = ( n7812 & n8117 ) | ( n7812 & n11035 ) | ( n8117 & n11035 ) ;
  assign n11037 = ( n7806 & ~n7809 ) | ( n7806 & n11036 ) | ( ~n7809 & n11036 ) ;
  assign n11038 = ( n7530 & ~n7270 ) | ( n7530 & n11037 ) | ( ~n7270 & n11037 ) ;
  assign n11039 = ( n7265 & n7267 ) | ( n7265 & n11038 ) | ( n7267 & n11038 ) ;
  assign n11040 = ( n7122 & ~n7125 ) | ( n7122 & n11039 ) | ( ~n7125 & n11039 ) ;
  assign n11041 = ( n6995 & ~n6547 ) | ( n6995 & n11040 ) | ( ~n6547 & n11040 ) ;
  assign n11042 = ( n6542 & n6544 ) | ( n6542 & n11041 ) | ( n6544 & n11041 ) ;
  assign n11043 = ( n6419 & ~n6181 ) | ( n6419 & n11042 ) | ( ~n6181 & n11042 ) ;
  assign n11044 = ( n6179 & ~n5986 ) | ( n6179 & n11043 ) | ( ~n5986 & n11043 ) ;
  assign n11045 = ( n5981 & n5983 ) | ( n5981 & n11044 ) | ( n5983 & n11044 ) ;
  assign n11046 = ( n5861 & ~n5773 ) | ( n5861 & n11045 ) | ( ~n5773 & n11045 ) ;
  assign n11047 = ( n5769 & ~n5353 ) | ( n5769 & n11046 ) | ( ~n5353 & n11046 ) ;
  assign n11048 = ( n5168 & n5350 ) | ( n5168 & n11047 ) | ( n5350 & n11047 ) ;
  assign n11049 = ( n5159 & n5165 ) | ( n5159 & n11048 ) | ( n5165 & n11048 ) ;
  assign n11050 = ( n5020 & n5075 ) | ( n5020 & n11049 ) | ( n5075 & n11049 ) ;
  assign n11051 = ( n4973 & n4999 ) | ( n4973 & n5017 ) | ( n4999 & n5017 ) ;
  assign n11052 = ( n4983 & n4986 ) | ( n4983 & n4996 ) | ( n4986 & n4996 ) ;
  assign n11053 = ( n4505 & ~n4638 ) | ( n4505 & n4648 ) | ( ~n4638 & n4648 ) ;
  assign n11054 = ( n4638 & ~n4649 ) | ( n4638 & n11053 ) | ( ~n4649 & n11053 ) ;
  assign n11058 = ~n863 & n4482 ;
  assign n11055 = n599 | n4962 ;
  assign n11056 = n702 | n4495 ;
  assign n11057 = n11055 &  n11056 ;
  assign n11059 = ( n863 & n11058 ) | ( n863 & n11057 ) | ( n11058 & n11057 ) ;
  assign n11060 = ( n4452 & ~n4478 ) | ( n4452 & n11059 ) | ( ~n4478 & n11059 ) ;
  assign n11061 = ~n4452 & n11060 ;
  assign n11062 = ( x26 & ~n11059 ) | ( x26 & n11061 ) | ( ~n11059 & n11061 ) ;
  assign n11063 = ( n11059 & ~x26 ) | ( n11059 & n11061 ) | ( ~x26 & n11061 ) ;
  assign n11064 = ( n11062 & ~n11061 ) | ( n11062 & n11063 ) | ( ~n11061 & n11063 ) ;
  assign n11065 = ( n11052 & ~n11054 ) | ( n11052 & n11064 ) | ( ~n11054 & n11064 ) ;
  assign n11066 = ( n11052 & ~n11064 ) | ( n11052 & n11054 ) | ( ~n11064 & n11054 ) ;
  assign n11067 = ( n11065 & ~n11052 ) | ( n11065 & n11066 ) | ( ~n11052 & n11066 ) ;
  assign n11068 = ( n11050 & n11051 ) | ( n11050 & n11067 ) | ( n11051 & n11067 ) ;
  assign n11069 = ( n11052 & n11054 ) | ( n11052 & n11064 ) | ( n11054 & n11064 ) ;
  assign n11070 = ( n4502 & ~n4649 ) | ( n4502 & n4652 ) | ( ~n4649 & n4652 ) ;
  assign n11071 = ( n4649 & ~n4653 ) | ( n4649 & n11070 ) | ( ~n4653 & n11070 ) ;
  assign n11072 = ( n11068 & n11069 ) | ( n11068 & n11071 ) | ( n11069 & n11071 ) ;
  assign n11073 = ( n4493 & n4653 ) | ( n4493 & n11072 ) | ( n4653 & n11072 ) ;
  assign n11074 = ( n4491 & ~n4461 ) | ( n4491 & n11073 ) | ( ~n4461 & n11073 ) ;
  assign n11075 = ( n4458 & ~n4053 ) | ( n4458 & n11074 ) | ( ~n4053 & n11074 ) ;
  assign n3944 = x29 | n3943 ;
  assign n3945 = x29 &  n3943 ;
  assign n3946 = ( n3944 & ~n3945 ) | ( n3944 & 1'b0 ) | ( ~n3945 & 1'b0 ) ;
  assign n4047 = ( n3946 & ~n3931 ) | ( n3946 & n4046 ) | ( ~n3931 & n4046 ) ;
  assign n11076 = ( n3928 & ~n11075 ) | ( n3928 & n4047 ) | ( ~n11075 & n4047 ) ;
  assign n11077 = ( n3928 & ~n4047 ) | ( n3928 & n11075 ) | ( ~n4047 & n11075 ) ;
  assign n11078 = ( n3928 & ~n11076 ) | ( n3928 & ~n11077 ) | ( ~n11076 & ~n11077 ) ;
  assign n11083 = ( n4053 & n4458 ) | ( n4053 & n11074 ) | ( n4458 & n11074 ) ;
  assign n11084 = ( n4053 & ~n4458 ) | ( n4053 & n11074 ) | ( ~n4458 & n11074 ) ;
  assign n11085 = ( ~n4458 & n11083 ) | ( ~n4458 & ~n11084 ) | ( n11083 & ~n11084 ) ;
  assign n11079 = ( n4461 & n4491 ) | ( n4461 & n11073 ) | ( n4491 & n11073 ) ;
  assign n11080 = ( n4461 & ~n4491 ) | ( n4461 & n11073 ) | ( ~n4491 & n11073 ) ;
  assign n11081 = ( ~n4491 & n11079 ) | ( ~n4491 & ~n11080 ) | ( n11079 & ~n11080 ) ;
  assign n11090 = ( n4493 & ~n4653 ) | ( n4493 & n11072 ) | ( ~n4653 & n11072 ) ;
  assign n11091 = ( n4653 & ~n11073 ) | ( n4653 & n11090 ) | ( ~n11073 & n11090 ) ;
  assign n11092 = ( n11068 & ~n11069 ) | ( n11068 & n11071 ) | ( ~n11069 & n11071 ) ;
  assign n11093 = ( n11069 & ~n11072 ) | ( n11069 & n11092 ) | ( ~n11072 & n11092 ) ;
  assign n11094 = ( n11050 & ~n11051 ) | ( n11050 & n11067 ) | ( ~n11051 & n11067 ) ;
  assign n11095 = ( n11051 & ~n11068 ) | ( n11051 & n11094 ) | ( ~n11068 & n11094 ) ;
  assign n11096 = ( n5075 & ~n5020 ) | ( n5075 & n11049 ) | ( ~n5020 & n11049 ) ;
  assign n11097 = ( n5020 & ~n11049 ) | ( n5020 & n5075 ) | ( ~n11049 & n5075 ) ;
  assign n11098 = ( ~n5075 & n11096 ) | ( ~n5075 & n11097 ) | ( n11096 & n11097 ) ;
  assign n11099 = ( n5159 & ~n11048 ) | ( n5159 & n5165 ) | ( ~n11048 & n5165 ) ;
  assign n11100 = ( n5165 & ~n5159 ) | ( n5165 & n11048 ) | ( ~n5159 & n11048 ) ;
  assign n11101 = ( ~n5165 & n11099 ) | ( ~n5165 & n11100 ) | ( n11099 & n11100 ) ;
  assign n11102 = ( n5350 & ~n5168 ) | ( n5350 & n11047 ) | ( ~n5168 & n11047 ) ;
  assign n11103 = ( n5168 & ~n11047 ) | ( n5168 & n5350 ) | ( ~n11047 & n5350 ) ;
  assign n11104 = ( n11102 & ~n5350 ) | ( n11102 & n11103 ) | ( ~n5350 & n11103 ) ;
  assign n11105 = ( n5353 & n5769 ) | ( n5353 & n11046 ) | ( n5769 & n11046 ) ;
  assign n11106 = ( n5353 & ~n5769 ) | ( n5353 & n11046 ) | ( ~n5769 & n11046 ) ;
  assign n11107 = ( n5769 & ~n11105 ) | ( n5769 & n11106 ) | ( ~n11105 & n11106 ) ;
  assign n11108 = ( n5773 & n5861 ) | ( n5773 & n11045 ) | ( n5861 & n11045 ) ;
  assign n11109 = ( n5773 & ~n5861 ) | ( n5773 & n11045 ) | ( ~n5861 & n11045 ) ;
  assign n11110 = ( ~n5861 & n11108 ) | ( ~n5861 & ~n11109 ) | ( n11108 & ~n11109 ) ;
  assign n11114 = ( n5986 & n6179 ) | ( n5986 & n11043 ) | ( n6179 & n11043 ) ;
  assign n11115 = ( n5986 & ~n6179 ) | ( n5986 & n11043 ) | ( ~n6179 & n11043 ) ;
  assign n11116 = ( n6179 & ~n11114 ) | ( n6179 & n11115 ) | ( ~n11114 & n11115 ) ;
  assign n11111 = ( n5981 & ~n11044 ) | ( n5981 & n5983 ) | ( ~n11044 & n5983 ) ;
  assign n11112 = ( n5983 & ~n5981 ) | ( n5983 & n11044 ) | ( ~n5981 & n11044 ) ;
  assign n11113 = ( n11111 & ~n5983 ) | ( n11111 & n11112 ) | ( ~n5983 & n11112 ) ;
  assign n11120 = ( n6542 & ~n11041 ) | ( n6542 & n6544 ) | ( ~n11041 & n6544 ) ;
  assign n11121 = ( n6544 & ~n6542 ) | ( n6544 & n11041 ) | ( ~n6542 & n11041 ) ;
  assign n11122 = ( ~n6544 & n11120 ) | ( ~n6544 & n11121 ) | ( n11120 & n11121 ) ;
  assign n11117 = ( n6181 & n6419 ) | ( n6181 & n11042 ) | ( n6419 & n11042 ) ;
  assign n11118 = ( n6181 & ~n6419 ) | ( n6181 & n11042 ) | ( ~n6419 & n11042 ) ;
  assign n11119 = ( n6419 & ~n11117 ) | ( n6419 & n11118 ) | ( ~n11117 & n11118 ) ;
  assign n11123 = ( n6547 & n6995 ) | ( n6547 & n11040 ) | ( n6995 & n11040 ) ;
  assign n11124 = ( n6547 & ~n6995 ) | ( n6547 & n11040 ) | ( ~n6995 & n11040 ) ;
  assign n11125 = ( n6995 & ~n11123 ) | ( n6995 & n11124 ) | ( ~n11123 & n11124 ) ;
  assign n11126 = ( n7125 & ~n7122 ) | ( n7125 & n11039 ) | ( ~n7122 & n11039 ) ;
  assign n11127 = ( n7122 & ~n11039 ) | ( n7122 & n7125 ) | ( ~n11039 & n7125 ) ;
  assign n11128 = ( n7125 & ~n11126 ) | ( n7125 & ~n11127 ) | ( ~n11126 & ~n11127 ) ;
  assign n11129 = ( n7265 & ~n11038 ) | ( n7265 & n7267 ) | ( ~n11038 & n7267 ) ;
  assign n11130 = ( n7267 & ~n7265 ) | ( n7267 & n11038 ) | ( ~n7265 & n11038 ) ;
  assign n11131 = ( n11129 & ~n7267 ) | ( n11129 & n11130 ) | ( ~n7267 & n11130 ) ;
  assign n11132 = ( n7270 & n7530 ) | ( n7270 & n11037 ) | ( n7530 & n11037 ) ;
  assign n11133 = ( n7270 & ~n7530 ) | ( n7270 & n11037 ) | ( ~n7530 & n11037 ) ;
  assign n11134 = ( n7530 & ~n11132 ) | ( n7530 & n11133 ) | ( ~n11132 & n11133 ) ;
  assign n11135 = ( n7809 & ~n7806 ) | ( n7809 & n11036 ) | ( ~n7806 & n11036 ) ;
  assign n11136 = ( n7806 & ~n11036 ) | ( n7806 & n7809 ) | ( ~n11036 & n7809 ) ;
  assign n11137 = ( n7809 & ~n11135 ) | ( n7809 & ~n11136 ) | ( ~n11135 & ~n11136 ) ;
  assign n11138 = ( n8117 & ~n7812 ) | ( n8117 & n11035 ) | ( ~n7812 & n11035 ) ;
  assign n11139 = ( n7812 & ~n11035 ) | ( n7812 & n8117 ) | ( ~n11035 & n8117 ) ;
  assign n11140 = ( ~n8117 & n11138 ) | ( ~n8117 & n11139 ) | ( n11138 & n11139 ) ;
  assign n11141 = ( n8120 & n8440 ) | ( n8120 & n11034 ) | ( n8440 & n11034 ) ;
  assign n11142 = ( n8120 & ~n8440 ) | ( n8120 & n11034 ) | ( ~n8440 & n11034 ) ;
  assign n11143 = ( ~n8440 & n11141 ) | ( ~n8440 & ~n11142 ) | ( n11141 & ~n11142 ) ;
  assign n11144 = ( n8790 & ~n8787 ) | ( n8790 & n11033 ) | ( ~n8787 & n11033 ) ;
  assign n11145 = ( n8787 & ~n11033 ) | ( n8787 & n8790 ) | ( ~n11033 & n8790 ) ;
  assign n11146 = ( n8790 & ~n11144 ) | ( n8790 & ~n11145 ) | ( ~n11144 & ~n11145 ) ;
  assign n11150 = ( n9174 & n9569 ) | ( n9174 & n11031 ) | ( n9569 & n11031 ) ;
  assign n11151 = ( n9174 & ~n9569 ) | ( n9174 & n11031 ) | ( ~n9569 & n11031 ) ;
  assign n11152 = ( n9569 & ~n11150 ) | ( n9569 & n11151 ) | ( ~n11150 & n11151 ) ;
  assign n11147 = ( n9172 & ~n9170 ) | ( n9172 & n11032 ) | ( ~n9170 & n11032 ) ;
  assign n11148 = ( n9170 & ~n11032 ) | ( n9170 & n9172 ) | ( ~n11032 & n9172 ) ;
  assign n11149 = ( n9172 & ~n11147 ) | ( n9172 & ~n11148 ) | ( ~n11147 & ~n11148 ) ;
  assign n11153 = ( n10010 & ~n10008 ) | ( n10010 & n11030 ) | ( ~n10008 & n11030 ) ;
  assign n11154 = ( n10008 & ~n11030 ) | ( n10008 & n10010 ) | ( ~n11030 & n10010 ) ;
  assign n11155 = ( n11153 & ~n10010 ) | ( n11153 & n11154 ) | ( ~n10010 & n11154 ) ;
  assign n11159 = ( n10482 & ~n10042 ) | ( n10482 & n11028 ) | ( ~n10042 & n11028 ) ;
  assign n11160 = ( n10042 & ~n11028 ) | ( n10042 & n10482 ) | ( ~n11028 & n10482 ) ;
  assign n11161 = ( ~n10482 & n11159 ) | ( ~n10482 & n11160 ) | ( n11159 & n11160 ) ;
  assign n11156 = ( n10040 & ~n10037 ) | ( n10040 & n11029 ) | ( ~n10037 & n11029 ) ;
  assign n11157 = ( n10037 & ~n11029 ) | ( n10037 & n10040 ) | ( ~n11029 & n10040 ) ;
  assign n11158 = ( n11156 & ~n10040 ) | ( n11156 & n11157 ) | ( ~n10040 & n11157 ) ;
  assign n11162 = ( n10496 & ~n10484 ) | ( n10496 & n11027 ) | ( ~n10484 & n11027 ) ;
  assign n11163 = ( n10484 & ~n10496 ) | ( n10484 & n11027 ) | ( ~n10496 & n11027 ) ;
  assign n11164 = ( n11162 & ~n11027 ) | ( n11162 & n11163 ) | ( ~n11027 & n11163 ) ;
  assign n11165 = ( n10498 & ~n11026 ) | ( n10498 & n10509 ) | ( ~n11026 & n10509 ) ;
  assign n11166 = ( n10509 & ~n11027 ) | ( n10509 & ~n11165 ) | ( ~n11027 & ~n11165 ) ;
  assign n11167 = ( n10511 & ~n10521 ) | ( n10511 & n11025 ) | ( ~n10521 & n11025 ) ;
  assign n11168 = ( n10521 & ~n11026 ) | ( n10521 & n11167 ) | ( ~n11026 & n11167 ) ;
  assign n11169 = ( n10535 & ~n11023 ) | ( n10535 & n10545 ) | ( ~n11023 & n10545 ) ;
  assign n11170 = ( n11024 & ~n10545 ) | ( n11024 & n11169 ) | ( ~n10545 & n11169 ) ;
  assign n11173 = n11170 &  n11168 ;
  assign n11171 = ( n10523 & ~n10533 ) | ( n10523 & n11024 ) | ( ~n10533 & n11024 ) ;
  assign n11172 = ( n10533 & ~n11025 ) | ( n10533 & n11171 ) | ( ~n11025 & n11171 ) ;
  assign n11174 = ( n11168 & ~n11173 ) | ( n11168 & n11172 ) | ( ~n11173 & n11172 ) ;
  assign n11175 = ( n11166 & n11168 ) | ( n11166 & n11174 ) | ( n11168 & n11174 ) ;
  assign n11176 = ( n11164 & n11166 ) | ( n11164 & n11175 ) | ( n11166 & n11175 ) ;
  assign n11177 = ( n11161 & n11164 ) | ( n11161 & n11176 ) | ( n11164 & n11176 ) ;
  assign n11178 = ( n11161 & ~n11158 ) | ( n11161 & n11177 ) | ( ~n11158 & n11177 ) ;
  assign n11179 = ( n11155 & ~n11178 ) | ( n11155 & n11158 ) | ( ~n11178 & n11158 ) ;
  assign n11180 = ( n11152 & n11155 ) | ( n11152 & n11179 ) | ( n11155 & n11179 ) ;
  assign n11181 = ( n11152 & ~n11149 ) | ( n11152 & n11180 ) | ( ~n11149 & n11180 ) ;
  assign n11182 = ( n11146 & ~n11181 ) | ( n11146 & n11149 ) | ( ~n11181 & n11149 ) ;
  assign n11183 = ( n11143 & n11146 ) | ( n11143 & n11182 ) | ( n11146 & n11182 ) ;
  assign n11184 = ( n11140 & n11143 ) | ( n11140 & n11183 ) | ( n11143 & n11183 ) ;
  assign n11185 = ( n11137 & n11140 ) | ( n11137 & n11184 ) | ( n11140 & n11184 ) ;
  assign n11186 = ( n11137 & ~n11134 ) | ( n11137 & n11185 ) | ( ~n11134 & n11185 ) ;
  assign n11187 = ( n11131 & ~n11134 ) | ( n11131 & n11186 ) | ( ~n11134 & n11186 ) ;
  assign n11188 = ( n11128 & n11131 ) | ( n11128 & n11187 ) | ( n11131 & n11187 ) ;
  assign n11189 = ( n11128 & ~n11125 ) | ( n11128 & n11188 ) | ( ~n11125 & n11188 ) ;
  assign n11190 = ( n11122 & ~n11125 ) | ( n11122 & n11189 ) | ( ~n11125 & n11189 ) ;
  assign n11191 = ( n11122 & ~n11119 ) | ( n11122 & n11190 ) | ( ~n11119 & n11190 ) ;
  assign n11192 = ( n11116 & ~n11191 ) | ( n11116 & n11119 ) | ( ~n11191 & n11119 ) ;
  assign n11193 = ( n11116 & ~n11113 ) | ( n11116 & n11192 ) | ( ~n11113 & n11192 ) ;
  assign n11194 = ( n11110 & ~n11193 ) | ( n11110 & n11113 ) | ( ~n11193 & n11113 ) ;
  assign n11195 = ( n11110 & ~n11107 ) | ( n11110 & n11194 ) | ( ~n11107 & n11194 ) ;
  assign n11196 = ( n11104 & ~n11107 ) | ( n11104 & n11195 ) | ( ~n11107 & n11195 ) ;
  assign n11197 = ( n11101 & n11104 ) | ( n11101 & n11196 ) | ( n11104 & n11196 ) ;
  assign n11198 = ( n11098 & n11101 ) | ( n11098 & n11197 ) | ( n11101 & n11197 ) ;
  assign n11199 = ( n11095 & n11098 ) | ( n11095 & n11198 ) | ( n11098 & n11198 ) ;
  assign n11200 = ( n11093 & n11095 ) | ( n11093 & n11199 ) | ( n11095 & n11199 ) ;
  assign n11201 = ( n11091 & n11093 ) | ( n11091 & n11200 ) | ( n11093 & n11200 ) ;
  assign n11202 = ( n11081 & n11091 ) | ( n11081 & n11201 ) | ( n11091 & n11201 ) ;
  assign n11203 = ( n11081 & n11085 ) | ( n11081 & n11202 ) | ( n11085 & n11202 ) ;
  assign n11205 = ( n11078 & n11085 ) | ( n11078 & n11203 ) | ( n11085 & n11203 ) ;
  assign n11204 = ( n11085 & ~n11078 ) | ( n11085 & n11203 ) | ( ~n11078 & n11203 ) ;
  assign n11206 = ( n11078 & ~n11205 ) | ( n11078 & n11204 ) | ( ~n11205 & n11204 ) ;
  assign n11082 = n10015 | n11081 ;
  assign n11086 = n10486 | n11085 ;
  assign n11087 = n11082 &  n11086 ;
  assign n11088 = n10499 &  n11078 ;
  assign n11089 = ( n11087 & ~n10499 ) | ( n11087 & n11088 ) | ( ~n10499 & n11088 ) ;
  assign n11207 = ( n11089 & ~n10017 ) | ( n11089 & n11206 ) | ( ~n10017 & n11206 ) ;
  assign n11208 = ~n11206 & n11207 ;
  assign n11210 = ( x2 & n11089 ) | ( x2 & n11208 ) | ( n11089 & n11208 ) ;
  assign n11209 = ( x2 & ~n11208 ) | ( x2 & n11089 ) | ( ~n11208 & n11089 ) ;
  assign n11211 = ( n11208 & ~n11210 ) | ( n11208 & n11209 ) | ( ~n11210 & n11209 ) ;
  assign n11217 = ( n11098 & ~n11101 ) | ( n11098 & n11197 ) | ( ~n11101 & n11197 ) ;
  assign n11218 = ( n11101 & ~n11198 ) | ( n11101 & n11217 ) | ( ~n11198 & n11217 ) ;
  assign n11212 = ( n8105 & ~n11104 ) | ( n8105 & 1'b0 ) | ( ~n11104 & 1'b0 ) ;
  assign n11213 = n8429 | n11101 ;
  assign n11214 = ~n11212 & n11213 ;
  assign n11215 = ~n8764 & n11098 ;
  assign n11216 = ( n8764 & n11214 ) | ( n8764 & n11215 ) | ( n11214 & n11215 ) ;
  assign n11219 = ( n11216 & ~n8107 ) | ( n11216 & n11218 ) | ( ~n8107 & n11218 ) ;
  assign n11220 = ~n11218 & n11219 ;
  assign n11222 = ( x8 & n11216 ) | ( x8 & n11220 ) | ( n11216 & n11220 ) ;
  assign n11221 = ( x8 & ~n11220 ) | ( x8 & n11216 ) | ( ~n11220 & n11216 ) ;
  assign n11223 = ( n11220 & ~n11222 ) | ( n11220 & n11221 ) | ( ~n11222 & n11221 ) ;
  assign n11227 = n11116 | n7097 ;
  assign n11224 = n6530 | n11122 ;
  assign n11225 = ~n6983 & n11119 ;
  assign n11226 = ( n11224 & ~n11225 ) | ( n11224 & 1'b0 ) | ( ~n11225 & 1'b0 ) ;
  assign n11228 = ( n7097 & ~n11227 ) | ( n7097 & n11226 ) | ( ~n11227 & n11226 ) ;
  assign n11229 = ( n11119 & ~n11116 ) | ( n11119 & n11191 ) | ( ~n11116 & n11191 ) ;
  assign n11230 = ( n11192 & ~n11119 ) | ( n11192 & n11229 ) | ( ~n11119 & n11229 ) ;
  assign n11231 = ( n11228 & ~n6532 ) | ( n11228 & n11230 ) | ( ~n6532 & n11230 ) ;
  assign n11232 = ~n11230 & n11231 ;
  assign n11233 = ( x14 & ~n11228 ) | ( x14 & n11232 ) | ( ~n11228 & n11232 ) ;
  assign n11234 = ( n11228 & ~x14 ) | ( n11228 & n11232 ) | ( ~x14 & n11232 ) ;
  assign n11235 = ( n11233 & ~n11232 ) | ( n11233 & n11234 ) | ( ~n11232 & n11234 ) ;
  assign n11241 = ( n11134 & ~n11185 ) | ( n11134 & n11137 ) | ( ~n11185 & n11137 ) ;
  assign n11242 = ( n11186 & ~n11137 ) | ( n11186 & n11241 ) | ( ~n11137 & n11241 ) ;
  assign n11239 = n11134 | n5837 ;
  assign n11236 = ( n5339 & ~n11140 ) | ( n5339 & 1'b0 ) | ( ~n11140 & 1'b0 ) ;
  assign n11237 = n5761 | n11137 ;
  assign n11238 = ~n11236 & n11237 ;
  assign n11240 = ( n5837 & ~n11239 ) | ( n5837 & n11238 ) | ( ~n11239 & n11238 ) ;
  assign n11243 = ( n5341 & ~n11240 ) | ( n5341 & n11242 ) | ( ~n11240 & n11242 ) ;
  assign n11244 = ( n11242 & ~n11243 ) | ( n11242 & 1'b0 ) | ( ~n11243 & 1'b0 ) ;
  assign n11246 = ( x20 & n11240 ) | ( x20 & n11244 ) | ( n11240 & n11244 ) ;
  assign n11245 = ( x20 & ~n11244 ) | ( x20 & n11240 ) | ( ~n11244 & n11240 ) ;
  assign n11247 = ( n11244 & ~n11246 ) | ( n11244 & n11245 ) | ( ~n11246 & n11245 ) ;
  assign n11251 = n11152 | n4962 ;
  assign n11248 = ~n4495 & n11155 ;
  assign n11249 = ~n4482 & n11158 ;
  assign n11250 = n11248 | n11249 ;
  assign n11252 = ( n11251 & ~n4962 ) | ( n11251 & n11250 ) | ( ~n4962 & n11250 ) ;
  assign n11253 = ( n11152 & ~n11155 ) | ( n11152 & n11179 ) | ( ~n11155 & n11179 ) ;
  assign n11254 = ( n11155 & ~n11180 ) | ( n11155 & n11253 ) | ( ~n11180 & n11253 ) ;
  assign n11255 = ( n4478 & n11252 ) | ( n4478 & n11254 ) | ( n11252 & n11254 ) ;
  assign n11256 = ( n11254 & ~n11255 ) | ( n11254 & 1'b0 ) | ( ~n11255 & 1'b0 ) ;
  assign n11257 = ( n11252 & ~x26 ) | ( n11252 & n11256 ) | ( ~x26 & n11256 ) ;
  assign n11258 = ( x26 & ~n11252 ) | ( x26 & n11256 ) | ( ~n11252 & n11256 ) ;
  assign n11259 = ( n11257 & ~n11256 ) | ( n11257 & n11258 ) | ( ~n11256 & n11258 ) ;
  assign n11354 = n2332 | n2548 ;
  assign n11355 = ( n3015 & ~n11354 ) | ( n3015 & n3243 ) | ( ~n11354 & n3243 ) ;
  assign n11356 = ~n3015 & n11355 ;
  assign n11357 = ( n11356 & ~n1017 ) | ( n11356 & n2914 ) | ( ~n1017 & n2914 ) ;
  assign n11358 = ( n11357 & ~n2914 ) | ( n11357 & 1'b0 ) | ( ~n2914 & 1'b0 ) ;
  assign n11359 = ( n2943 & ~n6770 ) | ( n2943 & n11358 ) | ( ~n6770 & n11358 ) ;
  assign n11360 = ( n11359 & ~n2943 ) | ( n11359 & 1'b0 ) | ( ~n2943 & 1'b0 ) ;
  assign n11331 = n363 | n2110 ;
  assign n11332 = ( n258 & ~n349 ) | ( n258 & n11331 ) | ( ~n349 & n11331 ) ;
  assign n11333 = n349 | n11332 ;
  assign n11334 = ( n281 & ~n745 ) | ( n281 & n11333 ) | ( ~n745 & n11333 ) ;
  assign n11335 = n745 | n11334 ;
  assign n11336 = n276 | n11335 ;
  assign n11342 = n791 | n1192 ;
  assign n11343 = ( n3888 & ~n883 ) | ( n3888 & n11342 ) | ( ~n883 & n11342 ) ;
  assign n11344 = n883 | n11343 ;
  assign n11337 = ( n624 & ~n1877 ) | ( n624 & 1'b0 ) | ( ~n1877 & 1'b0 ) ;
  assign n11338 = ( n130 & ~n408 ) | ( n130 & n11337 ) | ( ~n408 & n11337 ) ;
  assign n11339 = ~n130 & n11338 ;
  assign n11340 = ( n236 & ~n43 ) | ( n236 & n11339 ) | ( ~n43 & n11339 ) ;
  assign n11341 = ~n236 & n11340 ;
  assign n11345 = ( n189 & ~n11344 ) | ( n189 & n11341 ) | ( ~n11344 & n11341 ) ;
  assign n11346 = ~n189 & n11345 ;
  assign n11347 = ( n1072 & ~n11336 ) | ( n1072 & n11346 ) | ( ~n11336 & n11346 ) ;
  assign n11348 = ~n1072 & n11347 ;
  assign n11349 = ( n457 & ~n605 ) | ( n457 & n11348 ) | ( ~n605 & n11348 ) ;
  assign n11350 = ~n457 & n11349 ;
  assign n11351 = ( n664 & ~n269 ) | ( n664 & n11350 ) | ( ~n269 & n11350 ) ;
  assign n11352 = ~n664 & n11351 ;
  assign n11353 = ~n431 & n11352 ;
  assign n11361 = ( n570 & ~n11360 ) | ( n570 & n11353 ) | ( ~n11360 & n11353 ) ;
  assign n11362 = ( n789 & ~n11361 ) | ( n789 & n11353 ) | ( ~n11361 & n11353 ) ;
  assign n11363 = ~n789 & n11362 ;
  assign n11364 = ( n524 & ~n11363 ) | ( n524 & n734 ) | ( ~n11363 & n734 ) ;
  assign n11365 = ( n524 & ~n11364 ) | ( n524 & 1'b0 ) | ( ~n11364 & 1'b0 ) ;
  assign n11366 = ( n77 & ~n11365 ) | ( n77 & n484 ) | ( ~n11365 & n484 ) ;
  assign n11367 = ( n484 & ~n11366 ) | ( n484 & 1'b0 ) | ( ~n11366 & 1'b0 ) ;
  assign n11370 = n3653 | n11172 ;
  assign n11371 = n3657 &  n11170 ;
  assign n11372 = ( n11370 & ~n11371 ) | ( n11370 & 1'b0 ) | ( ~n11371 & 1'b0 ) ;
  assign n11320 = n11170 | n11172 ;
  assign n11368 = n11170 &  n11172 ;
  assign n11369 = ( n11320 & ~n11368 ) | ( n11320 & 1'b0 ) | ( ~n11368 & 1'b0 ) ;
  assign n11373 = ~n3644 & n11369 ;
  assign n11374 = ( n3644 & n11372 ) | ( n3644 & n11373 ) | ( n11372 & n11373 ) ;
  assign n11375 = n11367 | n11374 ;
  assign n11403 = ( n11367 & ~n11374 ) | ( n11367 & 1'b0 ) | ( ~n11374 & 1'b0 ) ;
  assign n11404 = ( n11375 & ~n11367 ) | ( n11375 & n11403 ) | ( ~n11367 & n11403 ) ;
  assign n11394 = ~n4430 & n11164 ;
  assign n11391 = n523 | n11168 ;
  assign n11392 = n3939 | n11166 ;
  assign n11393 = n11391 &  n11392 ;
  assign n11395 = ( n4430 & n11394 ) | ( n4430 & n11393 ) | ( n11394 & n11393 ) ;
  assign n11396 = ( n11164 & ~n11166 ) | ( n11164 & n11175 ) | ( ~n11166 & n11175 ) ;
  assign n11397 = ( n11166 & ~n11176 ) | ( n11166 & n11396 ) | ( ~n11176 & n11396 ) ;
  assign n11398 = n601 | n11397 ;
  assign n11399 = n11395 &  n11398 ;
  assign n11400 = x29 &  n11399 ;
  assign n11401 = x29 | n11399 ;
  assign n11402 = ~n11400 & n11401 ;
  assign n11405 = n3643 &  n11170 ;
  assign n11428 = ~n4430 & n11166 ;
  assign n11425 = n523 | n11172 ;
  assign n11426 = n3939 | n11168 ;
  assign n11427 = n11425 &  n11426 ;
  assign n11429 = ( n4430 & n11428 ) | ( n4430 & n11427 ) | ( n11428 & n11427 ) ;
  assign n11430 = ( n11166 & ~n11168 ) | ( n11166 & n11174 ) | ( ~n11168 & n11174 ) ;
  assign n11431 = ( n11168 & ~n11175 ) | ( n11168 & n11430 ) | ( ~n11175 & n11430 ) ;
  assign n11432 = n601 | n11431 ;
  assign n11433 = n11429 &  n11432 ;
  assign n11434 = x29 &  n11433 ;
  assign n11435 = x29 | n11433 ;
  assign n11436 = ~n11434 & n11435 ;
  assign n11409 = ~n601 & n11369 ;
  assign n11406 = ~n3939 & n11170 ;
  assign n11407 = n4430 | n11172 ;
  assign n11408 = ~n11406 & n11407 ;
  assign n11410 = ( n601 & n11409 ) | ( n601 & n11408 ) | ( n11409 & n11408 ) ;
  assign n11411 = n521 &  n11170 ;
  assign n11412 = ( x29 & ~n11410 ) | ( x29 & n11411 ) | ( ~n11410 & n11411 ) ;
  assign n11413 = ( x29 & ~n11412 ) | ( x29 & 1'b0 ) | ( ~n11412 & 1'b0 ) ;
  assign n11321 = ( n11168 & ~n11320 ) | ( n11168 & 1'b0 ) | ( ~n11320 & 1'b0 ) ;
  assign n11322 = ~n11168 & n11320 ;
  assign n11323 = n11321 | n11322 ;
  assign n11417 = ~n4430 & n11168 ;
  assign n11414 = ~n523 & n11170 ;
  assign n11415 = n3939 | n11172 ;
  assign n11416 = ~n11414 & n11415 ;
  assign n11418 = ( n4430 & n11417 ) | ( n4430 & n11416 ) | ( n11417 & n11416 ) ;
  assign n11419 = ( n601 & ~n11418 ) | ( n601 & n11323 ) | ( ~n11418 & n11323 ) ;
  assign n11420 = ( n11323 & ~n11419 ) | ( n11323 & 1'b0 ) | ( ~n11419 & 1'b0 ) ;
  assign n11422 = ( x29 & n11418 ) | ( x29 & n11420 ) | ( n11418 & n11420 ) ;
  assign n11421 = ( x29 & ~n11420 ) | ( x29 & n11418 ) | ( ~n11420 & n11418 ) ;
  assign n11423 = ( n11420 & ~n11422 ) | ( n11420 & n11421 ) | ( ~n11422 & n11421 ) ;
  assign n11424 = ( n11413 & ~n11423 ) | ( n11413 & 1'b0 ) | ( ~n11423 & 1'b0 ) ;
  assign n11437 = ( n11405 & ~n11436 ) | ( n11405 & n11424 ) | ( ~n11436 & n11424 ) ;
  assign n11442 = ( n11402 & n11404 ) | ( n11402 & n11437 ) | ( n11404 & n11437 ) ;
  assign n11443 = ( n11402 & ~n11404 ) | ( n11402 & n11437 ) | ( ~n11404 & n11437 ) ;
  assign n11444 = ( n11404 & ~n11442 ) | ( n11404 & n11443 ) | ( ~n11442 & n11443 ) ;
  assign n11448 = n11155 | n4962 ;
  assign n11445 = n4482 | n11161 ;
  assign n11446 = ~n4495 & n11158 ;
  assign n11447 = ( n11445 & ~n11446 ) | ( n11445 & 1'b0 ) | ( ~n11446 & 1'b0 ) ;
  assign n11449 = ( n4962 & ~n11448 ) | ( n4962 & n11447 ) | ( ~n11448 & n11447 ) ;
  assign n11450 = ( n11158 & ~n11155 ) | ( n11158 & n11178 ) | ( ~n11155 & n11178 ) ;
  assign n11451 = ( n11179 & ~n11158 ) | ( n11179 & n11450 ) | ( ~n11158 & n11450 ) ;
  assign n11452 = ( n11449 & ~n4478 ) | ( n11449 & n11451 ) | ( ~n4478 & n11451 ) ;
  assign n11453 = ~n11451 & n11452 ;
  assign n11454 = ( x26 & ~n11449 ) | ( x26 & n11453 ) | ( ~n11449 & n11453 ) ;
  assign n11455 = ( n11449 & ~x26 ) | ( n11449 & n11453 ) | ( ~x26 & n11453 ) ;
  assign n11456 = ( n11454 & ~n11453 ) | ( n11454 & n11455 ) | ( ~n11453 & n11455 ) ;
  assign n11457 = n4962 &  n11158 ;
  assign n11458 = n4495 | n11161 ;
  assign n11459 = n4482 | n11164 ;
  assign n11460 = n11458 &  n11459 ;
  assign n11461 = ( n11457 & ~n11158 ) | ( n11457 & n11460 ) | ( ~n11158 & n11460 ) ;
  assign n11462 = ( n11158 & ~n11177 ) | ( n11158 & n11161 ) | ( ~n11177 & n11161 ) ;
  assign n11463 = ( n11178 & ~n11161 ) | ( n11178 & n11462 ) | ( ~n11161 & n11462 ) ;
  assign n11464 = ~n4478 & n11463 ;
  assign n11465 = ( n11461 & ~n11464 ) | ( n11461 & 1'b0 ) | ( ~n11464 & 1'b0 ) ;
  assign n11466 = x26 &  n11465 ;
  assign n11467 = x26 | n11465 ;
  assign n11468 = ~n11466 & n11467 ;
  assign n11469 = ( n11424 & ~n11405 ) | ( n11424 & n11436 ) | ( ~n11405 & n11436 ) ;
  assign n11470 = ( n11405 & ~n11424 ) | ( n11405 & n11436 ) | ( ~n11424 & n11436 ) ;
  assign n11471 = ( n11469 & ~n11436 ) | ( n11469 & n11470 ) | ( ~n11436 & n11470 ) ;
  assign n11475 = ~n4962 & n11161 ;
  assign n11472 = n4482 | n11166 ;
  assign n11473 = n4495 | n11164 ;
  assign n11474 = n11472 &  n11473 ;
  assign n11476 = ( n4962 & n11475 ) | ( n4962 & n11474 ) | ( n11475 & n11474 ) ;
  assign n11384 = ( n11161 & ~n11164 ) | ( n11161 & n11176 ) | ( ~n11164 & n11176 ) ;
  assign n11385 = ( n11164 & ~n11177 ) | ( n11164 & n11384 ) | ( ~n11177 & n11384 ) ;
  assign n11477 = n4478 | n11385 ;
  assign n11478 = n11476 &  n11477 ;
  assign n11479 = x26 &  n11478 ;
  assign n11480 = x26 | n11478 ;
  assign n11481 = ~n11479 & n11480 ;
  assign n11482 = ~n11413 & n11423 ;
  assign n11483 = n11424 | n11482 ;
  assign n11484 = x29 &  n11411 ;
  assign n11485 = n11410 &  n11484 ;
  assign n11486 = n11410 | n11484 ;
  assign n11487 = ~n11485 & n11486 ;
  assign n11521 = ~n4962 & n11166 ;
  assign n11518 = n4482 | n11172 ;
  assign n11519 = n4495 | n11168 ;
  assign n11520 = n11518 &  n11519 ;
  assign n11522 = ( n4962 & n11521 ) | ( n4962 & n11520 ) | ( n11521 & n11520 ) ;
  assign n11523 = n4478 | n11431 ;
  assign n11524 = n11522 &  n11523 ;
  assign n11525 = x26 &  n11524 ;
  assign n11526 = x26 | n11524 ;
  assign n11527 = ~n11525 & n11526 ;
  assign n11501 = ~n4478 & n11369 ;
  assign n11498 = n4962 | n11172 ;
  assign n11499 = ~n4495 & n11170 ;
  assign n11500 = ( n11498 & ~n11499 ) | ( n11498 & 1'b0 ) | ( ~n11499 & 1'b0 ) ;
  assign n11502 = ( n4478 & n11501 ) | ( n4478 & n11500 ) | ( n11501 & n11500 ) ;
  assign n11503 = n4474 &  n11170 ;
  assign n11505 = ( x26 & ~n11502 ) | ( x26 & n11503 ) | ( ~n11502 & n11503 ) ;
  assign n11506 = ( x26 & ~n11505 ) | ( x26 & 1'b0 ) | ( ~n11505 & 1'b0 ) ;
  assign n11510 = ~n4962 & n11168 ;
  assign n11507 = ~n4482 & n11170 ;
  assign n11508 = n4495 | n11172 ;
  assign n11509 = ~n11507 & n11508 ;
  assign n11511 = ( n4962 & n11510 ) | ( n4962 & n11509 ) | ( n11510 & n11509 ) ;
  assign n11512 = ( n4478 & ~n11511 ) | ( n4478 & n11323 ) | ( ~n11511 & n11323 ) ;
  assign n11513 = ( n11323 & ~n11512 ) | ( n11323 & 1'b0 ) | ( ~n11512 & 1'b0 ) ;
  assign n11515 = ( x26 & n11511 ) | ( x26 & n11513 ) | ( n11511 & n11513 ) ;
  assign n11514 = ( x26 & ~n11513 ) | ( x26 & n11511 ) | ( ~n11513 & n11511 ) ;
  assign n11516 = ( n11513 & ~n11515 ) | ( n11513 & n11514 ) | ( ~n11515 & n11514 ) ;
  assign n11517 = ( n11506 & ~n11516 ) | ( n11506 & 1'b0 ) | ( ~n11516 & 1'b0 ) ;
  assign n11528 = ( n11411 & ~n11527 ) | ( n11411 & n11517 ) | ( ~n11527 & n11517 ) ;
  assign n11491 = ~n4962 & n11164 ;
  assign n11488 = n4482 | n11168 ;
  assign n11489 = n4495 | n11166 ;
  assign n11490 = n11488 &  n11489 ;
  assign n11492 = ( n4962 & n11491 ) | ( n4962 & n11490 ) | ( n11491 & n11490 ) ;
  assign n11493 = ( n11397 & ~n4478 ) | ( n11397 & n11492 ) | ( ~n4478 & n11492 ) ;
  assign n11494 = ~n11397 & n11493 ;
  assign n11495 = ( x26 & ~n11492 ) | ( x26 & n11494 ) | ( ~n11492 & n11494 ) ;
  assign n11496 = ( n11492 & ~x26 ) | ( n11492 & n11494 ) | ( ~x26 & n11494 ) ;
  assign n11497 = ( n11495 & ~n11494 ) | ( n11495 & n11496 ) | ( ~n11494 & n11496 ) ;
  assign n11529 = ( n11487 & ~n11528 ) | ( n11487 & n11497 ) | ( ~n11528 & n11497 ) ;
  assign n11530 = ( n11481 & n11483 ) | ( n11481 & n11529 ) | ( n11483 & n11529 ) ;
  assign n11531 = ( n11468 & n11471 ) | ( n11468 & n11530 ) | ( n11471 & n11530 ) ;
  assign n11532 = ( n11444 & n11456 ) | ( n11444 & n11531 ) | ( n11456 & n11531 ) ;
  assign n11260 = n52 | n237 ;
  assign n11261 = ( n670 & ~n86 ) | ( n670 & n11260 ) | ( ~n86 & n11260 ) ;
  assign n11262 = n86 | n11261 ;
  assign n11263 = n207 | n1626 ;
  assign n11264 = ( n192 & ~n411 ) | ( n192 & n11263 ) | ( ~n411 & n11263 ) ;
  assign n11265 = n411 | n11264 ;
  assign n11266 = n1196 | n2347 ;
  assign n11267 = ( n3442 & ~n11265 ) | ( n3442 & n11266 ) | ( ~n11265 & n11266 ) ;
  assign n11268 = ( n1167 & n11267 ) | ( n1167 & n11265 ) | ( n11267 & n11265 ) ;
  assign n11269 = ( n1167 & ~n11268 ) | ( n1167 & 1'b0 ) | ( ~n11268 & 1'b0 ) ;
  assign n11270 = ( n2862 & n11262 ) | ( n2862 & n11269 ) | ( n11262 & n11269 ) ;
  assign n11271 = ( n794 & ~n11262 ) | ( n794 & n11270 ) | ( ~n11262 & n11270 ) ;
  assign n11272 = ~n794 & n11271 ;
  assign n11273 = ( n605 & ~n1244 ) | ( n605 & n11272 ) | ( ~n1244 & n11272 ) ;
  assign n11274 = ~n605 & n11273 ;
  assign n11275 = ( n346 & ~n2309 ) | ( n346 & n11274 ) | ( ~n2309 & n11274 ) ;
  assign n11276 = ~n346 & n11275 ;
  assign n11277 = ( n69 & ~n127 ) | ( n69 & n11276 ) | ( ~n127 & n11276 ) ;
  assign n11278 = ~n69 & n11277 ;
  assign n11279 = ( n208 & ~n11278 ) | ( n208 & n354 ) | ( ~n11278 & n354 ) ;
  assign n11280 = ( n354 & ~n11279 ) | ( n354 & 1'b0 ) | ( ~n11279 & 1'b0 ) ;
  assign n11281 = ~n95 & n11280 ;
  assign n11302 = n1460 | n3961 ;
  assign n11303 = ( n795 & ~n1704 ) | ( n795 & n11302 ) | ( ~n1704 & n11302 ) ;
  assign n11304 = n1704 | n11303 ;
  assign n11282 = n679 | n796 ;
  assign n11283 = n403 | n11282 ;
  assign n11284 = ( n2332 & ~n2062 ) | ( n2332 & n11283 ) | ( ~n2062 & n11283 ) ;
  assign n11285 = n2062 | n11284 ;
  assign n11286 = ( n1877 & ~n1823 ) | ( n1877 & n11285 ) | ( ~n1823 & n11285 ) ;
  assign n11287 = n1823 | n11286 ;
  assign n11288 = ( n667 & ~n1762 ) | ( n667 & n11287 ) | ( ~n1762 & n11287 ) ;
  assign n11289 = n1762 | n11288 ;
  assign n11290 = ( n775 & ~n61 ) | ( n775 & n11289 ) | ( ~n61 & n11289 ) ;
  assign n11291 = n61 | n11290 ;
  assign n11292 = ( n338 & ~n196 ) | ( n338 & n11291 ) | ( ~n196 & n11291 ) ;
  assign n11293 = n196 | n11292 ;
  assign n11294 = n432 | n11293 ;
  assign n11295 = n260 | n1098 ;
  assign n11296 = ( n789 & ~n234 ) | ( n789 & n11295 ) | ( ~n234 & n11295 ) ;
  assign n11297 = n234 | n11296 ;
  assign n11298 = ( n217 & ~n245 ) | ( n217 & n11297 ) | ( ~n245 & n11297 ) ;
  assign n11299 = n245 | n11298 ;
  assign n11300 = ( n80 & ~n205 ) | ( n80 & n11299 ) | ( ~n205 & n11299 ) ;
  assign n11301 = n205 | n11300 ;
  assign n11305 = ( n11304 & ~n11294 ) | ( n11304 & n11301 ) | ( ~n11294 & n11301 ) ;
  assign n11306 = ( n11281 & n11305 ) | ( n11281 & n11294 ) | ( n11305 & n11294 ) ;
  assign n11307 = ( n11281 & ~n11306 ) | ( n11281 & 1'b0 ) | ( ~n11306 & 1'b0 ) ;
  assign n11308 = ( n2187 & ~n3741 ) | ( n2187 & n11307 ) | ( ~n3741 & n11307 ) ;
  assign n11309 = ~n2187 & n11308 ;
  assign n11310 = ( n602 & ~n409 ) | ( n602 & n11309 ) | ( ~n409 & n11309 ) ;
  assign n11311 = ~n602 & n11310 ;
  assign n11312 = ( n284 & ~n415 ) | ( n284 & n11311 ) | ( ~n415 & n11311 ) ;
  assign n11313 = ~n284 & n11312 ;
  assign n11314 = ( n734 & ~n188 ) | ( n734 & n11313 ) | ( ~n188 & n11313 ) ;
  assign n11315 = ~n734 & n11314 ;
  assign n11316 = ( n382 & ~n531 ) | ( n382 & n11315 ) | ( ~n531 & n11315 ) ;
  assign n11317 = ~n382 & n11316 ;
  assign n11318 = ( n225 & ~n77 ) | ( n225 & n11317 ) | ( ~n77 & n11317 ) ;
  assign n11319 = ~n225 & n11318 ;
  assign n11324 = ~n3644 & n11323 ;
  assign n11325 = n3652 &  n11170 ;
  assign n11326 = ( n3657 & ~n11172 ) | ( n3657 & 1'b0 ) | ( ~n11172 & 1'b0 ) ;
  assign n11327 = n11325 | n11326 ;
  assign n11328 = ~n3653 & n11168 ;
  assign n11329 = ( n3653 & ~n11327 ) | ( n3653 & n11328 ) | ( ~n11327 & n11328 ) ;
  assign n11330 = ~n11324 & n11329 ;
  assign n11376 = ( n11319 & n11330 ) | ( n11319 & n11375 ) | ( n11330 & n11375 ) ;
  assign n11377 = ( n11330 & ~n11319 ) | ( n11330 & n11375 ) | ( ~n11319 & n11375 ) ;
  assign n11378 = ( n11319 & ~n11376 ) | ( n11319 & n11377 ) | ( ~n11376 & n11377 ) ;
  assign n11382 = ~n4430 & n11161 ;
  assign n11379 = n523 | n11166 ;
  assign n11380 = n3939 | n11164 ;
  assign n11381 = n11379 &  n11380 ;
  assign n11383 = ( n4430 & n11382 ) | ( n4430 & n11381 ) | ( n11382 & n11381 ) ;
  assign n11386 = n601 | n11385 ;
  assign n11387 = n11383 &  n11386 ;
  assign n11388 = x29 &  n11387 ;
  assign n11389 = x29 | n11387 ;
  assign n11390 = ~n11388 & n11389 ;
  assign n11438 = ( n11404 & ~n11402 ) | ( n11404 & n11437 ) | ( ~n11402 & n11437 ) ;
  assign n11440 = ( n11378 & n11390 ) | ( n11378 & n11438 ) | ( n11390 & n11438 ) ;
  assign n11439 = ( n11390 & ~n11378 ) | ( n11390 & n11438 ) | ( ~n11378 & n11438 ) ;
  assign n11441 = ( n11378 & ~n11440 ) | ( n11378 & n11439 ) | ( ~n11440 & n11439 ) ;
  assign n11533 = ( n11259 & ~n11532 ) | ( n11259 & n11441 ) | ( ~n11532 & n11441 ) ;
  assign n11534 = ( n11259 & ~n11441 ) | ( n11259 & n11532 ) | ( ~n11441 & n11532 ) ;
  assign n11535 = ( n11533 & ~n11259 ) | ( n11533 & n11534 ) | ( ~n11259 & n11534 ) ;
  assign n11539 = ~n5135 & n11143 ;
  assign n11536 = n5010 | n11149 ;
  assign n11537 = n5067 | n11146 ;
  assign n11538 = n11536 &  n11537 ;
  assign n11540 = ( n5135 & n11539 ) | ( n5135 & n11538 ) | ( n11539 & n11538 ) ;
  assign n11541 = ( n11143 & ~n11146 ) | ( n11143 & n11182 ) | ( ~n11146 & n11182 ) ;
  assign n11542 = ( n11146 & ~n11183 ) | ( n11146 & n11541 ) | ( ~n11183 & n11541 ) ;
  assign n11543 = n5012 | n11542 ;
  assign n11544 = n11540 &  n11543 ;
  assign n11545 = x23 &  n11544 ;
  assign n11546 = x23 | n11544 ;
  assign n11547 = ~n11545 & n11546 ;
  assign n11551 = ~n5135 & n11146 ;
  assign n11548 = ~n5010 & n11152 ;
  assign n11549 = n5067 | n11149 ;
  assign n11550 = ~n11548 & n11549 ;
  assign n11552 = ( n5135 & n11551 ) | ( n5135 & n11550 ) | ( n11551 & n11550 ) ;
  assign n11553 = ( n11149 & ~n11146 ) | ( n11149 & n11181 ) | ( ~n11146 & n11181 ) ;
  assign n11554 = ( n11182 & ~n11149 ) | ( n11182 & n11553 ) | ( ~n11149 & n11553 ) ;
  assign n11555 = ~n5012 & n11554 ;
  assign n11556 = ( n11552 & ~n11555 ) | ( n11552 & 1'b0 ) | ( ~n11555 & 1'b0 ) ;
  assign n11557 = x23 &  n11556 ;
  assign n11558 = x23 | n11556 ;
  assign n11559 = ~n11557 & n11558 ;
  assign n11560 = ( n11456 & ~n11444 ) | ( n11456 & n11531 ) | ( ~n11444 & n11531 ) ;
  assign n11561 = ( n11444 & ~n11531 ) | ( n11444 & n11456 ) | ( ~n11531 & n11456 ) ;
  assign n11562 = ( n11560 & ~n11456 ) | ( n11560 & n11561 ) | ( ~n11456 & n11561 ) ;
  assign n11563 = ( n11468 & ~n11530 ) | ( n11468 & n11471 ) | ( ~n11530 & n11471 ) ;
  assign n11564 = ( n11471 & ~n11468 ) | ( n11471 & n11530 ) | ( ~n11468 & n11530 ) ;
  assign n11565 = ( n11563 & ~n11471 ) | ( n11563 & n11564 ) | ( ~n11471 & n11564 ) ;
  assign n11571 = ( n11149 & ~n11180 ) | ( n11149 & n11152 ) | ( ~n11180 & n11152 ) ;
  assign n11572 = ( n11181 & ~n11152 ) | ( n11181 & n11571 ) | ( ~n11152 & n11571 ) ;
  assign n11566 = ~n5010 & n11155 ;
  assign n11567 = ~n5067 & n11152 ;
  assign n11568 = n11566 | n11567 ;
  assign n11569 = ~n5135 & n11149 ;
  assign n11570 = ( n5135 & ~n11568 ) | ( n5135 & n11569 ) | ( ~n11568 & n11569 ) ;
  assign n11573 = ( n11570 & ~n5012 ) | ( n11570 & n11572 ) | ( ~n5012 & n11572 ) ;
  assign n11574 = ~n11572 & n11573 ;
  assign n11576 = ( x23 & n11570 ) | ( x23 & n11574 ) | ( n11570 & n11574 ) ;
  assign n11575 = ( x23 & ~n11574 ) | ( x23 & n11570 ) | ( ~n11574 & n11570 ) ;
  assign n11577 = ( n11574 & ~n11576 ) | ( n11574 & n11575 ) | ( ~n11576 & n11575 ) ;
  assign n11578 = ( n11481 & ~n11483 ) | ( n11481 & n11529 ) | ( ~n11483 & n11529 ) ;
  assign n11579 = ( n11483 & ~n11481 ) | ( n11483 & n11529 ) | ( ~n11481 & n11529 ) ;
  assign n11580 = ( n11578 & ~n11529 ) | ( n11578 & n11579 ) | ( ~n11529 & n11579 ) ;
  assign n11584 = n11152 | n5135 ;
  assign n11581 = ~n5010 & n11158 ;
  assign n11582 = ~n5067 & n11155 ;
  assign n11583 = n11581 | n11582 ;
  assign n11585 = ( n11584 & ~n5135 ) | ( n11584 & n11583 ) | ( ~n5135 & n11583 ) ;
  assign n11586 = ( n5012 & n11254 ) | ( n5012 & n11585 ) | ( n11254 & n11585 ) ;
  assign n11587 = ( n11254 & ~n11586 ) | ( n11254 & 1'b0 ) | ( ~n11586 & 1'b0 ) ;
  assign n11588 = ( n11585 & ~x23 ) | ( n11585 & n11587 ) | ( ~x23 & n11587 ) ;
  assign n11589 = ( x23 & ~n11585 ) | ( x23 & n11587 ) | ( ~n11585 & n11587 ) ;
  assign n11590 = ( n11588 & ~n11587 ) | ( n11588 & n11589 ) | ( ~n11587 & n11589 ) ;
  assign n11594 = n11155 | n5135 ;
  assign n11591 = n5010 | n11161 ;
  assign n11592 = ~n5067 & n11158 ;
  assign n11593 = ( n11591 & ~n11592 ) | ( n11591 & 1'b0 ) | ( ~n11592 & 1'b0 ) ;
  assign n11595 = ( n5135 & ~n11594 ) | ( n5135 & n11593 ) | ( ~n11594 & n11593 ) ;
  assign n11596 = n5012 | n11451 ;
  assign n11597 = n11595 &  n11596 ;
  assign n11598 = x23 &  n11597 ;
  assign n11599 = x23 | n11597 ;
  assign n11600 = ~n11598 & n11599 ;
  assign n11601 = ( n11497 & ~n11487 ) | ( n11497 & n11528 ) | ( ~n11487 & n11528 ) ;
  assign n11602 = ( n11529 & ~n11497 ) | ( n11529 & n11601 ) | ( ~n11497 & n11601 ) ;
  assign n11604 = ( n11411 & n11517 ) | ( n11411 & n11527 ) | ( n11517 & n11527 ) ;
  assign n11603 = ( n11411 & ~n11517 ) | ( n11411 & n11527 ) | ( ~n11517 & n11527 ) ;
  assign n11605 = ( n11517 & ~n11604 ) | ( n11517 & n11603 ) | ( ~n11604 & n11603 ) ;
  assign n11606 = n5135 &  n11158 ;
  assign n11607 = n5010 | n11164 ;
  assign n11608 = n5067 | n11161 ;
  assign n11609 = n11607 &  n11608 ;
  assign n11610 = ( n11606 & ~n11158 ) | ( n11606 & n11609 ) | ( ~n11158 & n11609 ) ;
  assign n11611 = ( n5012 & ~n11610 ) | ( n5012 & n11463 ) | ( ~n11610 & n11463 ) ;
  assign n11612 = ( n11463 & ~n11611 ) | ( n11463 & 1'b0 ) | ( ~n11611 & 1'b0 ) ;
  assign n11614 = ( x23 & n11610 ) | ( x23 & n11612 ) | ( n11610 & n11612 ) ;
  assign n11613 = ( x23 & ~n11612 ) | ( x23 & n11610 ) | ( ~n11612 & n11610 ) ;
  assign n11615 = ( n11612 & ~n11614 ) | ( n11612 & n11613 ) | ( ~n11614 & n11613 ) ;
  assign n11619 = ~n5135 & n11161 ;
  assign n11616 = n5010 | n11166 ;
  assign n11617 = n5067 | n11164 ;
  assign n11618 = n11616 &  n11617 ;
  assign n11620 = ( n5135 & n11619 ) | ( n5135 & n11618 ) | ( n11619 & n11618 ) ;
  assign n11621 = n5012 | n11385 ;
  assign n11622 = n11620 &  n11621 ;
  assign n11623 = x23 &  n11622 ;
  assign n11624 = x23 | n11622 ;
  assign n11625 = ~n11623 & n11624 ;
  assign n11626 = ~n11506 & n11516 ;
  assign n11627 = n11517 | n11626 ;
  assign n11504 = ( x26 & ~n11503 ) | ( x26 & 1'b0 ) | ( ~n11503 & 1'b0 ) ;
  assign n11628 = ( n11502 & ~x26 ) | ( n11502 & n11504 ) | ( ~x26 & n11504 ) ;
  assign n11629 = ( x26 & ~n11504 ) | ( x26 & n11502 ) | ( ~n11504 & n11502 ) ;
  assign n11630 = ( n11628 & ~n11502 ) | ( n11628 & n11629 ) | ( ~n11502 & n11629 ) ;
  assign n11660 = ~n5135 & n11166 ;
  assign n11657 = n5010 | n11172 ;
  assign n11658 = n5067 | n11168 ;
  assign n11659 = n11657 &  n11658 ;
  assign n11661 = ( n5135 & n11660 ) | ( n5135 & n11659 ) | ( n11660 & n11659 ) ;
  assign n11662 = n5012 | n11431 ;
  assign n11663 = n11661 &  n11662 ;
  assign n11664 = x23 &  n11663 ;
  assign n11665 = x23 | n11663 ;
  assign n11666 = ~n11664 & n11665 ;
  assign n11641 = n5005 &  n11170 ;
  assign n11645 = ~n5012 & n11369 ;
  assign n11642 = ~n5067 & n11170 ;
  assign n11643 = n5135 | n11172 ;
  assign n11644 = ~n11642 & n11643 ;
  assign n11646 = ( n5012 & n11645 ) | ( n5012 & n11644 ) | ( n11645 & n11644 ) ;
  assign n11652 = n11323 | n5012 ;
  assign n11650 = ~n5135 & n11168 ;
  assign n11647 = ~n5010 & n11170 ;
  assign n11648 = n5067 | n11172 ;
  assign n11649 = ~n11647 & n11648 ;
  assign n11651 = ( n5135 & n11650 ) | ( n5135 & n11649 ) | ( n11650 & n11649 ) ;
  assign n11653 = ( n5012 & ~n11652 ) | ( n5012 & n11651 ) | ( ~n11652 & n11651 ) ;
  assign n11654 = ( n11641 & n11646 ) | ( n11641 & n11653 ) | ( n11646 & n11653 ) ;
  assign n11655 = ( x23 & ~n11654 ) | ( x23 & n11641 ) | ( ~n11654 & n11641 ) ;
  assign n11656 = ( x23 & ~n11655 ) | ( x23 & 1'b0 ) | ( ~n11655 & 1'b0 ) ;
  assign n11667 = ( n11503 & ~n11666 ) | ( n11503 & n11656 ) | ( ~n11666 & n11656 ) ;
  assign n11634 = ~n5135 & n11164 ;
  assign n11631 = n5010 | n11168 ;
  assign n11632 = n5067 | n11166 ;
  assign n11633 = n11631 &  n11632 ;
  assign n11635 = ( n5135 & n11634 ) | ( n5135 & n11633 ) | ( n11634 & n11633 ) ;
  assign n11636 = ( n11397 & ~n5012 ) | ( n11397 & n11635 ) | ( ~n5012 & n11635 ) ;
  assign n11637 = ~n11397 & n11636 ;
  assign n11638 = ( x23 & ~n11635 ) | ( x23 & n11637 ) | ( ~n11635 & n11637 ) ;
  assign n11639 = ( n11635 & ~x23 ) | ( n11635 & n11637 ) | ( ~x23 & n11637 ) ;
  assign n11640 = ( n11638 & ~n11637 ) | ( n11638 & n11639 ) | ( ~n11637 & n11639 ) ;
  assign n11668 = ( n11630 & ~n11667 ) | ( n11630 & n11640 ) | ( ~n11667 & n11640 ) ;
  assign n11669 = ( n11625 & n11627 ) | ( n11625 & n11668 ) | ( n11627 & n11668 ) ;
  assign n11670 = ( n11605 & n11615 ) | ( n11605 & n11669 ) | ( n11615 & n11669 ) ;
  assign n11671 = ( n11600 & ~n11602 ) | ( n11600 & n11670 ) | ( ~n11602 & n11670 ) ;
  assign n11672 = ( n11580 & ~n11590 ) | ( n11580 & n11671 ) | ( ~n11590 & n11671 ) ;
  assign n11673 = ( n11565 & n11577 ) | ( n11565 & n11672 ) | ( n11577 & n11672 ) ;
  assign n11674 = ( n11559 & n11562 ) | ( n11559 & n11673 ) | ( n11562 & n11673 ) ;
  assign n11675 = ( n11535 & ~n11547 ) | ( n11535 & n11674 ) | ( ~n11547 & n11674 ) ;
  assign n11676 = ( n11535 & ~n11674 ) | ( n11535 & n11547 ) | ( ~n11674 & n11547 ) ;
  assign n11677 = ( n11675 & ~n11535 ) | ( n11675 & n11676 ) | ( ~n11535 & n11676 ) ;
  assign n11678 = ( n11562 & ~n11559 ) | ( n11562 & n11673 ) | ( ~n11559 & n11673 ) ;
  assign n11679 = ( n11559 & ~n11673 ) | ( n11559 & n11562 ) | ( ~n11673 & n11562 ) ;
  assign n11680 = ( n11678 & ~n11562 ) | ( n11678 & n11679 ) | ( ~n11562 & n11679 ) ;
  assign n11686 = ( n11137 & ~n11140 ) | ( n11137 & n11184 ) | ( ~n11140 & n11184 ) ;
  assign n11687 = ( n11140 & ~n11185 ) | ( n11140 & n11686 ) | ( ~n11185 & n11686 ) ;
  assign n11684 = ~n5837 & n11137 ;
  assign n11681 = ( n5339 & ~n11143 ) | ( n5339 & 1'b0 ) | ( ~n11143 & 1'b0 ) ;
  assign n11682 = n5761 | n11140 ;
  assign n11683 = ~n11681 & n11682 ;
  assign n11685 = ( n5837 & n11684 ) | ( n5837 & n11683 ) | ( n11684 & n11683 ) ;
  assign n11688 = ( n11685 & ~n5341 ) | ( n11685 & n11687 ) | ( ~n5341 & n11687 ) ;
  assign n11689 = ~n11687 & n11688 ;
  assign n11691 = ( x20 & n11685 ) | ( x20 & n11689 ) | ( n11685 & n11689 ) ;
  assign n11690 = ( x20 & ~n11689 ) | ( x20 & n11685 ) | ( ~n11689 & n11685 ) ;
  assign n11692 = ( n11689 & ~n11691 ) | ( n11689 & n11690 ) | ( ~n11691 & n11690 ) ;
  assign n11696 = ~n5837 & n11140 ;
  assign n11693 = ( n5339 & ~n11146 ) | ( n5339 & 1'b0 ) | ( ~n11146 & 1'b0 ) ;
  assign n11694 = n5761 | n11143 ;
  assign n11695 = ~n11693 & n11694 ;
  assign n11697 = ( n5837 & n11696 ) | ( n5837 & n11695 ) | ( n11696 & n11695 ) ;
  assign n11698 = ( n11140 & ~n11143 ) | ( n11140 & n11183 ) | ( ~n11143 & n11183 ) ;
  assign n11699 = ( n11143 & ~n11184 ) | ( n11143 & n11698 ) | ( ~n11184 & n11698 ) ;
  assign n11700 = n5341 | n11699 ;
  assign n11701 = n11697 &  n11700 ;
  assign n11702 = x20 &  n11701 ;
  assign n11703 = x20 | n11701 ;
  assign n11704 = ~n11702 & n11703 ;
  assign n11705 = ( n11565 & ~n11577 ) | ( n11565 & n11672 ) | ( ~n11577 & n11672 ) ;
  assign n11706 = ( n11577 & ~n11673 ) | ( n11577 & n11705 ) | ( ~n11673 & n11705 ) ;
  assign n11710 = ~n5837 & n11143 ;
  assign n11707 = ( n5339 & ~n11149 ) | ( n5339 & 1'b0 ) | ( ~n11149 & 1'b0 ) ;
  assign n11708 = n5761 | n11146 ;
  assign n11709 = ~n11707 & n11708 ;
  assign n11711 = ( n5837 & n11710 ) | ( n5837 & n11709 ) | ( n11710 & n11709 ) ;
  assign n11712 = n5341 | n11542 ;
  assign n11713 = n11711 &  n11712 ;
  assign n11714 = x20 &  n11713 ;
  assign n11715 = x20 | n11713 ;
  assign n11716 = ~n11714 & n11715 ;
  assign n11717 = ( n11580 & n11590 ) | ( n11580 & n11671 ) | ( n11590 & n11671 ) ;
  assign n11718 = ( n11590 & ~n11717 ) | ( n11590 & n11672 ) | ( ~n11717 & n11672 ) ;
  assign n11725 = ~n5837 & n11146 ;
  assign n11722 = n5339 &  n11152 ;
  assign n11723 = n5761 | n11149 ;
  assign n11724 = ~n11722 & n11723 ;
  assign n11726 = ( n5837 & n11725 ) | ( n5837 & n11724 ) | ( n11725 & n11724 ) ;
  assign n11727 = ( n5341 & ~n11726 ) | ( n5341 & n11554 ) | ( ~n11726 & n11554 ) ;
  assign n11728 = ( n11554 & ~n11727 ) | ( n11554 & 1'b0 ) | ( ~n11727 & 1'b0 ) ;
  assign n11729 = ( x20 & ~n11726 ) | ( x20 & n11728 ) | ( ~n11726 & n11728 ) ;
  assign n11730 = ( n11726 & ~x20 ) | ( n11726 & n11728 ) | ( ~x20 & n11728 ) ;
  assign n11731 = ( n11729 & ~n11728 ) | ( n11729 & n11730 ) | ( ~n11728 & n11730 ) ;
  assign n11719 = ( n11602 & ~n11600 ) | ( n11602 & n11670 ) | ( ~n11600 & n11670 ) ;
  assign n11720 = ( n11600 & ~n11670 ) | ( n11600 & n11602 ) | ( ~n11670 & n11602 ) ;
  assign n11721 = ( n11719 & ~n11602 ) | ( n11719 & n11720 ) | ( ~n11602 & n11720 ) ;
  assign n11732 = ( n11615 & ~n11605 ) | ( n11615 & n11669 ) | ( ~n11605 & n11669 ) ;
  assign n11733 = ( n11605 & ~n11669 ) | ( n11605 & n11615 ) | ( ~n11669 & n11615 ) ;
  assign n11734 = ( n11732 & ~n11615 ) | ( n11732 & n11733 ) | ( ~n11615 & n11733 ) ;
  assign n11735 = n5339 &  n11155 ;
  assign n11736 = ~n5761 & n11152 ;
  assign n11737 = n11735 | n11736 ;
  assign n11738 = ~n5837 & n11149 ;
  assign n11739 = ( n5837 & ~n11737 ) | ( n5837 & n11738 ) | ( ~n11737 & n11738 ) ;
  assign n11740 = ( n11572 & ~n5341 ) | ( n11572 & n11739 ) | ( ~n5341 & n11739 ) ;
  assign n11741 = ~n11572 & n11740 ;
  assign n11743 = ( x20 & n11739 ) | ( x20 & n11741 ) | ( n11739 & n11741 ) ;
  assign n11742 = ( x20 & ~n11741 ) | ( x20 & n11739 ) | ( ~n11741 & n11739 ) ;
  assign n11744 = ( n11741 & ~n11743 ) | ( n11741 & n11742 ) | ( ~n11743 & n11742 ) ;
  assign n11745 = ( n11625 & ~n11627 ) | ( n11625 & n11668 ) | ( ~n11627 & n11668 ) ;
  assign n11746 = ( n11627 & ~n11625 ) | ( n11627 & n11668 ) | ( ~n11625 & n11668 ) ;
  assign n11747 = ( n11745 & ~n11668 ) | ( n11745 & n11746 ) | ( ~n11668 & n11746 ) ;
  assign n11751 = n11152 | n5837 ;
  assign n11748 = n5339 &  n11158 ;
  assign n11749 = ~n5761 & n11155 ;
  assign n11750 = n11748 | n11749 ;
  assign n11752 = ( n11751 & ~n5837 ) | ( n11751 & n11750 ) | ( ~n5837 & n11750 ) ;
  assign n11753 = ( n5341 & n11254 ) | ( n5341 & n11752 ) | ( n11254 & n11752 ) ;
  assign n11754 = ( n11254 & ~n11753 ) | ( n11254 & 1'b0 ) | ( ~n11753 & 1'b0 ) ;
  assign n11755 = ( n11752 & ~x20 ) | ( n11752 & n11754 ) | ( ~x20 & n11754 ) ;
  assign n11756 = ( x20 & ~n11752 ) | ( x20 & n11754 ) | ( ~n11752 & n11754 ) ;
  assign n11757 = ( n11755 & ~n11754 ) | ( n11755 & n11756 ) | ( ~n11754 & n11756 ) ;
  assign n11761 = n11155 | n5837 ;
  assign n11758 = ( n5339 & ~n11161 ) | ( n5339 & 1'b0 ) | ( ~n11161 & 1'b0 ) ;
  assign n11759 = ~n5761 & n11158 ;
  assign n11760 = n11758 | n11759 ;
  assign n11762 = ( n11761 & ~n5837 ) | ( n11761 & n11760 ) | ( ~n5837 & n11760 ) ;
  assign n11763 = n5341 | n11451 ;
  assign n11764 = ~n11762 & n11763 ;
  assign n11765 = x20 &  n11764 ;
  assign n11766 = x20 | n11764 ;
  assign n11767 = ~n11765 & n11766 ;
  assign n11768 = ( n11630 & n11640 ) | ( n11630 & n11667 ) | ( n11640 & n11667 ) ;
  assign n11769 = ( n11630 & ~n11640 ) | ( n11630 & n11667 ) | ( ~n11640 & n11667 ) ;
  assign n11770 = ( n11640 & ~n11768 ) | ( n11640 & n11769 ) | ( ~n11768 & n11769 ) ;
  assign n11772 = ( n11503 & n11656 ) | ( n11503 & n11666 ) | ( n11656 & n11666 ) ;
  assign n11771 = ( n11503 & ~n11656 ) | ( n11503 & n11666 ) | ( ~n11656 & n11666 ) ;
  assign n11773 = ( n11656 & ~n11772 ) | ( n11656 & n11771 ) | ( ~n11772 & n11771 ) ;
  assign n11777 = n11158 | n5837 ;
  assign n11774 = ( n5339 & ~n11164 ) | ( n5339 & 1'b0 ) | ( ~n11164 & 1'b0 ) ;
  assign n11775 = n5761 | n11161 ;
  assign n11776 = ~n11774 & n11775 ;
  assign n11778 = ( n5837 & ~n11777 ) | ( n5837 & n11776 ) | ( ~n11777 & n11776 ) ;
  assign n11779 = ( n5341 & ~n11778 ) | ( n5341 & n11463 ) | ( ~n11778 & n11463 ) ;
  assign n11780 = ( n11463 & ~n11779 ) | ( n11463 & 1'b0 ) | ( ~n11779 & 1'b0 ) ;
  assign n11782 = ( x20 & n11778 ) | ( x20 & n11780 ) | ( n11778 & n11780 ) ;
  assign n11781 = ( x20 & ~n11780 ) | ( x20 & n11778 ) | ( ~n11780 & n11778 ) ;
  assign n11783 = ( n11780 & ~n11782 ) | ( n11780 & n11781 ) | ( ~n11782 & n11781 ) ;
  assign n11784 = ( n5339 & ~n11166 ) | ( n5339 & 1'b0 ) | ( ~n11166 & 1'b0 ) ;
  assign n11785 = n5761 | n11164 ;
  assign n11786 = ~n11784 & n11785 ;
  assign n11787 = ~n5837 & n11161 ;
  assign n11788 = ( n5837 & n11786 ) | ( n5837 & n11787 ) | ( n11786 & n11787 ) ;
  assign n11789 = n5341 | n11385 ;
  assign n11790 = n11788 &  n11789 ;
  assign n11791 = x20 &  n11790 ;
  assign n11792 = x20 | n11790 ;
  assign n11793 = ~n11791 & n11792 ;
  assign n11794 = ( x23 & n11641 ) | ( x23 & n11646 ) | ( n11641 & n11646 ) ;
  assign n11795 = ~n11641 & n11794 ;
  assign n11796 = ( n11653 & ~x23 ) | ( n11653 & n11795 ) | ( ~x23 & n11795 ) ;
  assign n11797 = ( x23 & ~n11653 ) | ( x23 & n11795 ) | ( ~n11653 & n11795 ) ;
  assign n11798 = ( n11796 & ~n11795 ) | ( n11796 & n11797 ) | ( ~n11795 & n11797 ) ;
  assign n11799 = x23 &  n11641 ;
  assign n11800 = n11646 &  n11799 ;
  assign n11801 = n11646 | n11799 ;
  assign n11802 = ~n11800 & n11801 ;
  assign n11832 = ~n5837 & n11166 ;
  assign n11829 = ( n5339 & ~n11172 ) | ( n5339 & 1'b0 ) | ( ~n11172 & 1'b0 ) ;
  assign n11830 = n5761 | n11168 ;
  assign n11831 = ~n11829 & n11830 ;
  assign n11833 = ( n5837 & n11832 ) | ( n5837 & n11831 ) | ( n11832 & n11831 ) ;
  assign n11834 = n5341 | n11431 ;
  assign n11835 = n11833 &  n11834 ;
  assign n11836 = x20 &  n11835 ;
  assign n11837 = x20 | n11835 ;
  assign n11838 = ~n11836 & n11837 ;
  assign n11813 = n5337 &  n11170 ;
  assign n11817 = ~n5341 & n11369 ;
  assign n11814 = ~n5761 & n11170 ;
  assign n11815 = n5837 | n11172 ;
  assign n11816 = ~n11814 & n11815 ;
  assign n11818 = ( n5341 & n11817 ) | ( n5341 & n11816 ) | ( n11817 & n11816 ) ;
  assign n11824 = n11323 | n5341 ;
  assign n11822 = ~n5837 & n11168 ;
  assign n11819 = n5339 &  n11170 ;
  assign n11820 = n5761 | n11172 ;
  assign n11821 = ~n11819 & n11820 ;
  assign n11823 = ( n5837 & n11822 ) | ( n5837 & n11821 ) | ( n11822 & n11821 ) ;
  assign n11825 = ( n5341 & ~n11824 ) | ( n5341 & n11823 ) | ( ~n11824 & n11823 ) ;
  assign n11826 = ( n11813 & n11818 ) | ( n11813 & n11825 ) | ( n11818 & n11825 ) ;
  assign n11827 = ( x20 & ~n11826 ) | ( x20 & n11813 ) | ( ~n11826 & n11813 ) ;
  assign n11828 = ( x20 & ~n11827 ) | ( x20 & 1'b0 ) | ( ~n11827 & 1'b0 ) ;
  assign n11839 = ( n11641 & ~n11838 ) | ( n11641 & n11828 ) | ( ~n11838 & n11828 ) ;
  assign n11806 = ~n5837 & n11164 ;
  assign n11803 = ( n5339 & ~n11168 ) | ( n5339 & 1'b0 ) | ( ~n11168 & 1'b0 ) ;
  assign n11804 = n5761 | n11166 ;
  assign n11805 = ~n11803 & n11804 ;
  assign n11807 = ( n5837 & n11806 ) | ( n5837 & n11805 ) | ( n11806 & n11805 ) ;
  assign n11808 = ( n11397 & ~n5341 ) | ( n11397 & n11807 ) | ( ~n5341 & n11807 ) ;
  assign n11809 = ~n11397 & n11808 ;
  assign n11810 = ( x20 & ~n11807 ) | ( x20 & n11809 ) | ( ~n11807 & n11809 ) ;
  assign n11811 = ( n11807 & ~x20 ) | ( n11807 & n11809 ) | ( ~x20 & n11809 ) ;
  assign n11812 = ( n11810 & ~n11809 ) | ( n11810 & n11811 ) | ( ~n11809 & n11811 ) ;
  assign n11840 = ( n11802 & ~n11839 ) | ( n11802 & n11812 ) | ( ~n11839 & n11812 ) ;
  assign n11841 = ( n11793 & n11798 ) | ( n11793 & n11840 ) | ( n11798 & n11840 ) ;
  assign n11842 = ( n11773 & n11783 ) | ( n11773 & n11841 ) | ( n11783 & n11841 ) ;
  assign n11843 = ( n11767 & ~n11770 ) | ( n11767 & n11842 ) | ( ~n11770 & n11842 ) ;
  assign n11844 = ( n11747 & ~n11757 ) | ( n11747 & n11843 ) | ( ~n11757 & n11843 ) ;
  assign n11845 = ( n11734 & n11744 ) | ( n11734 & n11844 ) | ( n11744 & n11844 ) ;
  assign n11846 = ( n11731 & ~n11721 ) | ( n11731 & n11845 ) | ( ~n11721 & n11845 ) ;
  assign n11847 = ( n11716 & ~n11718 ) | ( n11716 & n11846 ) | ( ~n11718 & n11846 ) ;
  assign n11848 = ( n11704 & n11706 ) | ( n11704 & n11847 ) | ( n11706 & n11847 ) ;
  assign n11849 = ( n11680 & n11692 ) | ( n11680 & n11848 ) | ( n11692 & n11848 ) ;
  assign n11850 = ( n11247 & n11677 ) | ( n11247 & n11849 ) | ( n11677 & n11849 ) ;
  assign n11851 = ( n11677 & ~n11247 ) | ( n11677 & n11849 ) | ( ~n11247 & n11849 ) ;
  assign n11852 = ( n11247 & ~n11850 ) | ( n11247 & n11851 ) | ( ~n11850 & n11851 ) ;
  assign n11853 = n6395 &  n11125 ;
  assign n11854 = n5970 | n11131 ;
  assign n11855 = n6170 | n11128 ;
  assign n11856 = n11854 &  n11855 ;
  assign n11857 = ( n11853 & ~n11125 ) | ( n11853 & n11856 ) | ( ~n11125 & n11856 ) ;
  assign n11858 = ( n11125 & ~n11188 ) | ( n11125 & n11128 ) | ( ~n11188 & n11128 ) ;
  assign n11859 = ( n11189 & ~n11128 ) | ( n11189 & n11858 ) | ( ~n11128 & n11858 ) ;
  assign n11860 = ~n5972 & n11859 ;
  assign n11861 = ( n11857 & ~n11860 ) | ( n11857 & 1'b0 ) | ( ~n11860 & 1'b0 ) ;
  assign n11862 = x17 &  n11861 ;
  assign n11863 = x17 | n11861 ;
  assign n11864 = ~n11862 & n11863 ;
  assign n11868 = ~n6395 & n11128 ;
  assign n11865 = ~n5970 & n11134 ;
  assign n11866 = n6170 | n11131 ;
  assign n11867 = ~n11865 & n11866 ;
  assign n11869 = ( n6395 & n11868 ) | ( n6395 & n11867 ) | ( n11868 & n11867 ) ;
  assign n11870 = ( n11128 & ~n11131 ) | ( n11128 & n11187 ) | ( ~n11131 & n11187 ) ;
  assign n11871 = ( n11131 & ~n11188 ) | ( n11131 & n11870 ) | ( ~n11188 & n11870 ) ;
  assign n11872 = n5972 | n11871 ;
  assign n11873 = n11869 &  n11872 ;
  assign n11874 = x17 &  n11873 ;
  assign n11875 = x17 | n11873 ;
  assign n11876 = ~n11874 & n11875 ;
  assign n11877 = ( n11680 & ~n11692 ) | ( n11680 & n11848 ) | ( ~n11692 & n11848 ) ;
  assign n11878 = ( n11692 & ~n11849 ) | ( n11692 & n11877 ) | ( ~n11849 & n11877 ) ;
  assign n11879 = ( n11704 & ~n11847 ) | ( n11704 & n11706 ) | ( ~n11847 & n11706 ) ;
  assign n11880 = ( n11706 & ~n11704 ) | ( n11706 & n11847 ) | ( ~n11704 & n11847 ) ;
  assign n11881 = ( n11879 & ~n11706 ) | ( n11879 & n11880 ) | ( ~n11706 & n11880 ) ;
  assign n11887 = ( n11131 & n11134 ) | ( n11131 & n11186 ) | ( n11134 & n11186 ) ;
  assign n11888 = ( n11134 & ~n11887 ) | ( n11134 & n11187 ) | ( ~n11887 & n11187 ) ;
  assign n11885 = ~n6395 & n11131 ;
  assign n11882 = n5970 | n11137 ;
  assign n11883 = ~n6170 & n11134 ;
  assign n11884 = ( n11882 & ~n11883 ) | ( n11882 & 1'b0 ) | ( ~n11883 & 1'b0 ) ;
  assign n11886 = ( n6395 & n11885 ) | ( n6395 & n11884 ) | ( n11885 & n11884 ) ;
  assign n11889 = ( n5972 & ~n11886 ) | ( n5972 & n11888 ) | ( ~n11886 & n11888 ) ;
  assign n11890 = ( n11888 & ~n11889 ) | ( n11888 & 1'b0 ) | ( ~n11889 & 1'b0 ) ;
  assign n11892 = ( x17 & n11886 ) | ( x17 & n11890 ) | ( n11886 & n11890 ) ;
  assign n11891 = ( x17 & ~n11890 ) | ( x17 & n11886 ) | ( ~n11890 & n11886 ) ;
  assign n11893 = ( n11890 & ~n11892 ) | ( n11890 & n11891 ) | ( ~n11892 & n11891 ) ;
  assign n11900 = n11134 | n6395 ;
  assign n11897 = n5970 | n11140 ;
  assign n11898 = n6170 | n11137 ;
  assign n11899 = n11897 &  n11898 ;
  assign n11901 = ( n6395 & ~n11900 ) | ( n6395 & n11899 ) | ( ~n11900 & n11899 ) ;
  assign n11902 = ( n5972 & ~n11901 ) | ( n5972 & n11242 ) | ( ~n11901 & n11242 ) ;
  assign n11903 = ( n11242 & ~n11902 ) | ( n11242 & 1'b0 ) | ( ~n11902 & 1'b0 ) ;
  assign n11905 = ( x17 & n11901 ) | ( x17 & n11903 ) | ( n11901 & n11903 ) ;
  assign n11904 = ( x17 & ~n11903 ) | ( x17 & n11901 ) | ( ~n11903 & n11901 ) ;
  assign n11906 = ( n11903 & ~n11905 ) | ( n11903 & n11904 ) | ( ~n11905 & n11904 ) ;
  assign n11894 = ( n11716 & ~n11846 ) | ( n11716 & n11718 ) | ( ~n11846 & n11718 ) ;
  assign n11895 = ( n11718 & ~n11716 ) | ( n11718 & n11846 ) | ( ~n11716 & n11846 ) ;
  assign n11896 = ( n11894 & ~n11718 ) | ( n11894 & n11895 ) | ( ~n11718 & n11895 ) ;
  assign n11910 = ~n6395 & n11137 ;
  assign n11907 = n5970 | n11143 ;
  assign n11908 = n6170 | n11140 ;
  assign n11909 = n11907 &  n11908 ;
  assign n11911 = ( n6395 & n11910 ) | ( n6395 & n11909 ) | ( n11910 & n11909 ) ;
  assign n11912 = n5972 | n11687 ;
  assign n11913 = n11911 &  n11912 ;
  assign n11914 = x17 &  n11913 ;
  assign n11915 = x17 | n11913 ;
  assign n11916 = ~n11914 & n11915 ;
  assign n11917 = ( n11721 & ~n11845 ) | ( n11721 & n11731 ) | ( ~n11845 & n11731 ) ;
  assign n11918 = ( n11846 & ~n11731 ) | ( n11846 & n11917 ) | ( ~n11731 & n11917 ) ;
  assign n11922 = ~n6395 & n11140 ;
  assign n11919 = n5970 | n11146 ;
  assign n11920 = n6170 | n11143 ;
  assign n11921 = n11919 &  n11920 ;
  assign n11923 = ( n6395 & n11922 ) | ( n6395 & n11921 ) | ( n11922 & n11921 ) ;
  assign n11924 = n5972 | n11699 ;
  assign n11925 = n11923 &  n11924 ;
  assign n11926 = x17 &  n11925 ;
  assign n11927 = x17 | n11925 ;
  assign n11928 = ~n11926 & n11927 ;
  assign n11929 = ( n11734 & ~n11744 ) | ( n11734 & n11844 ) | ( ~n11744 & n11844 ) ;
  assign n11930 = ( n11744 & ~n11845 ) | ( n11744 & n11929 ) | ( ~n11845 & n11929 ) ;
  assign n11934 = ~n6395 & n11143 ;
  assign n11931 = n5970 | n11149 ;
  assign n11932 = n6170 | n11146 ;
  assign n11933 = n11931 &  n11932 ;
  assign n11935 = ( n6395 & n11934 ) | ( n6395 & n11933 ) | ( n11934 & n11933 ) ;
  assign n11936 = n5972 | n11542 ;
  assign n11937 = n11935 &  n11936 ;
  assign n11938 = x17 &  n11937 ;
  assign n11939 = x17 | n11937 ;
  assign n11940 = ~n11938 & n11939 ;
  assign n11941 = ( n11747 & n11757 ) | ( n11747 & n11843 ) | ( n11757 & n11843 ) ;
  assign n11942 = ( n11757 & ~n11941 ) | ( n11757 & n11844 ) | ( ~n11941 & n11844 ) ;
  assign n11949 = ~n6395 & n11146 ;
  assign n11946 = ~n5970 & n11152 ;
  assign n11947 = n6170 | n11149 ;
  assign n11948 = ~n11946 & n11947 ;
  assign n11950 = ( n6395 & n11949 ) | ( n6395 & n11948 ) | ( n11949 & n11948 ) ;
  assign n11951 = ( n5972 & ~n11950 ) | ( n5972 & n11554 ) | ( ~n11950 & n11554 ) ;
  assign n11952 = ( n11554 & ~n11951 ) | ( n11554 & 1'b0 ) | ( ~n11951 & 1'b0 ) ;
  assign n11953 = ( x17 & ~n11950 ) | ( x17 & n11952 ) | ( ~n11950 & n11952 ) ;
  assign n11954 = ( n11950 & ~x17 ) | ( n11950 & n11952 ) | ( ~x17 & n11952 ) ;
  assign n11955 = ( n11953 & ~n11952 ) | ( n11953 & n11954 ) | ( ~n11952 & n11954 ) ;
  assign n11943 = ( n11770 & ~n11767 ) | ( n11770 & n11842 ) | ( ~n11767 & n11842 ) ;
  assign n11944 = ( n11767 & ~n11842 ) | ( n11767 & n11770 ) | ( ~n11842 & n11770 ) ;
  assign n11945 = ( n11943 & ~n11770 ) | ( n11943 & n11944 ) | ( ~n11770 & n11944 ) ;
  assign n11956 = ( n11783 & ~n11773 ) | ( n11783 & n11841 ) | ( ~n11773 & n11841 ) ;
  assign n11957 = ( n11773 & ~n11841 ) | ( n11773 & n11783 ) | ( ~n11841 & n11783 ) ;
  assign n11958 = ( n11956 & ~n11783 ) | ( n11956 & n11957 ) | ( ~n11783 & n11957 ) ;
  assign n11959 = ~n5970 & n11155 ;
  assign n11960 = ~n6170 & n11152 ;
  assign n11961 = n11959 | n11960 ;
  assign n11962 = ~n6395 & n11149 ;
  assign n11963 = ( n6395 & ~n11961 ) | ( n6395 & n11962 ) | ( ~n11961 & n11962 ) ;
  assign n11964 = ( n11572 & ~n5972 ) | ( n11572 & n11963 ) | ( ~n5972 & n11963 ) ;
  assign n11965 = ~n11572 & n11964 ;
  assign n11967 = ( x17 & n11963 ) | ( x17 & n11965 ) | ( n11963 & n11965 ) ;
  assign n11966 = ( x17 & ~n11965 ) | ( x17 & n11963 ) | ( ~n11965 & n11963 ) ;
  assign n11968 = ( n11965 & ~n11967 ) | ( n11965 & n11966 ) | ( ~n11967 & n11966 ) ;
  assign n11969 = ( n11793 & ~n11840 ) | ( n11793 & n11798 ) | ( ~n11840 & n11798 ) ;
  assign n11970 = ( n11798 & ~n11793 ) | ( n11798 & n11840 ) | ( ~n11793 & n11840 ) ;
  assign n11971 = ( n11969 & ~n11798 ) | ( n11969 & n11970 ) | ( ~n11798 & n11970 ) ;
  assign n11975 = n11152 | n6395 ;
  assign n11972 = ~n5970 & n11158 ;
  assign n11973 = ~n6170 & n11155 ;
  assign n11974 = n11972 | n11973 ;
  assign n11976 = ( n11975 & ~n6395 ) | ( n11975 & n11974 ) | ( ~n6395 & n11974 ) ;
  assign n11977 = ( n5972 & n11254 ) | ( n5972 & n11976 ) | ( n11254 & n11976 ) ;
  assign n11978 = ( n11254 & ~n11977 ) | ( n11254 & 1'b0 ) | ( ~n11977 & 1'b0 ) ;
  assign n11979 = ( n11976 & ~x17 ) | ( n11976 & n11978 ) | ( ~x17 & n11978 ) ;
  assign n11980 = ( x17 & ~n11976 ) | ( x17 & n11978 ) | ( ~n11976 & n11978 ) ;
  assign n11981 = ( n11979 & ~n11978 ) | ( n11979 & n11980 ) | ( ~n11978 & n11980 ) ;
  assign n11985 = n11155 | n6395 ;
  assign n11982 = n5970 | n11161 ;
  assign n11983 = ~n6170 & n11158 ;
  assign n11984 = ( n11982 & ~n11983 ) | ( n11982 & 1'b0 ) | ( ~n11983 & 1'b0 ) ;
  assign n11986 = ( n6395 & ~n11985 ) | ( n6395 & n11984 ) | ( ~n11985 & n11984 ) ;
  assign n11987 = n5972 | n11451 ;
  assign n11988 = n11986 &  n11987 ;
  assign n11989 = x17 &  n11988 ;
  assign n11990 = x17 | n11988 ;
  assign n11991 = ~n11989 & n11990 ;
  assign n11992 = ( n11812 & ~n11802 ) | ( n11812 & n11839 ) | ( ~n11802 & n11839 ) ;
  assign n11993 = ( n11840 & ~n11812 ) | ( n11840 & n11992 ) | ( ~n11812 & n11992 ) ;
  assign n11995 = ( n11641 & n11828 ) | ( n11641 & n11838 ) | ( n11828 & n11838 ) ;
  assign n11994 = ( n11641 & ~n11828 ) | ( n11641 & n11838 ) | ( ~n11828 & n11838 ) ;
  assign n11996 = ( n11828 & ~n11995 ) | ( n11828 & n11994 ) | ( ~n11995 & n11994 ) ;
  assign n11997 = n6395 &  n11158 ;
  assign n11998 = n5970 | n11164 ;
  assign n11999 = n6170 | n11161 ;
  assign n12000 = n11998 &  n11999 ;
  assign n12001 = ( n11997 & ~n11158 ) | ( n11997 & n12000 ) | ( ~n11158 & n12000 ) ;
  assign n12002 = ( n5972 & ~n12001 ) | ( n5972 & n11463 ) | ( ~n12001 & n11463 ) ;
  assign n12003 = ( n11463 & ~n12002 ) | ( n11463 & 1'b0 ) | ( ~n12002 & 1'b0 ) ;
  assign n12005 = ( x17 & n12001 ) | ( x17 & n12003 ) | ( n12001 & n12003 ) ;
  assign n12004 = ( x17 & ~n12003 ) | ( x17 & n12001 ) | ( ~n12003 & n12001 ) ;
  assign n12006 = ( n12003 & ~n12005 ) | ( n12003 & n12004 ) | ( ~n12005 & n12004 ) ;
  assign n12010 = ~n6395 & n11161 ;
  assign n12007 = n5970 | n11166 ;
  assign n12008 = n6170 | n11164 ;
  assign n12009 = n12007 &  n12008 ;
  assign n12011 = ( n6395 & n12010 ) | ( n6395 & n12009 ) | ( n12010 & n12009 ) ;
  assign n12012 = n5972 | n11385 ;
  assign n12013 = n12011 &  n12012 ;
  assign n12014 = x17 &  n12013 ;
  assign n12015 = x17 | n12013 ;
  assign n12016 = ~n12014 & n12015 ;
  assign n12017 = ( x20 & n11813 ) | ( x20 & n11818 ) | ( n11813 & n11818 ) ;
  assign n12018 = ~n11813 & n12017 ;
  assign n12019 = ( n11825 & ~x20 ) | ( n11825 & n12018 ) | ( ~x20 & n12018 ) ;
  assign n12020 = ( x20 & ~n11825 ) | ( x20 & n12018 ) | ( ~n11825 & n12018 ) ;
  assign n12021 = ( n12019 & ~n12018 ) | ( n12019 & n12020 ) | ( ~n12018 & n12020 ) ;
  assign n12022 = x20 &  n11813 ;
  assign n12023 = n11818 &  n12022 ;
  assign n12024 = n11818 | n12022 ;
  assign n12025 = ~n12023 & n12024 ;
  assign n12055 = ~n6395 & n11166 ;
  assign n12052 = n5970 | n11172 ;
  assign n12053 = n6170 | n11168 ;
  assign n12054 = n12052 &  n12053 ;
  assign n12056 = ( n6395 & n12055 ) | ( n6395 & n12054 ) | ( n12055 & n12054 ) ;
  assign n12057 = n5972 | n11431 ;
  assign n12058 = n12056 &  n12057 ;
  assign n12059 = x17 &  n12058 ;
  assign n12060 = x17 | n12058 ;
  assign n12061 = ~n12059 & n12060 ;
  assign n12036 = n5965 &  n11170 ;
  assign n12040 = ~n5972 & n11369 ;
  assign n12037 = ~n6170 & n11170 ;
  assign n12038 = n6395 | n11172 ;
  assign n12039 = ~n12037 & n12038 ;
  assign n12041 = ( n5972 & n12040 ) | ( n5972 & n12039 ) | ( n12040 & n12039 ) ;
  assign n12047 = n11323 | n5972 ;
  assign n12045 = ~n6395 & n11168 ;
  assign n12042 = ~n5970 & n11170 ;
  assign n12043 = n6170 | n11172 ;
  assign n12044 = ~n12042 & n12043 ;
  assign n12046 = ( n6395 & n12045 ) | ( n6395 & n12044 ) | ( n12045 & n12044 ) ;
  assign n12048 = ( n5972 & ~n12047 ) | ( n5972 & n12046 ) | ( ~n12047 & n12046 ) ;
  assign n12049 = ( n12036 & n12041 ) | ( n12036 & n12048 ) | ( n12041 & n12048 ) ;
  assign n12050 = ( x17 & ~n12049 ) | ( x17 & n12036 ) | ( ~n12049 & n12036 ) ;
  assign n12051 = ( x17 & ~n12050 ) | ( x17 & 1'b0 ) | ( ~n12050 & 1'b0 ) ;
  assign n12062 = ( n11813 & ~n12061 ) | ( n11813 & n12051 ) | ( ~n12061 & n12051 ) ;
  assign n12029 = ~n6395 & n11164 ;
  assign n12026 = n5970 | n11168 ;
  assign n12027 = n6170 | n11166 ;
  assign n12028 = n12026 &  n12027 ;
  assign n12030 = ( n6395 & n12029 ) | ( n6395 & n12028 ) | ( n12029 & n12028 ) ;
  assign n12031 = ( n11397 & ~n5972 ) | ( n11397 & n12030 ) | ( ~n5972 & n12030 ) ;
  assign n12032 = ~n11397 & n12031 ;
  assign n12033 = ( x17 & ~n12030 ) | ( x17 & n12032 ) | ( ~n12030 & n12032 ) ;
  assign n12034 = ( n12030 & ~x17 ) | ( n12030 & n12032 ) | ( ~x17 & n12032 ) ;
  assign n12035 = ( n12033 & ~n12032 ) | ( n12033 & n12034 ) | ( ~n12032 & n12034 ) ;
  assign n12063 = ( n12025 & ~n12062 ) | ( n12025 & n12035 ) | ( ~n12062 & n12035 ) ;
  assign n12064 = ( n12016 & n12021 ) | ( n12016 & n12063 ) | ( n12021 & n12063 ) ;
  assign n12065 = ( n11996 & n12006 ) | ( n11996 & n12064 ) | ( n12006 & n12064 ) ;
  assign n12066 = ( n11991 & ~n11993 ) | ( n11991 & n12065 ) | ( ~n11993 & n12065 ) ;
  assign n12067 = ( n11971 & ~n11981 ) | ( n11971 & n12066 ) | ( ~n11981 & n12066 ) ;
  assign n12068 = ( n11958 & n11968 ) | ( n11958 & n12067 ) | ( n11968 & n12067 ) ;
  assign n12069 = ( n11955 & ~n11945 ) | ( n11955 & n12068 ) | ( ~n11945 & n12068 ) ;
  assign n12070 = ( n11940 & ~n11942 ) | ( n11940 & n12069 ) | ( ~n11942 & n12069 ) ;
  assign n12071 = ( n11928 & n11930 ) | ( n11928 & n12070 ) | ( n11930 & n12070 ) ;
  assign n12072 = ( n11916 & ~n11918 ) | ( n11916 & n12071 ) | ( ~n11918 & n12071 ) ;
  assign n12073 = ( n11906 & ~n11896 ) | ( n11906 & n12072 ) | ( ~n11896 & n12072 ) ;
  assign n12074 = ( n11881 & n11893 ) | ( n11881 & n12073 ) | ( n11893 & n12073 ) ;
  assign n12075 = ( n11876 & n11878 ) | ( n11876 & n12074 ) | ( n11878 & n12074 ) ;
  assign n12076 = ( n11852 & ~n11864 ) | ( n11852 & n12075 ) | ( ~n11864 & n12075 ) ;
  assign n12077 = ( n11852 & ~n12075 ) | ( n11852 & n11864 ) | ( ~n12075 & n11864 ) ;
  assign n12078 = ( n12076 & ~n11852 ) | ( n12076 & n12077 ) | ( ~n11852 & n12077 ) ;
  assign n12079 = ( n11878 & ~n11876 ) | ( n11878 & n12074 ) | ( ~n11876 & n12074 ) ;
  assign n12080 = ( n11876 & ~n12074 ) | ( n11876 & n11878 ) | ( ~n12074 & n11878 ) ;
  assign n12081 = ( n12079 & ~n11878 ) | ( n12079 & n12080 ) | ( ~n11878 & n12080 ) ;
  assign n12082 = n7097 &  n11119 ;
  assign n12083 = ~n6530 & n11125 ;
  assign n12084 = n6983 | n11122 ;
  assign n12085 = ~n12083 & n12084 ;
  assign n12086 = ( n12082 & ~n11119 ) | ( n12082 & n12085 ) | ( ~n11119 & n12085 ) ;
  assign n12087 = ( n11119 & ~n11190 ) | ( n11119 & n11122 ) | ( ~n11190 & n11122 ) ;
  assign n12088 = ( n11191 & ~n11122 ) | ( n11191 & n12087 ) | ( ~n11122 & n12087 ) ;
  assign n12089 = ( n6532 & ~n12086 ) | ( n6532 & n12088 ) | ( ~n12086 & n12088 ) ;
  assign n12090 = ( n12088 & ~n12089 ) | ( n12088 & 1'b0 ) | ( ~n12089 & 1'b0 ) ;
  assign n12091 = ( x14 & ~n12086 ) | ( x14 & n12090 ) | ( ~n12086 & n12090 ) ;
  assign n12092 = ( n12086 & ~x14 ) | ( n12086 & n12090 ) | ( ~x14 & n12090 ) ;
  assign n12093 = ( n12091 & ~n12090 ) | ( n12091 & n12092 ) | ( ~n12090 & n12092 ) ;
  assign n12097 = ~n7097 & n11122 ;
  assign n12094 = n6530 | n11128 ;
  assign n12095 = ~n6983 & n11125 ;
  assign n12096 = ( n12094 & ~n12095 ) | ( n12094 & 1'b0 ) | ( ~n12095 & 1'b0 ) ;
  assign n12098 = ( n7097 & n12097 ) | ( n7097 & n12096 ) | ( n12097 & n12096 ) ;
  assign n12099 = ( n11122 & n11125 ) | ( n11122 & n11189 ) | ( n11125 & n11189 ) ;
  assign n12100 = ( n11125 & ~n12099 ) | ( n11125 & n11190 ) | ( ~n12099 & n11190 ) ;
  assign n12101 = ~n6532 & n12100 ;
  assign n12102 = ( n12098 & ~n12101 ) | ( n12098 & 1'b0 ) | ( ~n12101 & 1'b0 ) ;
  assign n12103 = x14 &  n12102 ;
  assign n12104 = x14 | n12102 ;
  assign n12105 = ~n12103 & n12104 ;
  assign n12106 = ( n11881 & ~n11893 ) | ( n11881 & n12073 ) | ( ~n11893 & n12073 ) ;
  assign n12107 = ( n11893 & ~n12074 ) | ( n11893 & n12106 ) | ( ~n12074 & n12106 ) ;
  assign n12108 = n7097 &  n11125 ;
  assign n12109 = n6530 | n11131 ;
  assign n12110 = n6983 | n11128 ;
  assign n12111 = n12109 &  n12110 ;
  assign n12112 = ( n12108 & ~n11125 ) | ( n12108 & n12111 ) | ( ~n11125 & n12111 ) ;
  assign n12113 = ~n6532 & n11859 ;
  assign n12114 = ( n12112 & ~n12113 ) | ( n12112 & 1'b0 ) | ( ~n12113 & 1'b0 ) ;
  assign n12115 = x14 &  n12114 ;
  assign n12116 = x14 | n12114 ;
  assign n12117 = ~n12115 & n12116 ;
  assign n12118 = ( n11896 & ~n12072 ) | ( n11896 & n11906 ) | ( ~n12072 & n11906 ) ;
  assign n12119 = ( n12073 & ~n11906 ) | ( n12073 & n12118 ) | ( ~n11906 & n12118 ) ;
  assign n12126 = ~n7097 & n11128 ;
  assign n12123 = ~n6530 & n11134 ;
  assign n12124 = n6983 | n11131 ;
  assign n12125 = ~n12123 & n12124 ;
  assign n12127 = ( n7097 & n12126 ) | ( n7097 & n12125 ) | ( n12126 & n12125 ) ;
  assign n12128 = ( n11871 & ~n6532 ) | ( n11871 & n12127 ) | ( ~n6532 & n12127 ) ;
  assign n12129 = ~n11871 & n12128 ;
  assign n12130 = ( x14 & ~n12127 ) | ( x14 & n12129 ) | ( ~n12127 & n12129 ) ;
  assign n12131 = ( n12127 & ~x14 ) | ( n12127 & n12129 ) | ( ~x14 & n12129 ) ;
  assign n12132 = ( n12130 & ~n12129 ) | ( n12130 & n12131 ) | ( ~n12129 & n12131 ) ;
  assign n12120 = ( n11918 & ~n11916 ) | ( n11918 & n12071 ) | ( ~n11916 & n12071 ) ;
  assign n12121 = ( n11916 & ~n12071 ) | ( n11916 & n11918 ) | ( ~n12071 & n11918 ) ;
  assign n12122 = ( n12120 & ~n11918 ) | ( n12120 & n12121 ) | ( ~n11918 & n12121 ) ;
  assign n12133 = ( n11930 & ~n11928 ) | ( n11930 & n12070 ) | ( ~n11928 & n12070 ) ;
  assign n12134 = ( n11928 & ~n12070 ) | ( n11928 & n11930 ) | ( ~n12070 & n11930 ) ;
  assign n12135 = ( n12133 & ~n11930 ) | ( n12133 & n12134 ) | ( ~n11930 & n12134 ) ;
  assign n12139 = ~n7097 & n11131 ;
  assign n12136 = n6530 | n11137 ;
  assign n12137 = ~n6983 & n11134 ;
  assign n12138 = ( n12136 & ~n12137 ) | ( n12136 & 1'b0 ) | ( ~n12137 & 1'b0 ) ;
  assign n12140 = ( n7097 & n12139 ) | ( n7097 & n12138 ) | ( n12139 & n12138 ) ;
  assign n12141 = ( n6532 & ~n12140 ) | ( n6532 & n11888 ) | ( ~n12140 & n11888 ) ;
  assign n12142 = ( n11888 & ~n12141 ) | ( n11888 & 1'b0 ) | ( ~n12141 & 1'b0 ) ;
  assign n12144 = ( x14 & n12140 ) | ( x14 & n12142 ) | ( n12140 & n12142 ) ;
  assign n12143 = ( x14 & ~n12142 ) | ( x14 & n12140 ) | ( ~n12142 & n12140 ) ;
  assign n12145 = ( n12142 & ~n12144 ) | ( n12142 & n12143 ) | ( ~n12144 & n12143 ) ;
  assign n12152 = n11134 | n7097 ;
  assign n12149 = n6530 | n11140 ;
  assign n12150 = n6983 | n11137 ;
  assign n12151 = n12149 &  n12150 ;
  assign n12153 = ( n7097 & ~n12152 ) | ( n7097 & n12151 ) | ( ~n12152 & n12151 ) ;
  assign n12154 = ( n6532 & ~n12153 ) | ( n6532 & n11242 ) | ( ~n12153 & n11242 ) ;
  assign n12155 = ( n11242 & ~n12154 ) | ( n11242 & 1'b0 ) | ( ~n12154 & 1'b0 ) ;
  assign n12157 = ( x14 & n12153 ) | ( x14 & n12155 ) | ( n12153 & n12155 ) ;
  assign n12156 = ( x14 & ~n12155 ) | ( x14 & n12153 ) | ( ~n12155 & n12153 ) ;
  assign n12158 = ( n12155 & ~n12157 ) | ( n12155 & n12156 ) | ( ~n12157 & n12156 ) ;
  assign n12146 = ( n11940 & ~n12069 ) | ( n11940 & n11942 ) | ( ~n12069 & n11942 ) ;
  assign n12147 = ( n11942 & ~n11940 ) | ( n11942 & n12069 ) | ( ~n11940 & n12069 ) ;
  assign n12148 = ( n12146 & ~n11942 ) | ( n12146 & n12147 ) | ( ~n11942 & n12147 ) ;
  assign n12162 = ~n7097 & n11137 ;
  assign n12159 = n6530 | n11143 ;
  assign n12160 = n6983 | n11140 ;
  assign n12161 = n12159 &  n12160 ;
  assign n12163 = ( n7097 & n12162 ) | ( n7097 & n12161 ) | ( n12162 & n12161 ) ;
  assign n12164 = n6532 | n11687 ;
  assign n12165 = n12163 &  n12164 ;
  assign n12166 = x14 &  n12165 ;
  assign n12167 = x14 | n12165 ;
  assign n12168 = ~n12166 & n12167 ;
  assign n12169 = ( n11945 & ~n12068 ) | ( n11945 & n11955 ) | ( ~n12068 & n11955 ) ;
  assign n12170 = ( n12069 & ~n11955 ) | ( n12069 & n12169 ) | ( ~n11955 & n12169 ) ;
  assign n12174 = ~n7097 & n11140 ;
  assign n12171 = n6530 | n11146 ;
  assign n12172 = n6983 | n11143 ;
  assign n12173 = n12171 &  n12172 ;
  assign n12175 = ( n7097 & n12174 ) | ( n7097 & n12173 ) | ( n12174 & n12173 ) ;
  assign n12176 = n6532 | n11699 ;
  assign n12177 = n12175 &  n12176 ;
  assign n12178 = x14 &  n12177 ;
  assign n12179 = x14 | n12177 ;
  assign n12180 = ~n12178 & n12179 ;
  assign n12181 = ( n11958 & ~n11968 ) | ( n11958 & n12067 ) | ( ~n11968 & n12067 ) ;
  assign n12182 = ( n11968 & ~n12068 ) | ( n11968 & n12181 ) | ( ~n12068 & n12181 ) ;
  assign n12186 = ~n7097 & n11143 ;
  assign n12183 = n6530 | n11149 ;
  assign n12184 = n6983 | n11146 ;
  assign n12185 = n12183 &  n12184 ;
  assign n12187 = ( n7097 & n12186 ) | ( n7097 & n12185 ) | ( n12186 & n12185 ) ;
  assign n12188 = n6532 | n11542 ;
  assign n12189 = n12187 &  n12188 ;
  assign n12190 = x14 &  n12189 ;
  assign n12191 = x14 | n12189 ;
  assign n12192 = ~n12190 & n12191 ;
  assign n12193 = ( n11971 & n11981 ) | ( n11971 & n12066 ) | ( n11981 & n12066 ) ;
  assign n12194 = ( n11981 & ~n12193 ) | ( n11981 & n12067 ) | ( ~n12193 & n12067 ) ;
  assign n12201 = ~n7097 & n11146 ;
  assign n12198 = ~n6530 & n11152 ;
  assign n12199 = n6983 | n11149 ;
  assign n12200 = ~n12198 & n12199 ;
  assign n12202 = ( n7097 & n12201 ) | ( n7097 & n12200 ) | ( n12201 & n12200 ) ;
  assign n12203 = ( n6532 & ~n12202 ) | ( n6532 & n11554 ) | ( ~n12202 & n11554 ) ;
  assign n12204 = ( n11554 & ~n12203 ) | ( n11554 & 1'b0 ) | ( ~n12203 & 1'b0 ) ;
  assign n12205 = ( x14 & ~n12202 ) | ( x14 & n12204 ) | ( ~n12202 & n12204 ) ;
  assign n12206 = ( n12202 & ~x14 ) | ( n12202 & n12204 ) | ( ~x14 & n12204 ) ;
  assign n12207 = ( n12205 & ~n12204 ) | ( n12205 & n12206 ) | ( ~n12204 & n12206 ) ;
  assign n12195 = ( n11993 & ~n11991 ) | ( n11993 & n12065 ) | ( ~n11991 & n12065 ) ;
  assign n12196 = ( n11991 & ~n12065 ) | ( n11991 & n11993 ) | ( ~n12065 & n11993 ) ;
  assign n12197 = ( n12195 & ~n11993 ) | ( n12195 & n12196 ) | ( ~n11993 & n12196 ) ;
  assign n12208 = ( n12006 & ~n11996 ) | ( n12006 & n12064 ) | ( ~n11996 & n12064 ) ;
  assign n12209 = ( n11996 & ~n12064 ) | ( n11996 & n12006 ) | ( ~n12064 & n12006 ) ;
  assign n12210 = ( n12208 & ~n12006 ) | ( n12208 & n12209 ) | ( ~n12006 & n12209 ) ;
  assign n12211 = ~n6530 & n11155 ;
  assign n12212 = ~n6983 & n11152 ;
  assign n12213 = n12211 | n12212 ;
  assign n12214 = ~n7097 & n11149 ;
  assign n12215 = ( n7097 & ~n12213 ) | ( n7097 & n12214 ) | ( ~n12213 & n12214 ) ;
  assign n12216 = ( n11572 & ~n6532 ) | ( n11572 & n12215 ) | ( ~n6532 & n12215 ) ;
  assign n12217 = ~n11572 & n12216 ;
  assign n12219 = ( x14 & n12215 ) | ( x14 & n12217 ) | ( n12215 & n12217 ) ;
  assign n12218 = ( x14 & ~n12217 ) | ( x14 & n12215 ) | ( ~n12217 & n12215 ) ;
  assign n12220 = ( n12217 & ~n12219 ) | ( n12217 & n12218 ) | ( ~n12219 & n12218 ) ;
  assign n12221 = ( n12016 & ~n12063 ) | ( n12016 & n12021 ) | ( ~n12063 & n12021 ) ;
  assign n12222 = ( n12021 & ~n12016 ) | ( n12021 & n12063 ) | ( ~n12016 & n12063 ) ;
  assign n12223 = ( n12221 & ~n12021 ) | ( n12221 & n12222 ) | ( ~n12021 & n12222 ) ;
  assign n12227 = n11152 | n7097 ;
  assign n12224 = ~n6530 & n11158 ;
  assign n12225 = ~n6983 & n11155 ;
  assign n12226 = n12224 | n12225 ;
  assign n12228 = ( n12227 & ~n7097 ) | ( n12227 & n12226 ) | ( ~n7097 & n12226 ) ;
  assign n12229 = ( n6532 & n11254 ) | ( n6532 & n12228 ) | ( n11254 & n12228 ) ;
  assign n12230 = ( n11254 & ~n12229 ) | ( n11254 & 1'b0 ) | ( ~n12229 & 1'b0 ) ;
  assign n12231 = ( n12228 & ~x14 ) | ( n12228 & n12230 ) | ( ~x14 & n12230 ) ;
  assign n12232 = ( x14 & ~n12228 ) | ( x14 & n12230 ) | ( ~n12228 & n12230 ) ;
  assign n12233 = ( n12231 & ~n12230 ) | ( n12231 & n12232 ) | ( ~n12230 & n12232 ) ;
  assign n12237 = n11155 | n7097 ;
  assign n12234 = n6530 | n11161 ;
  assign n12235 = ~n6983 & n11158 ;
  assign n12236 = ( n12234 & ~n12235 ) | ( n12234 & 1'b0 ) | ( ~n12235 & 1'b0 ) ;
  assign n12238 = ( n7097 & ~n12237 ) | ( n7097 & n12236 ) | ( ~n12237 & n12236 ) ;
  assign n12239 = n6532 | n11451 ;
  assign n12240 = n12238 &  n12239 ;
  assign n12241 = x14 &  n12240 ;
  assign n12242 = x14 | n12240 ;
  assign n12243 = ~n12241 & n12242 ;
  assign n12244 = ( n12035 & ~n12025 ) | ( n12035 & n12062 ) | ( ~n12025 & n12062 ) ;
  assign n12245 = ( n12063 & ~n12035 ) | ( n12063 & n12244 ) | ( ~n12035 & n12244 ) ;
  assign n12247 = ( n11813 & n12051 ) | ( n11813 & n12061 ) | ( n12051 & n12061 ) ;
  assign n12246 = ( n11813 & ~n12051 ) | ( n11813 & n12061 ) | ( ~n12051 & n12061 ) ;
  assign n12248 = ( n12051 & ~n12247 ) | ( n12051 & n12246 ) | ( ~n12247 & n12246 ) ;
  assign n12249 = n7097 &  n11158 ;
  assign n12250 = n6530 | n11164 ;
  assign n12251 = n6983 | n11161 ;
  assign n12252 = n12250 &  n12251 ;
  assign n12253 = ( n12249 & ~n11158 ) | ( n12249 & n12252 ) | ( ~n11158 & n12252 ) ;
  assign n12254 = ( n6532 & ~n12253 ) | ( n6532 & n11463 ) | ( ~n12253 & n11463 ) ;
  assign n12255 = ( n11463 & ~n12254 ) | ( n11463 & 1'b0 ) | ( ~n12254 & 1'b0 ) ;
  assign n12257 = ( x14 & n12253 ) | ( x14 & n12255 ) | ( n12253 & n12255 ) ;
  assign n12256 = ( x14 & ~n12255 ) | ( x14 & n12253 ) | ( ~n12255 & n12253 ) ;
  assign n12258 = ( n12255 & ~n12257 ) | ( n12255 & n12256 ) | ( ~n12257 & n12256 ) ;
  assign n12262 = ~n7097 & n11161 ;
  assign n12259 = n6530 | n11166 ;
  assign n12260 = n6983 | n11164 ;
  assign n12261 = n12259 &  n12260 ;
  assign n12263 = ( n7097 & n12262 ) | ( n7097 & n12261 ) | ( n12262 & n12261 ) ;
  assign n12264 = n6532 | n11385 ;
  assign n12265 = n12263 &  n12264 ;
  assign n12266 = x14 &  n12265 ;
  assign n12267 = x14 | n12265 ;
  assign n12268 = ~n12266 & n12267 ;
  assign n12269 = ( x17 & n12036 ) | ( x17 & n12041 ) | ( n12036 & n12041 ) ;
  assign n12270 = ~n12036 & n12269 ;
  assign n12271 = ( n12048 & ~x17 ) | ( n12048 & n12270 ) | ( ~x17 & n12270 ) ;
  assign n12272 = ( x17 & ~n12048 ) | ( x17 & n12270 ) | ( ~n12048 & n12270 ) ;
  assign n12273 = ( n12271 & ~n12270 ) | ( n12271 & n12272 ) | ( ~n12270 & n12272 ) ;
  assign n12274 = x17 &  n12036 ;
  assign n12275 = n12041 &  n12274 ;
  assign n12276 = n12041 | n12274 ;
  assign n12277 = ~n12275 & n12276 ;
  assign n12307 = ~n7097 & n11166 ;
  assign n12304 = n6530 | n11172 ;
  assign n12305 = n6983 | n11168 ;
  assign n12306 = n12304 &  n12305 ;
  assign n12308 = ( n7097 & n12307 ) | ( n7097 & n12306 ) | ( n12307 & n12306 ) ;
  assign n12309 = n6532 | n11431 ;
  assign n12310 = n12308 &  n12309 ;
  assign n12311 = x14 &  n12310 ;
  assign n12312 = x14 | n12310 ;
  assign n12313 = ~n12311 & n12312 ;
  assign n12288 = n6525 &  n11170 ;
  assign n12292 = ~n6532 & n11369 ;
  assign n12289 = ~n6983 & n11170 ;
  assign n12290 = n7097 | n11172 ;
  assign n12291 = ~n12289 & n12290 ;
  assign n12293 = ( n6532 & n12292 ) | ( n6532 & n12291 ) | ( n12292 & n12291 ) ;
  assign n12299 = n11323 | n6532 ;
  assign n12297 = ~n7097 & n11168 ;
  assign n12294 = ~n6530 & n11170 ;
  assign n12295 = n6983 | n11172 ;
  assign n12296 = ~n12294 & n12295 ;
  assign n12298 = ( n7097 & n12297 ) | ( n7097 & n12296 ) | ( n12297 & n12296 ) ;
  assign n12300 = ( n6532 & ~n12299 ) | ( n6532 & n12298 ) | ( ~n12299 & n12298 ) ;
  assign n12301 = ( n12288 & n12293 ) | ( n12288 & n12300 ) | ( n12293 & n12300 ) ;
  assign n12302 = ( x14 & ~n12301 ) | ( x14 & n12288 ) | ( ~n12301 & n12288 ) ;
  assign n12303 = ( x14 & ~n12302 ) | ( x14 & 1'b0 ) | ( ~n12302 & 1'b0 ) ;
  assign n12314 = ( n12036 & ~n12313 ) | ( n12036 & n12303 ) | ( ~n12313 & n12303 ) ;
  assign n12281 = ~n7097 & n11164 ;
  assign n12278 = n6530 | n11168 ;
  assign n12279 = n6983 | n11166 ;
  assign n12280 = n12278 &  n12279 ;
  assign n12282 = ( n7097 & n12281 ) | ( n7097 & n12280 ) | ( n12281 & n12280 ) ;
  assign n12283 = ( n11397 & ~n6532 ) | ( n11397 & n12282 ) | ( ~n6532 & n12282 ) ;
  assign n12284 = ~n11397 & n12283 ;
  assign n12285 = ( x14 & ~n12282 ) | ( x14 & n12284 ) | ( ~n12282 & n12284 ) ;
  assign n12286 = ( n12282 & ~x14 ) | ( n12282 & n12284 ) | ( ~x14 & n12284 ) ;
  assign n12287 = ( n12285 & ~n12284 ) | ( n12285 & n12286 ) | ( ~n12284 & n12286 ) ;
  assign n12315 = ( n12277 & ~n12314 ) | ( n12277 & n12287 ) | ( ~n12314 & n12287 ) ;
  assign n12316 = ( n12268 & n12273 ) | ( n12268 & n12315 ) | ( n12273 & n12315 ) ;
  assign n12317 = ( n12248 & n12258 ) | ( n12248 & n12316 ) | ( n12258 & n12316 ) ;
  assign n12318 = ( n12243 & ~n12245 ) | ( n12243 & n12317 ) | ( ~n12245 & n12317 ) ;
  assign n12319 = ( n12223 & ~n12233 ) | ( n12223 & n12318 ) | ( ~n12233 & n12318 ) ;
  assign n12320 = ( n12210 & n12220 ) | ( n12210 & n12319 ) | ( n12220 & n12319 ) ;
  assign n12321 = ( n12207 & ~n12197 ) | ( n12207 & n12320 ) | ( ~n12197 & n12320 ) ;
  assign n12322 = ( n12192 & ~n12194 ) | ( n12192 & n12321 ) | ( ~n12194 & n12321 ) ;
  assign n12323 = ( n12180 & n12182 ) | ( n12180 & n12322 ) | ( n12182 & n12322 ) ;
  assign n12324 = ( n12168 & ~n12170 ) | ( n12168 & n12323 ) | ( ~n12170 & n12323 ) ;
  assign n12325 = ( n12158 & ~n12148 ) | ( n12158 & n12324 ) | ( ~n12148 & n12324 ) ;
  assign n12326 = ( n12135 & n12145 ) | ( n12135 & n12325 ) | ( n12145 & n12325 ) ;
  assign n12327 = ( n12132 & ~n12122 ) | ( n12132 & n12326 ) | ( ~n12122 & n12326 ) ;
  assign n12328 = ( n12117 & ~n12119 ) | ( n12117 & n12327 ) | ( ~n12119 & n12327 ) ;
  assign n12329 = ( n12105 & n12107 ) | ( n12105 & n12328 ) | ( n12107 & n12328 ) ;
  assign n12330 = ( n12081 & n12093 ) | ( n12081 & n12329 ) | ( n12093 & n12329 ) ;
  assign n12331 = ( n11235 & n12078 ) | ( n11235 & n12330 ) | ( n12078 & n12330 ) ;
  assign n12332 = ( n12078 & ~n11235 ) | ( n12078 & n12330 ) | ( ~n11235 & n12330 ) ;
  assign n12333 = ( n11235 & ~n12331 ) | ( n11235 & n12332 ) | ( ~n12331 & n12332 ) ;
  assign n12337 = n11107 | n7783 ;
  assign n12334 = ( n7253 & ~n11113 ) | ( n7253 & 1'b0 ) | ( ~n11113 & 1'b0 ) ;
  assign n12335 = n7518 | n11110 ;
  assign n12336 = ~n12334 & n12335 ;
  assign n12338 = ( n7783 & ~n12337 ) | ( n7783 & n12336 ) | ( ~n12337 & n12336 ) ;
  assign n12339 = ( n11107 & n11110 ) | ( n11107 & n11194 ) | ( n11110 & n11194 ) ;
  assign n12340 = ( n11107 & ~n12339 ) | ( n11107 & n11195 ) | ( ~n12339 & n11195 ) ;
  assign n12341 = ~n7255 & n12340 ;
  assign n12342 = ( n12338 & ~n12341 ) | ( n12338 & 1'b0 ) | ( ~n12341 & 1'b0 ) ;
  assign n12343 = x11 &  n12342 ;
  assign n12344 = x11 | n12342 ;
  assign n12345 = ~n12343 & n12344 ;
  assign n12349 = ~n7783 & n11110 ;
  assign n12346 = n7253 &  n11116 ;
  assign n12347 = n7518 | n11113 ;
  assign n12348 = ~n12346 & n12347 ;
  assign n12350 = ( n7783 & n12349 ) | ( n7783 & n12348 ) | ( n12349 & n12348 ) ;
  assign n12351 = ( n11113 & ~n11110 ) | ( n11113 & n11193 ) | ( ~n11110 & n11193 ) ;
  assign n12352 = ( n11194 & ~n11113 ) | ( n11194 & n12351 ) | ( ~n11113 & n12351 ) ;
  assign n12353 = ~n7255 & n12352 ;
  assign n12354 = ( n12350 & ~n12353 ) | ( n12350 & 1'b0 ) | ( ~n12353 & 1'b0 ) ;
  assign n12355 = x11 &  n12354 ;
  assign n12356 = x11 | n12354 ;
  assign n12357 = ~n12355 & n12356 ;
  assign n12358 = ( n12081 & ~n12093 ) | ( n12081 & n12329 ) | ( ~n12093 & n12329 ) ;
  assign n12359 = ( n12093 & ~n12330 ) | ( n12093 & n12358 ) | ( ~n12330 & n12358 ) ;
  assign n12360 = ( n12105 & ~n12328 ) | ( n12105 & n12107 ) | ( ~n12328 & n12107 ) ;
  assign n12361 = ( n12107 & ~n12105 ) | ( n12107 & n12328 ) | ( ~n12105 & n12328 ) ;
  assign n12362 = ( n12360 & ~n12107 ) | ( n12360 & n12361 ) | ( ~n12107 & n12361 ) ;
  assign n12368 = ( n11113 & ~n11192 ) | ( n11113 & n11116 ) | ( ~n11192 & n11116 ) ;
  assign n12369 = ( n11193 & ~n11116 ) | ( n11193 & n12368 ) | ( ~n11116 & n12368 ) ;
  assign n12363 = n7253 &  n11119 ;
  assign n12364 = ~n7518 & n11116 ;
  assign n12365 = n12363 | n12364 ;
  assign n12366 = ~n7783 & n11113 ;
  assign n12367 = ( n7783 & ~n12365 ) | ( n7783 & n12366 ) | ( ~n12365 & n12366 ) ;
  assign n12370 = ( n12367 & ~n7255 ) | ( n12367 & n12369 ) | ( ~n7255 & n12369 ) ;
  assign n12371 = ~n12369 & n12370 ;
  assign n12373 = ( x11 & n12367 ) | ( x11 & n12371 ) | ( n12367 & n12371 ) ;
  assign n12372 = ( x11 & ~n12371 ) | ( x11 & n12367 ) | ( ~n12371 & n12367 ) ;
  assign n12374 = ( n12371 & ~n12373 ) | ( n12371 & n12372 ) | ( ~n12373 & n12372 ) ;
  assign n12381 = n11116 | n7783 ;
  assign n12378 = ( n7253 & ~n11122 ) | ( n7253 & 1'b0 ) | ( ~n11122 & 1'b0 ) ;
  assign n12379 = ~n7518 & n11119 ;
  assign n12380 = n12378 | n12379 ;
  assign n12382 = ( n12381 & ~n7783 ) | ( n12381 & n12380 ) | ( ~n7783 & n12380 ) ;
  assign n12383 = ( n7255 & ~n11230 ) | ( n7255 & n12382 ) | ( ~n11230 & n12382 ) ;
  assign n12384 = n11230 | n12383 ;
  assign n12386 = ( x11 & n12382 ) | ( x11 & n12384 ) | ( n12382 & n12384 ) ;
  assign n12385 = ( x11 & ~n12384 ) | ( x11 & n12382 ) | ( ~n12384 & n12382 ) ;
  assign n12387 = ( n12384 & ~n12386 ) | ( n12384 & n12385 ) | ( ~n12386 & n12385 ) ;
  assign n12375 = ( n12117 & ~n12327 ) | ( n12117 & n12119 ) | ( ~n12327 & n12119 ) ;
  assign n12376 = ( n12119 & ~n12117 ) | ( n12119 & n12327 ) | ( ~n12117 & n12327 ) ;
  assign n12377 = ( n12375 & ~n12119 ) | ( n12375 & n12376 ) | ( ~n12119 & n12376 ) ;
  assign n12391 = n7783 | n11119 ;
  assign n12388 = n7253 &  n11125 ;
  assign n12389 = n7518 | n11122 ;
  assign n12390 = ~n12388 & n12389 ;
  assign n12392 = ( n7783 & ~n12391 ) | ( n7783 & n12390 ) | ( ~n12391 & n12390 ) ;
  assign n12393 = ~n7255 & n12088 ;
  assign n12394 = ( n12392 & ~n12393 ) | ( n12392 & 1'b0 ) | ( ~n12393 & 1'b0 ) ;
  assign n12395 = x11 &  n12394 ;
  assign n12396 = x11 | n12394 ;
  assign n12397 = ~n12395 & n12396 ;
  assign n12398 = ( n12122 & ~n12326 ) | ( n12122 & n12132 ) | ( ~n12326 & n12132 ) ;
  assign n12399 = ( n12327 & ~n12132 ) | ( n12327 & n12398 ) | ( ~n12132 & n12398 ) ;
  assign n12400 = ( n7253 & ~n11128 ) | ( n7253 & 1'b0 ) | ( ~n11128 & 1'b0 ) ;
  assign n12401 = ~n7518 & n11125 ;
  assign n12402 = n12400 | n12401 ;
  assign n12403 = ~n7783 & n11122 ;
  assign n12404 = ( n7783 & ~n12402 ) | ( n7783 & n12403 ) | ( ~n12402 & n12403 ) ;
  assign n12405 = ~n7255 & n12100 ;
  assign n12406 = ( n12404 & ~n12405 ) | ( n12404 & 1'b0 ) | ( ~n12405 & 1'b0 ) ;
  assign n12407 = x11 &  n12406 ;
  assign n12408 = x11 | n12406 ;
  assign n12409 = ~n12407 & n12408 ;
  assign n12410 = ( n12135 & ~n12145 ) | ( n12135 & n12325 ) | ( ~n12145 & n12325 ) ;
  assign n12411 = ( n12145 & ~n12326 ) | ( n12145 & n12410 ) | ( ~n12326 & n12410 ) ;
  assign n12415 = n7783 | n11125 ;
  assign n12412 = ( n7253 & ~n11131 ) | ( n7253 & 1'b0 ) | ( ~n11131 & 1'b0 ) ;
  assign n12413 = n7518 | n11128 ;
  assign n12414 = ~n12412 & n12413 ;
  assign n12416 = ( n7783 & ~n12415 ) | ( n7783 & n12414 ) | ( ~n12415 & n12414 ) ;
  assign n12417 = ~n7255 & n11859 ;
  assign n12418 = ( n12416 & ~n12417 ) | ( n12416 & 1'b0 ) | ( ~n12417 & 1'b0 ) ;
  assign n12419 = x11 &  n12418 ;
  assign n12420 = x11 | n12418 ;
  assign n12421 = ~n12419 & n12420 ;
  assign n12422 = ( n12148 & ~n12324 ) | ( n12148 & n12158 ) | ( ~n12324 & n12158 ) ;
  assign n12423 = ( n12325 & ~n12158 ) | ( n12325 & n12422 ) | ( ~n12158 & n12422 ) ;
  assign n12430 = ~n7783 & n11128 ;
  assign n12427 = n7253 &  n11134 ;
  assign n12428 = n7518 | n11131 ;
  assign n12429 = ~n12427 & n12428 ;
  assign n12431 = ( n7783 & n12430 ) | ( n7783 & n12429 ) | ( n12430 & n12429 ) ;
  assign n12432 = ( n11871 & ~n7255 ) | ( n11871 & n12431 ) | ( ~n7255 & n12431 ) ;
  assign n12433 = ~n11871 & n12432 ;
  assign n12434 = ( x11 & ~n12431 ) | ( x11 & n12433 ) | ( ~n12431 & n12433 ) ;
  assign n12435 = ( n12431 & ~x11 ) | ( n12431 & n12433 ) | ( ~x11 & n12433 ) ;
  assign n12436 = ( n12434 & ~n12433 ) | ( n12434 & n12435 ) | ( ~n12433 & n12435 ) ;
  assign n12424 = ( n12170 & ~n12168 ) | ( n12170 & n12323 ) | ( ~n12168 & n12323 ) ;
  assign n12425 = ( n12168 & ~n12323 ) | ( n12168 & n12170 ) | ( ~n12323 & n12170 ) ;
  assign n12426 = ( n12424 & ~n12170 ) | ( n12424 & n12425 ) | ( ~n12170 & n12425 ) ;
  assign n12437 = ( n12182 & ~n12180 ) | ( n12182 & n12322 ) | ( ~n12180 & n12322 ) ;
  assign n12438 = ( n12180 & ~n12322 ) | ( n12180 & n12182 ) | ( ~n12322 & n12182 ) ;
  assign n12439 = ( n12437 & ~n12182 ) | ( n12437 & n12438 ) | ( ~n12182 & n12438 ) ;
  assign n12440 = ( n7253 & ~n11137 ) | ( n7253 & 1'b0 ) | ( ~n11137 & 1'b0 ) ;
  assign n12441 = ~n7518 & n11134 ;
  assign n12442 = n12440 | n12441 ;
  assign n12443 = ~n7783 & n11131 ;
  assign n12444 = ( n7783 & ~n12442 ) | ( n7783 & n12443 ) | ( ~n12442 & n12443 ) ;
  assign n12445 = ( n7255 & ~n12444 ) | ( n7255 & n11888 ) | ( ~n12444 & n11888 ) ;
  assign n12446 = ( n11888 & ~n12445 ) | ( n11888 & 1'b0 ) | ( ~n12445 & 1'b0 ) ;
  assign n12448 = ( x11 & n12444 ) | ( x11 & n12446 ) | ( n12444 & n12446 ) ;
  assign n12447 = ( x11 & ~n12446 ) | ( x11 & n12444 ) | ( ~n12446 & n12444 ) ;
  assign n12449 = ( n12446 & ~n12448 ) | ( n12446 & n12447 ) | ( ~n12448 & n12447 ) ;
  assign n12456 = n11134 | n7783 ;
  assign n12453 = ( n7253 & ~n11140 ) | ( n7253 & 1'b0 ) | ( ~n11140 & 1'b0 ) ;
  assign n12454 = n7518 | n11137 ;
  assign n12455 = ~n12453 & n12454 ;
  assign n12457 = ( n7783 & ~n12456 ) | ( n7783 & n12455 ) | ( ~n12456 & n12455 ) ;
  assign n12458 = ( n7255 & ~n12457 ) | ( n7255 & n11242 ) | ( ~n12457 & n11242 ) ;
  assign n12459 = ( n11242 & ~n12458 ) | ( n11242 & 1'b0 ) | ( ~n12458 & 1'b0 ) ;
  assign n12461 = ( x11 & n12457 ) | ( x11 & n12459 ) | ( n12457 & n12459 ) ;
  assign n12460 = ( x11 & ~n12459 ) | ( x11 & n12457 ) | ( ~n12459 & n12457 ) ;
  assign n12462 = ( n12459 & ~n12461 ) | ( n12459 & n12460 ) | ( ~n12461 & n12460 ) ;
  assign n12450 = ( n12192 & ~n12321 ) | ( n12192 & n12194 ) | ( ~n12321 & n12194 ) ;
  assign n12451 = ( n12194 & ~n12192 ) | ( n12194 & n12321 ) | ( ~n12192 & n12321 ) ;
  assign n12452 = ( n12450 & ~n12194 ) | ( n12450 & n12451 ) | ( ~n12194 & n12451 ) ;
  assign n12466 = ~n7783 & n11137 ;
  assign n12463 = ( n7253 & ~n11143 ) | ( n7253 & 1'b0 ) | ( ~n11143 & 1'b0 ) ;
  assign n12464 = n7518 | n11140 ;
  assign n12465 = ~n12463 & n12464 ;
  assign n12467 = ( n7783 & n12466 ) | ( n7783 & n12465 ) | ( n12466 & n12465 ) ;
  assign n12468 = n7255 | n11687 ;
  assign n12469 = n12467 &  n12468 ;
  assign n12470 = x11 &  n12469 ;
  assign n12471 = x11 | n12469 ;
  assign n12472 = ~n12470 & n12471 ;
  assign n12473 = ( n12197 & ~n12320 ) | ( n12197 & n12207 ) | ( ~n12320 & n12207 ) ;
  assign n12474 = ( n12321 & ~n12207 ) | ( n12321 & n12473 ) | ( ~n12207 & n12473 ) ;
  assign n12478 = ~n7783 & n11140 ;
  assign n12475 = ( n7253 & ~n11146 ) | ( n7253 & 1'b0 ) | ( ~n11146 & 1'b0 ) ;
  assign n12476 = n7518 | n11143 ;
  assign n12477 = ~n12475 & n12476 ;
  assign n12479 = ( n7783 & n12478 ) | ( n7783 & n12477 ) | ( n12478 & n12477 ) ;
  assign n12480 = n7255 | n11699 ;
  assign n12481 = n12479 &  n12480 ;
  assign n12482 = x11 &  n12481 ;
  assign n12483 = x11 | n12481 ;
  assign n12484 = ~n12482 & n12483 ;
  assign n12485 = ( n12210 & ~n12220 ) | ( n12210 & n12319 ) | ( ~n12220 & n12319 ) ;
  assign n12486 = ( n12220 & ~n12320 ) | ( n12220 & n12485 ) | ( ~n12320 & n12485 ) ;
  assign n12490 = ~n7783 & n11143 ;
  assign n12487 = ( n7253 & ~n11149 ) | ( n7253 & 1'b0 ) | ( ~n11149 & 1'b0 ) ;
  assign n12488 = n7518 | n11146 ;
  assign n12489 = ~n12487 & n12488 ;
  assign n12491 = ( n7783 & n12490 ) | ( n7783 & n12489 ) | ( n12490 & n12489 ) ;
  assign n12492 = n7255 | n11542 ;
  assign n12493 = n12491 &  n12492 ;
  assign n12494 = x11 &  n12493 ;
  assign n12495 = x11 | n12493 ;
  assign n12496 = ~n12494 & n12495 ;
  assign n12497 = ( n12223 & n12233 ) | ( n12223 & n12318 ) | ( n12233 & n12318 ) ;
  assign n12498 = ( n12233 & ~n12497 ) | ( n12233 & n12319 ) | ( ~n12497 & n12319 ) ;
  assign n12505 = ~n7783 & n11146 ;
  assign n12502 = n7253 &  n11152 ;
  assign n12503 = n7518 | n11149 ;
  assign n12504 = ~n12502 & n12503 ;
  assign n12506 = ( n7783 & n12505 ) | ( n7783 & n12504 ) | ( n12505 & n12504 ) ;
  assign n12507 = ( n7255 & ~n12506 ) | ( n7255 & n11554 ) | ( ~n12506 & n11554 ) ;
  assign n12508 = ( n11554 & ~n12507 ) | ( n11554 & 1'b0 ) | ( ~n12507 & 1'b0 ) ;
  assign n12509 = ( x11 & ~n12506 ) | ( x11 & n12508 ) | ( ~n12506 & n12508 ) ;
  assign n12510 = ( n12506 & ~x11 ) | ( n12506 & n12508 ) | ( ~x11 & n12508 ) ;
  assign n12511 = ( n12509 & ~n12508 ) | ( n12509 & n12510 ) | ( ~n12508 & n12510 ) ;
  assign n12499 = ( n12245 & ~n12243 ) | ( n12245 & n12317 ) | ( ~n12243 & n12317 ) ;
  assign n12500 = ( n12243 & ~n12317 ) | ( n12243 & n12245 ) | ( ~n12317 & n12245 ) ;
  assign n12501 = ( n12499 & ~n12245 ) | ( n12499 & n12500 ) | ( ~n12245 & n12500 ) ;
  assign n12512 = ( n12258 & ~n12248 ) | ( n12258 & n12316 ) | ( ~n12248 & n12316 ) ;
  assign n12513 = ( n12248 & ~n12316 ) | ( n12248 & n12258 ) | ( ~n12316 & n12258 ) ;
  assign n12514 = ( n12512 & ~n12258 ) | ( n12512 & n12513 ) | ( ~n12258 & n12513 ) ;
  assign n12515 = n7253 &  n11155 ;
  assign n12516 = ~n7518 & n11152 ;
  assign n12517 = n12515 | n12516 ;
  assign n12518 = ~n7783 & n11149 ;
  assign n12519 = ( n7783 & ~n12517 ) | ( n7783 & n12518 ) | ( ~n12517 & n12518 ) ;
  assign n12520 = ( n11572 & ~n7255 ) | ( n11572 & n12519 ) | ( ~n7255 & n12519 ) ;
  assign n12521 = ~n11572 & n12520 ;
  assign n12523 = ( x11 & n12519 ) | ( x11 & n12521 ) | ( n12519 & n12521 ) ;
  assign n12522 = ( x11 & ~n12521 ) | ( x11 & n12519 ) | ( ~n12521 & n12519 ) ;
  assign n12524 = ( n12521 & ~n12523 ) | ( n12521 & n12522 ) | ( ~n12523 & n12522 ) ;
  assign n12525 = ( n12268 & ~n12315 ) | ( n12268 & n12273 ) | ( ~n12315 & n12273 ) ;
  assign n12526 = ( n12273 & ~n12268 ) | ( n12273 & n12315 ) | ( ~n12268 & n12315 ) ;
  assign n12527 = ( n12525 & ~n12273 ) | ( n12525 & n12526 ) | ( ~n12273 & n12526 ) ;
  assign n12531 = n11152 | n7783 ;
  assign n12528 = n7253 &  n11158 ;
  assign n12529 = ~n7518 & n11155 ;
  assign n12530 = n12528 | n12529 ;
  assign n12532 = ( n12531 & ~n7783 ) | ( n12531 & n12530 ) | ( ~n7783 & n12530 ) ;
  assign n12533 = ( n7255 & n11254 ) | ( n7255 & n12532 ) | ( n11254 & n12532 ) ;
  assign n12534 = ( n11254 & ~n12533 ) | ( n11254 & 1'b0 ) | ( ~n12533 & 1'b0 ) ;
  assign n12535 = ( n12532 & ~x11 ) | ( n12532 & n12534 ) | ( ~x11 & n12534 ) ;
  assign n12536 = ( x11 & ~n12532 ) | ( x11 & n12534 ) | ( ~n12532 & n12534 ) ;
  assign n12537 = ( n12535 & ~n12534 ) | ( n12535 & n12536 ) | ( ~n12534 & n12536 ) ;
  assign n12541 = n11155 | n7783 ;
  assign n12538 = ( n7253 & ~n11161 ) | ( n7253 & 1'b0 ) | ( ~n11161 & 1'b0 ) ;
  assign n12539 = ~n7518 & n11158 ;
  assign n12540 = n12538 | n12539 ;
  assign n12542 = ( n12541 & ~n7783 ) | ( n12541 & n12540 ) | ( ~n7783 & n12540 ) ;
  assign n12543 = n7255 | n11451 ;
  assign n12544 = ~n12542 & n12543 ;
  assign n12545 = x11 &  n12544 ;
  assign n12546 = x11 | n12544 ;
  assign n12547 = ~n12545 & n12546 ;
  assign n12548 = ( n12287 & ~n12277 ) | ( n12287 & n12314 ) | ( ~n12277 & n12314 ) ;
  assign n12549 = ( n12315 & ~n12287 ) | ( n12315 & n12548 ) | ( ~n12287 & n12548 ) ;
  assign n12551 = ( n12036 & n12303 ) | ( n12036 & n12313 ) | ( n12303 & n12313 ) ;
  assign n12550 = ( n12036 & ~n12303 ) | ( n12036 & n12313 ) | ( ~n12303 & n12313 ) ;
  assign n12552 = ( n12303 & ~n12551 ) | ( n12303 & n12550 ) | ( ~n12551 & n12550 ) ;
  assign n12556 = n11158 | n7783 ;
  assign n12553 = ( n7253 & ~n11164 ) | ( n7253 & 1'b0 ) | ( ~n11164 & 1'b0 ) ;
  assign n12554 = n7518 | n11161 ;
  assign n12555 = ~n12553 & n12554 ;
  assign n12557 = ( n7783 & ~n12556 ) | ( n7783 & n12555 ) | ( ~n12556 & n12555 ) ;
  assign n12558 = ( n7255 & ~n12557 ) | ( n7255 & n11463 ) | ( ~n12557 & n11463 ) ;
  assign n12559 = ( n11463 & ~n12558 ) | ( n11463 & 1'b0 ) | ( ~n12558 & 1'b0 ) ;
  assign n12561 = ( x11 & n12557 ) | ( x11 & n12559 ) | ( n12557 & n12559 ) ;
  assign n12560 = ( x11 & ~n12559 ) | ( x11 & n12557 ) | ( ~n12559 & n12557 ) ;
  assign n12562 = ( n12559 & ~n12561 ) | ( n12559 & n12560 ) | ( ~n12561 & n12560 ) ;
  assign n12563 = ( n7253 & ~n11166 ) | ( n7253 & 1'b0 ) | ( ~n11166 & 1'b0 ) ;
  assign n12564 = n7518 | n11164 ;
  assign n12565 = ~n12563 & n12564 ;
  assign n12566 = ~n7783 & n11161 ;
  assign n12567 = ( n7783 & n12565 ) | ( n7783 & n12566 ) | ( n12565 & n12566 ) ;
  assign n12568 = n7255 | n11385 ;
  assign n12569 = n12567 &  n12568 ;
  assign n12570 = x11 &  n12569 ;
  assign n12571 = x11 | n12569 ;
  assign n12572 = ~n12570 & n12571 ;
  assign n12573 = ( x14 & n12288 ) | ( x14 & n12293 ) | ( n12288 & n12293 ) ;
  assign n12574 = ~n12288 & n12573 ;
  assign n12575 = ( n12300 & ~x14 ) | ( n12300 & n12574 ) | ( ~x14 & n12574 ) ;
  assign n12576 = ( x14 & ~n12300 ) | ( x14 & n12574 ) | ( ~n12300 & n12574 ) ;
  assign n12577 = ( n12575 & ~n12574 ) | ( n12575 & n12576 ) | ( ~n12574 & n12576 ) ;
  assign n12578 = x14 &  n12288 ;
  assign n12579 = n12293 &  n12578 ;
  assign n12580 = n12293 | n12578 ;
  assign n12581 = ~n12579 & n12580 ;
  assign n12611 = ~n7783 & n11166 ;
  assign n12608 = ( n7253 & ~n11172 ) | ( n7253 & 1'b0 ) | ( ~n11172 & 1'b0 ) ;
  assign n12609 = n7518 | n11168 ;
  assign n12610 = ~n12608 & n12609 ;
  assign n12612 = ( n7783 & n12611 ) | ( n7783 & n12610 ) | ( n12611 & n12610 ) ;
  assign n12613 = n7255 | n11431 ;
  assign n12614 = n12612 &  n12613 ;
  assign n12615 = x11 &  n12614 ;
  assign n12616 = x11 | n12614 ;
  assign n12617 = ~n12615 & n12616 ;
  assign n12592 = n7251 &  n11170 ;
  assign n12596 = ~n7255 & n11369 ;
  assign n12593 = ~n7518 & n11170 ;
  assign n12594 = n7783 | n11172 ;
  assign n12595 = ~n12593 & n12594 ;
  assign n12597 = ( n7255 & n12596 ) | ( n7255 & n12595 ) | ( n12596 & n12595 ) ;
  assign n12603 = n11323 | n7255 ;
  assign n12601 = ~n7783 & n11168 ;
  assign n12598 = n7253 &  n11170 ;
  assign n12599 = n7518 | n11172 ;
  assign n12600 = ~n12598 & n12599 ;
  assign n12602 = ( n7783 & n12601 ) | ( n7783 & n12600 ) | ( n12601 & n12600 ) ;
  assign n12604 = ( n7255 & ~n12603 ) | ( n7255 & n12602 ) | ( ~n12603 & n12602 ) ;
  assign n12605 = ( n12592 & n12597 ) | ( n12592 & n12604 ) | ( n12597 & n12604 ) ;
  assign n12606 = ( x11 & ~n12605 ) | ( x11 & n12592 ) | ( ~n12605 & n12592 ) ;
  assign n12607 = ( x11 & ~n12606 ) | ( x11 & 1'b0 ) | ( ~n12606 & 1'b0 ) ;
  assign n12618 = ( n12288 & ~n12617 ) | ( n12288 & n12607 ) | ( ~n12617 & n12607 ) ;
  assign n12585 = ~n7783 & n11164 ;
  assign n12582 = ( n7253 & ~n11168 ) | ( n7253 & 1'b0 ) | ( ~n11168 & 1'b0 ) ;
  assign n12583 = n7518 | n11166 ;
  assign n12584 = ~n12582 & n12583 ;
  assign n12586 = ( n7783 & n12585 ) | ( n7783 & n12584 ) | ( n12585 & n12584 ) ;
  assign n12587 = ( n11397 & ~n7255 ) | ( n11397 & n12586 ) | ( ~n7255 & n12586 ) ;
  assign n12588 = ~n11397 & n12587 ;
  assign n12589 = ( x11 & ~n12586 ) | ( x11 & n12588 ) | ( ~n12586 & n12588 ) ;
  assign n12590 = ( n12586 & ~x11 ) | ( n12586 & n12588 ) | ( ~x11 & n12588 ) ;
  assign n12591 = ( n12589 & ~n12588 ) | ( n12589 & n12590 ) | ( ~n12588 & n12590 ) ;
  assign n12619 = ( n12581 & ~n12618 ) | ( n12581 & n12591 ) | ( ~n12618 & n12591 ) ;
  assign n12620 = ( n12572 & n12577 ) | ( n12572 & n12619 ) | ( n12577 & n12619 ) ;
  assign n12621 = ( n12552 & n12562 ) | ( n12552 & n12620 ) | ( n12562 & n12620 ) ;
  assign n12622 = ( n12547 & ~n12549 ) | ( n12547 & n12621 ) | ( ~n12549 & n12621 ) ;
  assign n12623 = ( n12527 & ~n12537 ) | ( n12527 & n12622 ) | ( ~n12537 & n12622 ) ;
  assign n12624 = ( n12514 & n12524 ) | ( n12514 & n12623 ) | ( n12524 & n12623 ) ;
  assign n12625 = ( n12511 & ~n12501 ) | ( n12511 & n12624 ) | ( ~n12501 & n12624 ) ;
  assign n12626 = ( n12496 & ~n12498 ) | ( n12496 & n12625 ) | ( ~n12498 & n12625 ) ;
  assign n12627 = ( n12484 & n12486 ) | ( n12484 & n12626 ) | ( n12486 & n12626 ) ;
  assign n12628 = ( n12472 & ~n12474 ) | ( n12472 & n12627 ) | ( ~n12474 & n12627 ) ;
  assign n12629 = ( n12462 & ~n12452 ) | ( n12462 & n12628 ) | ( ~n12452 & n12628 ) ;
  assign n12630 = ( n12439 & n12449 ) | ( n12439 & n12629 ) | ( n12449 & n12629 ) ;
  assign n12631 = ( n12436 & ~n12426 ) | ( n12436 & n12630 ) | ( ~n12426 & n12630 ) ;
  assign n12632 = ( n12421 & ~n12423 ) | ( n12421 & n12631 ) | ( ~n12423 & n12631 ) ;
  assign n12633 = ( n12409 & n12411 ) | ( n12409 & n12632 ) | ( n12411 & n12632 ) ;
  assign n12634 = ( n12397 & ~n12399 ) | ( n12397 & n12633 ) | ( ~n12399 & n12633 ) ;
  assign n12635 = ( n12387 & ~n12377 ) | ( n12387 & n12634 ) | ( ~n12377 & n12634 ) ;
  assign n12636 = ( n12362 & n12374 ) | ( n12362 & n12635 ) | ( n12374 & n12635 ) ;
  assign n12637 = ( n12357 & n12359 ) | ( n12357 & n12636 ) | ( n12359 & n12636 ) ;
  assign n12638 = ( n12333 & ~n12345 ) | ( n12333 & n12637 ) | ( ~n12345 & n12637 ) ;
  assign n12639 = ( n12333 & ~n12637 ) | ( n12333 & n12345 ) | ( ~n12637 & n12345 ) ;
  assign n12640 = ( n12638 & ~n12333 ) | ( n12638 & n12639 ) | ( ~n12333 & n12639 ) ;
  assign n12641 = ( n12359 & ~n12357 ) | ( n12359 & n12636 ) | ( ~n12357 & n12636 ) ;
  assign n12642 = ( n12357 & ~n12636 ) | ( n12357 & n12359 ) | ( ~n12636 & n12359 ) ;
  assign n12643 = ( n12641 & ~n12359 ) | ( n12641 & n12642 ) | ( ~n12359 & n12642 ) ;
  assign n12649 = ( n11101 & ~n11104 ) | ( n11101 & n11196 ) | ( ~n11104 & n11196 ) ;
  assign n12650 = ( n11104 & ~n11197 ) | ( n11104 & n12649 ) | ( ~n11197 & n12649 ) ;
  assign n12647 = ~n8764 & n11101 ;
  assign n12644 = n8105 &  n11107 ;
  assign n12645 = n8429 | n11104 ;
  assign n12646 = ~n12644 & n12645 ;
  assign n12648 = ( n8764 & n12647 ) | ( n8764 & n12646 ) | ( n12647 & n12646 ) ;
  assign n12651 = ( n12648 & ~n8107 ) | ( n12648 & n12650 ) | ( ~n8107 & n12650 ) ;
  assign n12652 = ~n12650 & n12651 ;
  assign n12654 = ( x8 & n12648 ) | ( x8 & n12652 ) | ( n12648 & n12652 ) ;
  assign n12653 = ( x8 & ~n12652 ) | ( x8 & n12648 ) | ( ~n12652 & n12648 ) ;
  assign n12655 = ( n12652 & ~n12654 ) | ( n12652 & n12653 ) | ( ~n12654 & n12653 ) ;
  assign n12656 = ( n8105 & ~n11110 ) | ( n8105 & 1'b0 ) | ( ~n11110 & 1'b0 ) ;
  assign n12657 = ~n8429 & n11107 ;
  assign n12658 = n12656 | n12657 ;
  assign n12659 = ~n8764 & n11104 ;
  assign n12660 = ( n8764 & ~n12658 ) | ( n8764 & n12659 ) | ( ~n12658 & n12659 ) ;
  assign n12661 = ( n11104 & n11107 ) | ( n11104 & n11195 ) | ( n11107 & n11195 ) ;
  assign n12662 = ( n11107 & ~n12661 ) | ( n11107 & n11196 ) | ( ~n12661 & n11196 ) ;
  assign n12663 = ~n8107 & n12662 ;
  assign n12664 = ( n12660 & ~n12663 ) | ( n12660 & 1'b0 ) | ( ~n12663 & 1'b0 ) ;
  assign n12665 = x8 &  n12664 ;
  assign n12666 = x8 | n12664 ;
  assign n12667 = ~n12665 & n12666 ;
  assign n12668 = ( n12362 & ~n12374 ) | ( n12362 & n12635 ) | ( ~n12374 & n12635 ) ;
  assign n12669 = ( n12374 & ~n12636 ) | ( n12374 & n12668 ) | ( ~n12636 & n12668 ) ;
  assign n12673 = n11107 | n8764 ;
  assign n12670 = ( n8105 & ~n11113 ) | ( n8105 & 1'b0 ) | ( ~n11113 & 1'b0 ) ;
  assign n12671 = n8429 | n11110 ;
  assign n12672 = ~n12670 & n12671 ;
  assign n12674 = ( n8764 & ~n12673 ) | ( n8764 & n12672 ) | ( ~n12673 & n12672 ) ;
  assign n12675 = ~n8107 & n12340 ;
  assign n12676 = ( n12674 & ~n12675 ) | ( n12674 & 1'b0 ) | ( ~n12675 & 1'b0 ) ;
  assign n12677 = x8 &  n12676 ;
  assign n12678 = x8 | n12676 ;
  assign n12679 = ~n12677 & n12678 ;
  assign n12680 = ( n12377 & ~n12634 ) | ( n12377 & n12387 ) | ( ~n12634 & n12387 ) ;
  assign n12681 = ( n12635 & ~n12387 ) | ( n12635 & n12680 ) | ( ~n12387 & n12680 ) ;
  assign n12688 = ~n8764 & n11110 ;
  assign n12685 = n8105 &  n11116 ;
  assign n12686 = n8429 | n11113 ;
  assign n12687 = ~n12685 & n12686 ;
  assign n12689 = ( n8764 & n12688 ) | ( n8764 & n12687 ) | ( n12688 & n12687 ) ;
  assign n12690 = ( n8107 & ~n12689 ) | ( n8107 & n12352 ) | ( ~n12689 & n12352 ) ;
  assign n12691 = ( n12352 & ~n12690 ) | ( n12352 & 1'b0 ) | ( ~n12690 & 1'b0 ) ;
  assign n12693 = ( x8 & n12689 ) | ( x8 & n12691 ) | ( n12689 & n12691 ) ;
  assign n12692 = ( x8 & ~n12691 ) | ( x8 & n12689 ) | ( ~n12691 & n12689 ) ;
  assign n12694 = ( n12691 & ~n12693 ) | ( n12691 & n12692 ) | ( ~n12693 & n12692 ) ;
  assign n12682 = ( n12399 & ~n12397 ) | ( n12399 & n12633 ) | ( ~n12397 & n12633 ) ;
  assign n12683 = ( n12397 & ~n12633 ) | ( n12397 & n12399 ) | ( ~n12633 & n12399 ) ;
  assign n12684 = ( n12682 & ~n12399 ) | ( n12682 & n12683 ) | ( ~n12399 & n12683 ) ;
  assign n12695 = ( n12411 & ~n12409 ) | ( n12411 & n12632 ) | ( ~n12409 & n12632 ) ;
  assign n12696 = ( n12409 & ~n12632 ) | ( n12409 & n12411 ) | ( ~n12632 & n12411 ) ;
  assign n12697 = ( n12695 & ~n12411 ) | ( n12695 & n12696 ) | ( ~n12411 & n12696 ) ;
  assign n12698 = n8105 &  n11119 ;
  assign n12699 = ~n8429 & n11116 ;
  assign n12700 = n12698 | n12699 ;
  assign n12701 = ~n8764 & n11113 ;
  assign n12702 = ( n8764 & ~n12700 ) | ( n8764 & n12701 ) | ( ~n12700 & n12701 ) ;
  assign n12703 = ( n12369 & ~n8107 ) | ( n12369 & n12702 ) | ( ~n8107 & n12702 ) ;
  assign n12704 = ~n12369 & n12703 ;
  assign n12706 = ( x8 & n12702 ) | ( x8 & n12704 ) | ( n12702 & n12704 ) ;
  assign n12705 = ( x8 & ~n12704 ) | ( x8 & n12702 ) | ( ~n12704 & n12702 ) ;
  assign n12707 = ( n12704 & ~n12706 ) | ( n12704 & n12705 ) | ( ~n12706 & n12705 ) ;
  assign n12714 = n11116 | n8764 ;
  assign n12711 = ( n8105 & ~n11122 ) | ( n8105 & 1'b0 ) | ( ~n11122 & 1'b0 ) ;
  assign n12712 = ~n8429 & n11119 ;
  assign n12713 = n12711 | n12712 ;
  assign n12715 = ( n12714 & ~n8764 ) | ( n12714 & n12713 ) | ( ~n8764 & n12713 ) ;
  assign n12716 = ( n8107 & ~n11230 ) | ( n8107 & n12715 ) | ( ~n11230 & n12715 ) ;
  assign n12717 = n11230 | n12716 ;
  assign n12719 = ( x8 & n12715 ) | ( x8 & n12717 ) | ( n12715 & n12717 ) ;
  assign n12718 = ( x8 & ~n12717 ) | ( x8 & n12715 ) | ( ~n12717 & n12715 ) ;
  assign n12720 = ( n12717 & ~n12719 ) | ( n12717 & n12718 ) | ( ~n12719 & n12718 ) ;
  assign n12708 = ( n12421 & ~n12631 ) | ( n12421 & n12423 ) | ( ~n12631 & n12423 ) ;
  assign n12709 = ( n12423 & ~n12421 ) | ( n12423 & n12631 ) | ( ~n12421 & n12631 ) ;
  assign n12710 = ( n12708 & ~n12423 ) | ( n12708 & n12709 ) | ( ~n12423 & n12709 ) ;
  assign n12724 = n8764 | n11119 ;
  assign n12721 = n8105 &  n11125 ;
  assign n12722 = n8429 | n11122 ;
  assign n12723 = ~n12721 & n12722 ;
  assign n12725 = ( n8764 & ~n12724 ) | ( n8764 & n12723 ) | ( ~n12724 & n12723 ) ;
  assign n12726 = ~n8107 & n12088 ;
  assign n12727 = ( n12725 & ~n12726 ) | ( n12725 & 1'b0 ) | ( ~n12726 & 1'b0 ) ;
  assign n12728 = x8 &  n12727 ;
  assign n12729 = x8 | n12727 ;
  assign n12730 = ~n12728 & n12729 ;
  assign n12731 = ( n12426 & ~n12630 ) | ( n12426 & n12436 ) | ( ~n12630 & n12436 ) ;
  assign n12732 = ( n12631 & ~n12436 ) | ( n12631 & n12731 ) | ( ~n12436 & n12731 ) ;
  assign n12733 = ( n8105 & ~n11128 ) | ( n8105 & 1'b0 ) | ( ~n11128 & 1'b0 ) ;
  assign n12734 = ~n8429 & n11125 ;
  assign n12735 = n12733 | n12734 ;
  assign n12736 = ~n8764 & n11122 ;
  assign n12737 = ( n8764 & ~n12735 ) | ( n8764 & n12736 ) | ( ~n12735 & n12736 ) ;
  assign n12738 = ~n8107 & n12100 ;
  assign n12739 = ( n12737 & ~n12738 ) | ( n12737 & 1'b0 ) | ( ~n12738 & 1'b0 ) ;
  assign n12740 = x8 &  n12739 ;
  assign n12741 = x8 | n12739 ;
  assign n12742 = ~n12740 & n12741 ;
  assign n12743 = ( n12439 & ~n12449 ) | ( n12439 & n12629 ) | ( ~n12449 & n12629 ) ;
  assign n12744 = ( n12449 & ~n12630 ) | ( n12449 & n12743 ) | ( ~n12630 & n12743 ) ;
  assign n12748 = n8764 | n11125 ;
  assign n12745 = ( n8105 & ~n11131 ) | ( n8105 & 1'b0 ) | ( ~n11131 & 1'b0 ) ;
  assign n12746 = n8429 | n11128 ;
  assign n12747 = ~n12745 & n12746 ;
  assign n12749 = ( n8764 & ~n12748 ) | ( n8764 & n12747 ) | ( ~n12748 & n12747 ) ;
  assign n12750 = ~n8107 & n11859 ;
  assign n12751 = ( n12749 & ~n12750 ) | ( n12749 & 1'b0 ) | ( ~n12750 & 1'b0 ) ;
  assign n12752 = x8 &  n12751 ;
  assign n12753 = x8 | n12751 ;
  assign n12754 = ~n12752 & n12753 ;
  assign n12755 = ( n12452 & ~n12628 ) | ( n12452 & n12462 ) | ( ~n12628 & n12462 ) ;
  assign n12756 = ( n12629 & ~n12462 ) | ( n12629 & n12755 ) | ( ~n12462 & n12755 ) ;
  assign n12763 = ~n8764 & n11128 ;
  assign n12760 = n8105 &  n11134 ;
  assign n12761 = n8429 | n11131 ;
  assign n12762 = ~n12760 & n12761 ;
  assign n12764 = ( n8764 & n12763 ) | ( n8764 & n12762 ) | ( n12763 & n12762 ) ;
  assign n12765 = ( n11871 & ~n8107 ) | ( n11871 & n12764 ) | ( ~n8107 & n12764 ) ;
  assign n12766 = ~n11871 & n12765 ;
  assign n12767 = ( x8 & ~n12764 ) | ( x8 & n12766 ) | ( ~n12764 & n12766 ) ;
  assign n12768 = ( n12764 & ~x8 ) | ( n12764 & n12766 ) | ( ~x8 & n12766 ) ;
  assign n12769 = ( n12767 & ~n12766 ) | ( n12767 & n12768 ) | ( ~n12766 & n12768 ) ;
  assign n12757 = ( n12474 & ~n12472 ) | ( n12474 & n12627 ) | ( ~n12472 & n12627 ) ;
  assign n12758 = ( n12472 & ~n12627 ) | ( n12472 & n12474 ) | ( ~n12627 & n12474 ) ;
  assign n12759 = ( n12757 & ~n12474 ) | ( n12757 & n12758 ) | ( ~n12474 & n12758 ) ;
  assign n12770 = ( n12486 & ~n12484 ) | ( n12486 & n12626 ) | ( ~n12484 & n12626 ) ;
  assign n12771 = ( n12484 & ~n12626 ) | ( n12484 & n12486 ) | ( ~n12626 & n12486 ) ;
  assign n12772 = ( n12770 & ~n12486 ) | ( n12770 & n12771 ) | ( ~n12486 & n12771 ) ;
  assign n12773 = ( n8105 & ~n11137 ) | ( n8105 & 1'b0 ) | ( ~n11137 & 1'b0 ) ;
  assign n12774 = ~n8429 & n11134 ;
  assign n12775 = n12773 | n12774 ;
  assign n12776 = ~n8764 & n11131 ;
  assign n12777 = ( n8764 & ~n12775 ) | ( n8764 & n12776 ) | ( ~n12775 & n12776 ) ;
  assign n12778 = ( n8107 & ~n12777 ) | ( n8107 & n11888 ) | ( ~n12777 & n11888 ) ;
  assign n12779 = ( n11888 & ~n12778 ) | ( n11888 & 1'b0 ) | ( ~n12778 & 1'b0 ) ;
  assign n12781 = ( x8 & n12777 ) | ( x8 & n12779 ) | ( n12777 & n12779 ) ;
  assign n12780 = ( x8 & ~n12779 ) | ( x8 & n12777 ) | ( ~n12779 & n12777 ) ;
  assign n12782 = ( n12779 & ~n12781 ) | ( n12779 & n12780 ) | ( ~n12781 & n12780 ) ;
  assign n12789 = n11134 | n8764 ;
  assign n12786 = ( n8105 & ~n11140 ) | ( n8105 & 1'b0 ) | ( ~n11140 & 1'b0 ) ;
  assign n12787 = n8429 | n11137 ;
  assign n12788 = ~n12786 & n12787 ;
  assign n12790 = ( n8764 & ~n12789 ) | ( n8764 & n12788 ) | ( ~n12789 & n12788 ) ;
  assign n12791 = ( n8107 & ~n12790 ) | ( n8107 & n11242 ) | ( ~n12790 & n11242 ) ;
  assign n12792 = ( n11242 & ~n12791 ) | ( n11242 & 1'b0 ) | ( ~n12791 & 1'b0 ) ;
  assign n12794 = ( x8 & n12790 ) | ( x8 & n12792 ) | ( n12790 & n12792 ) ;
  assign n12793 = ( x8 & ~n12792 ) | ( x8 & n12790 ) | ( ~n12792 & n12790 ) ;
  assign n12795 = ( n12792 & ~n12794 ) | ( n12792 & n12793 ) | ( ~n12794 & n12793 ) ;
  assign n12783 = ( n12496 & ~n12625 ) | ( n12496 & n12498 ) | ( ~n12625 & n12498 ) ;
  assign n12784 = ( n12498 & ~n12496 ) | ( n12498 & n12625 ) | ( ~n12496 & n12625 ) ;
  assign n12785 = ( n12783 & ~n12498 ) | ( n12783 & n12784 ) | ( ~n12498 & n12784 ) ;
  assign n12799 = ~n8764 & n11137 ;
  assign n12796 = ( n8105 & ~n11143 ) | ( n8105 & 1'b0 ) | ( ~n11143 & 1'b0 ) ;
  assign n12797 = n8429 | n11140 ;
  assign n12798 = ~n12796 & n12797 ;
  assign n12800 = ( n8764 & n12799 ) | ( n8764 & n12798 ) | ( n12799 & n12798 ) ;
  assign n12801 = n8107 | n11687 ;
  assign n12802 = n12800 &  n12801 ;
  assign n12803 = x8 &  n12802 ;
  assign n12804 = x8 | n12802 ;
  assign n12805 = ~n12803 & n12804 ;
  assign n12806 = ( n12501 & ~n12624 ) | ( n12501 & n12511 ) | ( ~n12624 & n12511 ) ;
  assign n12807 = ( n12625 & ~n12511 ) | ( n12625 & n12806 ) | ( ~n12511 & n12806 ) ;
  assign n12811 = ~n8764 & n11140 ;
  assign n12808 = ( n8105 & ~n11146 ) | ( n8105 & 1'b0 ) | ( ~n11146 & 1'b0 ) ;
  assign n12809 = n8429 | n11143 ;
  assign n12810 = ~n12808 & n12809 ;
  assign n12812 = ( n8764 & n12811 ) | ( n8764 & n12810 ) | ( n12811 & n12810 ) ;
  assign n12813 = n8107 | n11699 ;
  assign n12814 = n12812 &  n12813 ;
  assign n12815 = x8 &  n12814 ;
  assign n12816 = x8 | n12814 ;
  assign n12817 = ~n12815 & n12816 ;
  assign n12818 = ( n12514 & ~n12524 ) | ( n12514 & n12623 ) | ( ~n12524 & n12623 ) ;
  assign n12819 = ( n12524 & ~n12624 ) | ( n12524 & n12818 ) | ( ~n12624 & n12818 ) ;
  assign n12823 = ~n8764 & n11143 ;
  assign n12820 = ( n8105 & ~n11149 ) | ( n8105 & 1'b0 ) | ( ~n11149 & 1'b0 ) ;
  assign n12821 = n8429 | n11146 ;
  assign n12822 = ~n12820 & n12821 ;
  assign n12824 = ( n8764 & n12823 ) | ( n8764 & n12822 ) | ( n12823 & n12822 ) ;
  assign n12825 = n8107 | n11542 ;
  assign n12826 = n12824 &  n12825 ;
  assign n12827 = x8 &  n12826 ;
  assign n12828 = x8 | n12826 ;
  assign n12829 = ~n12827 & n12828 ;
  assign n12830 = ( n12527 & n12537 ) | ( n12527 & n12622 ) | ( n12537 & n12622 ) ;
  assign n12831 = ( n12537 & ~n12830 ) | ( n12537 & n12623 ) | ( ~n12830 & n12623 ) ;
  assign n12838 = ~n8764 & n11146 ;
  assign n12835 = n8105 &  n11152 ;
  assign n12836 = n8429 | n11149 ;
  assign n12837 = ~n12835 & n12836 ;
  assign n12839 = ( n8764 & n12838 ) | ( n8764 & n12837 ) | ( n12838 & n12837 ) ;
  assign n12840 = ( n8107 & ~n12839 ) | ( n8107 & n11554 ) | ( ~n12839 & n11554 ) ;
  assign n12841 = ( n11554 & ~n12840 ) | ( n11554 & 1'b0 ) | ( ~n12840 & 1'b0 ) ;
  assign n12842 = ( x8 & ~n12839 ) | ( x8 & n12841 ) | ( ~n12839 & n12841 ) ;
  assign n12843 = ( n12839 & ~x8 ) | ( n12839 & n12841 ) | ( ~x8 & n12841 ) ;
  assign n12844 = ( n12842 & ~n12841 ) | ( n12842 & n12843 ) | ( ~n12841 & n12843 ) ;
  assign n12832 = ( n12549 & ~n12547 ) | ( n12549 & n12621 ) | ( ~n12547 & n12621 ) ;
  assign n12833 = ( n12547 & ~n12621 ) | ( n12547 & n12549 ) | ( ~n12621 & n12549 ) ;
  assign n12834 = ( n12832 & ~n12549 ) | ( n12832 & n12833 ) | ( ~n12549 & n12833 ) ;
  assign n12845 = ( n12562 & ~n12552 ) | ( n12562 & n12620 ) | ( ~n12552 & n12620 ) ;
  assign n12846 = ( n12552 & ~n12620 ) | ( n12552 & n12562 ) | ( ~n12620 & n12562 ) ;
  assign n12847 = ( n12845 & ~n12562 ) | ( n12845 & n12846 ) | ( ~n12562 & n12846 ) ;
  assign n12848 = n8105 &  n11155 ;
  assign n12849 = ~n8429 & n11152 ;
  assign n12850 = n12848 | n12849 ;
  assign n12851 = ~n8764 & n11149 ;
  assign n12852 = ( n8764 & ~n12850 ) | ( n8764 & n12851 ) | ( ~n12850 & n12851 ) ;
  assign n12853 = ( n11572 & ~n8107 ) | ( n11572 & n12852 ) | ( ~n8107 & n12852 ) ;
  assign n12854 = ~n11572 & n12853 ;
  assign n12856 = ( x8 & n12852 ) | ( x8 & n12854 ) | ( n12852 & n12854 ) ;
  assign n12855 = ( x8 & ~n12854 ) | ( x8 & n12852 ) | ( ~n12854 & n12852 ) ;
  assign n12857 = ( n12854 & ~n12856 ) | ( n12854 & n12855 ) | ( ~n12856 & n12855 ) ;
  assign n12858 = ( n12572 & ~n12619 ) | ( n12572 & n12577 ) | ( ~n12619 & n12577 ) ;
  assign n12859 = ( n12577 & ~n12572 ) | ( n12577 & n12619 ) | ( ~n12572 & n12619 ) ;
  assign n12860 = ( n12858 & ~n12577 ) | ( n12858 & n12859 ) | ( ~n12577 & n12859 ) ;
  assign n12864 = n11152 | n8764 ;
  assign n12861 = n8105 &  n11158 ;
  assign n12862 = ~n8429 & n11155 ;
  assign n12863 = n12861 | n12862 ;
  assign n12865 = ( n12864 & ~n8764 ) | ( n12864 & n12863 ) | ( ~n8764 & n12863 ) ;
  assign n12866 = ( n8107 & n11254 ) | ( n8107 & n12865 ) | ( n11254 & n12865 ) ;
  assign n12867 = ( n11254 & ~n12866 ) | ( n11254 & 1'b0 ) | ( ~n12866 & 1'b0 ) ;
  assign n12868 = ( n12865 & ~x8 ) | ( n12865 & n12867 ) | ( ~x8 & n12867 ) ;
  assign n12869 = ( x8 & ~n12865 ) | ( x8 & n12867 ) | ( ~n12865 & n12867 ) ;
  assign n12870 = ( n12868 & ~n12867 ) | ( n12868 & n12869 ) | ( ~n12867 & n12869 ) ;
  assign n12874 = n11155 | n8764 ;
  assign n12871 = ( n8105 & ~n11161 ) | ( n8105 & 1'b0 ) | ( ~n11161 & 1'b0 ) ;
  assign n12872 = ~n8429 & n11158 ;
  assign n12873 = n12871 | n12872 ;
  assign n12875 = ( n12874 & ~n8764 ) | ( n12874 & n12873 ) | ( ~n8764 & n12873 ) ;
  assign n12876 = n8107 | n11451 ;
  assign n12877 = ~n12875 & n12876 ;
  assign n12878 = x8 &  n12877 ;
  assign n12879 = x8 | n12877 ;
  assign n12880 = ~n12878 & n12879 ;
  assign n12881 = ( n12591 & ~n12581 ) | ( n12591 & n12618 ) | ( ~n12581 & n12618 ) ;
  assign n12882 = ( n12619 & ~n12591 ) | ( n12619 & n12881 ) | ( ~n12591 & n12881 ) ;
  assign n12884 = ( n12288 & n12607 ) | ( n12288 & n12617 ) | ( n12607 & n12617 ) ;
  assign n12883 = ( n12288 & ~n12607 ) | ( n12288 & n12617 ) | ( ~n12607 & n12617 ) ;
  assign n12885 = ( n12607 & ~n12884 ) | ( n12607 & n12883 ) | ( ~n12884 & n12883 ) ;
  assign n12889 = n11158 | n8764 ;
  assign n12886 = ( n8105 & ~n11164 ) | ( n8105 & 1'b0 ) | ( ~n11164 & 1'b0 ) ;
  assign n12887 = n8429 | n11161 ;
  assign n12888 = ~n12886 & n12887 ;
  assign n12890 = ( n8764 & ~n12889 ) | ( n8764 & n12888 ) | ( ~n12889 & n12888 ) ;
  assign n12891 = ( n8107 & ~n12890 ) | ( n8107 & n11463 ) | ( ~n12890 & n11463 ) ;
  assign n12892 = ( n11463 & ~n12891 ) | ( n11463 & 1'b0 ) | ( ~n12891 & 1'b0 ) ;
  assign n12894 = ( x8 & n12890 ) | ( x8 & n12892 ) | ( n12890 & n12892 ) ;
  assign n12893 = ( x8 & ~n12892 ) | ( x8 & n12890 ) | ( ~n12892 & n12890 ) ;
  assign n12895 = ( n12892 & ~n12894 ) | ( n12892 & n12893 ) | ( ~n12894 & n12893 ) ;
  assign n12896 = ( n8105 & ~n11166 ) | ( n8105 & 1'b0 ) | ( ~n11166 & 1'b0 ) ;
  assign n12897 = n8429 | n11164 ;
  assign n12898 = ~n12896 & n12897 ;
  assign n12899 = ~n8764 & n11161 ;
  assign n12900 = ( n8764 & n12898 ) | ( n8764 & n12899 ) | ( n12898 & n12899 ) ;
  assign n12901 = n8107 | n11385 ;
  assign n12902 = n12900 &  n12901 ;
  assign n12903 = x8 &  n12902 ;
  assign n12904 = x8 | n12902 ;
  assign n12905 = ~n12903 & n12904 ;
  assign n12906 = ( x11 & n12592 ) | ( x11 & n12597 ) | ( n12592 & n12597 ) ;
  assign n12907 = ~n12592 & n12906 ;
  assign n12908 = ( n12604 & ~x11 ) | ( n12604 & n12907 ) | ( ~x11 & n12907 ) ;
  assign n12909 = ( x11 & ~n12604 ) | ( x11 & n12907 ) | ( ~n12604 & n12907 ) ;
  assign n12910 = ( n12908 & ~n12907 ) | ( n12908 & n12909 ) | ( ~n12907 & n12909 ) ;
  assign n12911 = x11 &  n12592 ;
  assign n12912 = n12597 &  n12911 ;
  assign n12913 = n12597 | n12911 ;
  assign n12914 = ~n12912 & n12913 ;
  assign n12944 = ~n8764 & n11166 ;
  assign n12941 = ( n8105 & ~n11172 ) | ( n8105 & 1'b0 ) | ( ~n11172 & 1'b0 ) ;
  assign n12942 = n8429 | n11168 ;
  assign n12943 = ~n12941 & n12942 ;
  assign n12945 = ( n8764 & n12944 ) | ( n8764 & n12943 ) | ( n12944 & n12943 ) ;
  assign n12946 = n8107 | n11431 ;
  assign n12947 = n12945 &  n12946 ;
  assign n12948 = x8 &  n12947 ;
  assign n12949 = x8 | n12947 ;
  assign n12950 = ~n12948 & n12949 ;
  assign n12925 = n8103 &  n11170 ;
  assign n12929 = ~n8107 & n11369 ;
  assign n12926 = ~n8429 & n11170 ;
  assign n12927 = n8764 | n11172 ;
  assign n12928 = ~n12926 & n12927 ;
  assign n12930 = ( n8107 & n12929 ) | ( n8107 & n12928 ) | ( n12929 & n12928 ) ;
  assign n12936 = n11323 | n8107 ;
  assign n12934 = ~n8764 & n11168 ;
  assign n12931 = n8105 &  n11170 ;
  assign n12932 = n8429 | n11172 ;
  assign n12933 = ~n12931 & n12932 ;
  assign n12935 = ( n8764 & n12934 ) | ( n8764 & n12933 ) | ( n12934 & n12933 ) ;
  assign n12937 = ( n8107 & ~n12936 ) | ( n8107 & n12935 ) | ( ~n12936 & n12935 ) ;
  assign n12938 = ( n12925 & n12930 ) | ( n12925 & n12937 ) | ( n12930 & n12937 ) ;
  assign n12939 = ( x8 & ~n12938 ) | ( x8 & n12925 ) | ( ~n12938 & n12925 ) ;
  assign n12940 = ( x8 & ~n12939 ) | ( x8 & 1'b0 ) | ( ~n12939 & 1'b0 ) ;
  assign n12951 = ( n12592 & ~n12950 ) | ( n12592 & n12940 ) | ( ~n12950 & n12940 ) ;
  assign n12918 = ~n8764 & n11164 ;
  assign n12915 = ( n8105 & ~n11168 ) | ( n8105 & 1'b0 ) | ( ~n11168 & 1'b0 ) ;
  assign n12916 = n8429 | n11166 ;
  assign n12917 = ~n12915 & n12916 ;
  assign n12919 = ( n8764 & n12918 ) | ( n8764 & n12917 ) | ( n12918 & n12917 ) ;
  assign n12920 = ( n11397 & ~n8107 ) | ( n11397 & n12919 ) | ( ~n8107 & n12919 ) ;
  assign n12921 = ~n11397 & n12920 ;
  assign n12922 = ( x8 & ~n12919 ) | ( x8 & n12921 ) | ( ~n12919 & n12921 ) ;
  assign n12923 = ( n12919 & ~x8 ) | ( n12919 & n12921 ) | ( ~x8 & n12921 ) ;
  assign n12924 = ( n12922 & ~n12921 ) | ( n12922 & n12923 ) | ( ~n12921 & n12923 ) ;
  assign n12952 = ( n12914 & ~n12951 ) | ( n12914 & n12924 ) | ( ~n12951 & n12924 ) ;
  assign n12953 = ( n12905 & n12910 ) | ( n12905 & n12952 ) | ( n12910 & n12952 ) ;
  assign n12954 = ( n12885 & n12895 ) | ( n12885 & n12953 ) | ( n12895 & n12953 ) ;
  assign n12955 = ( n12880 & ~n12882 ) | ( n12880 & n12954 ) | ( ~n12882 & n12954 ) ;
  assign n12956 = ( n12860 & ~n12870 ) | ( n12860 & n12955 ) | ( ~n12870 & n12955 ) ;
  assign n12957 = ( n12847 & n12857 ) | ( n12847 & n12956 ) | ( n12857 & n12956 ) ;
  assign n12958 = ( n12844 & ~n12834 ) | ( n12844 & n12957 ) | ( ~n12834 & n12957 ) ;
  assign n12959 = ( n12829 & ~n12831 ) | ( n12829 & n12958 ) | ( ~n12831 & n12958 ) ;
  assign n12960 = ( n12817 & n12819 ) | ( n12817 & n12959 ) | ( n12819 & n12959 ) ;
  assign n12961 = ( n12805 & ~n12807 ) | ( n12805 & n12960 ) | ( ~n12807 & n12960 ) ;
  assign n12962 = ( n12795 & ~n12785 ) | ( n12795 & n12961 ) | ( ~n12785 & n12961 ) ;
  assign n12963 = ( n12772 & n12782 ) | ( n12772 & n12962 ) | ( n12782 & n12962 ) ;
  assign n12964 = ( n12769 & ~n12759 ) | ( n12769 & n12963 ) | ( ~n12759 & n12963 ) ;
  assign n12965 = ( n12754 & ~n12756 ) | ( n12754 & n12964 ) | ( ~n12756 & n12964 ) ;
  assign n12966 = ( n12742 & n12744 ) | ( n12742 & n12965 ) | ( n12744 & n12965 ) ;
  assign n12967 = ( n12730 & ~n12732 ) | ( n12730 & n12966 ) | ( ~n12732 & n12966 ) ;
  assign n12968 = ( n12720 & ~n12710 ) | ( n12720 & n12967 ) | ( ~n12710 & n12967 ) ;
  assign n12969 = ( n12697 & n12707 ) | ( n12697 & n12968 ) | ( n12707 & n12968 ) ;
  assign n12970 = ( n12694 & ~n12684 ) | ( n12694 & n12969 ) | ( ~n12684 & n12969 ) ;
  assign n12971 = ( n12679 & ~n12681 ) | ( n12679 & n12970 ) | ( ~n12681 & n12970 ) ;
  assign n12972 = ( n12667 & n12669 ) | ( n12667 & n12971 ) | ( n12669 & n12971 ) ;
  assign n12973 = ( n12643 & n12655 ) | ( n12643 & n12972 ) | ( n12655 & n12972 ) ;
  assign n12974 = ( n11223 & n12640 ) | ( n11223 & n12973 ) | ( n12640 & n12973 ) ;
  assign n12975 = ( n12640 & ~n11223 ) | ( n12640 & n12973 ) | ( ~n11223 & n12973 ) ;
  assign n12976 = ( n11223 & ~n12974 ) | ( n11223 & n12975 ) | ( ~n12974 & n12975 ) ;
  assign n12980 = ~n9997 & n11091 ;
  assign n12977 = n9160 | n11095 ;
  assign n12978 = n9558 | n11093 ;
  assign n12979 = n12977 &  n12978 ;
  assign n12981 = ( n9997 & n12980 ) | ( n9997 & n12979 ) | ( n12980 & n12979 ) ;
  assign n12982 = ( n11093 & ~n11091 ) | ( n11093 & n11200 ) | ( ~n11091 & n11200 ) ;
  assign n12983 = ( n11091 & ~n11093 ) | ( n11091 & n11200 ) | ( ~n11093 & n11200 ) ;
  assign n12984 = ( n12982 & ~n11200 ) | ( n12982 & n12983 ) | ( ~n11200 & n12983 ) ;
  assign n12985 = n9155 | n12984 ;
  assign n12986 = n12981 &  n12985 ;
  assign n12987 = x5 &  n12986 ;
  assign n12988 = x5 | n12986 ;
  assign n12989 = ~n12987 & n12988 ;
  assign n12993 = ~n9997 & n11093 ;
  assign n12990 = n9160 | n11098 ;
  assign n12991 = n9558 | n11095 ;
  assign n12992 = n12990 &  n12991 ;
  assign n12994 = ( n9997 & n12993 ) | ( n9997 & n12992 ) | ( n12993 & n12992 ) ;
  assign n12995 = ( n11095 & ~n11093 ) | ( n11095 & n11199 ) | ( ~n11093 & n11199 ) ;
  assign n12996 = ( n11093 & ~n11095 ) | ( n11093 & n11199 ) | ( ~n11095 & n11199 ) ;
  assign n12997 = ( n12995 & ~n11199 ) | ( n12995 & n12996 ) | ( ~n11199 & n12996 ) ;
  assign n12998 = n9155 | n12997 ;
  assign n12999 = n12994 &  n12998 ;
  assign n13000 = x5 &  n12999 ;
  assign n13001 = x5 | n12999 ;
  assign n13002 = ~n13000 & n13001 ;
  assign n13003 = ( n12643 & ~n12655 ) | ( n12643 & n12972 ) | ( ~n12655 & n12972 ) ;
  assign n13004 = ( n12655 & ~n12973 ) | ( n12655 & n13003 ) | ( ~n12973 & n13003 ) ;
  assign n13005 = ( n12667 & ~n12971 ) | ( n12667 & n12669 ) | ( ~n12971 & n12669 ) ;
  assign n13006 = ( n12669 & ~n12667 ) | ( n12669 & n12971 ) | ( ~n12667 & n12971 ) ;
  assign n13007 = ( n13005 & ~n12669 ) | ( n13005 & n13006 ) | ( ~n12669 & n13006 ) ;
  assign n13013 = ( n11098 & ~n11095 ) | ( n11098 & n11198 ) | ( ~n11095 & n11198 ) ;
  assign n13014 = ( n11095 & ~n11199 ) | ( n11095 & n13013 ) | ( ~n11199 & n13013 ) ;
  assign n13011 = ~n9997 & n11095 ;
  assign n13008 = n9160 | n11101 ;
  assign n13009 = n9558 | n11098 ;
  assign n13010 = n13008 &  n13009 ;
  assign n13012 = ( n9997 & n13011 ) | ( n9997 & n13010 ) | ( n13011 & n13010 ) ;
  assign n13015 = ( n13012 & ~n9155 ) | ( n13012 & n13014 ) | ( ~n9155 & n13014 ) ;
  assign n13016 = ~n13014 & n13015 ;
  assign n13018 = ( x5 & n13012 ) | ( x5 & n13016 ) | ( n13012 & n13016 ) ;
  assign n13017 = ( x5 & ~n13016 ) | ( x5 & n13012 ) | ( ~n13016 & n13012 ) ;
  assign n13019 = ( n13016 & ~n13018 ) | ( n13016 & n13017 ) | ( ~n13018 & n13017 ) ;
  assign n13026 = ~n9997 & n11098 ;
  assign n13023 = n9160 | n11104 ;
  assign n13024 = n9558 | n11101 ;
  assign n13025 = n13023 &  n13024 ;
  assign n13027 = ( n9997 & n13026 ) | ( n9997 & n13025 ) | ( n13026 & n13025 ) ;
  assign n13028 = ( n11218 & ~n9155 ) | ( n11218 & n13027 ) | ( ~n9155 & n13027 ) ;
  assign n13029 = ~n11218 & n13028 ;
  assign n13031 = ( x5 & n13027 ) | ( x5 & n13029 ) | ( n13027 & n13029 ) ;
  assign n13030 = ( x5 & ~n13029 ) | ( x5 & n13027 ) | ( ~n13029 & n13027 ) ;
  assign n13032 = ( n13029 & ~n13031 ) | ( n13029 & n13030 ) | ( ~n13031 & n13030 ) ;
  assign n13020 = ( n12679 & ~n12970 ) | ( n12679 & n12681 ) | ( ~n12970 & n12681 ) ;
  assign n13021 = ( n12681 & ~n12679 ) | ( n12681 & n12970 ) | ( ~n12679 & n12970 ) ;
  assign n13022 = ( n13020 & ~n12681 ) | ( n13020 & n13021 ) | ( ~n12681 & n13021 ) ;
  assign n13036 = ~n9997 & n11101 ;
  assign n13033 = ~n9160 & n11107 ;
  assign n13034 = n9558 | n11104 ;
  assign n13035 = ~n13033 & n13034 ;
  assign n13037 = ( n9997 & n13036 ) | ( n9997 & n13035 ) | ( n13036 & n13035 ) ;
  assign n13038 = n9155 | n12650 ;
  assign n13039 = n13037 &  n13038 ;
  assign n13040 = x5 &  n13039 ;
  assign n13041 = x5 | n13039 ;
  assign n13042 = ~n13040 & n13041 ;
  assign n13043 = ( n12684 & ~n12969 ) | ( n12684 & n12694 ) | ( ~n12969 & n12694 ) ;
  assign n13044 = ( n12970 & ~n12694 ) | ( n12970 & n13043 ) | ( ~n12694 & n13043 ) ;
  assign n13048 = ~n9997 & n11104 ;
  assign n13045 = n9160 | n11110 ;
  assign n13046 = ~n9558 & n11107 ;
  assign n13047 = ( n13045 & ~n13046 ) | ( n13045 & 1'b0 ) | ( ~n13046 & 1'b0 ) ;
  assign n13049 = ( n9997 & n13048 ) | ( n9997 & n13047 ) | ( n13048 & n13047 ) ;
  assign n13050 = ~n9155 & n12662 ;
  assign n13051 = ( n13049 & ~n13050 ) | ( n13049 & 1'b0 ) | ( ~n13050 & 1'b0 ) ;
  assign n13052 = x5 &  n13051 ;
  assign n13053 = x5 | n13051 ;
  assign n13054 = ~n13052 & n13053 ;
  assign n13055 = ( n12697 & ~n12707 ) | ( n12697 & n12968 ) | ( ~n12707 & n12968 ) ;
  assign n13056 = ( n12707 & ~n12969 ) | ( n12707 & n13055 ) | ( ~n12969 & n13055 ) ;
  assign n13060 = n11107 | n9997 ;
  assign n13057 = n9160 | n11113 ;
  assign n13058 = n9558 | n11110 ;
  assign n13059 = n13057 &  n13058 ;
  assign n13061 = ( n9997 & ~n13060 ) | ( n9997 & n13059 ) | ( ~n13060 & n13059 ) ;
  assign n13062 = ~n9155 & n12340 ;
  assign n13063 = ( n13061 & ~n13062 ) | ( n13061 & 1'b0 ) | ( ~n13062 & 1'b0 ) ;
  assign n13064 = x5 &  n13063 ;
  assign n13065 = x5 | n13063 ;
  assign n13066 = ~n13064 & n13065 ;
  assign n13067 = ( n12710 & ~n12967 ) | ( n12710 & n12720 ) | ( ~n12967 & n12720 ) ;
  assign n13068 = ( n12968 & ~n12720 ) | ( n12968 & n13067 ) | ( ~n12720 & n13067 ) ;
  assign n13075 = ~n9997 & n11110 ;
  assign n13072 = ~n9160 & n11116 ;
  assign n13073 = n9558 | n11113 ;
  assign n13074 = ~n13072 & n13073 ;
  assign n13076 = ( n9997 & n13075 ) | ( n9997 & n13074 ) | ( n13075 & n13074 ) ;
  assign n13077 = ( n9155 & ~n13076 ) | ( n9155 & n12352 ) | ( ~n13076 & n12352 ) ;
  assign n13078 = ( n12352 & ~n13077 ) | ( n12352 & 1'b0 ) | ( ~n13077 & 1'b0 ) ;
  assign n13080 = ( x5 & n13076 ) | ( x5 & n13078 ) | ( n13076 & n13078 ) ;
  assign n13079 = ( x5 & ~n13078 ) | ( x5 & n13076 ) | ( ~n13078 & n13076 ) ;
  assign n13081 = ( n13078 & ~n13080 ) | ( n13078 & n13079 ) | ( ~n13080 & n13079 ) ;
  assign n13069 = ( n12732 & ~n12730 ) | ( n12732 & n12966 ) | ( ~n12730 & n12966 ) ;
  assign n13070 = ( n12730 & ~n12966 ) | ( n12730 & n12732 ) | ( ~n12966 & n12732 ) ;
  assign n13071 = ( n13069 & ~n12732 ) | ( n13069 & n13070 ) | ( ~n12732 & n13070 ) ;
  assign n13082 = ( n12744 & ~n12742 ) | ( n12744 & n12965 ) | ( ~n12742 & n12965 ) ;
  assign n13083 = ( n12742 & ~n12965 ) | ( n12742 & n12744 ) | ( ~n12965 & n12744 ) ;
  assign n13084 = ( n13082 & ~n12744 ) | ( n13082 & n13083 ) | ( ~n12744 & n13083 ) ;
  assign n13086 = ~n9160 & n11119 ;
  assign n13087 = ~n9558 & n11116 ;
  assign n13088 = n13086 | n13087 ;
  assign n13085 = ( n9997 & ~n11113 ) | ( n9997 & 1'b0 ) | ( ~n11113 & 1'b0 ) ;
  assign n13089 = ( n11113 & ~n13088 ) | ( n11113 & n13085 ) | ( ~n13088 & n13085 ) ;
  assign n13090 = ( n12369 & ~n9155 ) | ( n12369 & n13089 ) | ( ~n9155 & n13089 ) ;
  assign n13091 = ~n12369 & n13090 ;
  assign n13093 = ( x5 & n13089 ) | ( x5 & n13091 ) | ( n13089 & n13091 ) ;
  assign n13092 = ( x5 & ~n13091 ) | ( x5 & n13089 ) | ( ~n13091 & n13089 ) ;
  assign n13094 = ( n13091 & ~n13093 ) | ( n13091 & n13092 ) | ( ~n13093 & n13092 ) ;
  assign n13101 = n11116 | n9997 ;
  assign n13098 = n9160 | n11122 ;
  assign n13099 = ~n9558 & n11119 ;
  assign n13100 = ( n13098 & ~n13099 ) | ( n13098 & 1'b0 ) | ( ~n13099 & 1'b0 ) ;
  assign n13102 = ( n9997 & ~n13101 ) | ( n9997 & n13100 ) | ( ~n13101 & n13100 ) ;
  assign n13103 = ( n11230 & ~n9155 ) | ( n11230 & n13102 ) | ( ~n9155 & n13102 ) ;
  assign n13104 = ~n11230 & n13103 ;
  assign n13105 = ( x5 & ~n13102 ) | ( x5 & n13104 ) | ( ~n13102 & n13104 ) ;
  assign n13106 = ( n13102 & ~x5 ) | ( n13102 & n13104 ) | ( ~x5 & n13104 ) ;
  assign n13107 = ( n13105 & ~n13104 ) | ( n13105 & n13106 ) | ( ~n13104 & n13106 ) ;
  assign n13095 = ( n12754 & ~n12964 ) | ( n12754 & n12756 ) | ( ~n12964 & n12756 ) ;
  assign n13096 = ( n12756 & ~n12754 ) | ( n12756 & n12964 ) | ( ~n12754 & n12964 ) ;
  assign n13097 = ( n13095 & ~n12756 ) | ( n13095 & n13096 ) | ( ~n12756 & n13096 ) ;
  assign n13108 = n9997 &  n11119 ;
  assign n13109 = ~n9160 & n11125 ;
  assign n13110 = n9558 | n11122 ;
  assign n13111 = ~n13109 & n13110 ;
  assign n13112 = ( n13108 & ~n11119 ) | ( n13108 & n13111 ) | ( ~n11119 & n13111 ) ;
  assign n13113 = ~n9155 & n12088 ;
  assign n13114 = ( n13112 & ~n13113 ) | ( n13112 & 1'b0 ) | ( ~n13113 & 1'b0 ) ;
  assign n13115 = x5 &  n13114 ;
  assign n13116 = x5 | n13114 ;
  assign n13117 = ~n13115 & n13116 ;
  assign n13118 = ( n12759 & ~n12963 ) | ( n12759 & n12769 ) | ( ~n12963 & n12769 ) ;
  assign n13119 = ( n12964 & ~n12769 ) | ( n12964 & n13118 ) | ( ~n12769 & n13118 ) ;
  assign n13123 = ~n9997 & n11122 ;
  assign n13120 = n9160 | n11128 ;
  assign n13121 = ~n9558 & n11125 ;
  assign n13122 = ( n13120 & ~n13121 ) | ( n13120 & 1'b0 ) | ( ~n13121 & 1'b0 ) ;
  assign n13124 = ( n9997 & n13123 ) | ( n9997 & n13122 ) | ( n13123 & n13122 ) ;
  assign n13125 = ~n9155 & n12100 ;
  assign n13126 = ( n13124 & ~n13125 ) | ( n13124 & 1'b0 ) | ( ~n13125 & 1'b0 ) ;
  assign n13127 = x5 &  n13126 ;
  assign n13128 = x5 | n13126 ;
  assign n13129 = ~n13127 & n13128 ;
  assign n13130 = ( n12772 & ~n12782 ) | ( n12772 & n12962 ) | ( ~n12782 & n12962 ) ;
  assign n13131 = ( n12782 & ~n12963 ) | ( n12782 & n13130 ) | ( ~n12963 & n13130 ) ;
  assign n13132 = n9997 &  n11125 ;
  assign n13133 = n9160 | n11131 ;
  assign n13134 = n9558 | n11128 ;
  assign n13135 = n13133 &  n13134 ;
  assign n13136 = ( n13132 & ~n11125 ) | ( n13132 & n13135 ) | ( ~n11125 & n13135 ) ;
  assign n13137 = ~n9155 & n11859 ;
  assign n13138 = ( n13136 & ~n13137 ) | ( n13136 & 1'b0 ) | ( ~n13137 & 1'b0 ) ;
  assign n13139 = x5 &  n13138 ;
  assign n13140 = x5 | n13138 ;
  assign n13141 = ~n13139 & n13140 ;
  assign n13142 = ( n12785 & ~n12961 ) | ( n12785 & n12795 ) | ( ~n12961 & n12795 ) ;
  assign n13143 = ( n12962 & ~n12795 ) | ( n12962 & n13142 ) | ( ~n12795 & n13142 ) ;
  assign n13150 = ~n9997 & n11128 ;
  assign n13147 = ~n9160 & n11134 ;
  assign n13148 = n9558 | n11131 ;
  assign n13149 = ~n13147 & n13148 ;
  assign n13151 = ( n9997 & n13150 ) | ( n9997 & n13149 ) | ( n13150 & n13149 ) ;
  assign n13152 = ( n11871 & ~n9155 ) | ( n11871 & n13151 ) | ( ~n9155 & n13151 ) ;
  assign n13153 = ~n11871 & n13152 ;
  assign n13154 = ( x5 & ~n13151 ) | ( x5 & n13153 ) | ( ~n13151 & n13153 ) ;
  assign n13155 = ( n13151 & ~x5 ) | ( n13151 & n13153 ) | ( ~x5 & n13153 ) ;
  assign n13156 = ( n13154 & ~n13153 ) | ( n13154 & n13155 ) | ( ~n13153 & n13155 ) ;
  assign n13144 = ( n12807 & ~n12805 ) | ( n12807 & n12960 ) | ( ~n12805 & n12960 ) ;
  assign n13145 = ( n12805 & ~n12960 ) | ( n12805 & n12807 ) | ( ~n12960 & n12807 ) ;
  assign n13146 = ( n13144 & ~n12807 ) | ( n13144 & n13145 ) | ( ~n12807 & n13145 ) ;
  assign n13157 = ( n12819 & ~n12817 ) | ( n12819 & n12959 ) | ( ~n12817 & n12959 ) ;
  assign n13158 = ( n12817 & ~n12959 ) | ( n12817 & n12819 ) | ( ~n12959 & n12819 ) ;
  assign n13159 = ( n13157 & ~n12819 ) | ( n13157 & n13158 ) | ( ~n12819 & n13158 ) ;
  assign n13163 = ~n9997 & n11131 ;
  assign n13160 = n9160 | n11137 ;
  assign n13161 = ~n9558 & n11134 ;
  assign n13162 = ( n13160 & ~n13161 ) | ( n13160 & 1'b0 ) | ( ~n13161 & 1'b0 ) ;
  assign n13164 = ( n9997 & n13163 ) | ( n9997 & n13162 ) | ( n13163 & n13162 ) ;
  assign n13165 = ( n9155 & ~n13164 ) | ( n9155 & n11888 ) | ( ~n13164 & n11888 ) ;
  assign n13166 = ( n11888 & ~n13165 ) | ( n11888 & 1'b0 ) | ( ~n13165 & 1'b0 ) ;
  assign n13168 = ( x5 & n13164 ) | ( x5 & n13166 ) | ( n13164 & n13166 ) ;
  assign n13167 = ( x5 & ~n13166 ) | ( x5 & n13164 ) | ( ~n13166 & n13164 ) ;
  assign n13169 = ( n13166 & ~n13168 ) | ( n13166 & n13167 ) | ( ~n13168 & n13167 ) ;
  assign n13176 = n11134 | n9997 ;
  assign n13173 = n9160 | n11140 ;
  assign n13174 = n9558 | n11137 ;
  assign n13175 = n13173 &  n13174 ;
  assign n13177 = ( n9997 & ~n13176 ) | ( n9997 & n13175 ) | ( ~n13176 & n13175 ) ;
  assign n13178 = ( n9155 & ~n13177 ) | ( n9155 & n11242 ) | ( ~n13177 & n11242 ) ;
  assign n13179 = ( n11242 & ~n13178 ) | ( n11242 & 1'b0 ) | ( ~n13178 & 1'b0 ) ;
  assign n13181 = ( x5 & n13177 ) | ( x5 & n13179 ) | ( n13177 & n13179 ) ;
  assign n13180 = ( x5 & ~n13179 ) | ( x5 & n13177 ) | ( ~n13179 & n13177 ) ;
  assign n13182 = ( n13179 & ~n13181 ) | ( n13179 & n13180 ) | ( ~n13181 & n13180 ) ;
  assign n13170 = ( n12829 & ~n12958 ) | ( n12829 & n12831 ) | ( ~n12958 & n12831 ) ;
  assign n13171 = ( n12831 & ~n12829 ) | ( n12831 & n12958 ) | ( ~n12829 & n12958 ) ;
  assign n13172 = ( n13170 & ~n12831 ) | ( n13170 & n13171 ) | ( ~n12831 & n13171 ) ;
  assign n13186 = ~n9997 & n11137 ;
  assign n13183 = n9160 | n11143 ;
  assign n13184 = n9558 | n11140 ;
  assign n13185 = n13183 &  n13184 ;
  assign n13187 = ( n9997 & n13186 ) | ( n9997 & n13185 ) | ( n13186 & n13185 ) ;
  assign n13188 = n9155 | n11687 ;
  assign n13189 = n13187 &  n13188 ;
  assign n13190 = x5 &  n13189 ;
  assign n13191 = x5 | n13189 ;
  assign n13192 = ~n13190 & n13191 ;
  assign n13193 = ( n12834 & ~n12957 ) | ( n12834 & n12844 ) | ( ~n12957 & n12844 ) ;
  assign n13194 = ( n12958 & ~n12844 ) | ( n12958 & n13193 ) | ( ~n12844 & n13193 ) ;
  assign n13198 = ~n9997 & n11140 ;
  assign n13195 = n9160 | n11146 ;
  assign n13196 = n9558 | n11143 ;
  assign n13197 = n13195 &  n13196 ;
  assign n13199 = ( n9997 & n13198 ) | ( n9997 & n13197 ) | ( n13198 & n13197 ) ;
  assign n13200 = n9155 | n11699 ;
  assign n13201 = n13199 &  n13200 ;
  assign n13202 = x5 &  n13201 ;
  assign n13203 = x5 | n13201 ;
  assign n13204 = ~n13202 & n13203 ;
  assign n13205 = ( n12847 & ~n12857 ) | ( n12847 & n12956 ) | ( ~n12857 & n12956 ) ;
  assign n13206 = ( n12857 & ~n12957 ) | ( n12857 & n13205 ) | ( ~n12957 & n13205 ) ;
  assign n13210 = ~n9997 & n11143 ;
  assign n13207 = n9160 | n11149 ;
  assign n13208 = n9558 | n11146 ;
  assign n13209 = n13207 &  n13208 ;
  assign n13211 = ( n9997 & n13210 ) | ( n9997 & n13209 ) | ( n13210 & n13209 ) ;
  assign n13212 = n9155 | n11542 ;
  assign n13213 = n13211 &  n13212 ;
  assign n13214 = x5 &  n13213 ;
  assign n13215 = x5 | n13213 ;
  assign n13216 = ~n13214 & n13215 ;
  assign n13217 = ( n12860 & n12870 ) | ( n12860 & n12955 ) | ( n12870 & n12955 ) ;
  assign n13218 = ( n12870 & ~n13217 ) | ( n12870 & n12956 ) | ( ~n13217 & n12956 ) ;
  assign n13225 = ~n9997 & n11146 ;
  assign n13222 = ~n9160 & n11152 ;
  assign n13223 = n9558 | n11149 ;
  assign n13224 = ~n13222 & n13223 ;
  assign n13226 = ( n9997 & n13225 ) | ( n9997 & n13224 ) | ( n13225 & n13224 ) ;
  assign n13227 = ( n9155 & ~n13226 ) | ( n9155 & n11554 ) | ( ~n13226 & n11554 ) ;
  assign n13228 = ( n11554 & ~n13227 ) | ( n11554 & 1'b0 ) | ( ~n13227 & 1'b0 ) ;
  assign n13229 = ( x5 & ~n13226 ) | ( x5 & n13228 ) | ( ~n13226 & n13228 ) ;
  assign n13230 = ( n13226 & ~x5 ) | ( n13226 & n13228 ) | ( ~x5 & n13228 ) ;
  assign n13231 = ( n13229 & ~n13228 ) | ( n13229 & n13230 ) | ( ~n13228 & n13230 ) ;
  assign n13219 = ( n12882 & ~n12880 ) | ( n12882 & n12954 ) | ( ~n12880 & n12954 ) ;
  assign n13220 = ( n12880 & ~n12954 ) | ( n12880 & n12882 ) | ( ~n12954 & n12882 ) ;
  assign n13221 = ( n13219 & ~n12882 ) | ( n13219 & n13220 ) | ( ~n12882 & n13220 ) ;
  assign n13232 = ( n12895 & ~n12885 ) | ( n12895 & n12953 ) | ( ~n12885 & n12953 ) ;
  assign n13233 = ( n12885 & ~n12953 ) | ( n12885 & n12895 ) | ( ~n12953 & n12895 ) ;
  assign n13234 = ( n13232 & ~n12895 ) | ( n13232 & n13233 ) | ( ~n12895 & n13233 ) ;
  assign n13235 = ~n9160 & n11155 ;
  assign n13236 = ~n9558 & n11152 ;
  assign n13237 = n13235 | n13236 ;
  assign n13238 = ~n9997 & n11149 ;
  assign n13239 = ( n9997 & ~n13237 ) | ( n9997 & n13238 ) | ( ~n13237 & n13238 ) ;
  assign n13240 = ( n11572 & ~n9155 ) | ( n11572 & n13239 ) | ( ~n9155 & n13239 ) ;
  assign n13241 = ~n11572 & n13240 ;
  assign n13243 = ( x5 & n13239 ) | ( x5 & n13241 ) | ( n13239 & n13241 ) ;
  assign n13242 = ( x5 & ~n13241 ) | ( x5 & n13239 ) | ( ~n13241 & n13239 ) ;
  assign n13244 = ( n13241 & ~n13243 ) | ( n13241 & n13242 ) | ( ~n13243 & n13242 ) ;
  assign n13245 = ( n12905 & ~n12952 ) | ( n12905 & n12910 ) | ( ~n12952 & n12910 ) ;
  assign n13246 = ( n12910 & ~n12905 ) | ( n12910 & n12952 ) | ( ~n12905 & n12952 ) ;
  assign n13247 = ( n13245 & ~n12910 ) | ( n13245 & n13246 ) | ( ~n12910 & n13246 ) ;
  assign n13251 = n11152 | n9997 ;
  assign n13248 = ~n9160 & n11158 ;
  assign n13249 = ~n9558 & n11155 ;
  assign n13250 = n13248 | n13249 ;
  assign n13252 = ( n13251 & ~n9997 ) | ( n13251 & n13250 ) | ( ~n9997 & n13250 ) ;
  assign n13253 = ( n9155 & n11254 ) | ( n9155 & n13252 ) | ( n11254 & n13252 ) ;
  assign n13254 = ( n11254 & ~n13253 ) | ( n11254 & 1'b0 ) | ( ~n13253 & 1'b0 ) ;
  assign n13255 = ( n13252 & ~x5 ) | ( n13252 & n13254 ) | ( ~x5 & n13254 ) ;
  assign n13256 = ( x5 & ~n13252 ) | ( x5 & n13254 ) | ( ~n13252 & n13254 ) ;
  assign n13257 = ( n13255 & ~n13254 ) | ( n13255 & n13256 ) | ( ~n13254 & n13256 ) ;
  assign n13261 = n11155 | n9997 ;
  assign n13258 = n9160 | n11161 ;
  assign n13259 = ~n9558 & n11158 ;
  assign n13260 = ( n13258 & ~n13259 ) | ( n13258 & 1'b0 ) | ( ~n13259 & 1'b0 ) ;
  assign n13262 = ( n9997 & ~n13261 ) | ( n9997 & n13260 ) | ( ~n13261 & n13260 ) ;
  assign n13263 = n9155 | n11451 ;
  assign n13264 = n13262 &  n13263 ;
  assign n13265 = x5 &  n13264 ;
  assign n13266 = x5 | n13264 ;
  assign n13267 = ~n13265 & n13266 ;
  assign n13268 = ( n12924 & ~n12914 ) | ( n12924 & n12951 ) | ( ~n12914 & n12951 ) ;
  assign n13269 = ( n12952 & ~n12924 ) | ( n12952 & n13268 ) | ( ~n12924 & n13268 ) ;
  assign n13271 = ( n12592 & n12940 ) | ( n12592 & n12950 ) | ( n12940 & n12950 ) ;
  assign n13270 = ( n12592 & ~n12940 ) | ( n12592 & n12950 ) | ( ~n12940 & n12950 ) ;
  assign n13272 = ( n12940 & ~n13271 ) | ( n12940 & n13270 ) | ( ~n13271 & n13270 ) ;
  assign n13273 = n9997 &  n11158 ;
  assign n13274 = n9160 | n11164 ;
  assign n13275 = n9558 | n11161 ;
  assign n13276 = n13274 &  n13275 ;
  assign n13277 = ( n13273 & ~n11158 ) | ( n13273 & n13276 ) | ( ~n11158 & n13276 ) ;
  assign n13278 = ( n9155 & ~n13277 ) | ( n9155 & n11463 ) | ( ~n13277 & n11463 ) ;
  assign n13279 = ( n11463 & ~n13278 ) | ( n11463 & 1'b0 ) | ( ~n13278 & 1'b0 ) ;
  assign n13281 = ( x5 & n13277 ) | ( x5 & n13279 ) | ( n13277 & n13279 ) ;
  assign n13280 = ( x5 & ~n13279 ) | ( x5 & n13277 ) | ( ~n13279 & n13277 ) ;
  assign n13282 = ( n13279 & ~n13281 ) | ( n13279 & n13280 ) | ( ~n13281 & n13280 ) ;
  assign n13286 = ~n9997 & n11161 ;
  assign n13283 = n9160 | n11166 ;
  assign n13284 = n9558 | n11164 ;
  assign n13285 = n13283 &  n13284 ;
  assign n13287 = ( n9997 & n13286 ) | ( n9997 & n13285 ) | ( n13286 & n13285 ) ;
  assign n13288 = n9155 | n11385 ;
  assign n13289 = n13287 &  n13288 ;
  assign n13290 = x5 &  n13289 ;
  assign n13291 = x5 | n13289 ;
  assign n13292 = ~n13290 & n13291 ;
  assign n13293 = ( x8 & n12925 ) | ( x8 & n12930 ) | ( n12925 & n12930 ) ;
  assign n13294 = ~n12925 & n13293 ;
  assign n13295 = ( n12937 & ~x8 ) | ( n12937 & n13294 ) | ( ~x8 & n13294 ) ;
  assign n13296 = ( x8 & ~n12937 ) | ( x8 & n13294 ) | ( ~n12937 & n13294 ) ;
  assign n13297 = ( n13295 & ~n13294 ) | ( n13295 & n13296 ) | ( ~n13294 & n13296 ) ;
  assign n13298 = x8 &  n12925 ;
  assign n13299 = n12930 &  n13298 ;
  assign n13300 = n12930 | n13298 ;
  assign n13301 = ~n13299 & n13300 ;
  assign n13331 = ~n9997 & n11166 ;
  assign n13328 = n9160 | n11172 ;
  assign n13329 = n9558 | n11168 ;
  assign n13330 = n13328 &  n13329 ;
  assign n13332 = ( n9997 & n13331 ) | ( n9997 & n13330 ) | ( n13331 & n13330 ) ;
  assign n13333 = n9155 | n11431 ;
  assign n13334 = n13332 &  n13333 ;
  assign n13335 = x5 &  n13334 ;
  assign n13336 = x5 | n13334 ;
  assign n13337 = ~n13335 & n13336 ;
  assign n13312 = n9154 &  n11170 ;
  assign n13316 = ~n9155 & n11369 ;
  assign n13313 = ~n9558 & n11170 ;
  assign n13314 = n9997 | n11172 ;
  assign n13315 = ~n13313 & n13314 ;
  assign n13317 = ( n9155 & n13316 ) | ( n9155 & n13315 ) | ( n13316 & n13315 ) ;
  assign n13323 = n11323 | n9155 ;
  assign n13321 = ~n9997 & n11168 ;
  assign n13318 = ~n9160 & n11170 ;
  assign n13319 = n9558 | n11172 ;
  assign n13320 = ~n13318 & n13319 ;
  assign n13322 = ( n9997 & n13321 ) | ( n9997 & n13320 ) | ( n13321 & n13320 ) ;
  assign n13324 = ( n9155 & ~n13323 ) | ( n9155 & n13322 ) | ( ~n13323 & n13322 ) ;
  assign n13325 = ( n13312 & n13317 ) | ( n13312 & n13324 ) | ( n13317 & n13324 ) ;
  assign n13326 = ( x5 & ~n13325 ) | ( x5 & n13312 ) | ( ~n13325 & n13312 ) ;
  assign n13327 = ( x5 & ~n13326 ) | ( x5 & 1'b0 ) | ( ~n13326 & 1'b0 ) ;
  assign n13338 = ( n12925 & ~n13337 ) | ( n12925 & n13327 ) | ( ~n13337 & n13327 ) ;
  assign n13305 = ~n9997 & n11164 ;
  assign n13302 = n9160 | n11168 ;
  assign n13303 = n9558 | n11166 ;
  assign n13304 = n13302 &  n13303 ;
  assign n13306 = ( n9997 & n13305 ) | ( n9997 & n13304 ) | ( n13305 & n13304 ) ;
  assign n13307 = ( n11397 & ~n9155 ) | ( n11397 & n13306 ) | ( ~n9155 & n13306 ) ;
  assign n13308 = ~n11397 & n13307 ;
  assign n13309 = ( x5 & ~n13306 ) | ( x5 & n13308 ) | ( ~n13306 & n13308 ) ;
  assign n13310 = ( n13306 & ~x5 ) | ( n13306 & n13308 ) | ( ~x5 & n13308 ) ;
  assign n13311 = ( n13309 & ~n13308 ) | ( n13309 & n13310 ) | ( ~n13308 & n13310 ) ;
  assign n13339 = ( n13301 & ~n13338 ) | ( n13301 & n13311 ) | ( ~n13338 & n13311 ) ;
  assign n13340 = ( n13292 & n13297 ) | ( n13292 & n13339 ) | ( n13297 & n13339 ) ;
  assign n13341 = ( n13272 & n13282 ) | ( n13272 & n13340 ) | ( n13282 & n13340 ) ;
  assign n13342 = ( n13267 & ~n13269 ) | ( n13267 & n13341 ) | ( ~n13269 & n13341 ) ;
  assign n13343 = ( n13247 & ~n13257 ) | ( n13247 & n13342 ) | ( ~n13257 & n13342 ) ;
  assign n13344 = ( n13234 & n13244 ) | ( n13234 & n13343 ) | ( n13244 & n13343 ) ;
  assign n13345 = ( n13231 & ~n13221 ) | ( n13231 & n13344 ) | ( ~n13221 & n13344 ) ;
  assign n13346 = ( n13216 & ~n13218 ) | ( n13216 & n13345 ) | ( ~n13218 & n13345 ) ;
  assign n13347 = ( n13204 & n13206 ) | ( n13204 & n13346 ) | ( n13206 & n13346 ) ;
  assign n13348 = ( n13192 & ~n13194 ) | ( n13192 & n13347 ) | ( ~n13194 & n13347 ) ;
  assign n13349 = ( n13182 & ~n13172 ) | ( n13182 & n13348 ) | ( ~n13172 & n13348 ) ;
  assign n13350 = ( n13159 & n13169 ) | ( n13159 & n13349 ) | ( n13169 & n13349 ) ;
  assign n13351 = ( n13156 & ~n13146 ) | ( n13156 & n13350 ) | ( ~n13146 & n13350 ) ;
  assign n13352 = ( n13141 & ~n13143 ) | ( n13141 & n13351 ) | ( ~n13143 & n13351 ) ;
  assign n13353 = ( n13129 & n13131 ) | ( n13129 & n13352 ) | ( n13131 & n13352 ) ;
  assign n13354 = ( n13117 & ~n13119 ) | ( n13117 & n13353 ) | ( ~n13119 & n13353 ) ;
  assign n13355 = ( n13107 & ~n13097 ) | ( n13107 & n13354 ) | ( ~n13097 & n13354 ) ;
  assign n13356 = ( n13084 & n13094 ) | ( n13084 & n13355 ) | ( n13094 & n13355 ) ;
  assign n13357 = ( n13081 & ~n13071 ) | ( n13081 & n13356 ) | ( ~n13071 & n13356 ) ;
  assign n13358 = ( n13066 & ~n13068 ) | ( n13066 & n13357 ) | ( ~n13068 & n13357 ) ;
  assign n13359 = ( n13054 & n13056 ) | ( n13054 & n13358 ) | ( n13056 & n13358 ) ;
  assign n13360 = ( n13042 & ~n13044 ) | ( n13042 & n13359 ) | ( ~n13044 & n13359 ) ;
  assign n13361 = ( n13032 & ~n13022 ) | ( n13032 & n13360 ) | ( ~n13022 & n13360 ) ;
  assign n13362 = ( n13007 & n13019 ) | ( n13007 & n13361 ) | ( n13019 & n13361 ) ;
  assign n13363 = ( n13002 & n13004 ) | ( n13002 & n13362 ) | ( n13004 & n13362 ) ;
  assign n13364 = ( n12976 & ~n12989 ) | ( n12976 & n13363 ) | ( ~n12989 & n13363 ) ;
  assign n13365 = ( n12976 & ~n13363 ) | ( n12976 & n12989 ) | ( ~n13363 & n12989 ) ;
  assign n13366 = ( n13364 & ~n12976 ) | ( n13364 & n13365 ) | ( ~n12976 & n13365 ) ;
  assign n13367 = ( n13004 & ~n13002 ) | ( n13004 & n13362 ) | ( ~n13002 & n13362 ) ;
  assign n13368 = ( n13002 & ~n13362 ) | ( n13002 & n13004 ) | ( ~n13362 & n13004 ) ;
  assign n13369 = ( n13367 & ~n13004 ) | ( n13367 & n13368 ) | ( ~n13004 & n13368 ) ;
  assign n13370 = n10015 | n11091 ;
  assign n13371 = n10486 | n11081 ;
  assign n13372 = n13370 &  n13371 ;
  assign n13373 = n10499 &  n11085 ;
  assign n13374 = ( n13372 & ~n10499 ) | ( n13372 & n13373 ) | ( ~n10499 & n13373 ) ;
  assign n13375 = ( n11081 & ~n11085 ) | ( n11081 & n11202 ) | ( ~n11085 & n11202 ) ;
  assign n13376 = ( n11085 & ~n11081 ) | ( n11085 & n11202 ) | ( ~n11081 & n11202 ) ;
  assign n13377 = ( n13375 & ~n11202 ) | ( n13375 & n13376 ) | ( ~n11202 & n13376 ) ;
  assign n13378 = ( n13374 & ~n10017 ) | ( n13374 & n13377 ) | ( ~n10017 & n13377 ) ;
  assign n13379 = ~n13377 & n13378 ;
  assign n13380 = ( x2 & ~n13374 ) | ( x2 & n13379 ) | ( ~n13374 & n13379 ) ;
  assign n13381 = ( n13374 & ~x2 ) | ( n13374 & n13379 ) | ( ~x2 & n13379 ) ;
  assign n13382 = ( n13380 & ~n13379 ) | ( n13380 & n13381 ) | ( ~n13379 & n13381 ) ;
  assign n13383 = ( n13007 & ~n13019 ) | ( n13007 & n13361 ) | ( ~n13019 & n13361 ) ;
  assign n13384 = ( n13019 & ~n13362 ) | ( n13019 & n13383 ) | ( ~n13362 & n13383 ) ;
  assign n13393 = ( x5 & n13312 ) | ( x5 & n13317 ) | ( n13312 & n13317 ) ;
  assign n13394 = ~n13312 & n13393 ;
  assign n13395 = ( n13324 & ~x5 ) | ( n13324 & n13394 ) | ( ~x5 & n13394 ) ;
  assign n13396 = ( x5 & ~n13324 ) | ( x5 & n13394 ) | ( ~n13324 & n13394 ) ;
  assign n13397 = ( n13395 & ~n13394 ) | ( n13395 & n13396 ) | ( ~n13394 & n13396 ) ;
  assign n13426 = n10015 | n11168 ;
  assign n13427 = n10486 | n11166 ;
  assign n13428 = n13426 &  n13427 ;
  assign n13429 = n10499 &  n11164 ;
  assign n13430 = ( n13428 & ~n10499 ) | ( n13428 & n13429 ) | ( ~n10499 & n13429 ) ;
  assign n13431 = ( n11397 & ~n10017 ) | ( n11397 & n13430 ) | ( ~n10017 & n13430 ) ;
  assign n13432 = ~n11397 & n13431 ;
  assign n13433 = ( x2 & ~n13430 ) | ( x2 & n13432 ) | ( ~n13430 & n13432 ) ;
  assign n13434 = ( n13430 & ~x2 ) | ( n13430 & n13432 ) | ( ~x2 & n13432 ) ;
  assign n13435 = ( n13433 & ~n13432 ) | ( n13433 & n13434 ) | ( ~n13432 & n13434 ) ;
  assign n13418 = n11166 &  n10499 ;
  assign n13415 = n10015 | n11172 ;
  assign n13416 = n10486 | n11168 ;
  assign n13417 = n13415 &  n13416 ;
  assign n13419 = ( n13418 & ~n10499 ) | ( n13418 & n13417 ) | ( ~n10499 & n13417 ) ;
  assign n13420 = n10017 | n11431 ;
  assign n13421 = n13419 &  n13420 ;
  assign n13422 = x2 &  n13421 ;
  assign n13423 = x2 | n13421 ;
  assign n13424 = ~n13422 & n13423 ;
  assign n13398 = n10567 &  n11323 ;
  assign n13404 = ( n10567 & ~n11369 ) | ( n10567 & 1'b0 ) | ( ~n11369 & 1'b0 ) ;
  assign n13405 = n10574 &  n11170 ;
  assign n13406 = ( x2 & ~n13405 ) | ( x2 & 1'b0 ) | ( ~n13405 & 1'b0 ) ;
  assign n13407 = n10499 &  n11172 ;
  assign n13408 = ( n13406 & ~n10499 ) | ( n13406 & n13407 ) | ( ~n10499 & n13407 ) ;
  assign n13409 = ~n13404 & n13408 ;
  assign n13399 = ~n10015 & n11170 ;
  assign n13400 = n10486 | n11172 ;
  assign n13401 = ~n13399 & n13400 ;
  assign n13402 = n10499 &  n11168 ;
  assign n13403 = ( n13401 & ~n10499 ) | ( n13401 & n13402 ) | ( ~n10499 & n13402 ) ;
  assign n13410 = x2 &  n13403 ;
  assign n13411 = ( n13409 & ~x2 ) | ( n13409 & n13410 ) | ( ~x2 & n13410 ) ;
  assign n13412 = ~n13398 & n13411 ;
  assign n13413 = ( x0 & ~n11170 ) | ( x0 & 1'b0 ) | ( ~n11170 & 1'b0 ) ;
  assign n13414 = ( n13412 & ~x0 ) | ( n13412 & n13413 ) | ( ~x0 & n13413 ) ;
  assign n13425 = ( n13312 & ~n13424 ) | ( n13312 & n13414 ) | ( ~n13424 & n13414 ) ;
  assign n13436 = x5 &  n13312 ;
  assign n13437 = n13317 &  n13436 ;
  assign n13438 = n13317 | n13436 ;
  assign n13439 = ~n13437 & n13438 ;
  assign n13440 = ( n13435 & ~n13425 ) | ( n13435 & n13439 ) | ( ~n13425 & n13439 ) ;
  assign n13444 = n11161 &  n10499 ;
  assign n13441 = n10015 | n11166 ;
  assign n13442 = n10486 | n11164 ;
  assign n13443 = n13441 &  n13442 ;
  assign n13445 = ( n13444 & ~n10499 ) | ( n13444 & n13443 ) | ( ~n10499 & n13443 ) ;
  assign n13446 = n10017 | n11385 ;
  assign n13447 = n13445 &  n13446 ;
  assign n13448 = x2 &  n13447 ;
  assign n13449 = x2 | n13447 ;
  assign n13450 = ~n13448 & n13449 ;
  assign n13451 = ( n13397 & n13440 ) | ( n13397 & n13450 ) | ( n13440 & n13450 ) ;
  assign n13455 = ~n11158 & n10499 ;
  assign n13452 = n10015 | n11164 ;
  assign n13453 = n10486 | n11161 ;
  assign n13454 = n13452 &  n13453 ;
  assign n13456 = ( n13455 & ~n10499 ) | ( n13455 & n13454 ) | ( ~n10499 & n13454 ) ;
  assign n13457 = ( n10017 & ~n13456 ) | ( n10017 & n11463 ) | ( ~n13456 & n11463 ) ;
  assign n13458 = ( n11463 & ~n13457 ) | ( n11463 & 1'b0 ) | ( ~n13457 & 1'b0 ) ;
  assign n13460 = ( x2 & n13456 ) | ( x2 & n13458 ) | ( n13456 & n13458 ) ;
  assign n13459 = ( x2 & ~n13458 ) | ( x2 & n13456 ) | ( ~n13458 & n13456 ) ;
  assign n13461 = ( n13458 & ~n13460 ) | ( n13458 & n13459 ) | ( ~n13460 & n13459 ) ;
  assign n13463 = ( n12925 & n13327 ) | ( n12925 & n13337 ) | ( n13327 & n13337 ) ;
  assign n13462 = ( n12925 & ~n13327 ) | ( n12925 & n13337 ) | ( ~n13327 & n13337 ) ;
  assign n13464 = ( n13327 & ~n13463 ) | ( n13327 & n13462 ) | ( ~n13463 & n13462 ) ;
  assign n13465 = ( n13451 & n13461 ) | ( n13451 & n13464 ) | ( n13461 & n13464 ) ;
  assign n13391 = ( n13311 & ~n13301 ) | ( n13311 & n13338 ) | ( ~n13301 & n13338 ) ;
  assign n13392 = ( n13339 & ~n13311 ) | ( n13339 & n13391 ) | ( ~n13311 & n13391 ) ;
  assign n13466 = n10015 | n11161 ;
  assign n13467 = ~n10486 & n11158 ;
  assign n13468 = ( n13466 & ~n13467 ) | ( n13466 & 1'b0 ) | ( ~n13467 & 1'b0 ) ;
  assign n13469 = ( n10499 & ~n11155 ) | ( n10499 & 1'b0 ) | ( ~n11155 & 1'b0 ) ;
  assign n13470 = ( n13468 & ~n10499 ) | ( n13468 & n13469 ) | ( ~n10499 & n13469 ) ;
  assign n13471 = n10017 | n11451 ;
  assign n13472 = n13470 &  n13471 ;
  assign n13473 = x2 &  n13472 ;
  assign n13474 = x2 | n13472 ;
  assign n13475 = ~n13473 & n13474 ;
  assign n13476 = ( n13465 & ~n13392 ) | ( n13465 & n13475 ) | ( ~n13392 & n13475 ) ;
  assign n13480 = ( n10499 & ~n11152 ) | ( n10499 & 1'b0 ) | ( ~n11152 & 1'b0 ) ;
  assign n13477 = ~n10015 & n11158 ;
  assign n13478 = ~n10486 & n11155 ;
  assign n13479 = n13477 | n13478 ;
  assign n13481 = ( n10499 & ~n13480 ) | ( n10499 & n13479 ) | ( ~n13480 & n13479 ) ;
  assign n13482 = ( n10017 & n11254 ) | ( n10017 & n13481 ) | ( n11254 & n13481 ) ;
  assign n13483 = ( n11254 & ~n13482 ) | ( n11254 & 1'b0 ) | ( ~n13482 & 1'b0 ) ;
  assign n13484 = ( n13481 & ~x2 ) | ( n13481 & n13483 ) | ( ~x2 & n13483 ) ;
  assign n13485 = ( x2 & ~n13481 ) | ( x2 & n13483 ) | ( ~n13481 & n13483 ) ;
  assign n13486 = ( n13484 & ~n13483 ) | ( n13484 & n13485 ) | ( ~n13483 & n13485 ) ;
  assign n13487 = ( n13292 & ~n13339 ) | ( n13292 & n13297 ) | ( ~n13339 & n13297 ) ;
  assign n13488 = ( n13297 & ~n13292 ) | ( n13297 & n13339 ) | ( ~n13292 & n13339 ) ;
  assign n13489 = ( n13487 & ~n13297 ) | ( n13487 & n13488 ) | ( ~n13297 & n13488 ) ;
  assign n13490 = ( n13476 & ~n13486 ) | ( n13476 & n13489 ) | ( ~n13486 & n13489 ) ;
  assign n13494 = n11149 &  n10499 ;
  assign n13491 = ~n10015 & n11155 ;
  assign n13492 = ~n10486 & n11152 ;
  assign n13493 = n13491 | n13492 ;
  assign n13495 = ( n10499 & ~n13494 ) | ( n10499 & n13493 ) | ( ~n13494 & n13493 ) ;
  assign n13496 = ( n10017 & ~n11572 ) | ( n10017 & n13495 ) | ( ~n11572 & n13495 ) ;
  assign n13497 = n11572 | n13496 ;
  assign n13498 = ( x2 & ~n13495 ) | ( x2 & n13497 ) | ( ~n13495 & n13497 ) ;
  assign n13499 = ( n13495 & ~x2 ) | ( n13495 & n13497 ) | ( ~x2 & n13497 ) ;
  assign n13500 = ( n13498 & ~n13497 ) | ( n13498 & n13499 ) | ( ~n13497 & n13499 ) ;
  assign n13501 = ( n13282 & ~n13272 ) | ( n13282 & n13340 ) | ( ~n13272 & n13340 ) ;
  assign n13502 = ( n13272 & ~n13340 ) | ( n13272 & n13282 ) | ( ~n13340 & n13282 ) ;
  assign n13503 = ( n13501 & ~n13282 ) | ( n13501 & n13502 ) | ( ~n13282 & n13502 ) ;
  assign n13504 = ( n13490 & n13500 ) | ( n13490 & n13503 ) | ( n13500 & n13503 ) ;
  assign n13515 = ( n13269 & ~n13267 ) | ( n13269 & n13341 ) | ( ~n13267 & n13341 ) ;
  assign n13516 = ( n13267 & ~n13341 ) | ( n13267 & n13269 ) | ( ~n13341 & n13269 ) ;
  assign n13517 = ( n13515 & ~n13269 ) | ( n13515 & n13516 ) | ( ~n13269 & n13516 ) ;
  assign n13505 = ~n10015 & n11152 ;
  assign n13506 = n10486 | n11149 ;
  assign n13507 = ~n13505 & n13506 ;
  assign n13508 = n10499 &  n11146 ;
  assign n13509 = ( n13507 & ~n10499 ) | ( n13507 & n13508 ) | ( ~n10499 & n13508 ) ;
  assign n13510 = ( n10017 & ~n13509 ) | ( n10017 & n11554 ) | ( ~n13509 & n11554 ) ;
  assign n13511 = ( n11554 & ~n13510 ) | ( n11554 & 1'b0 ) | ( ~n13510 & 1'b0 ) ;
  assign n13512 = ( x2 & ~n13509 ) | ( x2 & n13511 ) | ( ~n13509 & n13511 ) ;
  assign n13513 = ( n13509 & ~x2 ) | ( n13509 & n13511 ) | ( ~x2 & n13511 ) ;
  assign n13514 = ( n13512 & ~n13511 ) | ( n13512 & n13513 ) | ( ~n13511 & n13513 ) ;
  assign n13518 = ( n13504 & ~n13517 ) | ( n13504 & n13514 ) | ( ~n13517 & n13514 ) ;
  assign n13519 = ( n13247 & n13257 ) | ( n13247 & n13342 ) | ( n13257 & n13342 ) ;
  assign n13520 = ( n13257 & ~n13519 ) | ( n13257 & n13343 ) | ( ~n13519 & n13343 ) ;
  assign n13521 = n10015 | n11149 ;
  assign n13522 = n10486 | n11146 ;
  assign n13523 = n13521 &  n13522 ;
  assign n13524 = n10499 &  n11143 ;
  assign n13525 = ( n13523 & ~n10499 ) | ( n13523 & n13524 ) | ( ~n10499 & n13524 ) ;
  assign n13526 = n10017 | n11542 ;
  assign n13527 = n13525 &  n13526 ;
  assign n13528 = x2 &  n13527 ;
  assign n13529 = x2 | n13527 ;
  assign n13530 = ~n13528 & n13529 ;
  assign n13531 = ( n13518 & ~n13520 ) | ( n13518 & n13530 ) | ( ~n13520 & n13530 ) ;
  assign n13532 = ( n13234 & ~n13244 ) | ( n13234 & n13343 ) | ( ~n13244 & n13343 ) ;
  assign n13533 = ( n13244 & ~n13344 ) | ( n13244 & n13532 ) | ( ~n13344 & n13532 ) ;
  assign n13537 = n11140 &  n10499 ;
  assign n13534 = n10015 | n11146 ;
  assign n13535 = n10486 | n11143 ;
  assign n13536 = n13534 &  n13535 ;
  assign n13538 = ( n13537 & ~n10499 ) | ( n13537 & n13536 ) | ( ~n10499 & n13536 ) ;
  assign n13539 = n10017 | n11699 ;
  assign n13540 = n13538 &  n13539 ;
  assign n13541 = x2 &  n13540 ;
  assign n13542 = x2 | n13540 ;
  assign n13543 = ~n13541 & n13542 ;
  assign n13544 = ( n13531 & n13533 ) | ( n13531 & n13543 ) | ( n13533 & n13543 ) ;
  assign n13389 = ( n13221 & ~n13344 ) | ( n13221 & n13231 ) | ( ~n13344 & n13231 ) ;
  assign n13390 = ( n13345 & ~n13231 ) | ( n13345 & n13389 ) | ( ~n13231 & n13389 ) ;
  assign n13545 = n10015 | n11143 ;
  assign n13546 = n10486 | n11140 ;
  assign n13547 = n13545 &  n13546 ;
  assign n13548 = n10499 &  n11137 ;
  assign n13549 = ( n13547 & ~n10499 ) | ( n13547 & n13548 ) | ( ~n10499 & n13548 ) ;
  assign n13550 = n10017 | n11687 ;
  assign n13551 = n13549 &  n13550 ;
  assign n13552 = x2 &  n13551 ;
  assign n13553 = x2 | n13551 ;
  assign n13554 = ~n13552 & n13553 ;
  assign n13555 = ( n13544 & ~n13390 ) | ( n13544 & n13554 ) | ( ~n13390 & n13554 ) ;
  assign n13566 = ( n13216 & ~n13345 ) | ( n13216 & n13218 ) | ( ~n13345 & n13218 ) ;
  assign n13567 = ( n13218 & ~n13216 ) | ( n13218 & n13345 ) | ( ~n13216 & n13345 ) ;
  assign n13568 = ( n13566 & ~n13218 ) | ( n13566 & n13567 ) | ( ~n13218 & n13567 ) ;
  assign n13556 = n10015 | n11140 ;
  assign n13557 = n10486 | n11137 ;
  assign n13558 = n13556 &  n13557 ;
  assign n13559 = ( n10499 & ~n11134 ) | ( n10499 & 1'b0 ) | ( ~n11134 & 1'b0 ) ;
  assign n13560 = ( n13558 & ~n10499 ) | ( n13558 & n13559 ) | ( ~n10499 & n13559 ) ;
  assign n13561 = ( n10017 & ~n13560 ) | ( n10017 & n11242 ) | ( ~n13560 & n11242 ) ;
  assign n13562 = ( n11242 & ~n13561 ) | ( n11242 & 1'b0 ) | ( ~n13561 & 1'b0 ) ;
  assign n13564 = ( x2 & n13560 ) | ( x2 & n13562 ) | ( n13560 & n13562 ) ;
  assign n13563 = ( x2 & ~n13562 ) | ( x2 & n13560 ) | ( ~n13562 & n13560 ) ;
  assign n13565 = ( n13562 & ~n13564 ) | ( n13562 & n13563 ) | ( ~n13564 & n13563 ) ;
  assign n13569 = ( n13555 & ~n13568 ) | ( n13555 & n13565 ) | ( ~n13568 & n13565 ) ;
  assign n13570 = n10015 | n11137 ;
  assign n13571 = ~n10486 & n11134 ;
  assign n13572 = ( n13570 & ~n13571 ) | ( n13570 & 1'b0 ) | ( ~n13571 & 1'b0 ) ;
  assign n13573 = n10499 &  n11131 ;
  assign n13574 = ( n13572 & ~n10499 ) | ( n13572 & n13573 ) | ( ~n10499 & n13573 ) ;
  assign n13575 = ( n10017 & ~n13574 ) | ( n10017 & n11888 ) | ( ~n13574 & n11888 ) ;
  assign n13576 = ( n11888 & ~n13575 ) | ( n11888 & 1'b0 ) | ( ~n13575 & 1'b0 ) ;
  assign n13578 = ( x2 & n13574 ) | ( x2 & n13576 ) | ( n13574 & n13576 ) ;
  assign n13577 = ( x2 & ~n13576 ) | ( x2 & n13574 ) | ( ~n13576 & n13574 ) ;
  assign n13579 = ( n13576 & ~n13578 ) | ( n13576 & n13577 ) | ( ~n13578 & n13577 ) ;
  assign n13580 = ( n13206 & ~n13204 ) | ( n13206 & n13346 ) | ( ~n13204 & n13346 ) ;
  assign n13581 = ( n13204 & ~n13346 ) | ( n13204 & n13206 ) | ( ~n13346 & n13206 ) ;
  assign n13582 = ( n13580 & ~n13206 ) | ( n13580 & n13581 ) | ( ~n13206 & n13581 ) ;
  assign n13583 = ( n13569 & n13579 ) | ( n13569 & n13582 ) | ( n13579 & n13582 ) ;
  assign n13594 = ( n13194 & ~n13192 ) | ( n13194 & n13347 ) | ( ~n13192 & n13347 ) ;
  assign n13595 = ( n13192 & ~n13347 ) | ( n13192 & n13194 ) | ( ~n13347 & n13194 ) ;
  assign n13596 = ( n13594 & ~n13194 ) | ( n13594 & n13595 ) | ( ~n13194 & n13595 ) ;
  assign n13584 = ~n10015 & n11134 ;
  assign n13585 = n10486 | n11131 ;
  assign n13586 = ~n13584 & n13585 ;
  assign n13587 = n10499 &  n11128 ;
  assign n13588 = ( n13586 & ~n10499 ) | ( n13586 & n13587 ) | ( ~n10499 & n13587 ) ;
  assign n13589 = ( n11871 & ~n10017 ) | ( n11871 & n13588 ) | ( ~n10017 & n13588 ) ;
  assign n13590 = ~n11871 & n13589 ;
  assign n13591 = ( x2 & ~n13588 ) | ( x2 & n13590 ) | ( ~n13588 & n13590 ) ;
  assign n13592 = ( n13588 & ~x2 ) | ( n13588 & n13590 ) | ( ~x2 & n13590 ) ;
  assign n13593 = ( n13591 & ~n13590 ) | ( n13591 & n13592 ) | ( ~n13590 & n13592 ) ;
  assign n13597 = ( n13583 & ~n13596 ) | ( n13583 & n13593 ) | ( ~n13596 & n13593 ) ;
  assign n13598 = ( n13172 & ~n13348 ) | ( n13172 & n13182 ) | ( ~n13348 & n13182 ) ;
  assign n13599 = ( n13349 & ~n13182 ) | ( n13349 & n13598 ) | ( ~n13182 & n13598 ) ;
  assign n13603 = ~n11125 & n10499 ;
  assign n13600 = n10015 | n11131 ;
  assign n13601 = n10486 | n11128 ;
  assign n13602 = n13600 &  n13601 ;
  assign n13604 = ( n13603 & ~n10499 ) | ( n13603 & n13602 ) | ( ~n10499 & n13602 ) ;
  assign n13605 = ~n10017 & n11859 ;
  assign n13606 = ( n13604 & ~n13605 ) | ( n13604 & 1'b0 ) | ( ~n13605 & 1'b0 ) ;
  assign n13607 = x2 &  n13606 ;
  assign n13608 = x2 | n13606 ;
  assign n13609 = ~n13607 & n13608 ;
  assign n13610 = ( n13597 & ~n13599 ) | ( n13597 & n13609 ) | ( ~n13599 & n13609 ) ;
  assign n13611 = ( n13159 & ~n13169 ) | ( n13159 & n13349 ) | ( ~n13169 & n13349 ) ;
  assign n13612 = ( n13169 & ~n13350 ) | ( n13169 & n13611 ) | ( ~n13350 & n13611 ) ;
  assign n13613 = n10015 | n11128 ;
  assign n13614 = ~n10486 & n11125 ;
  assign n13615 = ( n13613 & ~n13614 ) | ( n13613 & 1'b0 ) | ( ~n13614 & 1'b0 ) ;
  assign n13616 = n10499 &  n11122 ;
  assign n13617 = ( n13615 & ~n10499 ) | ( n13615 & n13616 ) | ( ~n10499 & n13616 ) ;
  assign n13618 = ~n10017 & n12100 ;
  assign n13619 = ( n13617 & ~n13618 ) | ( n13617 & 1'b0 ) | ( ~n13618 & 1'b0 ) ;
  assign n13620 = x2 &  n13619 ;
  assign n13621 = x2 | n13619 ;
  assign n13622 = ~n13620 & n13621 ;
  assign n13623 = ( n13610 & n13612 ) | ( n13610 & n13622 ) | ( n13612 & n13622 ) ;
  assign n13387 = ( n13146 & ~n13350 ) | ( n13146 & n13156 ) | ( ~n13350 & n13156 ) ;
  assign n13388 = ( n13351 & ~n13156 ) | ( n13351 & n13387 ) | ( ~n13156 & n13387 ) ;
  assign n13627 = ~n11119 & n10499 ;
  assign n13624 = ~n10015 & n11125 ;
  assign n13625 = n10486 | n11122 ;
  assign n13626 = ~n13624 & n13625 ;
  assign n13628 = ( n13627 & ~n10499 ) | ( n13627 & n13626 ) | ( ~n10499 & n13626 ) ;
  assign n13629 = ~n10017 & n12088 ;
  assign n13630 = ( n13628 & ~n13629 ) | ( n13628 & 1'b0 ) | ( ~n13629 & 1'b0 ) ;
  assign n13631 = x2 &  n13630 ;
  assign n13632 = x2 | n13630 ;
  assign n13633 = ~n13631 & n13632 ;
  assign n13634 = ( n13623 & ~n13388 ) | ( n13623 & n13633 ) | ( ~n13388 & n13633 ) ;
  assign n13645 = ( n13141 & ~n13351 ) | ( n13141 & n13143 ) | ( ~n13351 & n13143 ) ;
  assign n13646 = ( n13143 & ~n13141 ) | ( n13143 & n13351 ) | ( ~n13141 & n13351 ) ;
  assign n13647 = ( n13645 & ~n13143 ) | ( n13645 & n13646 ) | ( ~n13143 & n13646 ) ;
  assign n13635 = n10015 | n11122 ;
  assign n13636 = ~n10486 & n11119 ;
  assign n13637 = ( n13635 & ~n13636 ) | ( n13635 & 1'b0 ) | ( ~n13636 & 1'b0 ) ;
  assign n13638 = ( n10499 & ~n11116 ) | ( n10499 & 1'b0 ) | ( ~n11116 & 1'b0 ) ;
  assign n13639 = ( n13637 & ~n10499 ) | ( n13637 & n13638 ) | ( ~n10499 & n13638 ) ;
  assign n13640 = ( n11230 & ~n10017 ) | ( n11230 & n13639 ) | ( ~n10017 & n13639 ) ;
  assign n13641 = ~n11230 & n13640 ;
  assign n13642 = ( x2 & ~n13639 ) | ( x2 & n13641 ) | ( ~n13639 & n13641 ) ;
  assign n13643 = ( n13639 & ~x2 ) | ( n13639 & n13641 ) | ( ~x2 & n13641 ) ;
  assign n13644 = ( n13642 & ~n13641 ) | ( n13642 & n13643 ) | ( ~n13641 & n13643 ) ;
  assign n13648 = ( n13634 & ~n13647 ) | ( n13634 & n13644 ) | ( ~n13647 & n13644 ) ;
  assign n13652 = n11113 &  n10499 ;
  assign n13649 = ~n10015 & n11119 ;
  assign n13650 = ~n10486 & n11116 ;
  assign n13651 = n13649 | n13650 ;
  assign n13653 = ( n10499 & ~n13652 ) | ( n10499 & n13651 ) | ( ~n13652 & n13651 ) ;
  assign n13654 = ( n10017 & ~n12369 ) | ( n10017 & n13653 ) | ( ~n12369 & n13653 ) ;
  assign n13655 = n12369 | n13654 ;
  assign n13656 = ( x2 & ~n13653 ) | ( x2 & n13655 ) | ( ~n13653 & n13655 ) ;
  assign n13657 = ( n13653 & ~x2 ) | ( n13653 & n13655 ) | ( ~x2 & n13655 ) ;
  assign n13658 = ( n13656 & ~n13655 ) | ( n13656 & n13657 ) | ( ~n13655 & n13657 ) ;
  assign n13659 = ( n13131 & ~n13129 ) | ( n13131 & n13352 ) | ( ~n13129 & n13352 ) ;
  assign n13660 = ( n13129 & ~n13352 ) | ( n13129 & n13131 ) | ( ~n13352 & n13131 ) ;
  assign n13661 = ( n13659 & ~n13131 ) | ( n13659 & n13660 ) | ( ~n13131 & n13660 ) ;
  assign n13662 = ( n13648 & n13658 ) | ( n13648 & n13661 ) | ( n13658 & n13661 ) ;
  assign n13673 = ( n13119 & ~n13117 ) | ( n13119 & n13353 ) | ( ~n13117 & n13353 ) ;
  assign n13674 = ( n13117 & ~n13353 ) | ( n13117 & n13119 ) | ( ~n13353 & n13119 ) ;
  assign n13675 = ( n13673 & ~n13119 ) | ( n13673 & n13674 ) | ( ~n13119 & n13674 ) ;
  assign n13663 = ~n10015 & n11116 ;
  assign n13664 = n10486 | n11113 ;
  assign n13665 = ~n13663 & n13664 ;
  assign n13666 = n10499 &  n11110 ;
  assign n13667 = ( n13665 & ~n10499 ) | ( n13665 & n13666 ) | ( ~n10499 & n13666 ) ;
  assign n13668 = ( n10017 & ~n13667 ) | ( n10017 & n12352 ) | ( ~n13667 & n12352 ) ;
  assign n13669 = ( n12352 & ~n13668 ) | ( n12352 & 1'b0 ) | ( ~n13668 & 1'b0 ) ;
  assign n13671 = ( x2 & n13667 ) | ( x2 & n13669 ) | ( n13667 & n13669 ) ;
  assign n13670 = ( x2 & ~n13669 ) | ( x2 & n13667 ) | ( ~n13669 & n13667 ) ;
  assign n13672 = ( n13669 & ~n13671 ) | ( n13669 & n13670 ) | ( ~n13671 & n13670 ) ;
  assign n13676 = ( n13662 & ~n13675 ) | ( n13662 & n13672 ) | ( ~n13675 & n13672 ) ;
  assign n13677 = ( n13097 & ~n13354 ) | ( n13097 & n13107 ) | ( ~n13354 & n13107 ) ;
  assign n13678 = ( n13355 & ~n13107 ) | ( n13355 & n13677 ) | ( ~n13107 & n13677 ) ;
  assign n13679 = n10015 | n11113 ;
  assign n13680 = n10486 | n11110 ;
  assign n13681 = n13679 &  n13680 ;
  assign n13682 = ( n10499 & ~n11107 ) | ( n10499 & 1'b0 ) | ( ~n11107 & 1'b0 ) ;
  assign n13683 = ( n13681 & ~n10499 ) | ( n13681 & n13682 ) | ( ~n10499 & n13682 ) ;
  assign n13684 = ~n10017 & n12340 ;
  assign n13685 = ( n13683 & ~n13684 ) | ( n13683 & 1'b0 ) | ( ~n13684 & 1'b0 ) ;
  assign n13686 = x2 &  n13685 ;
  assign n13687 = x2 | n13685 ;
  assign n13688 = ~n13686 & n13687 ;
  assign n13689 = ( n13676 & ~n13678 ) | ( n13676 & n13688 ) | ( ~n13678 & n13688 ) ;
  assign n13690 = ( n13084 & ~n13094 ) | ( n13084 & n13355 ) | ( ~n13094 & n13355 ) ;
  assign n13691 = ( n13094 & ~n13356 ) | ( n13094 & n13690 ) | ( ~n13356 & n13690 ) ;
  assign n13692 = n10015 | n11110 ;
  assign n13693 = ~n10486 & n11107 ;
  assign n13694 = ( n13692 & ~n13693 ) | ( n13692 & 1'b0 ) | ( ~n13693 & 1'b0 ) ;
  assign n13695 = n10499 &  n11104 ;
  assign n13696 = ( n13694 & ~n10499 ) | ( n13694 & n13695 ) | ( ~n10499 & n13695 ) ;
  assign n13697 = ~n10017 & n12662 ;
  assign n13698 = ( n13696 & ~n13697 ) | ( n13696 & 1'b0 ) | ( ~n13697 & 1'b0 ) ;
  assign n13699 = x2 &  n13698 ;
  assign n13700 = x2 | n13698 ;
  assign n13701 = ~n13699 & n13700 ;
  assign n13702 = ( n13689 & n13691 ) | ( n13689 & n13701 ) | ( n13691 & n13701 ) ;
  assign n13385 = ( n13071 & ~n13356 ) | ( n13071 & n13081 ) | ( ~n13356 & n13081 ) ;
  assign n13386 = ( n13357 & ~n13081 ) | ( n13357 & n13385 ) | ( ~n13081 & n13385 ) ;
  assign n13703 = ~n10015 & n11107 ;
  assign n13704 = n10486 | n11104 ;
  assign n13705 = ~n13703 & n13704 ;
  assign n13706 = n10499 &  n11101 ;
  assign n13707 = ( n13705 & ~n10499 ) | ( n13705 & n13706 ) | ( ~n10499 & n13706 ) ;
  assign n13708 = n10017 | n12650 ;
  assign n13709 = n13707 &  n13708 ;
  assign n13710 = x2 &  n13709 ;
  assign n13711 = x2 | n13709 ;
  assign n13712 = ~n13710 & n13711 ;
  assign n13713 = ( n13702 & ~n13386 ) | ( n13702 & n13712 ) | ( ~n13386 & n13712 ) ;
  assign n13724 = ( n13066 & ~n13357 ) | ( n13066 & n13068 ) | ( ~n13357 & n13068 ) ;
  assign n13725 = ( n13068 & ~n13066 ) | ( n13068 & n13357 ) | ( ~n13066 & n13357 ) ;
  assign n13726 = ( n13724 & ~n13068 ) | ( n13724 & n13725 ) | ( ~n13068 & n13725 ) ;
  assign n13717 = n11098 &  n10499 ;
  assign n13714 = n10015 | n11104 ;
  assign n13715 = n10486 | n11101 ;
  assign n13716 = n13714 &  n13715 ;
  assign n13718 = ( n13717 & ~n10499 ) | ( n13717 & n13716 ) | ( ~n10499 & n13716 ) ;
  assign n13719 = ( n11218 & ~n10017 ) | ( n11218 & n13718 ) | ( ~n10017 & n13718 ) ;
  assign n13720 = ~n11218 & n13719 ;
  assign n13722 = ( x2 & n13718 ) | ( x2 & n13720 ) | ( n13718 & n13720 ) ;
  assign n13721 = ( x2 & ~n13720 ) | ( x2 & n13718 ) | ( ~n13720 & n13718 ) ;
  assign n13723 = ( n13720 & ~n13722 ) | ( n13720 & n13721 ) | ( ~n13722 & n13721 ) ;
  assign n13727 = ( n13713 & ~n13726 ) | ( n13713 & n13723 ) | ( ~n13726 & n13723 ) ;
  assign n13728 = n10015 | n11101 ;
  assign n13729 = n10486 | n11098 ;
  assign n13730 = n13728 &  n13729 ;
  assign n13731 = n10499 &  n11095 ;
  assign n13732 = ( n13730 & ~n10499 ) | ( n13730 & n13731 ) | ( ~n10499 & n13731 ) ;
  assign n13733 = ( n13014 & ~n10017 ) | ( n13014 & n13732 ) | ( ~n10017 & n13732 ) ;
  assign n13734 = ~n13014 & n13733 ;
  assign n13736 = ( x2 & n13732 ) | ( x2 & n13734 ) | ( n13732 & n13734 ) ;
  assign n13735 = ( x2 & ~n13734 ) | ( x2 & n13732 ) | ( ~n13734 & n13732 ) ;
  assign n13737 = ( n13734 & ~n13736 ) | ( n13734 & n13735 ) | ( ~n13736 & n13735 ) ;
  assign n13738 = ( n13056 & ~n13054 ) | ( n13056 & n13358 ) | ( ~n13054 & n13358 ) ;
  assign n13739 = ( n13054 & ~n13358 ) | ( n13054 & n13056 ) | ( ~n13358 & n13056 ) ;
  assign n13740 = ( n13738 & ~n13056 ) | ( n13738 & n13739 ) | ( ~n13056 & n13739 ) ;
  assign n13741 = ( n13727 & n13737 ) | ( n13727 & n13740 ) | ( n13737 & n13740 ) ;
  assign n13752 = ( n13044 & ~n13042 ) | ( n13044 & n13359 ) | ( ~n13042 & n13359 ) ;
  assign n13753 = ( n13042 & ~n13359 ) | ( n13042 & n13044 ) | ( ~n13359 & n13044 ) ;
  assign n13754 = ( n13752 & ~n13044 ) | ( n13752 & n13753 ) | ( ~n13044 & n13753 ) ;
  assign n13742 = n10015 | n11098 ;
  assign n13743 = n10486 | n11095 ;
  assign n13744 = n13742 &  n13743 ;
  assign n13745 = n10499 &  n11093 ;
  assign n13746 = ( n13744 & ~n10499 ) | ( n13744 & n13745 ) | ( ~n10499 & n13745 ) ;
  assign n13747 = ( n12997 & ~n10017 ) | ( n12997 & n13746 ) | ( ~n10017 & n13746 ) ;
  assign n13748 = ~n12997 & n13747 ;
  assign n13749 = ( x2 & ~n13746 ) | ( x2 & n13748 ) | ( ~n13746 & n13748 ) ;
  assign n13750 = ( n13746 & ~x2 ) | ( n13746 & n13748 ) | ( ~x2 & n13748 ) ;
  assign n13751 = ( n13749 & ~n13748 ) | ( n13749 & n13750 ) | ( ~n13748 & n13750 ) ;
  assign n13755 = ( n13741 & ~n13754 ) | ( n13741 & n13751 ) | ( ~n13754 & n13751 ) ;
  assign n13756 = ( n13022 & ~n13360 ) | ( n13022 & n13032 ) | ( ~n13360 & n13032 ) ;
  assign n13757 = ( n13361 & ~n13032 ) | ( n13361 & n13756 ) | ( ~n13032 & n13756 ) ;
  assign n13758 = n10015 | n11095 ;
  assign n13759 = n10486 | n11093 ;
  assign n13760 = n13758 &  n13759 ;
  assign n13761 = n10499 &  n11091 ;
  assign n13762 = ( n13760 & ~n10499 ) | ( n13760 & n13761 ) | ( ~n10499 & n13761 ) ;
  assign n13763 = n10017 | n12984 ;
  assign n13764 = n13762 &  n13763 ;
  assign n13765 = x2 &  n13764 ;
  assign n13766 = x2 | n13764 ;
  assign n13767 = ~n13765 & n13766 ;
  assign n13768 = ( n13755 & ~n13757 ) | ( n13755 & n13767 ) | ( ~n13757 & n13767 ) ;
  assign n13769 = n10015 | n11093 ;
  assign n13770 = n10486 | n11091 ;
  assign n13771 = n13769 &  n13770 ;
  assign n13772 = n10499 &  n11081 ;
  assign n13773 = ( n13771 & ~n10499 ) | ( n13771 & n13772 ) | ( ~n10499 & n13772 ) ;
  assign n13774 = ( n11091 & ~n11081 ) | ( n11091 & n11201 ) | ( ~n11081 & n11201 ) ;
  assign n13775 = ( n11081 & ~n11202 ) | ( n11081 & n13774 ) | ( ~n11202 & n13774 ) ;
  assign n13776 = n10017 | n13775 ;
  assign n13777 = n13773 &  n13776 ;
  assign n13778 = x2 &  n13777 ;
  assign n13779 = x2 | n13777 ;
  assign n13780 = ~n13778 & n13779 ;
  assign n13781 = ( n13384 & n13768 ) | ( n13384 & n13780 ) | ( n13768 & n13780 ) ;
  assign n13782 = ( n13369 & n13382 ) | ( n13369 & n13781 ) | ( n13382 & n13781 ) ;
  assign n13783 = ( n11211 & n13366 ) | ( n11211 & n13782 ) | ( n13366 & n13782 ) ;
  assign n13784 = ( n13366 & ~n11211 ) | ( n13366 & n13782 ) | ( ~n11211 & n13782 ) ;
  assign n13785 = ( n11211 & ~n13783 ) | ( n11211 & n13784 ) | ( ~n13783 & n13784 ) ;
  assign n13786 = ( n13369 & ~n13382 ) | ( n13369 & n13781 ) | ( ~n13382 & n13781 ) ;
  assign n13787 = ( n13382 & ~n13782 ) | ( n13382 & n13786 ) | ( ~n13782 & n13786 ) ;
  assign n13788 = ~n13785 & n13787 ;
  assign n13789 = ( n13785 & ~n13787 ) | ( n13785 & 1'b0 ) | ( ~n13787 & 1'b0 ) ;
  assign n13790 = n13788 | n13789 ;
  assign n13794 = n13790 | n3644 ;
  assign n13791 = n3653 | n13785 ;
  assign n13792 = ( n3657 & ~n13787 ) | ( n3657 & 1'b0 ) | ( ~n13787 & 1'b0 ) ;
  assign n13793 = ( n13791 & ~n13792 ) | ( n13791 & 1'b0 ) | ( ~n13792 & 1'b0 ) ;
  assign n13795 = ( n3644 & ~n13794 ) | ( n3644 & n13793 ) | ( ~n13794 & n13793 ) ;
  assign n13796 = n514 | n13795 ;
  assign n13797 = n1327 | n2666 ;
  assign n13798 = ( n785 & ~n403 ) | ( n785 & n13797 ) | ( ~n403 & n13797 ) ;
  assign n13799 = n403 | n13798 ;
  assign n13800 = n212 | n13799 ;
  assign n13801 = ( n928 & ~n5454 ) | ( n928 & 1'b0 ) | ( ~n5454 & 1'b0 ) ;
  assign n13802 = ( n299 & ~n461 ) | ( n299 & n13801 ) | ( ~n461 & n13801 ) ;
  assign n13803 = ~n299 & n13802 ;
  assign n13804 = n541 | n669 ;
  assign n13805 = ( n13804 & ~n528 ) | ( n13804 & n665 ) | ( ~n528 & n665 ) ;
  assign n13806 = n528 | n13805 ;
  assign n13807 = n526 | n13806 ;
  assign n13808 = n2347 | n2633 ;
  assign n13809 = ( n13803 & n13807 ) | ( n13803 & n13808 ) | ( n13807 & n13808 ) ;
  assign n13810 = ( n2188 & ~n13803 ) | ( n2188 & n13809 ) | ( ~n13803 & n13809 ) ;
  assign n13811 = ( n2188 & ~n13810 ) | ( n2188 & 1'b0 ) | ( ~n13810 & 1'b0 ) ;
  assign n13812 = ( n810 & ~n13800 ) | ( n810 & n13811 ) | ( ~n13800 & n13811 ) ;
  assign n13813 = ( n13812 & ~n810 ) | ( n13812 & 1'b0 ) | ( ~n810 & 1'b0 ) ;
  assign n13814 = ( n163 & ~n733 ) | ( n163 & n13813 ) | ( ~n733 & n13813 ) ;
  assign n13815 = ~n163 & n13814 ;
  assign n13816 = ( n628 & ~n529 ) | ( n628 & n13815 ) | ( ~n529 & n13815 ) ;
  assign n13817 = ~n628 & n13816 ;
  assign n13818 = ~n196 & n13817 ;
  assign n13819 = ( x29 & n3776 ) | ( x29 & n13818 ) | ( n3776 & n13818 ) ;
  assign n13820 = ( x29 & ~n3776 ) | ( x29 & n13818 ) | ( ~n3776 & n13818 ) ;
  assign n13821 = ( n3776 & ~n13819 ) | ( n3776 & n13820 ) | ( ~n13819 & n13820 ) ;
  assign n13822 = n3644 | n4452 ;
  assign n13826 = n863 | n3652 ;
  assign n13823 = n599 | n3653 ;
  assign n13824 = ~n702 & n3657 ;
  assign n13825 = ( n13823 & ~n13824 ) | ( n13823 & 1'b0 ) | ( ~n13824 & 1'b0 ) ;
  assign n13827 = ( n863 & ~n13826 ) | ( n863 & n13825 ) | ( ~n13826 & n13825 ) ;
  assign n13828 = n13822 &  n13827 ;
  assign n13829 = ( n13821 & ~n3923 ) | ( n13821 & n13828 ) | ( ~n3923 & n13828 ) ;
  assign n13830 = ( n3923 & ~n13828 ) | ( n3923 & n13821 ) | ( ~n13828 & n13821 ) ;
  assign n13831 = ( n13829 & ~n13821 ) | ( n13829 & n13830 ) | ( ~n13821 & n13830 ) ;
  assign n13833 = ( n4047 & ~n3928 ) | ( n4047 & n11075 ) | ( ~n3928 & n11075 ) ;
  assign n13832 = ( n3642 & ~n3925 ) | ( n3642 & n3662 ) | ( ~n3925 & n3662 ) ;
  assign n13834 = ( n13831 & ~n13833 ) | ( n13831 & n13832 ) | ( ~n13833 & n13832 ) ;
  assign n13835 = ( n13831 & ~n13832 ) | ( n13831 & n13833 ) | ( ~n13832 & n13833 ) ;
  assign n13836 = ( ~n13831 & n13834 ) | ( ~n13831 & n13835 ) | ( n13834 & n13835 ) ;
  assign n13840 = n13836 &  n10499 ;
  assign n13837 = n10015 | n11085 ;
  assign n13838 = n10486 | n11078 ;
  assign n13839 = n13837 &  n13838 ;
  assign n13841 = ( n13840 & ~n10499 ) | ( n13840 & n13839 ) | ( ~n10499 & n13839 ) ;
  assign n13843 = ( n11078 & n11205 ) | ( n11078 & n13836 ) | ( n11205 & n13836 ) ;
  assign n13842 = ( n11205 & ~n11078 ) | ( n11205 & n13836 ) | ( ~n11078 & n13836 ) ;
  assign n13844 = ( n11078 & ~n13843 ) | ( n11078 & n13842 ) | ( ~n13843 & n13842 ) ;
  assign n13845 = ( n13841 & ~n10017 ) | ( n13841 & n13844 ) | ( ~n10017 & n13844 ) ;
  assign n13846 = ~n13844 & n13845 ;
  assign n13847 = ( x2 & ~n13841 ) | ( x2 & n13846 ) | ( ~n13841 & n13846 ) ;
  assign n13848 = ( n13841 & ~x2 ) | ( n13841 & n13846 ) | ( ~x2 & n13846 ) ;
  assign n13849 = ( n13847 & ~n13846 ) | ( n13847 & n13848 ) | ( ~n13846 & n13848 ) ;
  assign n13880 = ~n4482 & n11155 ;
  assign n13881 = ~n4495 & n11152 ;
  assign n13882 = n13880 | n13881 ;
  assign n13883 = ~n4962 & n11149 ;
  assign n13884 = ( n4962 & ~n13882 ) | ( n4962 & n13883 ) | ( ~n13882 & n13883 ) ;
  assign n13885 = ( n11572 & ~n4478 ) | ( n11572 & n13884 ) | ( ~n4478 & n13884 ) ;
  assign n13886 = ~n11572 & n13885 ;
  assign n13888 = ( x26 & n13884 ) | ( x26 & n13886 ) | ( n13884 & n13886 ) ;
  assign n13887 = ( x26 & ~n13886 ) | ( x26 & n13884 ) | ( ~n13886 & n13884 ) ;
  assign n13889 = ( n13886 & ~n13888 ) | ( n13886 & n13887 ) | ( ~n13888 & n13887 ) ;
  assign n13890 = n108 | n3419 ;
  assign n13891 = ( n13890 & ~n1672 ) | ( n13890 & n6679 ) | ( ~n1672 & n6679 ) ;
  assign n13892 = n1672 | n13891 ;
  assign n13893 = n5682 | n13892 ;
  assign n13894 = ( n3708 & ~n3753 ) | ( n3708 & n13893 ) | ( ~n3753 & n13893 ) ;
  assign n13895 = ( n4384 & ~n3708 ) | ( n4384 & n13894 ) | ( ~n3708 & n13894 ) ;
  assign n13896 = ( n4384 & ~n13895 ) | ( n4384 & 1'b0 ) | ( ~n13895 & 1'b0 ) ;
  assign n13897 = ( n747 & n820 ) | ( n747 & n13896 ) | ( n820 & n13896 ) ;
  assign n13898 = ~n747 & n13897 ;
  assign n13899 = ( n13898 & ~n495 ) | ( n13898 & n796 ) | ( ~n495 & n796 ) ;
  assign n13900 = ( n13899 & ~n796 ) | ( n13899 & 1'b0 ) | ( ~n796 & 1'b0 ) ;
  assign n13901 = ( n13900 & ~n531 ) | ( n13900 & n569 ) | ( ~n531 & n569 ) ;
  assign n13902 = ( n13901 & ~n569 ) | ( n13901 & 1'b0 ) | ( ~n569 & 1'b0 ) ;
  assign n13903 = ~n342 & n13902 ;
  assign n13909 = ~n3644 & n11431 ;
  assign n13904 = n3653 | n11166 ;
  assign n13905 = ( n3657 & ~n11168 ) | ( n3657 & 1'b0 ) | ( ~n11168 & 1'b0 ) ;
  assign n13906 = ( n3652 & ~n11172 ) | ( n3652 & 1'b0 ) | ( ~n11172 & 1'b0 ) ;
  assign n13907 = n13905 | n13906 ;
  assign n13908 = ( n13904 & ~n13907 ) | ( n13904 & 1'b0 ) | ( ~n13907 & 1'b0 ) ;
  assign n13910 = ( n3644 & n13909 ) | ( n3644 & n13908 ) | ( n13909 & n13908 ) ;
  assign n13911 = ( n11376 & ~n13903 ) | ( n11376 & n13910 ) | ( ~n13903 & n13910 ) ;
  assign n13912 = ( n11376 & ~n13910 ) | ( n11376 & n13903 ) | ( ~n13910 & n13903 ) ;
  assign n13913 = ( n13911 & ~n11376 ) | ( n13911 & n13912 ) | ( ~n11376 & n13912 ) ;
  assign n13914 = n4430 &  n11158 ;
  assign n13915 = n523 | n11164 ;
  assign n13916 = n3939 | n11161 ;
  assign n13917 = n13915 &  n13916 ;
  assign n13918 = ( n13914 & ~n11158 ) | ( n13914 & n13917 ) | ( ~n11158 & n13917 ) ;
  assign n13919 = ~n601 & n11463 ;
  assign n13920 = ( n13918 & ~n13919 ) | ( n13918 & 1'b0 ) | ( ~n13919 & 1'b0 ) ;
  assign n13921 = x29 &  n13920 ;
  assign n13922 = x29 | n13920 ;
  assign n13923 = ~n13921 & n13922 ;
  assign n13924 = ( n11378 & ~n11438 ) | ( n11378 & n11390 ) | ( ~n11438 & n11390 ) ;
  assign n13925 = ( n13913 & ~n13923 ) | ( n13913 & n13924 ) | ( ~n13923 & n13924 ) ;
  assign n13926 = ( n13913 & ~n13924 ) | ( n13913 & n13923 ) | ( ~n13924 & n13923 ) ;
  assign n13927 = ( n13925 & ~n13913 ) | ( n13925 & n13926 ) | ( ~n13913 & n13926 ) ;
  assign n13928 = ( n13889 & ~n11533 ) | ( n13889 & n13927 ) | ( ~n11533 & n13927 ) ;
  assign n13929 = ( n11533 & ~n13927 ) | ( n11533 & n13889 ) | ( ~n13927 & n13889 ) ;
  assign n13930 = ( n13928 & ~n13889 ) | ( n13928 & n13929 ) | ( ~n13889 & n13929 ) ;
  assign n13941 = ( n11535 & n11547 ) | ( n11535 & n11674 ) | ( n11547 & n11674 ) ;
  assign n13934 = ~n5135 & n11140 ;
  assign n13931 = n5010 | n11146 ;
  assign n13932 = n5067 | n11143 ;
  assign n13933 = n13931 &  n13932 ;
  assign n13935 = ( n5135 & n13934 ) | ( n5135 & n13933 ) | ( n13934 & n13933 ) ;
  assign n13936 = n5012 | n11699 ;
  assign n13937 = n13935 &  n13936 ;
  assign n13938 = x23 &  n13937 ;
  assign n13939 = x23 | n13937 ;
  assign n13940 = ~n13938 & n13939 ;
  assign n13942 = ( n13930 & ~n13941 ) | ( n13930 & n13940 ) | ( ~n13941 & n13940 ) ;
  assign n13943 = ( n13930 & ~n13940 ) | ( n13930 & n13941 ) | ( ~n13940 & n13941 ) ;
  assign n13944 = ( n13942 & ~n13930 ) | ( n13942 & n13943 ) | ( ~n13930 & n13943 ) ;
  assign n13870 = ( n5339 & ~n11137 ) | ( n5339 & 1'b0 ) | ( ~n11137 & 1'b0 ) ;
  assign n13871 = ~n5761 & n11134 ;
  assign n13872 = n13870 | n13871 ;
  assign n13873 = ~n5837 & n11131 ;
  assign n13874 = ( n5837 & ~n13872 ) | ( n5837 & n13873 ) | ( ~n13872 & n13873 ) ;
  assign n13875 = ( n5341 & ~n13874 ) | ( n5341 & n11888 ) | ( ~n13874 & n11888 ) ;
  assign n13876 = ( n11888 & ~n13875 ) | ( n11888 & 1'b0 ) | ( ~n13875 & 1'b0 ) ;
  assign n13878 = ( x20 & n13874 ) | ( x20 & n13876 ) | ( n13874 & n13876 ) ;
  assign n13877 = ( x20 & ~n13876 ) | ( x20 & n13874 ) | ( ~n13876 & n13874 ) ;
  assign n13879 = ( n13876 & ~n13878 ) | ( n13876 & n13877 ) | ( ~n13878 & n13877 ) ;
  assign n13945 = ( n11850 & ~n13944 ) | ( n11850 & n13879 ) | ( ~n13944 & n13879 ) ;
  assign n13946 = ( n13879 & ~n11850 ) | ( n13879 & n13944 ) | ( ~n11850 & n13944 ) ;
  assign n13947 = ( n13945 & ~n13879 ) | ( n13945 & n13946 ) | ( ~n13879 & n13946 ) ;
  assign n13958 = ( n11852 & n11864 ) | ( n11852 & n12075 ) | ( n11864 & n12075 ) ;
  assign n13951 = ~n6395 & n11122 ;
  assign n13948 = n5970 | n11128 ;
  assign n13949 = ~n6170 & n11125 ;
  assign n13950 = ( n13948 & ~n13949 ) | ( n13948 & 1'b0 ) | ( ~n13949 & 1'b0 ) ;
  assign n13952 = ( n6395 & n13951 ) | ( n6395 & n13950 ) | ( n13951 & n13950 ) ;
  assign n13953 = ~n5972 & n12100 ;
  assign n13954 = ( n13952 & ~n13953 ) | ( n13952 & 1'b0 ) | ( ~n13953 & 1'b0 ) ;
  assign n13955 = x17 &  n13954 ;
  assign n13956 = x17 | n13954 ;
  assign n13957 = ~n13955 & n13956 ;
  assign n13959 = ( n13947 & ~n13958 ) | ( n13947 & n13957 ) | ( ~n13958 & n13957 ) ;
  assign n13960 = ( n13947 & ~n13957 ) | ( n13947 & n13958 ) | ( ~n13957 & n13958 ) ;
  assign n13961 = ( n13959 & ~n13947 ) | ( n13959 & n13960 ) | ( ~n13947 & n13960 ) ;
  assign n13861 = ~n6530 & n11119 ;
  assign n13862 = ~n6983 & n11116 ;
  assign n13863 = n13861 | n13862 ;
  assign n13860 = ( n7097 & ~n11113 ) | ( n7097 & 1'b0 ) | ( ~n11113 & 1'b0 ) ;
  assign n13864 = ( n11113 & ~n13863 ) | ( n11113 & n13860 ) | ( ~n13863 & n13860 ) ;
  assign n13865 = ( n12369 & ~n6532 ) | ( n12369 & n13864 ) | ( ~n6532 & n13864 ) ;
  assign n13866 = ~n12369 & n13865 ;
  assign n13868 = ( x14 & n13864 ) | ( x14 & n13866 ) | ( n13864 & n13866 ) ;
  assign n13867 = ( x14 & ~n13866 ) | ( x14 & n13864 ) | ( ~n13866 & n13864 ) ;
  assign n13869 = ( n13866 & ~n13868 ) | ( n13866 & n13867 ) | ( ~n13868 & n13867 ) ;
  assign n13962 = ( n12331 & ~n13961 ) | ( n12331 & n13869 ) | ( ~n13961 & n13869 ) ;
  assign n13963 = ( n13869 & ~n12331 ) | ( n13869 & n13961 ) | ( ~n12331 & n13961 ) ;
  assign n13964 = ( n13962 & ~n13869 ) | ( n13962 & n13963 ) | ( ~n13869 & n13963 ) ;
  assign n13975 = ( n12333 & n12345 ) | ( n12333 & n12637 ) | ( n12345 & n12637 ) ;
  assign n13965 = ( n7253 & ~n11110 ) | ( n7253 & 1'b0 ) | ( ~n11110 & 1'b0 ) ;
  assign n13966 = ~n7518 & n11107 ;
  assign n13967 = n13965 | n13966 ;
  assign n13968 = ~n7783 & n11104 ;
  assign n13969 = ( n7783 & ~n13967 ) | ( n7783 & n13968 ) | ( ~n13967 & n13968 ) ;
  assign n13970 = ~n7255 & n12662 ;
  assign n13971 = ( n13969 & ~n13970 ) | ( n13969 & 1'b0 ) | ( ~n13970 & 1'b0 ) ;
  assign n13972 = x11 &  n13971 ;
  assign n13973 = x11 | n13971 ;
  assign n13974 = ~n13972 & n13973 ;
  assign n13976 = ( n13964 & ~n13975 ) | ( n13964 & n13974 ) | ( ~n13975 & n13974 ) ;
  assign n13977 = ( n13964 & ~n13974 ) | ( n13964 & n13975 ) | ( ~n13974 & n13975 ) ;
  assign n13978 = ( n13976 & ~n13964 ) | ( n13976 & n13977 ) | ( ~n13964 & n13977 ) ;
  assign n13853 = ~n8764 & n11095 ;
  assign n13850 = ( n8105 & ~n11101 ) | ( n8105 & 1'b0 ) | ( ~n11101 & 1'b0 ) ;
  assign n13851 = n8429 | n11098 ;
  assign n13852 = ~n13850 & n13851 ;
  assign n13854 = ( n8764 & n13853 ) | ( n8764 & n13852 ) | ( n13853 & n13852 ) ;
  assign n13855 = ( n13014 & ~n8107 ) | ( n13014 & n13854 ) | ( ~n8107 & n13854 ) ;
  assign n13856 = ~n13014 & n13855 ;
  assign n13858 = ( x8 & n13854 ) | ( x8 & n13856 ) | ( n13854 & n13856 ) ;
  assign n13857 = ( x8 & ~n13856 ) | ( x8 & n13854 ) | ( ~n13856 & n13854 ) ;
  assign n13859 = ( n13856 & ~n13858 ) | ( n13856 & n13857 ) | ( ~n13858 & n13857 ) ;
  assign n13979 = ( n12974 & ~n13978 ) | ( n12974 & n13859 ) | ( ~n13978 & n13859 ) ;
  assign n13980 = ( n13859 & ~n12974 ) | ( n13859 & n13978 ) | ( ~n12974 & n13978 ) ;
  assign n13981 = ( n13979 & ~n13859 ) | ( n13979 & n13980 ) | ( ~n13859 & n13980 ) ;
  assign n13992 = ( n12976 & n12989 ) | ( n12976 & n13363 ) | ( n12989 & n13363 ) ;
  assign n13985 = ~n9997 & n11081 ;
  assign n13982 = n9160 | n11093 ;
  assign n13983 = n9558 | n11091 ;
  assign n13984 = n13982 &  n13983 ;
  assign n13986 = ( n9997 & n13985 ) | ( n9997 & n13984 ) | ( n13985 & n13984 ) ;
  assign n13987 = n9155 | n13775 ;
  assign n13988 = n13986 &  n13987 ;
  assign n13989 = x5 &  n13988 ;
  assign n13990 = x5 | n13988 ;
  assign n13991 = ~n13989 & n13990 ;
  assign n13993 = ( n13981 & ~n13992 ) | ( n13981 & n13991 ) | ( ~n13992 & n13991 ) ;
  assign n13994 = ( n13981 & ~n13991 ) | ( n13981 & n13992 ) | ( ~n13991 & n13992 ) ;
  assign n13995 = ( n13993 & ~n13981 ) | ( n13993 & n13994 ) | ( ~n13981 & n13994 ) ;
  assign n13996 = ( n13783 & ~n13995 ) | ( n13783 & n13849 ) | ( ~n13995 & n13849 ) ;
  assign n13997 = ( n13849 & ~n13783 ) | ( n13849 & n13995 ) | ( ~n13783 & n13995 ) ;
  assign n13998 = ( n13849 & ~n13996 ) | ( n13849 & ~n13997 ) | ( ~n13996 & ~n13997 ) ;
  assign n13999 = n13788 &  n13998 ;
  assign n14000 = n13788 | n13998 ;
  assign n14001 = ~n13999 & n14000 ;
  assign n14002 = n3644 | n14001 ;
  assign n14003 = ( n3652 & ~n13787 ) | ( n3652 & 1'b0 ) | ( ~n13787 & 1'b0 ) ;
  assign n14004 = ( n3657 & ~n13785 ) | ( n3657 & 1'b0 ) | ( ~n13785 & 1'b0 ) ;
  assign n14005 = n14003 | n14004 ;
  assign n14006 = ~n3653 & n13998 ;
  assign n14007 = ( n3653 & ~n14005 ) | ( n3653 & n14006 ) | ( ~n14005 & n14006 ) ;
  assign n14008 = n14002 &  n14007 ;
  assign n14009 = n213 | n720 ;
  assign n14010 = n459 | n14009 ;
  assign n14011 = ( n301 & ~n889 ) | ( n301 & n14010 ) | ( ~n889 & n14010 ) ;
  assign n14012 = n889 | n14011 ;
  assign n14013 = ( n4138 & ~n632 ) | ( n4138 & n14012 ) | ( ~n632 & n14012 ) ;
  assign n14014 = n632 | n14013 ;
  assign n14015 = ( n4533 & ~n6732 ) | ( n4533 & n14014 ) | ( ~n6732 & n14014 ) ;
  assign n14016 = ( n4533 & ~n14015 ) | ( n4533 & 1'b0 ) | ( ~n14015 & 1'b0 ) ;
  assign n14017 = ( n1954 & n5576 ) | ( n1954 & n14016 ) | ( n5576 & n14016 ) ;
  assign n14018 = ~n1954 & n14017 ;
  assign n14019 = ( n1512 & ~n2082 ) | ( n1512 & n14018 ) | ( ~n2082 & n14018 ) ;
  assign n14020 = ~n1512 & n14019 ;
  assign n14021 = ( n402 & n1762 ) | ( n402 & n14020 ) | ( n1762 & n14020 ) ;
  assign n14022 = ~n1762 & n14021 ;
  assign n14023 = ( n14022 & ~n712 ) | ( n14022 & n800 ) | ( ~n712 & n800 ) ;
  assign n14024 = ( n14023 & ~n800 ) | ( n14023 & 1'b0 ) | ( ~n800 & 1'b0 ) ;
  assign n14025 = ( n453 & ~n452 ) | ( n453 & n14024 ) | ( ~n452 & n14024 ) ;
  assign n14026 = ~n453 & n14025 ;
  assign n14027 = ( n529 & ~n568 ) | ( n529 & n14026 ) | ( ~n568 & n14026 ) ;
  assign n14028 = ~n529 & n14027 ;
  assign n14029 = ( n13796 & n14008 ) | ( n13796 & n14028 ) | ( n14008 & n14028 ) ;
  assign n14030 = n62 | n415 ;
  assign n14031 = n721 | n14030 ;
  assign n14032 = ( n3663 & ~n5413 ) | ( n3663 & n14031 ) | ( ~n5413 & n14031 ) ;
  assign n14033 = ( n2889 & n5413 ) | ( n2889 & n14032 ) | ( n5413 & n14032 ) ;
  assign n14034 = ( n2889 & ~n14033 ) | ( n2889 & 1'b0 ) | ( ~n14033 & 1'b0 ) ;
  assign n14035 = ( n2525 & ~n5674 ) | ( n2525 & n14034 ) | ( ~n5674 & n14034 ) ;
  assign n14036 = ( n14035 & ~n2525 ) | ( n14035 & 1'b0 ) | ( ~n2525 & 1'b0 ) ;
  assign n14037 = ( n4513 & ~n14036 ) | ( n4513 & n1904 ) | ( ~n14036 & n1904 ) ;
  assign n14038 = ( n1904 & ~n14037 ) | ( n1904 & 1'b0 ) | ( ~n14037 & 1'b0 ) ;
  assign n14039 = ( n1093 & ~n570 ) | ( n1093 & n14038 ) | ( ~n570 & n14038 ) ;
  assign n14040 = ~n1093 & n14039 ;
  assign n14041 = ( n604 & ~n647 ) | ( n604 & n14040 ) | ( ~n647 & n14040 ) ;
  assign n14042 = ~n604 & n14041 ;
  assign n14043 = ( n761 & ~n864 ) | ( n761 & n14042 ) | ( ~n864 & n14042 ) ;
  assign n14044 = ~n761 & n14043 ;
  assign n14045 = ( n456 & ~n266 ) | ( n456 & n14044 ) | ( ~n266 & n14044 ) ;
  assign n14046 = ~n456 & n14045 ;
  assign n14047 = ~n236 & n14046 ;
  assign n14048 = ( n3923 & n13821 ) | ( n3923 & n13828 ) | ( n13821 & n13828 ) ;
  assign n14049 = ( n626 & ~n913 ) | ( n626 & 1'b0 ) | ( ~n913 & 1'b0 ) ;
  assign n14050 = ( n1243 & ~n5617 ) | ( n1243 & n14049 ) | ( ~n5617 & n14049 ) ;
  assign n14051 = ~n1243 & n14050 ;
  assign n14052 = ( n586 & n13800 ) | ( n586 & n14051 ) | ( n13800 & n14051 ) ;
  assign n14053 = ( n774 & ~n14052 ) | ( n774 & n13800 ) | ( ~n14052 & n13800 ) ;
  assign n14054 = ( n774 & ~n14053 ) | ( n774 & 1'b0 ) | ( ~n14053 & 1'b0 ) ;
  assign n14055 = ( n128 & ~n616 ) | ( n128 & n14054 ) | ( ~n616 & n14054 ) ;
  assign n14056 = ~n128 & n14055 ;
  assign n14057 = ( n72 & ~n865 ) | ( n72 & n14056 ) | ( ~n865 & n14056 ) ;
  assign n14058 = ~n72 & n14057 ;
  assign n14059 = ~n787 & n14058 ;
  assign n14063 = n3937 | n3644 ;
  assign n14060 = ~n702 & n3652 ;
  assign n14061 = ~n599 & n3657 ;
  assign n14062 = n14060 | n14061 ;
  assign n14064 = ( n14063 & ~n3644 ) | ( n14063 & n14062 ) | ( ~n3644 & n14062 ) ;
  assign n14065 = ( n13819 & ~n14059 ) | ( n13819 & n14064 ) | ( ~n14059 & n14064 ) ;
  assign n14066 = ( n13819 & ~n14064 ) | ( n13819 & n14059 ) | ( ~n14064 & n14059 ) ;
  assign n14067 = ( n14065 & ~n13819 ) | ( n14065 & n14066 ) | ( ~n13819 & n14066 ) ;
  assign n14068 = ( n13831 & n13832 ) | ( n13831 & n13833 ) | ( n13832 & n13833 ) ;
  assign n14069 = ( n14048 & ~n14067 ) | ( n14048 & n14068 ) | ( ~n14067 & n14068 ) ;
  assign n14070 = ( n14048 & ~n14068 ) | ( n14048 & n14067 ) | ( ~n14068 & n14067 ) ;
  assign n14071 = ( n14069 & ~n14048 ) | ( n14069 & n14070 ) | ( ~n14048 & n14070 ) ;
  assign n14078 = ( n13836 & n13843 ) | ( n13836 & n14071 ) | ( n13843 & n14071 ) ;
  assign n14077 = ( n13836 & ~n14071 ) | ( n13836 & n13843 ) | ( ~n14071 & n13843 ) ;
  assign n14079 = ( n14071 & ~n14078 ) | ( n14071 & n14077 ) | ( ~n14078 & n14077 ) ;
  assign n14072 = n10015 | n11078 ;
  assign n14073 = n10486 | n13836 ;
  assign n14074 = n14072 &  n14073 ;
  assign n14075 = n10499 &  n14071 ;
  assign n14076 = ( n14074 & ~n10499 ) | ( n14074 & n14075 ) | ( ~n10499 & n14075 ) ;
  assign n14080 = ( n14076 & ~n10017 ) | ( n14076 & n14079 ) | ( ~n10017 & n14079 ) ;
  assign n14081 = ~n14079 & n14080 ;
  assign n14083 = ( x2 & n14076 ) | ( x2 & n14081 ) | ( n14076 & n14081 ) ;
  assign n14082 = ( x2 & ~n14081 ) | ( x2 & n14076 ) | ( ~n14081 & n14076 ) ;
  assign n14084 = ( n14081 & ~n14083 ) | ( n14081 & n14082 ) | ( ~n14083 & n14082 ) ;
  assign n14085 = ( n8105 & ~n11098 ) | ( n8105 & 1'b0 ) | ( ~n11098 & 1'b0 ) ;
  assign n14086 = n8429 | n11095 ;
  assign n14087 = ~n14085 & n14086 ;
  assign n14088 = ~n8764 & n11093 ;
  assign n14089 = ( n8764 & n14087 ) | ( n8764 & n14088 ) | ( n14087 & n14088 ) ;
  assign n14090 = ( n12997 & ~n8107 ) | ( n12997 & n14089 ) | ( ~n8107 & n14089 ) ;
  assign n14091 = ~n12997 & n14090 ;
  assign n14092 = ( x8 & ~n14089 ) | ( x8 & n14091 ) | ( ~n14089 & n14091 ) ;
  assign n14093 = ( n14089 & ~x8 ) | ( n14089 & n14091 ) | ( ~x8 & n14091 ) ;
  assign n14094 = ( n14092 & ~n14091 ) | ( n14092 & n14093 ) | ( ~n14091 & n14093 ) ;
  assign n14098 = ~n7097 & n11110 ;
  assign n14095 = ~n6530 & n11116 ;
  assign n14096 = n6983 | n11113 ;
  assign n14097 = ~n14095 & n14096 ;
  assign n14099 = ( n7097 & n14098 ) | ( n7097 & n14097 ) | ( n14098 & n14097 ) ;
  assign n14100 = ( n6532 & ~n14099 ) | ( n6532 & n12352 ) | ( ~n14099 & n12352 ) ;
  assign n14101 = ( n12352 & ~n14100 ) | ( n12352 & 1'b0 ) | ( ~n14100 & 1'b0 ) ;
  assign n14103 = ( x14 & n14099 ) | ( x14 & n14101 ) | ( n14099 & n14101 ) ;
  assign n14102 = ( x14 & ~n14101 ) | ( x14 & n14099 ) | ( ~n14101 & n14099 ) ;
  assign n14104 = ( n14101 & ~n14103 ) | ( n14101 & n14102 ) | ( ~n14103 & n14102 ) ;
  assign n14108 = ~n5837 & n11128 ;
  assign n14105 = n5339 &  n11134 ;
  assign n14106 = n5761 | n11131 ;
  assign n14107 = ~n14105 & n14106 ;
  assign n14109 = ( n5837 & n14108 ) | ( n5837 & n14107 ) | ( n14108 & n14107 ) ;
  assign n14110 = ( n11871 & ~n5341 ) | ( n11871 & n14109 ) | ( ~n5341 & n14109 ) ;
  assign n14111 = ~n11871 & n14110 ;
  assign n14112 = ( x20 & ~n14109 ) | ( x20 & n14111 ) | ( ~n14109 & n14111 ) ;
  assign n14113 = ( n14109 & ~x20 ) | ( n14109 & n14111 ) | ( ~x20 & n14111 ) ;
  assign n14114 = ( n14112 & ~n14111 ) | ( n14112 & n14113 ) | ( ~n14111 & n14113 ) ;
  assign n14118 = ~n4962 & n11146 ;
  assign n14115 = ~n4482 & n11152 ;
  assign n14116 = n4495 | n11149 ;
  assign n14117 = ~n14115 & n14116 ;
  assign n14119 = ( n4962 & n14118 ) | ( n4962 & n14117 ) | ( n14118 & n14117 ) ;
  assign n14120 = ( n4478 & ~n14119 ) | ( n4478 & n11554 ) | ( ~n14119 & n11554 ) ;
  assign n14121 = ( n11554 & ~n14120 ) | ( n11554 & 1'b0 ) | ( ~n14120 & 1'b0 ) ;
  assign n14122 = ( x26 & ~n14119 ) | ( x26 & n14121 ) | ( ~n14119 & n14121 ) ;
  assign n14123 = ( n14119 & ~x26 ) | ( n14119 & n14121 ) | ( ~x26 & n14121 ) ;
  assign n14124 = ( n14122 & ~n14121 ) | ( n14122 & n14123 ) | ( ~n14121 & n14123 ) ;
  assign n14166 = n3653 | n11164 ;
  assign n14167 = ( n3657 & ~n11166 ) | ( n3657 & 1'b0 ) | ( ~n11166 & 1'b0 ) ;
  assign n14168 = ( n3652 & ~n11168 ) | ( n3652 & 1'b0 ) | ( ~n11168 & 1'b0 ) ;
  assign n14169 = n14167 | n14168 ;
  assign n14170 = ( n14166 & ~n14169 ) | ( n14166 & 1'b0 ) | ( ~n14169 & 1'b0 ) ;
  assign n14171 = ~n3644 & n11397 ;
  assign n14172 = ( n3644 & n14170 ) | ( n3644 & n14171 ) | ( n14170 & n14171 ) ;
  assign n14125 = ~n254 & n1106 ;
  assign n14126 = ( n224 & ~n425 ) | ( n224 & n14125 ) | ( ~n425 & n14125 ) ;
  assign n14127 = ~n224 & n14126 ;
  assign n14128 = ~n549 & n14127 ;
  assign n14129 = n852 | n2996 ;
  assign n14130 = ( n530 & ~n259 ) | ( n530 & n14129 ) | ( ~n259 & n14129 ) ;
  assign n14131 = n259 | n14130 ;
  assign n14132 = ( n235 & ~n493 ) | ( n235 & n14131 ) | ( ~n493 & n14131 ) ;
  assign n14133 = n493 | n14132 ;
  assign n14134 = ( n404 & ~n372 ) | ( n404 & n14133 ) | ( ~n372 & n14133 ) ;
  assign n14135 = n372 | n14134 ;
  assign n14136 = ( n132 & ~n556 ) | ( n132 & n14135 ) | ( ~n556 & n14135 ) ;
  assign n14137 = n556 | n14136 ;
  assign n14138 = ( n14128 & ~n489 ) | ( n14128 & n14137 ) | ( ~n489 & n14137 ) ;
  assign n14139 = ( n604 & ~n14138 ) | ( n604 & n14128 ) | ( ~n14138 & n14128 ) ;
  assign n14140 = ~n604 & n14139 ;
  assign n14141 = ( n1461 & ~n3245 ) | ( n1461 & n14140 ) | ( ~n3245 & n14140 ) ;
  assign n14142 = ~n1461 & n14141 ;
  assign n14143 = ( n789 & ~n605 ) | ( n789 & n14142 ) | ( ~n605 & n14142 ) ;
  assign n14144 = ~n789 & n14143 ;
  assign n14145 = ( n275 & ~n494 ) | ( n275 & n14144 ) | ( ~n494 & n14144 ) ;
  assign n14146 = ~n275 & n14145 ;
  assign n14147 = ( n554 & ~n909 ) | ( n554 & n14146 ) | ( ~n909 & n14146 ) ;
  assign n14148 = ~n554 & n14147 ;
  assign n14149 = ( n89 & ~n618 ) | ( n89 & n14148 ) | ( ~n618 & n14148 ) ;
  assign n14150 = ~n89 & n14149 ;
  assign n14151 = ~n83 & n14150 ;
  assign n14152 = n576 | n3031 ;
  assign n14153 = ( n2594 & ~n5220 ) | ( n2594 & n14152 ) | ( ~n5220 & n14152 ) ;
  assign n14154 = ( n2594 & ~n14153 ) | ( n2594 & 1'b0 ) | ( ~n14153 & 1'b0 ) ;
  assign n14155 = ( n1599 & n2451 ) | ( n1599 & n14154 ) | ( n2451 & n14154 ) ;
  assign n14156 = ~n1599 & n14155 ;
  assign n14157 = ( n3170 & ~n14156 ) | ( n3170 & n2084 ) | ( ~n14156 & n2084 ) ;
  assign n14158 = ( n2084 & ~n14157 ) | ( n2084 & 1'b0 ) | ( ~n14157 & 1'b0 ) ;
  assign n14159 = ( n2192 & n14151 ) | ( n2192 & n14158 ) | ( n14151 & n14158 ) ;
  assign n14160 = ~n2192 & n14159 ;
  assign n14161 = ( n280 & ~n797 ) | ( n280 & n14160 ) | ( ~n797 & n14160 ) ;
  assign n14162 = ~n280 & n14161 ;
  assign n14163 = ( n191 & ~n139 ) | ( n191 & n14162 ) | ( ~n139 & n14162 ) ;
  assign n14164 = ~n191 & n14163 ;
  assign n14165 = ~n559 & n14164 ;
  assign n14173 = ( n11376 & n13903 ) | ( n11376 & n13910 ) | ( n13903 & n13910 ) ;
  assign n14174 = ( n14172 & ~n14165 ) | ( n14172 & n14173 ) | ( ~n14165 & n14173 ) ;
  assign n14175 = ( n14165 & ~n14172 ) | ( n14165 & n14173 ) | ( ~n14172 & n14173 ) ;
  assign n14176 = ( n14174 & ~n14173 ) | ( n14174 & n14175 ) | ( ~n14173 & n14175 ) ;
  assign n14180 = n11155 | n4430 ;
  assign n14177 = n523 | n11161 ;
  assign n14178 = ~n3939 & n11158 ;
  assign n14179 = ( n14177 & ~n14178 ) | ( n14177 & 1'b0 ) | ( ~n14178 & 1'b0 ) ;
  assign n14181 = ( n4430 & ~n14180 ) | ( n4430 & n14179 ) | ( ~n14180 & n14179 ) ;
  assign n14182 = n601 | n11451 ;
  assign n14183 = n14181 &  n14182 ;
  assign n14184 = x29 &  n14183 ;
  assign n14185 = x29 | n14183 ;
  assign n14186 = ~n14184 & n14185 ;
  assign n14187 = ( n13913 & n13923 ) | ( n13913 & n13924 ) | ( n13923 & n13924 ) ;
  assign n14188 = ( n14176 & ~n14186 ) | ( n14176 & n14187 ) | ( ~n14186 & n14187 ) ;
  assign n14189 = ( n14176 & ~n14187 ) | ( n14176 & n14186 ) | ( ~n14187 & n14186 ) ;
  assign n14190 = ( n14188 & ~n14176 ) | ( n14188 & n14189 ) | ( ~n14176 & n14189 ) ;
  assign n14191 = ( n13928 & n14124 ) | ( n13928 & n14190 ) | ( n14124 & n14190 ) ;
  assign n14192 = ( n13928 & ~n14124 ) | ( n13928 & n14190 ) | ( ~n14124 & n14190 ) ;
  assign n14193 = ( n14124 & ~n14191 ) | ( n14124 & n14192 ) | ( ~n14191 & n14192 ) ;
  assign n14197 = ~n5135 & n11137 ;
  assign n14194 = n5010 | n11143 ;
  assign n14195 = n5067 | n11140 ;
  assign n14196 = n14194 &  n14195 ;
  assign n14198 = ( n5135 & n14197 ) | ( n5135 & n14196 ) | ( n14197 & n14196 ) ;
  assign n14199 = n5012 | n11687 ;
  assign n14200 = n14198 &  n14199 ;
  assign n14201 = x23 &  n14200 ;
  assign n14202 = x23 | n14200 ;
  assign n14203 = ~n14201 & n14202 ;
  assign n14204 = ( n13940 & ~n13930 ) | ( n13940 & n13941 ) | ( ~n13930 & n13941 ) ;
  assign n14205 = ( n14193 & ~n14203 ) | ( n14193 & n14204 ) | ( ~n14203 & n14204 ) ;
  assign n14206 = ( n14193 & ~n14204 ) | ( n14193 & n14203 ) | ( ~n14204 & n14203 ) ;
  assign n14207 = ( n14205 & ~n14193 ) | ( n14205 & n14206 ) | ( ~n14193 & n14206 ) ;
  assign n14208 = ( n13945 & n14114 ) | ( n13945 & n14207 ) | ( n14114 & n14207 ) ;
  assign n14209 = ( n13945 & ~n14114 ) | ( n13945 & n14207 ) | ( ~n14114 & n14207 ) ;
  assign n14210 = ( n14114 & ~n14208 ) | ( n14114 & n14209 ) | ( ~n14208 & n14209 ) ;
  assign n14214 = n11119 | n6395 ;
  assign n14211 = ~n5970 & n11125 ;
  assign n14212 = n6170 | n11122 ;
  assign n14213 = ~n14211 & n14212 ;
  assign n14215 = ( n6395 & ~n14214 ) | ( n6395 & n14213 ) | ( ~n14214 & n14213 ) ;
  assign n14216 = ~n5972 & n12088 ;
  assign n14217 = ( n14215 & ~n14216 ) | ( n14215 & 1'b0 ) | ( ~n14216 & 1'b0 ) ;
  assign n14218 = x17 &  n14217 ;
  assign n14219 = x17 | n14217 ;
  assign n14220 = ~n14218 & n14219 ;
  assign n14221 = ( n13957 & ~n13947 ) | ( n13957 & n13958 ) | ( ~n13947 & n13958 ) ;
  assign n14222 = ( n14210 & ~n14220 ) | ( n14210 & n14221 ) | ( ~n14220 & n14221 ) ;
  assign n14223 = ( n14210 & ~n14221 ) | ( n14210 & n14220 ) | ( ~n14221 & n14220 ) ;
  assign n14224 = ( n14222 & ~n14210 ) | ( n14222 & n14223 ) | ( ~n14210 & n14223 ) ;
  assign n14225 = ( n13962 & n14104 ) | ( n13962 & n14224 ) | ( n14104 & n14224 ) ;
  assign n14226 = ( n13962 & ~n14104 ) | ( n13962 & n14224 ) | ( ~n14104 & n14224 ) ;
  assign n14227 = ( n14104 & ~n14225 ) | ( n14104 & n14226 ) | ( ~n14225 & n14226 ) ;
  assign n14231 = ~n7783 & n11101 ;
  assign n14228 = n7253 &  n11107 ;
  assign n14229 = n7518 | n11104 ;
  assign n14230 = ~n14228 & n14229 ;
  assign n14232 = ( n7783 & n14231 ) | ( n7783 & n14230 ) | ( n14231 & n14230 ) ;
  assign n14233 = n7255 | n12650 ;
  assign n14234 = n14232 &  n14233 ;
  assign n14235 = x11 &  n14234 ;
  assign n14236 = x11 | n14234 ;
  assign n14237 = ~n14235 & n14236 ;
  assign n14238 = ( n13974 & ~n13964 ) | ( n13974 & n13975 ) | ( ~n13964 & n13975 ) ;
  assign n14239 = ( n14227 & ~n14237 ) | ( n14227 & n14238 ) | ( ~n14237 & n14238 ) ;
  assign n14240 = ( n14227 & ~n14238 ) | ( n14227 & n14237 ) | ( ~n14238 & n14237 ) ;
  assign n14241 = ( n14239 & ~n14227 ) | ( n14239 & n14240 ) | ( ~n14227 & n14240 ) ;
  assign n14242 = ( n13979 & n14094 ) | ( n13979 & n14241 ) | ( n14094 & n14241 ) ;
  assign n14243 = ( n13979 & ~n14094 ) | ( n13979 & n14241 ) | ( ~n14094 & n14241 ) ;
  assign n14244 = ( n14094 & ~n14242 ) | ( n14094 & n14243 ) | ( ~n14242 & n14243 ) ;
  assign n14248 = ~n9997 & n11085 ;
  assign n14245 = n9160 | n11091 ;
  assign n14246 = n9558 | n11081 ;
  assign n14247 = n14245 &  n14246 ;
  assign n14249 = ( n9997 & n14248 ) | ( n9997 & n14247 ) | ( n14248 & n14247 ) ;
  assign n14250 = n9155 | n13377 ;
  assign n14251 = n14249 &  n14250 ;
  assign n14252 = x5 &  n14251 ;
  assign n14253 = x5 | n14251 ;
  assign n14254 = ~n14252 & n14253 ;
  assign n14255 = ( n13991 & ~n13981 ) | ( n13991 & n13992 ) | ( ~n13981 & n13992 ) ;
  assign n14256 = ( n14244 & ~n14254 ) | ( n14244 & n14255 ) | ( ~n14254 & n14255 ) ;
  assign n14257 = ( n14244 & ~n14255 ) | ( n14244 & n14254 ) | ( ~n14255 & n14254 ) ;
  assign n14258 = ( n14256 & ~n14244 ) | ( n14256 & n14257 ) | ( ~n14244 & n14257 ) ;
  assign n14259 = ( n13996 & n14084 ) | ( n13996 & n14258 ) | ( n14084 & n14258 ) ;
  assign n14260 = ( n13996 & ~n14084 ) | ( n13996 & n14258 ) | ( ~n14084 & n14258 ) ;
  assign n14261 = ( n14084 & ~n14259 ) | ( n14084 & n14260 ) | ( ~n14259 & n14260 ) ;
  assign n14263 = ~n13787 & n13998 ;
  assign n14264 = ( n13785 & ~n14263 ) | ( n13785 & n13998 ) | ( ~n14263 & n13998 ) ;
  assign n14266 = ( n13998 & n14261 ) | ( n13998 & n14264 ) | ( n14261 & n14264 ) ;
  assign n14265 = ( n14261 & ~n13998 ) | ( n14261 & n14264 ) | ( ~n13998 & n14264 ) ;
  assign n14267 = ( n13998 & ~n14266 ) | ( n13998 & n14265 ) | ( ~n14266 & n14265 ) ;
  assign n14272 = ~n3644 & n14267 ;
  assign n14262 = n3653 | n14261 ;
  assign n14268 = ( n3657 & ~n13998 ) | ( n3657 & 1'b0 ) | ( ~n13998 & 1'b0 ) ;
  assign n14269 = ( n3652 & ~n13785 ) | ( n3652 & 1'b0 ) | ( ~n13785 & 1'b0 ) ;
  assign n14270 = n14268 | n14269 ;
  assign n14271 = ( n14262 & ~n14270 ) | ( n14262 & 1'b0 ) | ( ~n14270 & 1'b0 ) ;
  assign n14273 = ( n3644 & n14272 ) | ( n3644 & n14271 ) | ( n14272 & n14271 ) ;
  assign n14274 = ( n14029 & n14047 ) | ( n14029 & n14273 ) | ( n14047 & n14273 ) ;
  assign n14282 = n3856 | n3998 ;
  assign n14275 = n2596 &  n2798 ;
  assign n14276 = ( n339 & ~n278 ) | ( n339 & n14275 ) | ( ~n278 & n14275 ) ;
  assign n14277 = ~n339 & n14276 ;
  assign n14278 = ( n255 & ~n14277 ) | ( n255 & n786 ) | ( ~n14277 & n786 ) ;
  assign n14279 = ( n786 & ~n14278 ) | ( n786 & 1'b0 ) | ( ~n14278 & 1'b0 ) ;
  assign n14280 = ( n228 & ~n139 ) | ( n228 & n14279 ) | ( ~n139 & n14279 ) ;
  assign n14281 = ~n228 & n14280 ;
  assign n14283 = ( n1046 & ~n14282 ) | ( n1046 & n14281 ) | ( ~n14282 & n14281 ) ;
  assign n14284 = ~n1046 & n14283 ;
  assign n14285 = ( n1679 & n2201 ) | ( n1679 & n14284 ) | ( n2201 & n14284 ) ;
  assign n14286 = ~n1679 & n14285 ;
  assign n14287 = ( n2029 & ~n2128 ) | ( n2029 & n14286 ) | ( ~n2128 & n14286 ) ;
  assign n14288 = ~n2029 & n14287 ;
  assign n14289 = ( n2666 & ~n102 ) | ( n2666 & n14288 ) | ( ~n102 & n14288 ) ;
  assign n14290 = ~n2666 & n14289 ;
  assign n14291 = ( n672 & ~n412 ) | ( n672 & n14290 ) | ( ~n412 & n14290 ) ;
  assign n14292 = ~n672 & n14291 ;
  assign n14293 = ( n384 & ~n266 ) | ( n384 & n14292 ) | ( ~n266 & n14292 ) ;
  assign n14294 = ~n384 & n14293 ;
  assign n14295 = ~n239 & n14294 ;
  assign n14296 = ( n45 & ~n48 ) | ( n45 & n103 ) | ( ~n48 & n103 ) ;
  assign n14297 = n48 | n14296 ;
  assign n14298 = ( n235 & ~n244 ) | ( n235 & n362 ) | ( ~n244 & n362 ) ;
  assign n14299 = n244 | n14298 ;
  assign n14300 = ( n52 & ~n271 ) | ( n52 & n14299 ) | ( ~n271 & n14299 ) ;
  assign n14301 = n271 | n14300 ;
  assign n14302 = ( n14297 & ~n45 ) | ( n14297 & n14301 ) | ( ~n45 & n14301 ) ;
  assign n14303 = n556 | n14302 ;
  assign n14304 = ( n2784 & ~n2687 ) | ( n2784 & n6633 ) | ( ~n2687 & n6633 ) ;
  assign n14305 = n2687 | n14304 ;
  assign n14306 = ( n72 & ~n61 ) | ( n72 & n14305 ) | ( ~n61 & n14305 ) ;
  assign n14307 = n61 | n14306 ;
  assign n14308 = ( n775 & ~n284 ) | ( n775 & n14307 ) | ( ~n284 & n14307 ) ;
  assign n14309 = n284 | n14308 ;
  assign n14310 = ( n382 & ~n459 ) | ( n382 & n14309 ) | ( ~n459 & n14309 ) ;
  assign n14311 = n459 | n14310 ;
  assign n14312 = ( n1030 & ~n3973 ) | ( n1030 & 1'b0 ) | ( ~n3973 & 1'b0 ) ;
  assign n14313 = ( n1991 & ~n3171 ) | ( n1991 & n14312 ) | ( ~n3171 & n14312 ) ;
  assign n14314 = ~n1991 & n14313 ;
  assign n14315 = ( n1511 & ~n1184 ) | ( n1511 & n14314 ) | ( ~n1184 & n14314 ) ;
  assign n14316 = ~n1511 & n14315 ;
  assign n14317 = ( n812 & ~n718 ) | ( n812 & n14316 ) | ( ~n718 & n14316 ) ;
  assign n14318 = ~n812 & n14317 ;
  assign n14319 = ( n149 & ~n274 ) | ( n149 & n14318 ) | ( ~n274 & n14318 ) ;
  assign n14320 = ~n149 & n14319 ;
  assign n14321 = ( n95 & ~n141 ) | ( n95 & n14320 ) | ( ~n141 & n14320 ) ;
  assign n14322 = ~n95 & n14321 ;
  assign n14323 = n2515 | n6059 ;
  assign n14324 = ( n14323 & ~n1729 ) | ( n14323 & n4808 ) | ( ~n1729 & n4808 ) ;
  assign n14325 = n1729 | n14324 ;
  assign n14326 = ( n1168 & ~n14322 ) | ( n1168 & n14325 ) | ( ~n14322 & n14325 ) ;
  assign n14327 = ( n1168 & ~n14326 ) | ( n1168 & 1'b0 ) | ( ~n14326 & 1'b0 ) ;
  assign n14328 = ( n14303 & ~n14311 ) | ( n14303 & n14327 ) | ( ~n14311 & n14327 ) ;
  assign n14329 = ~n14303 & n14328 ;
  assign n14330 = ( n906 & n14295 ) | ( n906 & n14329 ) | ( n14295 & n14329 ) ;
  assign n14331 = ~n906 & n14330 ;
  assign n14332 = ( n280 & ~n208 ) | ( n280 & n14331 ) | ( ~n208 & n14331 ) ;
  assign n14333 = ~n280 & n14332 ;
  assign n14334 = ( n214 & ~n192 ) | ( n214 & n14333 ) | ( ~n192 & n14333 ) ;
  assign n14335 = ~n214 & n14334 ;
  assign n14336 = ~n236 & n14335 ;
  assign n14356 = n10015 | n13836 ;
  assign n14357 = n10486 | n14071 ;
  assign n14358 = n14356 &  n14357 ;
  assign n14337 = ( n14059 & ~n13819 ) | ( n14059 & n14064 ) | ( ~n13819 & n14064 ) ;
  assign n14338 = ( n567 & ~n13807 ) | ( n567 & n931 ) | ( ~n13807 & n931 ) ;
  assign n14339 = ( n567 & ~n14338 ) | ( n567 & n662 ) | ( ~n14338 & n662 ) ;
  assign n14340 = ( n662 & ~n14339 ) | ( n662 & 1'b0 ) | ( ~n14339 & 1'b0 ) ;
  assign n14341 = ( n530 & ~n555 ) | ( n530 & n14340 ) | ( ~n555 & n14340 ) ;
  assign n14342 = ~n530 & n14341 ;
  assign n14343 = ( n237 & ~n568 ) | ( n237 & n14342 ) | ( ~n568 & n14342 ) ;
  assign n14344 = ~n237 & n14343 ;
  assign n14345 = ~n151 & n14344 ;
  assign n14346 = n3637 | n3644 ;
  assign n14347 = ~n599 & n3652 ;
  assign n14348 = ( n14346 & ~n14347 ) | ( n14346 & 1'b0 ) | ( ~n14347 & 1'b0 ) ;
  assign n14349 = ( n14345 & ~n14059 ) | ( n14345 & n14348 ) | ( ~n14059 & n14348 ) ;
  assign n14350 = ( n14059 & ~n14345 ) | ( n14059 & n14348 ) | ( ~n14345 & n14348 ) ;
  assign n14351 = ( n14349 & ~n14348 ) | ( n14349 & n14350 ) | ( ~n14348 & n14350 ) ;
  assign n14352 = ( n14048 & n14067 ) | ( n14048 & n14068 ) | ( n14067 & n14068 ) ;
  assign n14354 = ( n14337 & n14351 ) | ( n14337 & n14352 ) | ( n14351 & n14352 ) ;
  assign n14353 = ( n14351 & ~n14337 ) | ( n14351 & n14352 ) | ( ~n14337 & n14352 ) ;
  assign n14355 = ( n14337 & ~n14354 ) | ( n14337 & n14353 ) | ( ~n14354 & n14353 ) ;
  assign n14359 = n10499 &  n14355 ;
  assign n14360 = ( n14358 & ~n10499 ) | ( n14358 & n14359 ) | ( ~n10499 & n14359 ) ;
  assign n14361 = ( n14071 & ~n14355 ) | ( n14071 & n14078 ) | ( ~n14355 & n14078 ) ;
  assign n14362 = ( n14078 & ~n14071 ) | ( n14078 & n14355 ) | ( ~n14071 & n14355 ) ;
  assign n14363 = ( n14361 & ~n14078 ) | ( n14361 & n14362 ) | ( ~n14078 & n14362 ) ;
  assign n14364 = ( n14360 & ~n10017 ) | ( n14360 & n14363 ) | ( ~n10017 & n14363 ) ;
  assign n14365 = ~n14363 & n14364 ;
  assign n14366 = ( x2 & ~n14360 ) | ( x2 & n14365 ) | ( ~n14360 & n14365 ) ;
  assign n14367 = ( n14360 & ~x2 ) | ( n14360 & n14365 ) | ( ~x2 & n14365 ) ;
  assign n14368 = ( n14366 & ~n14365 ) | ( n14366 & n14367 ) | ( ~n14365 & n14367 ) ;
  assign n14438 = ~n3644 & n11385 ;
  assign n14433 = n3653 | n11161 ;
  assign n14434 = ( n3657 & ~n11164 ) | ( n3657 & 1'b0 ) | ( ~n11164 & 1'b0 ) ;
  assign n14435 = ( n3652 & ~n11166 ) | ( n3652 & 1'b0 ) | ( ~n11166 & 1'b0 ) ;
  assign n14436 = n14434 | n14435 ;
  assign n14437 = ( n14433 & ~n14436 ) | ( n14433 & 1'b0 ) | ( ~n14436 & 1'b0 ) ;
  assign n14439 = ( n3644 & n14438 ) | ( n3644 & n14437 ) | ( n14438 & n14437 ) ;
  assign n14409 = n1381 | n4716 ;
  assign n14410 = ( n1885 & ~n1268 ) | ( n1885 & n14409 ) | ( ~n1268 & n14409 ) ;
  assign n14411 = n1268 | n14410 ;
  assign n14412 = ( n490 & ~n272 ) | ( n490 & n14411 ) | ( ~n272 & n14411 ) ;
  assign n14413 = n272 | n14412 ;
  assign n14414 = ( n123 & ~n191 ) | ( n123 & n14413 ) | ( ~n191 & n14413 ) ;
  assign n14415 = n191 | n14414 ;
  assign n14416 = ( n353 & ~n561 ) | ( n353 & n14415 ) | ( ~n561 & n14415 ) ;
  assign n14417 = n561 | n14416 ;
  assign n14418 = n196 | n14417 ;
  assign n14419 = n2670 | n3244 ;
  assign n14420 = ( n1343 & n3996 ) | ( n1343 & n14419 ) | ( n3996 & n14419 ) ;
  assign n14421 = ( n1343 & ~n14420 ) | ( n1343 & 1'b0 ) | ( ~n14420 & 1'b0 ) ;
  assign n14422 = ( n14418 & ~n14421 ) | ( n14418 & n14295 ) | ( ~n14421 & n14295 ) ;
  assign n14423 = ( n1762 & ~n14422 ) | ( n1762 & n14295 ) | ( ~n14422 & n14295 ) ;
  assign n14424 = ~n1762 & n14423 ;
  assign n14425 = ( n157 & ~n912 ) | ( n157 & n14424 ) | ( ~n912 & n14424 ) ;
  assign n14426 = ~n157 & n14425 ;
  assign n14427 = ( n257 & ~n127 ) | ( n257 & n14426 ) | ( ~n127 & n14426 ) ;
  assign n14428 = ~n257 & n14427 ;
  assign n14429 = ( n222 & ~n14428 ) | ( n222 & n524 ) | ( ~n14428 & n524 ) ;
  assign n14430 = ( n524 & ~n14429 ) | ( n524 & 1'b0 ) | ( ~n14429 & 1'b0 ) ;
  assign n14431 = ( n14430 & ~n405 ) | ( n14430 & n454 ) | ( ~n405 & n454 ) ;
  assign n14432 = ( n14431 & ~n454 ) | ( n14431 & 1'b0 ) | ( ~n454 & 1'b0 ) ;
  assign n14440 = ( n14165 & n14172 ) | ( n14165 & n14173 ) | ( n14172 & n14173 ) ;
  assign n14441 = ( n14439 & ~n14432 ) | ( n14439 & n14440 ) | ( ~n14432 & n14440 ) ;
  assign n14442 = ( n14432 & ~n14439 ) | ( n14432 & n14440 ) | ( ~n14439 & n14440 ) ;
  assign n14443 = ( n14441 & ~n14440 ) | ( n14441 & n14442 ) | ( ~n14440 & n14442 ) ;
  assign n14447 = n11152 | n4430 ;
  assign n14444 = ~n523 & n11158 ;
  assign n14445 = ~n3939 & n11155 ;
  assign n14446 = n14444 | n14445 ;
  assign n14448 = ( n14447 & ~n4430 ) | ( n14447 & n14446 ) | ( ~n4430 & n14446 ) ;
  assign n14449 = ~n601 & n11254 ;
  assign n14450 = n14448 | n14449 ;
  assign n14451 = ( x29 & ~n14450 ) | ( x29 & 1'b0 ) | ( ~n14450 & 1'b0 ) ;
  assign n14452 = ~x29 & n14450 ;
  assign n14453 = n14451 | n14452 ;
  assign n14454 = ( n14176 & n14186 ) | ( n14176 & n14187 ) | ( n14186 & n14187 ) ;
  assign n14455 = ( n14443 & n14453 ) | ( n14443 & n14454 ) | ( n14453 & n14454 ) ;
  assign n14456 = ( n14453 & ~n14443 ) | ( n14453 & n14454 ) | ( ~n14443 & n14454 ) ;
  assign n14457 = ( n14443 & ~n14455 ) | ( n14443 & n14456 ) | ( ~n14455 & n14456 ) ;
  assign n14402 = ~n4962 & n11143 ;
  assign n14399 = n4482 | n11149 ;
  assign n14400 = n4495 | n11146 ;
  assign n14401 = n14399 &  n14400 ;
  assign n14403 = ( n4962 & n14402 ) | ( n4962 & n14401 ) | ( n14402 & n14401 ) ;
  assign n14404 = ( n11542 & ~n4478 ) | ( n11542 & n14403 ) | ( ~n4478 & n14403 ) ;
  assign n14405 = ~n11542 & n14404 ;
  assign n14407 = ( x26 & n14403 ) | ( x26 & n14405 ) | ( n14403 & n14405 ) ;
  assign n14406 = ( x26 & ~n14405 ) | ( x26 & n14403 ) | ( ~n14405 & n14403 ) ;
  assign n14408 = ( n14405 & ~n14407 ) | ( n14405 & n14406 ) | ( ~n14407 & n14406 ) ;
  assign n14458 = ( n14191 & ~n14457 ) | ( n14191 & n14408 ) | ( ~n14457 & n14408 ) ;
  assign n14459 = ( n14408 & ~n14191 ) | ( n14408 & n14457 ) | ( ~n14191 & n14457 ) ;
  assign n14460 = ( n14458 & ~n14408 ) | ( n14458 & n14459 ) | ( ~n14408 & n14459 ) ;
  assign n14471 = ( n14193 & n14203 ) | ( n14193 & n14204 ) | ( n14203 & n14204 ) ;
  assign n14464 = n11134 | n5135 ;
  assign n14461 = n5010 | n11140 ;
  assign n14462 = n5067 | n11137 ;
  assign n14463 = n14461 &  n14462 ;
  assign n14465 = ( n5135 & ~n14464 ) | ( n5135 & n14463 ) | ( ~n14464 & n14463 ) ;
  assign n14466 = ~n5012 & n11242 ;
  assign n14467 = ( n14465 & ~n14466 ) | ( n14465 & 1'b0 ) | ( ~n14466 & 1'b0 ) ;
  assign n14468 = x23 &  n14467 ;
  assign n14469 = x23 | n14467 ;
  assign n14470 = ~n14468 & n14469 ;
  assign n14472 = ( n14460 & ~n14471 ) | ( n14460 & n14470 ) | ( ~n14471 & n14470 ) ;
  assign n14473 = ( n14460 & ~n14470 ) | ( n14460 & n14471 ) | ( ~n14470 & n14471 ) ;
  assign n14474 = ( n14472 & ~n14460 ) | ( n14472 & n14473 ) | ( ~n14460 & n14473 ) ;
  assign n14392 = n5837 | n11125 ;
  assign n14389 = ( n5339 & ~n11131 ) | ( n5339 & 1'b0 ) | ( ~n11131 & 1'b0 ) ;
  assign n14390 = n5761 | n11128 ;
  assign n14391 = ~n14389 & n14390 ;
  assign n14393 = ( n5837 & ~n14392 ) | ( n5837 & n14391 ) | ( ~n14392 & n14391 ) ;
  assign n14394 = ( n5341 & ~n14393 ) | ( n5341 & n11859 ) | ( ~n14393 & n11859 ) ;
  assign n14395 = ( n11859 & ~n14394 ) | ( n11859 & 1'b0 ) | ( ~n14394 & 1'b0 ) ;
  assign n14397 = ( x20 & n14393 ) | ( x20 & n14395 ) | ( n14393 & n14395 ) ;
  assign n14396 = ( x20 & ~n14395 ) | ( x20 & n14393 ) | ( ~n14395 & n14393 ) ;
  assign n14398 = ( n14395 & ~n14397 ) | ( n14395 & n14396 ) | ( ~n14397 & n14396 ) ;
  assign n14475 = ( n14208 & ~n14474 ) | ( n14208 & n14398 ) | ( ~n14474 & n14398 ) ;
  assign n14476 = ( n14398 & ~n14208 ) | ( n14398 & n14474 ) | ( ~n14208 & n14474 ) ;
  assign n14477 = ( n14475 & ~n14398 ) | ( n14475 & n14476 ) | ( ~n14398 & n14476 ) ;
  assign n14488 = ( n14210 & n14220 ) | ( n14210 & n14221 ) | ( n14220 & n14221 ) ;
  assign n14481 = n11116 | n6395 ;
  assign n14478 = n5970 | n11122 ;
  assign n14479 = ~n6170 & n11119 ;
  assign n14480 = ( n14478 & ~n14479 ) | ( n14478 & 1'b0 ) | ( ~n14479 & 1'b0 ) ;
  assign n14482 = ( n6395 & ~n14481 ) | ( n6395 & n14480 ) | ( ~n14481 & n14480 ) ;
  assign n14483 = n5972 | n11230 ;
  assign n14484 = n14482 &  n14483 ;
  assign n14485 = x17 &  n14484 ;
  assign n14486 = x17 | n14484 ;
  assign n14487 = ~n14485 & n14486 ;
  assign n14489 = ( n14477 & ~n14488 ) | ( n14477 & n14487 ) | ( ~n14488 & n14487 ) ;
  assign n14490 = ( n14477 & ~n14487 ) | ( n14477 & n14488 ) | ( ~n14487 & n14488 ) ;
  assign n14491 = ( n14489 & ~n14477 ) | ( n14489 & n14490 ) | ( ~n14477 & n14490 ) ;
  assign n14382 = n11107 | n7097 ;
  assign n14379 = n6530 | n11113 ;
  assign n14380 = n6983 | n11110 ;
  assign n14381 = n14379 &  n14380 ;
  assign n14383 = ( n7097 & ~n14382 ) | ( n7097 & n14381 ) | ( ~n14382 & n14381 ) ;
  assign n14384 = ( n6532 & ~n14383 ) | ( n6532 & n12340 ) | ( ~n14383 & n12340 ) ;
  assign n14385 = ( n12340 & ~n14384 ) | ( n12340 & 1'b0 ) | ( ~n14384 & 1'b0 ) ;
  assign n14386 = ( x14 & ~n14383 ) | ( x14 & n14385 ) | ( ~n14383 & n14385 ) ;
  assign n14387 = ( n14383 & ~x14 ) | ( n14383 & n14385 ) | ( ~x14 & n14385 ) ;
  assign n14388 = ( n14386 & ~n14385 ) | ( n14386 & n14387 ) | ( ~n14385 & n14387 ) ;
  assign n14492 = ( n14225 & ~n14491 ) | ( n14225 & n14388 ) | ( ~n14491 & n14388 ) ;
  assign n14493 = ( n14388 & ~n14225 ) | ( n14388 & n14491 ) | ( ~n14225 & n14491 ) ;
  assign n14494 = ( n14492 & ~n14388 ) | ( n14492 & n14493 ) | ( ~n14388 & n14493 ) ;
  assign n14505 = ( n14227 & n14237 ) | ( n14227 & n14238 ) | ( n14237 & n14238 ) ;
  assign n14495 = ( n7253 & ~n11104 ) | ( n7253 & 1'b0 ) | ( ~n11104 & 1'b0 ) ;
  assign n14496 = n7518 | n11101 ;
  assign n14497 = ~n14495 & n14496 ;
  assign n14498 = ~n7783 & n11098 ;
  assign n14499 = ( n7783 & n14497 ) | ( n7783 & n14498 ) | ( n14497 & n14498 ) ;
  assign n14500 = n7255 | n11218 ;
  assign n14501 = n14499 &  n14500 ;
  assign n14502 = x11 &  n14501 ;
  assign n14503 = x11 | n14501 ;
  assign n14504 = ~n14502 & n14503 ;
  assign n14506 = ( n14494 & ~n14505 ) | ( n14494 & n14504 ) | ( ~n14505 & n14504 ) ;
  assign n14507 = ( n14494 & ~n14504 ) | ( n14494 & n14505 ) | ( ~n14504 & n14505 ) ;
  assign n14508 = ( n14506 & ~n14494 ) | ( n14506 & n14507 ) | ( ~n14494 & n14507 ) ;
  assign n14372 = ~n8764 & n11091 ;
  assign n14369 = ( n8105 & ~n11095 ) | ( n8105 & 1'b0 ) | ( ~n11095 & 1'b0 ) ;
  assign n14370 = n8429 | n11093 ;
  assign n14371 = ~n14369 & n14370 ;
  assign n14373 = ( n8764 & n14372 ) | ( n8764 & n14371 ) | ( n14372 & n14371 ) ;
  assign n14374 = ( n12984 & ~n8107 ) | ( n12984 & n14373 ) | ( ~n8107 & n14373 ) ;
  assign n14375 = ~n12984 & n14374 ;
  assign n14376 = ( x8 & ~n14373 ) | ( x8 & n14375 ) | ( ~n14373 & n14375 ) ;
  assign n14377 = ( n14373 & ~x8 ) | ( n14373 & n14375 ) | ( ~x8 & n14375 ) ;
  assign n14378 = ( n14376 & ~n14375 ) | ( n14376 & n14377 ) | ( ~n14375 & n14377 ) ;
  assign n14509 = ( n14242 & ~n14508 ) | ( n14242 & n14378 ) | ( ~n14508 & n14378 ) ;
  assign n14510 = ( n14378 & ~n14242 ) | ( n14378 & n14508 ) | ( ~n14242 & n14508 ) ;
  assign n14511 = ( n14509 & ~n14378 ) | ( n14509 & n14510 ) | ( ~n14378 & n14510 ) ;
  assign n14522 = ( n14244 & n14254 ) | ( n14244 & n14255 ) | ( n14254 & n14255 ) ;
  assign n14515 = ~n9997 & n11078 ;
  assign n14512 = n9160 | n11081 ;
  assign n14513 = n9558 | n11085 ;
  assign n14514 = n14512 &  n14513 ;
  assign n14516 = ( n9997 & n14515 ) | ( n9997 & n14514 ) | ( n14515 & n14514 ) ;
  assign n14517 = n9155 | n11206 ;
  assign n14518 = n14516 &  n14517 ;
  assign n14519 = x5 &  n14518 ;
  assign n14520 = x5 | n14518 ;
  assign n14521 = ~n14519 & n14520 ;
  assign n14523 = ( n14511 & ~n14522 ) | ( n14511 & n14521 ) | ( ~n14522 & n14521 ) ;
  assign n14524 = ( n14511 & ~n14521 ) | ( n14511 & n14522 ) | ( ~n14521 & n14522 ) ;
  assign n14525 = ( n14523 & ~n14511 ) | ( n14523 & n14524 ) | ( ~n14511 & n14524 ) ;
  assign n14526 = ( n14259 & ~n14525 ) | ( n14259 & n14368 ) | ( ~n14525 & n14368 ) ;
  assign n14527 = ( n14368 & ~n14259 ) | ( n14368 & n14525 ) | ( ~n14259 & n14525 ) ;
  assign n14528 = ( n14368 & ~n14526 ) | ( n14368 & ~n14527 ) | ( ~n14526 & ~n14527 ) ;
  assign n14531 = ( n14261 & n14266 ) | ( n14261 & n14528 ) | ( n14266 & n14528 ) ;
  assign n14530 = ( n14266 & ~n14261 ) | ( n14266 & n14528 ) | ( ~n14261 & n14528 ) ;
  assign n14532 = ( n14261 & ~n14531 ) | ( n14261 & n14530 ) | ( ~n14531 & n14530 ) ;
  assign n14537 = ~n3644 & n14532 ;
  assign n14529 = n3653 | n14528 ;
  assign n14533 = ( n3657 & ~n14261 ) | ( n3657 & 1'b0 ) | ( ~n14261 & 1'b0 ) ;
  assign n14534 = ( n3652 & ~n13998 ) | ( n3652 & 1'b0 ) | ( ~n13998 & 1'b0 ) ;
  assign n14535 = n14533 | n14534 ;
  assign n14536 = ( n14529 & ~n14535 ) | ( n14529 & 1'b0 ) | ( ~n14535 & 1'b0 ) ;
  assign n14538 = ( n3644 & n14537 ) | ( n3644 & n14536 ) | ( n14537 & n14536 ) ;
  assign n14539 = ( n14274 & n14336 ) | ( n14274 & n14538 ) | ( n14336 & n14538 ) ;
  assign n14608 = ~n523 & n11155 ;
  assign n14609 = ~n3939 & n11152 ;
  assign n14610 = n14608 | n14609 ;
  assign n14611 = ~n4430 & n11149 ;
  assign n14612 = ( n4430 & ~n14610 ) | ( n4430 & n14611 ) | ( ~n14610 & n14611 ) ;
  assign n14613 = ( n11572 & ~n601 ) | ( n11572 & n14612 ) | ( ~n601 & n14612 ) ;
  assign n14614 = ~n11572 & n14613 ;
  assign n14616 = ( x29 & n14612 ) | ( x29 & n14614 ) | ( n14612 & n14614 ) ;
  assign n14615 = ( x29 & ~n14614 ) | ( x29 & n14612 ) | ( ~n14614 & n14612 ) ;
  assign n14617 = ( n14614 & ~n14616 ) | ( n14614 & n14615 ) | ( ~n14616 & n14615 ) ;
  assign n14667 = ( n14432 & n14439 ) | ( n14432 & n14440 ) | ( n14439 & n14440 ) ;
  assign n14618 = n527 | n761 ;
  assign n14619 = n561 | n14618 ;
  assign n14620 = n3042 | n14619 ;
  assign n14621 = ( n5599 & ~n768 ) | ( n5599 & n14620 ) | ( ~n768 & n14620 ) ;
  assign n14622 = n768 | n14621 ;
  assign n14623 = ( n743 & ~n14622 ) | ( n743 & n3681 ) | ( ~n14622 & n3681 ) ;
  assign n14624 = ( n14623 & ~n743 ) | ( n14623 & 1'b0 ) | ( ~n743 & 1'b0 ) ;
  assign n14625 = ( n947 & ~n654 ) | ( n947 & n14624 ) | ( ~n654 & n14624 ) ;
  assign n14626 = ~n947 & n14625 ;
  assign n14627 = ( n477 & ~n14626 ) | ( n477 & n525 ) | ( ~n14626 & n525 ) ;
  assign n14628 = ( n525 & ~n14627 ) | ( n525 & 1'b0 ) | ( ~n14627 & 1'b0 ) ;
  assign n14629 = ( n787 & ~n568 ) | ( n787 & n14628 ) | ( ~n568 & n14628 ) ;
  assign n14630 = ~n787 & n14629 ;
  assign n14631 = ( n93 & ~n166 ) | ( n93 & n14630 ) | ( ~n166 & n14630 ) ;
  assign n14632 = ~n93 & n14631 ;
  assign n14641 = n270 | n3827 ;
  assign n14642 = n664 | n14641 ;
  assign n14643 = n2210 | n3464 ;
  assign n14644 = ( n14642 & ~n6630 ) | ( n14642 & n14643 ) | ( ~n6630 & n14643 ) ;
  assign n14645 = n6630 | n14644 ;
  assign n14633 = n1009 | n4344 ;
  assign n14634 = ( n888 & ~n14633 ) | ( n888 & n1991 ) | ( ~n14633 & n1991 ) ;
  assign n14635 = ~n1991 & n14634 ;
  assign n14636 = ( n425 & ~n2687 ) | ( n425 & n14635 ) | ( ~n2687 & n14635 ) ;
  assign n14637 = ~n425 & n14636 ;
  assign n14638 = ( n214 & ~n194 ) | ( n214 & n14637 ) | ( ~n194 & n14637 ) ;
  assign n14639 = ~n214 & n14638 ;
  assign n14640 = ~n556 & n14639 ;
  assign n14646 = ( n727 & ~n14645 ) | ( n727 & n14640 ) | ( ~n14645 & n14640 ) ;
  assign n14647 = ~n727 & n14646 ;
  assign n14648 = ( n2840 & n14632 ) | ( n2840 & n14647 ) | ( n14632 & n14647 ) ;
  assign n14649 = ~n2840 & n14648 ;
  assign n14650 = ( n2082 & ~n865 ) | ( n2082 & n14649 ) | ( ~n865 & n14649 ) ;
  assign n14651 = ~n2082 & n14650 ;
  assign n14652 = ( n402 & ~n14651 ) | ( n402 & n674 ) | ( ~n14651 & n674 ) ;
  assign n14653 = ( n624 & ~n402 ) | ( n624 & n14652 ) | ( ~n402 & n14652 ) ;
  assign n14654 = ( n624 & ~n14653 ) | ( n624 & 1'b0 ) | ( ~n14653 & 1'b0 ) ;
  assign n14655 = ( n233 & ~n14654 ) | ( n233 & n786 ) | ( ~n14654 & n786 ) ;
  assign n14656 = ( n786 & ~n14655 ) | ( n786 & 1'b0 ) | ( ~n14655 & 1'b0 ) ;
  assign n14657 = ( n571 & ~n492 ) | ( n571 & n14656 ) | ( ~n492 & n14656 ) ;
  assign n14658 = ~n571 & n14657 ;
  assign n14659 = ~n630 & n14658 ;
  assign n14660 = ~n3653 & n11158 ;
  assign n14661 = ( n3657 & ~n11161 ) | ( n3657 & 1'b0 ) | ( ~n11161 & 1'b0 ) ;
  assign n14662 = ( n3652 & ~n11164 ) | ( n3652 & 1'b0 ) | ( ~n11164 & 1'b0 ) ;
  assign n14663 = n14661 | n14662 ;
  assign n14664 = n14660 | n14663 ;
  assign n14665 = n3644 | n11463 ;
  assign n14666 = ( n14664 & ~n3644 ) | ( n14664 & n14665 ) | ( ~n3644 & n14665 ) ;
  assign n14669 = ( n14659 & n14666 ) | ( n14659 & n14667 ) | ( n14666 & n14667 ) ;
  assign n14668 = ( n14659 & ~n14667 ) | ( n14659 & n14666 ) | ( ~n14667 & n14666 ) ;
  assign n14670 = ( n14667 & ~n14669 ) | ( n14667 & n14668 ) | ( ~n14669 & n14668 ) ;
  assign n14671 = ( n14443 & ~n14453 ) | ( n14443 & n14454 ) | ( ~n14453 & n14454 ) ;
  assign n14672 = ( n14617 & n14670 ) | ( n14617 & n14671 ) | ( n14670 & n14671 ) ;
  assign n14673 = ( n14670 & ~n14617 ) | ( n14670 & n14671 ) | ( ~n14617 & n14671 ) ;
  assign n14674 = ( n14617 & ~n14672 ) | ( n14617 & n14673 ) | ( ~n14672 & n14673 ) ;
  assign n14601 = ~n4962 & n11140 ;
  assign n14598 = n4482 | n11146 ;
  assign n14599 = n4495 | n11143 ;
  assign n14600 = n14598 &  n14599 ;
  assign n14602 = ( n4962 & n14601 ) | ( n4962 & n14600 ) | ( n14601 & n14600 ) ;
  assign n14603 = ( n11699 & ~n4478 ) | ( n11699 & n14602 ) | ( ~n4478 & n14602 ) ;
  assign n14604 = ~n11699 & n14603 ;
  assign n14605 = ( x26 & ~n14602 ) | ( x26 & n14604 ) | ( ~n14602 & n14604 ) ;
  assign n14606 = ( n14602 & ~x26 ) | ( n14602 & n14604 ) | ( ~x26 & n14604 ) ;
  assign n14607 = ( n14605 & ~n14604 ) | ( n14605 & n14606 ) | ( ~n14604 & n14606 ) ;
  assign n14675 = ( n14458 & ~n14674 ) | ( n14458 & n14607 ) | ( ~n14674 & n14607 ) ;
  assign n14676 = ( n14607 & ~n14458 ) | ( n14607 & n14674 ) | ( ~n14458 & n14674 ) ;
  assign n14677 = ( n14675 & ~n14607 ) | ( n14675 & n14676 ) | ( ~n14607 & n14676 ) ;
  assign n14688 = ( n14470 & ~n14460 ) | ( n14470 & n14471 ) | ( ~n14460 & n14471 ) ;
  assign n14681 = ~n5135 & n11131 ;
  assign n14678 = n5010 | n11137 ;
  assign n14679 = ~n5067 & n11134 ;
  assign n14680 = ( n14678 & ~n14679 ) | ( n14678 & 1'b0 ) | ( ~n14679 & 1'b0 ) ;
  assign n14682 = ( n5135 & n14681 ) | ( n5135 & n14680 ) | ( n14681 & n14680 ) ;
  assign n14683 = ~n5012 & n11888 ;
  assign n14684 = ( n14682 & ~n14683 ) | ( n14682 & 1'b0 ) | ( ~n14683 & 1'b0 ) ;
  assign n14685 = x23 &  n14684 ;
  assign n14686 = x23 | n14684 ;
  assign n14687 = ~n14685 & n14686 ;
  assign n14689 = ( n14677 & ~n14688 ) | ( n14677 & n14687 ) | ( ~n14688 & n14687 ) ;
  assign n14690 = ( n14677 & ~n14687 ) | ( n14677 & n14688 ) | ( ~n14687 & n14688 ) ;
  assign n14691 = ( n14689 & ~n14677 ) | ( n14689 & n14690 ) | ( ~n14677 & n14690 ) ;
  assign n14588 = ( n5339 & ~n11128 ) | ( n5339 & 1'b0 ) | ( ~n11128 & 1'b0 ) ;
  assign n14589 = ~n5761 & n11125 ;
  assign n14590 = n14588 | n14589 ;
  assign n14591 = ~n5837 & n11122 ;
  assign n14592 = ( n5837 & ~n14590 ) | ( n5837 & n14591 ) | ( ~n14590 & n14591 ) ;
  assign n14593 = ( n5341 & ~n14592 ) | ( n5341 & n12100 ) | ( ~n14592 & n12100 ) ;
  assign n14594 = ( n12100 & ~n14593 ) | ( n12100 & 1'b0 ) | ( ~n14593 & 1'b0 ) ;
  assign n14595 = ( x20 & ~n14592 ) | ( x20 & n14594 ) | ( ~n14592 & n14594 ) ;
  assign n14596 = ( n14592 & ~x20 ) | ( n14592 & n14594 ) | ( ~x20 & n14594 ) ;
  assign n14597 = ( n14595 & ~n14594 ) | ( n14595 & n14596 ) | ( ~n14594 & n14596 ) ;
  assign n14692 = ( n14475 & ~n14691 ) | ( n14475 & n14597 ) | ( ~n14691 & n14597 ) ;
  assign n14693 = ( n14597 & ~n14475 ) | ( n14597 & n14691 ) | ( ~n14475 & n14691 ) ;
  assign n14694 = ( n14692 & ~n14597 ) | ( n14692 & n14693 ) | ( ~n14597 & n14693 ) ;
  assign n14705 = ( n14487 & ~n14477 ) | ( n14487 & n14488 ) | ( ~n14477 & n14488 ) ;
  assign n14695 = ~n5970 & n11119 ;
  assign n14696 = ~n6170 & n11116 ;
  assign n14697 = n14695 | n14696 ;
  assign n14698 = ~n6395 & n11113 ;
  assign n14699 = ( n6395 & ~n14697 ) | ( n6395 & n14698 ) | ( ~n14697 & n14698 ) ;
  assign n14700 = n5972 | n12369 ;
  assign n14701 = n14699 &  n14700 ;
  assign n14702 = x17 &  n14701 ;
  assign n14703 = x17 | n14701 ;
  assign n14704 = ~n14702 & n14703 ;
  assign n14706 = ( n14694 & ~n14705 ) | ( n14694 & n14704 ) | ( ~n14705 & n14704 ) ;
  assign n14707 = ( n14694 & ~n14704 ) | ( n14694 & n14705 ) | ( ~n14704 & n14705 ) ;
  assign n14708 = ( n14706 & ~n14694 ) | ( n14706 & n14707 ) | ( ~n14694 & n14707 ) ;
  assign n14581 = ~n7097 & n11104 ;
  assign n14578 = n6530 | n11110 ;
  assign n14579 = ~n6983 & n11107 ;
  assign n14580 = ( n14578 & ~n14579 ) | ( n14578 & 1'b0 ) | ( ~n14579 & 1'b0 ) ;
  assign n14582 = ( n7097 & n14581 ) | ( n7097 & n14580 ) | ( n14581 & n14580 ) ;
  assign n14583 = ( n6532 & ~n14582 ) | ( n6532 & n12662 ) | ( ~n14582 & n12662 ) ;
  assign n14584 = ( n12662 & ~n14583 ) | ( n12662 & 1'b0 ) | ( ~n14583 & 1'b0 ) ;
  assign n14585 = ( x14 & ~n14582 ) | ( x14 & n14584 ) | ( ~n14582 & n14584 ) ;
  assign n14586 = ( n14582 & ~x14 ) | ( n14582 & n14584 ) | ( ~x14 & n14584 ) ;
  assign n14587 = ( n14585 & ~n14584 ) | ( n14585 & n14586 ) | ( ~n14584 & n14586 ) ;
  assign n14709 = ( n14492 & ~n14708 ) | ( n14492 & n14587 ) | ( ~n14708 & n14587 ) ;
  assign n14710 = ( n14587 & ~n14492 ) | ( n14587 & n14708 ) | ( ~n14492 & n14708 ) ;
  assign n14711 = ( n14709 & ~n14587 ) | ( n14709 & n14710 ) | ( ~n14587 & n14710 ) ;
  assign n14722 = ( n14504 & ~n14494 ) | ( n14504 & n14505 ) | ( ~n14494 & n14505 ) ;
  assign n14715 = ~n7783 & n11095 ;
  assign n14712 = ( n7253 & ~n11101 ) | ( n7253 & 1'b0 ) | ( ~n11101 & 1'b0 ) ;
  assign n14713 = n7518 | n11098 ;
  assign n14714 = ~n14712 & n14713 ;
  assign n14716 = ( n7783 & n14715 ) | ( n7783 & n14714 ) | ( n14715 & n14714 ) ;
  assign n14717 = n7255 | n13014 ;
  assign n14718 = n14716 &  n14717 ;
  assign n14719 = x11 &  n14718 ;
  assign n14720 = x11 | n14718 ;
  assign n14721 = ~n14719 & n14720 ;
  assign n14723 = ( n14711 & ~n14722 ) | ( n14711 & n14721 ) | ( ~n14722 & n14721 ) ;
  assign n14724 = ( n14711 & ~n14721 ) | ( n14711 & n14722 ) | ( ~n14721 & n14722 ) ;
  assign n14725 = ( n14723 & ~n14711 ) | ( n14723 & n14724 ) | ( ~n14711 & n14724 ) ;
  assign n14571 = ~n8764 & n11081 ;
  assign n14568 = ( n8105 & ~n11093 ) | ( n8105 & 1'b0 ) | ( ~n11093 & 1'b0 ) ;
  assign n14569 = n8429 | n11091 ;
  assign n14570 = ~n14568 & n14569 ;
  assign n14572 = ( n8764 & n14571 ) | ( n8764 & n14570 ) | ( n14571 & n14570 ) ;
  assign n14573 = ( n13775 & ~n8107 ) | ( n13775 & n14572 ) | ( ~n8107 & n14572 ) ;
  assign n14574 = ~n13775 & n14573 ;
  assign n14576 = ( x8 & n14572 ) | ( x8 & n14574 ) | ( n14572 & n14574 ) ;
  assign n14575 = ( x8 & ~n14574 ) | ( x8 & n14572 ) | ( ~n14574 & n14572 ) ;
  assign n14577 = ( n14574 & ~n14576 ) | ( n14574 & n14575 ) | ( ~n14576 & n14575 ) ;
  assign n14726 = ( n14509 & ~n14725 ) | ( n14509 & n14577 ) | ( ~n14725 & n14577 ) ;
  assign n14727 = ( n14577 & ~n14509 ) | ( n14577 & n14725 ) | ( ~n14509 & n14725 ) ;
  assign n14728 = ( n14726 & ~n14577 ) | ( n14726 & n14727 ) | ( ~n14577 & n14727 ) ;
  assign n14739 = ( n14521 & ~n14511 ) | ( n14521 & n14522 ) | ( ~n14511 & n14522 ) ;
  assign n14732 = ~n9997 & n13836 ;
  assign n14729 = n9160 | n11085 ;
  assign n14730 = n9558 | n11078 ;
  assign n14731 = n14729 &  n14730 ;
  assign n14733 = ( n9997 & n14732 ) | ( n9997 & n14731 ) | ( n14732 & n14731 ) ;
  assign n14734 = n9155 | n13844 ;
  assign n14735 = n14733 &  n14734 ;
  assign n14736 = x5 &  n14735 ;
  assign n14737 = x5 | n14735 ;
  assign n14738 = ~n14736 & n14737 ;
  assign n14740 = ( n14728 & ~n14739 ) | ( n14728 & n14738 ) | ( ~n14739 & n14738 ) ;
  assign n14741 = ( n14728 & ~n14738 ) | ( n14728 & n14739 ) | ( ~n14738 & n14739 ) ;
  assign n14742 = ( n14740 & ~n14728 ) | ( n14740 & n14741 ) | ( ~n14728 & n14741 ) ;
  assign n14550 = ( n14337 & ~n14352 ) | ( n14337 & n14351 ) | ( ~n14352 & n14351 ) ;
  assign n14540 = n913 | n1231 ;
  assign n14541 = ~n541 & n841 ;
  assign n14542 = ( n694 & ~n14540 ) | ( n694 & n14541 ) | ( ~n14540 & n14541 ) ;
  assign n14543 = ~n694 & n14542 ;
  assign n14544 = ( n602 & ~n136 ) | ( n602 & n14543 ) | ( ~n136 & n14543 ) ;
  assign n14545 = ~n602 & n14544 ;
  assign n14546 = ~n529 & n14545 ;
  assign n14547 = n14059 &  n14546 ;
  assign n14548 = n14059 | n14546 ;
  assign n14549 = ~n14547 & n14548 ;
  assign n14552 = ( n14349 & n14549 ) | ( n14349 & n14550 ) | ( n14549 & n14550 ) ;
  assign n14551 = ( n14349 & ~n14550 ) | ( n14349 & n14549 ) | ( ~n14550 & n14549 ) ;
  assign n14553 = ( n14550 & ~n14552 ) | ( n14550 & n14551 ) | ( ~n14552 & n14551 ) ;
  assign n14557 = ~n14553 & n10499 ;
  assign n14554 = n10015 | n14071 ;
  assign n14555 = n10486 | n14355 ;
  assign n14556 = n14554 &  n14555 ;
  assign n14558 = ( n14557 & ~n10499 ) | ( n14557 & n14556 ) | ( ~n10499 & n14556 ) ;
  assign n14559 = ( n14071 & n14078 ) | ( n14071 & n14355 ) | ( n14078 & n14355 ) ;
  assign n14560 = ( n14355 & n14553 ) | ( n14355 & n14559 ) | ( n14553 & n14559 ) ;
  assign n14561 = ( n14355 & ~n14553 ) | ( n14355 & n14559 ) | ( ~n14553 & n14559 ) ;
  assign n14562 = ( n14553 & ~n14560 ) | ( n14553 & n14561 ) | ( ~n14560 & n14561 ) ;
  assign n14563 = ( n10017 & ~n14558 ) | ( n10017 & n14562 ) | ( ~n14558 & n14562 ) ;
  assign n14564 = ( n14562 & ~n14563 ) | ( n14562 & 1'b0 ) | ( ~n14563 & 1'b0 ) ;
  assign n14565 = ( x2 & ~n14558 ) | ( x2 & n14564 ) | ( ~n14558 & n14564 ) ;
  assign n14566 = ( n14558 & ~x2 ) | ( n14558 & n14564 ) | ( ~x2 & n14564 ) ;
  assign n14567 = ( n14565 & ~n14564 ) | ( n14565 & n14566 ) | ( ~n14564 & n14566 ) ;
  assign n14743 = ( n14526 & ~n14742 ) | ( n14526 & n14567 ) | ( ~n14742 & n14567 ) ;
  assign n14744 = ( n14567 & ~n14526 ) | ( n14567 & n14742 ) | ( ~n14526 & n14742 ) ;
  assign n14745 = ( n14743 & ~n14567 ) | ( n14743 & n14744 ) | ( ~n14567 & n14744 ) ;
  assign n14746 = ~n3653 & n14745 ;
  assign n14750 = ( n3657 & ~n14528 ) | ( n3657 & 1'b0 ) | ( ~n14528 & 1'b0 ) ;
  assign n14751 = ( n3652 & ~n14261 ) | ( n3652 & 1'b0 ) | ( ~n14261 & 1'b0 ) ;
  assign n14752 = n14750 | n14751 ;
  assign n14753 = n14746 | n14752 ;
  assign n14747 = ( n14528 & ~n14531 ) | ( n14528 & n14745 ) | ( ~n14531 & n14745 ) ;
  assign n14748 = ( n14528 & ~n14745 ) | ( n14528 & n14531 ) | ( ~n14745 & n14531 ) ;
  assign n14749 = ( n14747 & ~n14528 ) | ( n14747 & n14748 ) | ( ~n14528 & n14748 ) ;
  assign n14754 = n3644 | n14749 ;
  assign n14755 = ( n14753 & ~n3644 ) | ( n14753 & n14754 ) | ( ~n3644 & n14754 ) ;
  assign n14757 = ( n331 & n14539 ) | ( n331 & n14755 ) | ( n14539 & n14755 ) ;
  assign n14756 = ( n14539 & ~n331 ) | ( n14539 & n14755 ) | ( ~n331 & n14755 ) ;
  assign n14758 = ( n331 & ~n14757 ) | ( n331 & n14756 ) | ( ~n14757 & n14756 ) ;
  assign n14759 = n493 | n1494 ;
  assign n14760 = ( n721 & ~n140 ) | ( n721 & n14759 ) | ( ~n140 & n14759 ) ;
  assign n14761 = n140 | n14760 ;
  assign n14762 = n194 | n674 ;
  assign n14763 = n269 | n14762 ;
  assign n14764 = n384 | n711 ;
  assign n14765 = n43 | n14764 ;
  assign n14766 = ( n2594 & n14763 ) | ( n2594 & n14765 ) | ( n14763 & n14765 ) ;
  assign n14767 = ( n2594 & ~n14766 ) | ( n2594 & 1'b0 ) | ( ~n14766 & 1'b0 ) ;
  assign n14768 = ( n3971 & n14761 ) | ( n3971 & n14767 ) | ( n14761 & n14767 ) ;
  assign n14769 = ( n2426 & ~n14768 ) | ( n2426 & n14761 ) | ( ~n14768 & n14761 ) ;
  assign n14770 = ( n2426 & ~n14769 ) | ( n2426 & 1'b0 ) | ( ~n14769 & 1'b0 ) ;
  assign n14771 = ( n3304 & n3496 ) | ( n3304 & n14770 ) | ( n3496 & n14770 ) ;
  assign n14772 = ~n3304 & n14771 ;
  assign n14773 = ( n716 & ~n2702 ) | ( n716 & n14772 ) | ( ~n2702 & n14772 ) ;
  assign n14774 = ~n716 & n14773 ;
  assign n14775 = ( n208 & ~n374 ) | ( n208 & n14774 ) | ( ~n374 & n14774 ) ;
  assign n14776 = ~n208 & n14775 ;
  assign n14777 = ( n230 & ~n58 ) | ( n230 & n14776 ) | ( ~n58 & n14776 ) ;
  assign n14778 = ~n230 & n14777 ;
  assign n14779 = ( n77 & ~n120 ) | ( n77 & n14778 ) | ( ~n120 & n14778 ) ;
  assign n14780 = ~n77 & n14779 ;
  assign n14781 = n2801 | n6772 ;
  assign n14782 = ( n6717 & ~n1284 ) | ( n6717 & n14781 ) | ( ~n1284 & n14781 ) ;
  assign n14783 = n1284 | n14782 ;
  assign n14784 = ( n14418 & ~n14783 ) | ( n14418 & n4014 ) | ( ~n14783 & n4014 ) ;
  assign n14785 = ( n2461 & ~n14418 ) | ( n2461 & n14784 ) | ( ~n14418 & n14784 ) ;
  assign n14786 = ~n2461 & n14785 ;
  assign n14787 = ( n1270 & n14780 ) | ( n1270 & n14786 ) | ( n14780 & n14786 ) ;
  assign n14788 = ~n1270 & n14787 ;
  assign n14789 = ( n1093 & ~n2091 ) | ( n1093 & n14788 ) | ( ~n2091 & n14788 ) ;
  assign n14790 = ( n14789 & ~n1093 ) | ( n14789 & 1'b0 ) | ( ~n1093 & 1'b0 ) ;
  assign n14791 = ( n1824 & ~n218 ) | ( n1824 & n14790 ) | ( ~n218 & n14790 ) ;
  assign n14792 = ~n1824 & n14791 ;
  assign n14793 = ( n335 & ~n793 ) | ( n335 & n14792 ) | ( ~n793 & n14792 ) ;
  assign n14794 = ~n335 & n14793 ;
  assign n14795 = ~n156 & n14794 ;
  assign n14796 = ( n539 & ~n14795 ) | ( n539 & n525 ) | ( ~n14795 & n525 ) ;
  assign n14797 = ( n525 & ~n14796 ) | ( n525 & 1'b0 ) | ( ~n14796 & 1'b0 ) ;
  assign n14798 = ~n281 & n14797 ;
  assign n14799 = ( n14551 & ~n14547 ) | ( n14551 & n14798 ) | ( ~n14547 & n14798 ) ;
  assign n14800 = n14547 | n14799 ;
  assign n14805 = ( n14547 & ~n14798 ) | ( n14547 & n14551 ) | ( ~n14798 & n14551 ) ;
  assign n14806 = n14798 &  n14805 ;
  assign n14807 = ( n14800 & ~n14806 ) | ( n14800 & 1'b0 ) | ( ~n14806 & 1'b0 ) ;
  assign n15290 = ~n14807 & n10499 ;
  assign n15287 = ~n10015 & n14553 ;
  assign n14801 = ( n14547 & n14551 ) | ( n14547 & n14798 ) | ( n14551 & n14798 ) ;
  assign n14802 = ( n14547 & ~n14551 ) | ( n14547 & n14798 ) | ( ~n14551 & n14798 ) ;
  assign n14803 = ( ~n14551 & n14801 ) | ( ~n14551 & ~n14802 ) | ( n14801 & ~n14802 ) ;
  assign n15288 = n10486 | n14803 ;
  assign n15289 = ~n15287 & n15288 ;
  assign n15291 = ( n15290 & ~n10499 ) | ( n15290 & n15289 ) | ( ~n10499 & n15289 ) ;
  assign n14812 = ( n14561 & ~n14553 ) | ( n14561 & n14803 ) | ( ~n14553 & n14803 ) ;
  assign n15292 = ( n14803 & n14807 ) | ( n14803 & n14812 ) | ( n14807 & n14812 ) ;
  assign n15293 = ( n14807 & ~n14803 ) | ( n14807 & n14812 ) | ( ~n14803 & n14812 ) ;
  assign n15294 = ( n14803 & ~n15292 ) | ( n14803 & n15293 ) | ( ~n15292 & n15293 ) ;
  assign n15295 = ( n10017 & ~n15291 ) | ( n10017 & n15294 ) | ( ~n15291 & n15294 ) ;
  assign n15296 = ( n15294 & ~n15295 ) | ( n15294 & 1'b0 ) | ( ~n15295 & 1'b0 ) ;
  assign n15297 = ( x2 & ~n15291 ) | ( x2 & n15296 ) | ( ~n15291 & n15296 ) ;
  assign n15298 = ( n15291 & ~x2 ) | ( n15291 & n15296 ) | ( ~x2 & n15296 ) ;
  assign n15299 = ( n15297 & ~n15296 ) | ( n15297 & n15298 ) | ( ~n15296 & n15298 ) ;
  assign n15257 = ~n9997 & n14355 ;
  assign n15254 = n9160 | n13836 ;
  assign n15255 = n9558 | n14071 ;
  assign n15256 = n15254 &  n15255 ;
  assign n15258 = ( n9997 & n15257 ) | ( n9997 & n15256 ) | ( n15257 & n15256 ) ;
  assign n15259 = n9155 | n14363 ;
  assign n15260 = n15258 &  n15259 ;
  assign n15261 = x5 &  n15260 ;
  assign n15262 = x5 | n15260 ;
  assign n15263 = ~n15261 & n15262 ;
  assign n15269 = ~n9997 & n14071 ;
  assign n15266 = n9160 | n11078 ;
  assign n15267 = n9558 | n13836 ;
  assign n15268 = n15266 &  n15267 ;
  assign n15270 = ( n9997 & n15269 ) | ( n9997 & n15268 ) | ( n15269 & n15268 ) ;
  assign n15271 = n9155 | n14079 ;
  assign n15272 = n15270 &  n15271 ;
  assign n15273 = x5 &  n15272 ;
  assign n15274 = x5 | n15272 ;
  assign n15275 = ~n15273 & n15274 ;
  assign n15232 = ~n8764 & n11085 ;
  assign n15229 = ( n8105 & ~n11091 ) | ( n8105 & 1'b0 ) | ( ~n11091 & 1'b0 ) ;
  assign n15230 = n8429 | n11081 ;
  assign n15231 = ~n15229 & n15230 ;
  assign n15233 = ( n8764 & n15232 ) | ( n8764 & n15231 ) | ( n15232 & n15231 ) ;
  assign n15234 = ( n13377 & ~n8107 ) | ( n13377 & n15233 ) | ( ~n8107 & n15233 ) ;
  assign n15235 = ~n13377 & n15234 ;
  assign n15236 = ( x8 & ~n15233 ) | ( x8 & n15235 ) | ( ~n15233 & n15235 ) ;
  assign n15237 = ( n15233 & ~x8 ) | ( n15233 & n15235 ) | ( ~x8 & n15235 ) ;
  assign n15238 = ( n15236 & ~n15235 ) | ( n15236 & n15237 ) | ( ~n15235 & n15237 ) ;
  assign n15161 = ~n7097 & n11101 ;
  assign n15158 = ~n6530 & n11107 ;
  assign n15159 = n6983 | n11104 ;
  assign n15160 = ~n15158 & n15159 ;
  assign n15162 = ( n7097 & n15161 ) | ( n7097 & n15160 ) | ( n15161 & n15160 ) ;
  assign n15163 = ( n12650 & ~n6532 ) | ( n12650 & n15162 ) | ( ~n6532 & n15162 ) ;
  assign n15164 = ~n12650 & n15163 ;
  assign n15166 = ( x14 & n15162 ) | ( x14 & n15164 ) | ( n15162 & n15164 ) ;
  assign n15165 = ( x14 & ~n15164 ) | ( x14 & n15162 ) | ( ~n15164 & n15162 ) ;
  assign n15167 = ( n15164 & ~n15166 ) | ( n15164 & n15165 ) | ( ~n15166 & n15165 ) ;
  assign n15090 = n5837 | n11119 ;
  assign n15087 = n5339 &  n11125 ;
  assign n15088 = n5761 | n11122 ;
  assign n15089 = ~n15087 & n15088 ;
  assign n15091 = ( n5837 & ~n15090 ) | ( n5837 & n15089 ) | ( ~n15090 & n15089 ) ;
  assign n15092 = ( n5341 & ~n15091 ) | ( n5341 & n12088 ) | ( ~n15091 & n12088 ) ;
  assign n15093 = ( n12088 & ~n15092 ) | ( n12088 & 1'b0 ) | ( ~n15092 & 1'b0 ) ;
  assign n15094 = ( x20 & ~n15091 ) | ( x20 & n15093 ) | ( ~n15091 & n15093 ) ;
  assign n15095 = ( n15091 & ~x20 ) | ( n15091 & n15093 ) | ( ~x20 & n15093 ) ;
  assign n15096 = ( n15094 & ~n15093 ) | ( n15094 & n15095 ) | ( ~n15093 & n15095 ) ;
  assign n15019 = ~n4962 & n11137 ;
  assign n15016 = n4482 | n11143 ;
  assign n15017 = n4495 | n11140 ;
  assign n15018 = n15016 &  n15017 ;
  assign n15020 = ( n4962 & n15019 ) | ( n4962 & n15018 ) | ( n15019 & n15018 ) ;
  assign n15021 = ( n11687 & ~n4478 ) | ( n11687 & n15020 ) | ( ~n4478 & n15020 ) ;
  assign n15022 = ~n11687 & n15021 ;
  assign n15024 = ( x26 & n15020 ) | ( x26 & n15022 ) | ( n15020 & n15022 ) ;
  assign n15023 = ( x26 & ~n15022 ) | ( x26 & n15020 ) | ( ~n15022 & n15020 ) ;
  assign n15025 = ( n15022 & ~n15024 ) | ( n15022 & n15023 ) | ( ~n15024 & n15023 ) ;
  assign n14987 = ~n4430 & n11146 ;
  assign n14984 = ~n523 & n11152 ;
  assign n14985 = n3939 | n11149 ;
  assign n14986 = ~n14984 & n14985 ;
  assign n14988 = ( n4430 & n14987 ) | ( n4430 & n14986 ) | ( n14987 & n14986 ) ;
  assign n14989 = ( n601 & ~n14988 ) | ( n601 & n11554 ) | ( ~n14988 & n11554 ) ;
  assign n14990 = ( n11554 & ~n14989 ) | ( n11554 & 1'b0 ) | ( ~n14989 & 1'b0 ) ;
  assign n14991 = ( x29 & ~n14988 ) | ( x29 & n14990 ) | ( ~n14988 & n14990 ) ;
  assign n14992 = ( n14988 & ~x29 ) | ( n14988 & n14990 ) | ( ~x29 & n14990 ) ;
  assign n14993 = ( n14991 & ~n14990 ) | ( n14991 & n14992 ) | ( ~n14990 & n14992 ) ;
  assign n14956 = ~n3653 & n11155 ;
  assign n14957 = n3657 &  n11158 ;
  assign n14958 = ( n3652 & ~n11161 ) | ( n3652 & 1'b0 ) | ( ~n11161 & 1'b0 ) ;
  assign n14959 = n14957 | n14958 ;
  assign n14960 = n14956 | n14959 ;
  assign n14961 = ~n3644 & n11451 ;
  assign n14962 = ( n3644 & ~n14960 ) | ( n3644 & n14961 ) | ( ~n14960 & n14961 ) ;
  assign n14940 = n1356 | n2206 ;
  assign n14941 = ( n4197 & ~n4397 ) | ( n4197 & n14940 ) | ( ~n4397 & n14940 ) ;
  assign n14942 = n4397 | n14941 ;
  assign n14943 = ( n1070 & ~n4166 ) | ( n1070 & n14942 ) | ( ~n4166 & n14942 ) ;
  assign n14944 = ( n1070 & ~n14943 ) | ( n1070 & 1'b0 ) | ( ~n14943 & 1'b0 ) ;
  assign n14945 = ( n747 & n3681 ) | ( n747 & n14944 ) | ( n3681 & n14944 ) ;
  assign n14946 = ~n747 & n14945 ;
  assign n14947 = ( n2394 & ~n647 ) | ( n2394 & n14946 ) | ( ~n647 & n14946 ) ;
  assign n14948 = ~n2394 & n14947 ;
  assign n14949 = ( n788 & n11341 ) | ( n788 & n14948 ) | ( n11341 & n14948 ) ;
  assign n14950 = ~n788 & n14949 ;
  assign n14951 = ( n241 & ~n216 ) | ( n241 & n14950 ) | ( ~n216 & n14950 ) ;
  assign n14952 = ~n241 & n14951 ;
  assign n14953 = ( n151 & ~n384 ) | ( n151 & n14952 ) | ( ~n384 & n14952 ) ;
  assign n14954 = ~n151 & n14953 ;
  assign n14955 = ~n356 & n14954 ;
  assign n14963 = ( n14659 & ~n14666 ) | ( n14659 & n14667 ) | ( ~n14666 & n14667 ) ;
  assign n14981 = ( n14962 & ~n14955 ) | ( n14962 & n14963 ) | ( ~n14955 & n14963 ) ;
  assign n14982 = ( n14955 & ~n14962 ) | ( n14955 & n14963 ) | ( ~n14962 & n14963 ) ;
  assign n14983 = ( n14981 & ~n14963 ) | ( n14981 & n14982 ) | ( ~n14963 & n14982 ) ;
  assign n14994 = ( n14617 & ~n14670 ) | ( n14617 & n14671 ) | ( ~n14670 & n14671 ) ;
  assign n15013 = ( n14993 & ~n14983 ) | ( n14993 & n14994 ) | ( ~n14983 & n14994 ) ;
  assign n15014 = ( n14983 & ~n14994 ) | ( n14983 & n14993 ) | ( ~n14994 & n14993 ) ;
  assign n15015 = ( n15013 & ~n14993 ) | ( n15013 & n15014 ) | ( ~n14993 & n15014 ) ;
  assign n15026 = ( n14675 & n15015 ) | ( n14675 & n15025 ) | ( n15015 & n15025 ) ;
  assign n15063 = ( n14675 & ~n15025 ) | ( n14675 & n15015 ) | ( ~n15025 & n15015 ) ;
  assign n15064 = ( n15025 & ~n15026 ) | ( n15025 & n15063 ) | ( ~n15026 & n15063 ) ;
  assign n15056 = ~n5135 & n11128 ;
  assign n15053 = ~n5010 & n11134 ;
  assign n15054 = n5067 | n11131 ;
  assign n15055 = ~n15053 & n15054 ;
  assign n15057 = ( n5135 & n15056 ) | ( n5135 & n15055 ) | ( n15056 & n15055 ) ;
  assign n15058 = n5012 | n11871 ;
  assign n15059 = n15057 &  n15058 ;
  assign n15060 = x23 &  n15059 ;
  assign n15061 = x23 | n15059 ;
  assign n15062 = ~n15060 & n15061 ;
  assign n15065 = ( n14687 & ~n14677 ) | ( n14687 & n14688 ) | ( ~n14677 & n14688 ) ;
  assign n15084 = ( n15064 & ~n15062 ) | ( n15064 & n15065 ) | ( ~n15062 & n15065 ) ;
  assign n15085 = ( n15062 & ~n15065 ) | ( n15062 & n15064 ) | ( ~n15065 & n15064 ) ;
  assign n15086 = ( n15084 & ~n15064 ) | ( n15084 & n15085 ) | ( ~n15064 & n15085 ) ;
  assign n15097 = ( n14692 & n15086 ) | ( n14692 & n15096 ) | ( n15086 & n15096 ) ;
  assign n15134 = ( n14692 & ~n15096 ) | ( n14692 & n15086 ) | ( ~n15096 & n15086 ) ;
  assign n15135 = ( n15096 & ~n15097 ) | ( n15096 & n15134 ) | ( ~n15097 & n15134 ) ;
  assign n15127 = ~n6395 & n11110 ;
  assign n15124 = ~n5970 & n11116 ;
  assign n15125 = n6170 | n11113 ;
  assign n15126 = ~n15124 & n15125 ;
  assign n15128 = ( n6395 & n15127 ) | ( n6395 & n15126 ) | ( n15127 & n15126 ) ;
  assign n15129 = ~n5972 & n12352 ;
  assign n15130 = ( n15128 & ~n15129 ) | ( n15128 & 1'b0 ) | ( ~n15129 & 1'b0 ) ;
  assign n15131 = x17 &  n15130 ;
  assign n15132 = x17 | n15130 ;
  assign n15133 = ~n15131 & n15132 ;
  assign n15136 = ( n14704 & ~n14694 ) | ( n14704 & n14705 ) | ( ~n14694 & n14705 ) ;
  assign n15155 = ( n15135 & ~n15133 ) | ( n15135 & n15136 ) | ( ~n15133 & n15136 ) ;
  assign n15156 = ( n15133 & ~n15136 ) | ( n15133 & n15135 ) | ( ~n15136 & n15135 ) ;
  assign n15157 = ( n15155 & ~n15135 ) | ( n15155 & n15156 ) | ( ~n15135 & n15156 ) ;
  assign n15168 = ( n14709 & n15157 ) | ( n14709 & n15167 ) | ( n15157 & n15167 ) ;
  assign n15205 = ( n14709 & ~n15167 ) | ( n14709 & n15157 ) | ( ~n15167 & n15157 ) ;
  assign n15206 = ( n15167 & ~n15168 ) | ( n15167 & n15205 ) | ( ~n15168 & n15205 ) ;
  assign n15195 = ( n7253 & ~n11098 ) | ( n7253 & 1'b0 ) | ( ~n11098 & 1'b0 ) ;
  assign n15196 = n7518 | n11095 ;
  assign n15197 = ~n15195 & n15196 ;
  assign n15198 = ~n7783 & n11093 ;
  assign n15199 = ( n7783 & n15197 ) | ( n7783 & n15198 ) | ( n15197 & n15198 ) ;
  assign n15200 = n7255 | n12997 ;
  assign n15201 = n15199 &  n15200 ;
  assign n15202 = x11 &  n15201 ;
  assign n15203 = x11 | n15201 ;
  assign n15204 = ~n15202 & n15203 ;
  assign n15207 = ( n14721 & ~n14711 ) | ( n14721 & n14722 ) | ( ~n14711 & n14722 ) ;
  assign n15226 = ( n15206 & ~n15204 ) | ( n15206 & n15207 ) | ( ~n15204 & n15207 ) ;
  assign n15227 = ( n15204 & ~n15207 ) | ( n15204 & n15206 ) | ( ~n15207 & n15206 ) ;
  assign n15228 = ( n15226 & ~n15206 ) | ( n15226 & n15227 ) | ( ~n15206 & n15227 ) ;
  assign n15239 = ( n14726 & n15228 ) | ( n14726 & n15238 ) | ( n15228 & n15238 ) ;
  assign n15276 = ( n14726 & ~n15238 ) | ( n14726 & n15228 ) | ( ~n15238 & n15228 ) ;
  assign n15277 = ( n15238 & ~n15239 ) | ( n15238 & n15276 ) | ( ~n15239 & n15276 ) ;
  assign n15278 = ( n14738 & ~n14728 ) | ( n14738 & n14739 ) | ( ~n14728 & n14739 ) ;
  assign n15279 = ( n15275 & n15277 ) | ( n15275 & n15278 ) | ( n15277 & n15278 ) ;
  assign n15219 = ~n8764 & n11078 ;
  assign n15216 = ( n8105 & ~n11081 ) | ( n8105 & 1'b0 ) | ( ~n11081 & 1'b0 ) ;
  assign n15217 = n8429 | n11085 ;
  assign n15218 = ~n15216 & n15217 ;
  assign n15220 = ( n8764 & n15219 ) | ( n8764 & n15218 ) | ( n15219 & n15218 ) ;
  assign n15221 = ( n11206 & ~n8107 ) | ( n11206 & n15220 ) | ( ~n8107 & n15220 ) ;
  assign n15222 = ~n11206 & n15221 ;
  assign n15224 = ( x8 & n15220 ) | ( x8 & n15222 ) | ( n15220 & n15222 ) ;
  assign n15223 = ( x8 & ~n15222 ) | ( x8 & n15220 ) | ( ~n15222 & n15220 ) ;
  assign n15225 = ( n15222 & ~n15224 ) | ( n15222 & n15223 ) | ( ~n15224 & n15223 ) ;
  assign n15186 = ~n7783 & n11091 ;
  assign n15183 = ( n7253 & ~n11095 ) | ( n7253 & 1'b0 ) | ( ~n11095 & 1'b0 ) ;
  assign n15184 = n7518 | n11093 ;
  assign n15185 = ~n15183 & n15184 ;
  assign n15187 = ( n7783 & n15186 ) | ( n7783 & n15185 ) | ( n15186 & n15185 ) ;
  assign n15188 = n7255 | n12984 ;
  assign n15189 = n15187 &  n15188 ;
  assign n15190 = x11 &  n15189 ;
  assign n15191 = x11 | n15189 ;
  assign n15192 = ~n15190 & n15191 ;
  assign n15208 = ( n15204 & n15206 ) | ( n15204 & n15207 ) | ( n15206 & n15207 ) ;
  assign n15148 = ~n7097 & n11098 ;
  assign n15145 = n6530 | n11104 ;
  assign n15146 = n6983 | n11101 ;
  assign n15147 = n15145 &  n15146 ;
  assign n15149 = ( n7097 & n15148 ) | ( n7097 & n15147 ) | ( n15148 & n15147 ) ;
  assign n15150 = ( n11218 & ~n6532 ) | ( n11218 & n15149 ) | ( ~n6532 & n15149 ) ;
  assign n15151 = ~n11218 & n15150 ;
  assign n15153 = ( x14 & n15149 ) | ( x14 & n15151 ) | ( n15149 & n15151 ) ;
  assign n15152 = ( x14 & ~n15151 ) | ( x14 & n15149 ) | ( ~n15151 & n15149 ) ;
  assign n15154 = ( n15151 & ~n15153 ) | ( n15151 & n15152 ) | ( ~n15153 & n15152 ) ;
  assign n15115 = n11107 | n6395 ;
  assign n15112 = n5970 | n11113 ;
  assign n15113 = n6170 | n11110 ;
  assign n15114 = n15112 &  n15113 ;
  assign n15116 = ( n6395 & ~n15115 ) | ( n6395 & n15114 ) | ( ~n15115 & n15114 ) ;
  assign n15117 = ~n5972 & n12340 ;
  assign n15118 = ( n15116 & ~n15117 ) | ( n15116 & 1'b0 ) | ( ~n15117 & 1'b0 ) ;
  assign n15119 = x17 &  n15118 ;
  assign n15120 = x17 | n15118 ;
  assign n15121 = ~n15119 & n15120 ;
  assign n15137 = ( n15133 & n15135 ) | ( n15133 & n15136 ) | ( n15135 & n15136 ) ;
  assign n15077 = n11116 | n5837 ;
  assign n15074 = ( n5339 & ~n11122 ) | ( n5339 & 1'b0 ) | ( ~n11122 & 1'b0 ) ;
  assign n15075 = ~n5761 & n11119 ;
  assign n15076 = n15074 | n15075 ;
  assign n15078 = ( n15077 & ~n5837 ) | ( n15077 & n15076 ) | ( ~n5837 & n15076 ) ;
  assign n15079 = ( n5341 & ~n11230 ) | ( n5341 & n15078 ) | ( ~n11230 & n15078 ) ;
  assign n15080 = n11230 | n15079 ;
  assign n15082 = ( x20 & n15078 ) | ( x20 & n15080 ) | ( n15078 & n15080 ) ;
  assign n15081 = ( x20 & ~n15080 ) | ( x20 & n15078 ) | ( ~n15080 & n15078 ) ;
  assign n15083 = ( n15080 & ~n15082 ) | ( n15080 & n15081 ) | ( ~n15082 & n15081 ) ;
  assign n15041 = n5135 &  n11125 ;
  assign n15042 = n5010 | n11131 ;
  assign n15043 = n5067 | n11128 ;
  assign n15044 = n15042 &  n15043 ;
  assign n15045 = ( n15041 & ~n11125 ) | ( n15041 & n15044 ) | ( ~n11125 & n15044 ) ;
  assign n15046 = ~n5012 & n11859 ;
  assign n15047 = ( n15045 & ~n15046 ) | ( n15045 & 1'b0 ) | ( ~n15046 & 1'b0 ) ;
  assign n15048 = x23 &  n15047 ;
  assign n15049 = x23 | n15047 ;
  assign n15050 = ~n15048 & n15049 ;
  assign n15066 = ( n15062 & n15064 ) | ( n15062 & n15065 ) | ( n15064 & n15065 ) ;
  assign n15006 = n11134 | n4962 ;
  assign n15003 = n4482 | n11140 ;
  assign n15004 = n4495 | n11137 ;
  assign n15005 = n15003 &  n15004 ;
  assign n15007 = ( n4962 & ~n15006 ) | ( n4962 & n15005 ) | ( ~n15006 & n15005 ) ;
  assign n15008 = ( n4478 & ~n15007 ) | ( n4478 & n11242 ) | ( ~n15007 & n11242 ) ;
  assign n15009 = ( n11242 & ~n15008 ) | ( n11242 & 1'b0 ) | ( ~n15008 & 1'b0 ) ;
  assign n15011 = ( x26 & n15007 ) | ( x26 & n15009 ) | ( n15007 & n15009 ) ;
  assign n15010 = ( x26 & ~n15009 ) | ( x26 & n15007 ) | ( ~n15009 & n15007 ) ;
  assign n15012 = ( n15009 & ~n15011 ) | ( n15009 & n15010 ) | ( ~n15011 & n15010 ) ;
  assign n14974 = ~n4430 & n11143 ;
  assign n14971 = n523 | n11149 ;
  assign n14972 = n3939 | n11146 ;
  assign n14973 = n14971 &  n14972 ;
  assign n14975 = ( n4430 & n14974 ) | ( n4430 & n14973 ) | ( n14974 & n14973 ) ;
  assign n14976 = ( n11542 & ~n601 ) | ( n11542 & n14975 ) | ( ~n601 & n14975 ) ;
  assign n14977 = ~n11542 & n14976 ;
  assign n14979 = ( x29 & n14975 ) | ( x29 & n14977 ) | ( n14975 & n14977 ) ;
  assign n14978 = ( x29 & ~n14977 ) | ( x29 & n14975 ) | ( ~n14977 & n14975 ) ;
  assign n14980 = ( n14977 & ~n14979 ) | ( n14977 & n14978 ) | ( ~n14979 & n14978 ) ;
  assign n14938 = n11254 | n3644 ;
  assign n14933 = ~n3653 & n11152 ;
  assign n14934 = n3657 &  n11155 ;
  assign n14935 = n3652 &  n11158 ;
  assign n14936 = n14934 | n14935 ;
  assign n14937 = n14933 | n14936 ;
  assign n14939 = ( n14938 & ~n3644 ) | ( n14938 & n14937 ) | ( ~n3644 & n14937 ) ;
  assign n14895 = n2468 | n3042 ;
  assign n14896 = ( n712 & ~n208 ) | ( n712 & n14895 ) | ( ~n208 & n14895 ) ;
  assign n14897 = n208 | n14896 ;
  assign n14898 = ( n403 & ~n232 ) | ( n403 & n14897 ) | ( ~n232 & n14897 ) ;
  assign n14899 = n232 | n14898 ;
  assign n14900 = n476 | n14899 ;
  assign n14901 = n1546 | n2263 ;
  assign n14902 = ( n4176 & ~n3267 ) | ( n4176 & n14901 ) | ( ~n3267 & n14901 ) ;
  assign n14903 = n3267 | n14902 ;
  assign n14904 = ( n2575 & n3741 ) | ( n2575 & n14903 ) | ( n3741 & n14903 ) ;
  assign n14905 = ( n2575 & ~n14904 ) | ( n2575 & 1'b0 ) | ( ~n14904 & 1'b0 ) ;
  assign n14906 = ( n570 & ~n14900 ) | ( n570 & n14905 ) | ( ~n14900 & n14905 ) ;
  assign n14907 = ( n14906 & ~n570 ) | ( n14906 & 1'b0 ) | ( ~n570 & 1'b0 ) ;
  assign n14908 = ( n765 & ~n14907 ) | ( n765 & n786 ) | ( ~n14907 & n786 ) ;
  assign n14909 = ( n786 & ~n14908 ) | ( n786 & 1'b0 ) | ( ~n14908 & 1'b0 ) ;
  assign n14910 = ( n534 & ~n221 ) | ( n534 & n14909 ) | ( ~n221 & n14909 ) ;
  assign n14911 = ~n534 & n14910 ;
  assign n14912 = ~n618 & n14911 ;
  assign n14913 = ( n277 & ~n2593 ) | ( n277 & n14912 ) | ( ~n2593 & n14912 ) ;
  assign n14914 = ~n277 & n14913 ;
  assign n14915 = ( n224 & ~n460 ) | ( n224 & n14914 ) | ( ~n460 & n14914 ) ;
  assign n14916 = ~n224 & n14915 ;
  assign n14917 = ( n256 & ~n492 ) | ( n256 & n14916 ) | ( ~n492 & n14916 ) ;
  assign n14918 = ~n256 & n14917 ;
  assign n14919 = n740 | n3394 ;
  assign n14920 = ( n2508 & ~n14919 ) | ( n2508 & n2647 ) | ( ~n14919 & n2647 ) ;
  assign n14921 = ~n2508 & n14920 ;
  assign n14922 = ( n3337 & n14918 ) | ( n3337 & n14921 ) | ( n14918 & n14921 ) ;
  assign n14923 = ~n3337 & n14922 ;
  assign n14924 = ( n1883 & ~n2394 ) | ( n1883 & n14923 ) | ( ~n2394 & n14923 ) ;
  assign n14925 = ~n1883 & n14924 ;
  assign n14926 = ( n479 & ~n134 ) | ( n479 & n14925 ) | ( ~n134 & n14925 ) ;
  assign n14927 = ~n479 & n14926 ;
  assign n14928 = ( n678 & ~n797 ) | ( n678 & n14927 ) | ( ~n797 & n14927 ) ;
  assign n14929 = ~n678 & n14928 ;
  assign n14930 = ( n14929 & ~n340 ) | ( n14929 & n454 ) | ( ~n340 & n454 ) ;
  assign n14931 = ( n14930 & ~n454 ) | ( n14930 & 1'b0 ) | ( ~n454 & 1'b0 ) ;
  assign n14932 = ~n358 & n14931 ;
  assign n14964 = ( n14955 & n14962 ) | ( n14955 & n14963 ) | ( n14962 & n14963 ) ;
  assign n14969 = ( n14932 & n14939 ) | ( n14932 & n14964 ) | ( n14939 & n14964 ) ;
  assign n14965 = ( n14932 & ~n14939 ) | ( n14932 & n14964 ) | ( ~n14939 & n14964 ) ;
  assign n14970 = ( n14939 & ~n14969 ) | ( n14939 & n14965 ) | ( ~n14969 & n14965 ) ;
  assign n14995 = ( n14983 & n14993 ) | ( n14983 & n14994 ) | ( n14993 & n14994 ) ;
  assign n15000 = ( n14970 & n14980 ) | ( n14970 & n14995 ) | ( n14980 & n14995 ) ;
  assign n15001 = ( n14970 & ~n14980 ) | ( n14970 & n14995 ) | ( ~n14980 & n14995 ) ;
  assign n15002 = ( n14980 & ~n15000 ) | ( n14980 & n15001 ) | ( ~n15000 & n15001 ) ;
  assign n15027 = ( n15012 & ~n15002 ) | ( n15012 & n15026 ) | ( ~n15002 & n15026 ) ;
  assign n15051 = ( n15002 & ~n15026 ) | ( n15002 & n15012 ) | ( ~n15026 & n15012 ) ;
  assign n15052 = ( n15027 & ~n15012 ) | ( n15027 & n15051 ) | ( ~n15012 & n15051 ) ;
  assign n15071 = ( n15050 & ~n15066 ) | ( n15050 & n15052 ) | ( ~n15066 & n15052 ) ;
  assign n15072 = ( n15052 & ~n15050 ) | ( n15052 & n15066 ) | ( ~n15050 & n15066 ) ;
  assign n15073 = ( n15071 & ~n15052 ) | ( n15071 & n15072 ) | ( ~n15052 & n15072 ) ;
  assign n15098 = ( n15083 & ~n15073 ) | ( n15083 & n15097 ) | ( ~n15073 & n15097 ) ;
  assign n15122 = ( n15073 & ~n15097 ) | ( n15073 & n15083 ) | ( ~n15097 & n15083 ) ;
  assign n15123 = ( n15098 & ~n15083 ) | ( n15098 & n15122 ) | ( ~n15083 & n15122 ) ;
  assign n15142 = ( n15121 & ~n15137 ) | ( n15121 & n15123 ) | ( ~n15137 & n15123 ) ;
  assign n15143 = ( n15123 & ~n15121 ) | ( n15123 & n15137 ) | ( ~n15121 & n15137 ) ;
  assign n15144 = ( n15142 & ~n15123 ) | ( n15142 & n15143 ) | ( ~n15123 & n15143 ) ;
  assign n15169 = ( n15154 & ~n15144 ) | ( n15154 & n15168 ) | ( ~n15144 & n15168 ) ;
  assign n15193 = ( n15144 & ~n15168 ) | ( n15144 & n15154 ) | ( ~n15168 & n15154 ) ;
  assign n15194 = ( n15169 & ~n15154 ) | ( n15169 & n15193 ) | ( ~n15154 & n15193 ) ;
  assign n15213 = ( n15192 & ~n15208 ) | ( n15192 & n15194 ) | ( ~n15208 & n15194 ) ;
  assign n15214 = ( n15194 & ~n15192 ) | ( n15194 & n15208 ) | ( ~n15192 & n15208 ) ;
  assign n15215 = ( n15213 & ~n15194 ) | ( n15213 & n15214 ) | ( ~n15194 & n15214 ) ;
  assign n15240 = ( n15225 & ~n15215 ) | ( n15225 & n15239 ) | ( ~n15215 & n15239 ) ;
  assign n15264 = ( n15215 & ~n15239 ) | ( n15215 & n15225 ) | ( ~n15239 & n15225 ) ;
  assign n15265 = ( n15240 & ~n15225 ) | ( n15240 & n15264 ) | ( ~n15225 & n15264 ) ;
  assign n15284 = ( n15263 & ~n15279 ) | ( n15263 & n15265 ) | ( ~n15279 & n15265 ) ;
  assign n15285 = ( n15265 & ~n15263 ) | ( n15265 & n15279 ) | ( ~n15263 & n15279 ) ;
  assign n15286 = ( n15284 & ~n15265 ) | ( n15284 & n15285 ) | ( ~n15265 & n15285 ) ;
  assign n15300 = ( n15277 & ~n15275 ) | ( n15277 & n15278 ) | ( ~n15275 & n15278 ) ;
  assign n15301 = ( n15275 & ~n15278 ) | ( n15275 & n15277 ) | ( ~n15278 & n15277 ) ;
  assign n15302 = ( n15300 & ~n15277 ) | ( n15300 & n15301 ) | ( ~n15277 & n15301 ) ;
  assign n15308 = ( n14553 & ~n14803 ) | ( n14553 & n14561 ) | ( ~n14803 & n14561 ) ;
  assign n15309 = ( n14553 & ~n14561 ) | ( n14553 & n14803 ) | ( ~n14561 & n14803 ) ;
  assign n15310 = ( n15308 & ~n14553 ) | ( n15308 & n15309 ) | ( ~n14553 & n15309 ) ;
  assign n15303 = n10015 | n14355 ;
  assign n15304 = ~n10486 & n14553 ;
  assign n15305 = ( n15303 & ~n15304 ) | ( n15303 & 1'b0 ) | ( ~n15304 & 1'b0 ) ;
  assign n15306 = n10499 &  n14803 ;
  assign n15307 = ( n15305 & ~n10499 ) | ( n15305 & n15306 ) | ( ~n10499 & n15306 ) ;
  assign n15311 = ( n10017 & ~n15307 ) | ( n10017 & n15310 ) | ( ~n15307 & n15310 ) ;
  assign n15312 = ( n15310 & ~n15311 ) | ( n15310 & 1'b0 ) | ( ~n15311 & 1'b0 ) ;
  assign n15314 = ( x2 & n15307 ) | ( x2 & n15312 ) | ( n15307 & n15312 ) ;
  assign n15313 = ( x2 & ~n15312 ) | ( x2 & n15307 ) | ( ~n15312 & n15307 ) ;
  assign n15315 = ( n15312 & ~n15314 ) | ( n15312 & n15313 ) | ( ~n15314 & n15313 ) ;
  assign n15316 = ( n14743 & n15302 ) | ( n14743 & n15315 ) | ( n15302 & n15315 ) ;
  assign n15317 = ( n15299 & ~n15286 ) | ( n15299 & n15316 ) | ( ~n15286 & n15316 ) ;
  assign n15324 = ( n15286 & ~n15316 ) | ( n15286 & n15299 ) | ( ~n15316 & n15299 ) ;
  assign n15325 = ( n15299 & ~n15317 ) | ( n15299 & ~n15324 ) | ( ~n15317 & ~n15324 ) ;
  assign n15343 = ~n4430 & n15325 ;
  assign n15340 = ~n523 & n14745 ;
  assign n15321 = ( n14743 & ~n15315 ) | ( n14743 & n15302 ) | ( ~n15315 & n15302 ) ;
  assign n15322 = ( n15315 & ~n15316 ) | ( n15315 & n15321 ) | ( ~n15316 & n15321 ) ;
  assign n15341 = n3939 | n15322 ;
  assign n15342 = ~n15340 & n15341 ;
  assign n15344 = ( n4430 & n15343 ) | ( n4430 & n15342 ) | ( n15343 & n15342 ) ;
  assign n15330 = ( n14748 & ~n14745 ) | ( n14748 & n15322 ) | ( ~n14745 & n15322 ) ;
  assign n15331 = ( n15322 & n15325 ) | ( n15322 & n15330 ) | ( n15325 & n15330 ) ;
  assign n15345 = ( n15325 & ~n15322 ) | ( n15325 & n15330 ) | ( ~n15322 & n15330 ) ;
  assign n15346 = ( n15322 & ~n15331 ) | ( n15322 & n15345 ) | ( ~n15331 & n15345 ) ;
  assign n15347 = n601 | n15346 ;
  assign n15348 = n15344 &  n15347 ;
  assign n15349 = x29 &  n15348 ;
  assign n15350 = x29 | n15348 ;
  assign n15351 = ~n15349 & n15350 ;
  assign n15352 = ( n14336 & ~n14274 ) | ( n14336 & n14538 ) | ( ~n14274 & n14538 ) ;
  assign n15353 = ( n14274 & ~n14538 ) | ( n14274 & n14336 ) | ( ~n14538 & n14336 ) ;
  assign n15354 = ( n15352 & ~n14336 ) | ( n15352 & n15353 ) | ( ~n14336 & n15353 ) ;
  assign n15358 = ~n4430 & n15322 ;
  assign n15355 = n523 | n14528 ;
  assign n15356 = ~n3939 & n14745 ;
  assign n15357 = ( n15355 & ~n15356 ) | ( n15355 & 1'b0 ) | ( ~n15356 & 1'b0 ) ;
  assign n15359 = ( n4430 & n15358 ) | ( n4430 & n15357 ) | ( n15358 & n15357 ) ;
  assign n15360 = ( n14745 & n14748 ) | ( n14745 & n15322 ) | ( n14748 & n15322 ) ;
  assign n15361 = ( n14745 & ~n15360 ) | ( n14745 & n15330 ) | ( ~n15360 & n15330 ) ;
  assign n15362 = ~n601 & n15361 ;
  assign n15363 = ( n15359 & ~n15362 ) | ( n15359 & 1'b0 ) | ( ~n15362 & 1'b0 ) ;
  assign n15364 = x29 &  n15363 ;
  assign n15365 = x29 | n15363 ;
  assign n15366 = ~n15364 & n15365 ;
  assign n15367 = ( n14047 & ~n14029 ) | ( n14047 & n14273 ) | ( ~n14029 & n14273 ) ;
  assign n15368 = ( n14029 & ~n14273 ) | ( n14029 & n14047 ) | ( ~n14273 & n14047 ) ;
  assign n15369 = ( n15367 & ~n14047 ) | ( n15367 & n15368 ) | ( ~n14047 & n15368 ) ;
  assign n15373 = n14745 | n4430 ;
  assign n15370 = n523 | n14261 ;
  assign n15371 = n3939 | n14528 ;
  assign n15372 = n15370 &  n15371 ;
  assign n15374 = ( n4430 & ~n15373 ) | ( n4430 & n15372 ) | ( ~n15373 & n15372 ) ;
  assign n15375 = ~n601 & n14749 ;
  assign n15376 = ( n15374 & ~n15375 ) | ( n15374 & 1'b0 ) | ( ~n15375 & 1'b0 ) ;
  assign n15377 = x29 &  n15376 ;
  assign n15378 = x29 | n15376 ;
  assign n15379 = ~n15377 & n15378 ;
  assign n15395 = n13790 | n601 ;
  assign n15392 = n3939 | n13787 ;
  assign n15393 = n4430 | n13785 ;
  assign n15394 = n15392 &  n15393 ;
  assign n15396 = ( n601 & ~n15395 ) | ( n601 & n15394 ) | ( ~n15395 & n15394 ) ;
  assign n15403 = ~n601 & n14001 ;
  assign n15401 = ~n4430 & n13998 ;
  assign n15398 = n523 | n13787 ;
  assign n15399 = n3939 | n13785 ;
  assign n15400 = n15398 &  n15399 ;
  assign n15402 = ( n4430 & n15401 ) | ( n4430 & n15400 ) | ( n15401 & n15400 ) ;
  assign n15404 = ( n601 & n15403 ) | ( n601 & n15402 ) | ( n15403 & n15402 ) ;
  assign n15397 = ( n521 & ~n13787 ) | ( n521 & 1'b0 ) | ( ~n13787 & 1'b0 ) ;
  assign n15405 = ( n15396 & ~n15404 ) | ( n15396 & n15397 ) | ( ~n15404 & n15397 ) ;
  assign n15406 = ( x29 & ~n15396 ) | ( x29 & n15405 ) | ( ~n15396 & n15405 ) ;
  assign n15407 = ( x29 & ~n15406 ) | ( x29 & 1'b0 ) | ( ~n15406 & 1'b0 ) ;
  assign n15385 = ~n4430 & n14261 ;
  assign n15382 = n523 | n13785 ;
  assign n15383 = n3939 | n13998 ;
  assign n15384 = n15382 &  n15383 ;
  assign n15386 = ( n4430 & n15385 ) | ( n4430 & n15384 ) | ( n15385 & n15384 ) ;
  assign n15387 = ( n601 & ~n14267 ) | ( n601 & n15386 ) | ( ~n14267 & n15386 ) ;
  assign n15388 = ~n601 & n15387 ;
  assign n15389 = ( x29 & ~n15386 ) | ( x29 & n15388 ) | ( ~n15386 & n15388 ) ;
  assign n15390 = ( n15386 & ~x29 ) | ( n15386 & n15388 ) | ( ~x29 & n15388 ) ;
  assign n15391 = ( n15389 & ~n15388 ) | ( n15389 & n15390 ) | ( ~n15388 & n15390 ) ;
  assign n15408 = ( n3643 & ~n13787 ) | ( n3643 & 1'b0 ) | ( ~n13787 & 1'b0 ) ;
  assign n15409 = ( n15407 & ~n15391 ) | ( n15407 & n15408 ) | ( ~n15391 & n15408 ) ;
  assign n15416 = ~n4430 & n14528 ;
  assign n15413 = n523 | n13998 ;
  assign n15414 = n3939 | n14261 ;
  assign n15415 = n15413 &  n15414 ;
  assign n15417 = ( n4430 & n15416 ) | ( n4430 & n15415 ) | ( n15416 & n15415 ) ;
  assign n15418 = n601 | n14532 ;
  assign n15419 = n15417 &  n15418 ;
  assign n15420 = x29 &  n15419 ;
  assign n15421 = x29 | n15419 ;
  assign n15422 = ~n15420 & n15421 ;
  assign n15410 = ~n514 & n13795 ;
  assign n15411 = ( n514 & ~n13795 ) | ( n514 & 1'b0 ) | ( ~n13795 & 1'b0 ) ;
  assign n15412 = n15410 | n15411 ;
  assign n15423 = ( n15409 & ~n15422 ) | ( n15409 & n15412 ) | ( ~n15422 & n15412 ) ;
  assign n15380 = ( n13796 & ~n14008 ) | ( n13796 & n14028 ) | ( ~n14008 & n14028 ) ;
  assign n15381 = ( n14008 & ~n14029 ) | ( n14008 & n15380 ) | ( ~n14029 & n15380 ) ;
  assign n15424 = ( n15379 & ~n15423 ) | ( n15379 & n15381 ) | ( ~n15423 & n15381 ) ;
  assign n15425 = ( n15366 & n15369 ) | ( n15366 & n15424 ) | ( n15369 & n15424 ) ;
  assign n15426 = ( n15351 & n15354 ) | ( n15351 & n15425 ) | ( n15354 & n15425 ) ;
  assign n14810 = ~n14800 & n10499 ;
  assign n14804 = n10015 | n14803 ;
  assign n14808 = ~n10486 & n14807 ;
  assign n14809 = ( n14804 & ~n14808 ) | ( n14804 & 1'b0 ) | ( ~n14808 & 1'b0 ) ;
  assign n14811 = ( n14810 & ~n10499 ) | ( n14810 & n14809 ) | ( ~n10499 & n14809 ) ;
  assign n14813 = ( n14803 & ~n14807 ) | ( n14803 & n14812 ) | ( ~n14807 & n14812 ) ;
  assign n14814 = ( n14806 & ~n14813 ) | ( n14806 & 1'b0 ) | ( ~n14813 & 1'b0 ) ;
  assign n14815 = ~n14806 & n14813 ;
  assign n14816 = n14814 | n14815 ;
  assign n14817 = ( n14811 & ~n10017 ) | ( n14811 & n14816 ) | ( ~n10017 & n14816 ) ;
  assign n14818 = ~n14816 & n14817 ;
  assign n14819 = ( x2 & ~n14811 ) | ( x2 & n14818 ) | ( ~n14811 & n14818 ) ;
  assign n14820 = ( n14811 & ~x2 ) | ( n14811 & n14818 ) | ( ~x2 & n14818 ) ;
  assign n14821 = ( n14819 & ~n14818 ) | ( n14819 & n14820 ) | ( ~n14818 & n14820 ) ;
  assign n14825 = ~n8764 & n13836 ;
  assign n14822 = ( n8105 & ~n11085 ) | ( n8105 & 1'b0 ) | ( ~n11085 & 1'b0 ) ;
  assign n14823 = n8429 | n11078 ;
  assign n14824 = ~n14822 & n14823 ;
  assign n14826 = ( n8764 & n14825 ) | ( n8764 & n14824 ) | ( n14825 & n14824 ) ;
  assign n14827 = ( n13844 & ~n8107 ) | ( n13844 & n14826 ) | ( ~n8107 & n14826 ) ;
  assign n14828 = ~n13844 & n14827 ;
  assign n14829 = ( x8 & ~n14826 ) | ( x8 & n14828 ) | ( ~n14826 & n14828 ) ;
  assign n14830 = ( n14826 & ~x8 ) | ( n14826 & n14828 ) | ( ~x8 & n14828 ) ;
  assign n14831 = ( n14829 & ~n14828 ) | ( n14829 & n14830 ) | ( ~n14828 & n14830 ) ;
  assign n14835 = ~n7097 & n11095 ;
  assign n14832 = n6530 | n11101 ;
  assign n14833 = n6983 | n11098 ;
  assign n14834 = n14832 &  n14833 ;
  assign n14836 = ( n7097 & n14835 ) | ( n7097 & n14834 ) | ( n14835 & n14834 ) ;
  assign n14837 = ( n13014 & ~n6532 ) | ( n13014 & n14836 ) | ( ~n6532 & n14836 ) ;
  assign n14838 = ~n13014 & n14837 ;
  assign n14840 = ( x14 & n14836 ) | ( x14 & n14838 ) | ( n14836 & n14838 ) ;
  assign n14839 = ( x14 & ~n14838 ) | ( x14 & n14836 ) | ( ~n14838 & n14836 ) ;
  assign n14841 = ( n14838 & ~n14840 ) | ( n14838 & n14839 ) | ( ~n14840 & n14839 ) ;
  assign n14842 = n5339 &  n11119 ;
  assign n14843 = ~n5761 & n11116 ;
  assign n14844 = n14842 | n14843 ;
  assign n14845 = ~n5837 & n11113 ;
  assign n14846 = ( n5837 & ~n14844 ) | ( n5837 & n14845 ) | ( ~n14844 & n14845 ) ;
  assign n14847 = ( n12369 & ~n5341 ) | ( n12369 & n14846 ) | ( ~n5341 & n14846 ) ;
  assign n14848 = ~n12369 & n14847 ;
  assign n14850 = ( x20 & n14846 ) | ( x20 & n14848 ) | ( n14846 & n14848 ) ;
  assign n14849 = ( x20 & ~n14848 ) | ( x20 & n14846 ) | ( ~n14848 & n14846 ) ;
  assign n14851 = ( n14848 & ~n14850 ) | ( n14848 & n14849 ) | ( ~n14850 & n14849 ) ;
  assign n14855 = ~n4962 & n11131 ;
  assign n14852 = n4482 | n11137 ;
  assign n14853 = ~n4495 & n11134 ;
  assign n14854 = ( n14852 & ~n14853 ) | ( n14852 & 1'b0 ) | ( ~n14853 & 1'b0 ) ;
  assign n14856 = ( n4962 & n14855 ) | ( n4962 & n14854 ) | ( n14855 & n14854 ) ;
  assign n14857 = ( n4478 & ~n14856 ) | ( n4478 & n11888 ) | ( ~n14856 & n11888 ) ;
  assign n14858 = ( n11888 & ~n14857 ) | ( n11888 & 1'b0 ) | ( ~n14857 & 1'b0 ) ;
  assign n14860 = ( x26 & n14856 ) | ( x26 & n14858 ) | ( n14856 & n14858 ) ;
  assign n14859 = ( x26 & ~n14858 ) | ( x26 & n14856 ) | ( ~n14858 & n14856 ) ;
  assign n14861 = ( n14858 & ~n14860 ) | ( n14858 & n14859 ) | ( ~n14860 & n14859 ) ;
  assign n14865 = ~n4430 & n11140 ;
  assign n14862 = n523 | n11146 ;
  assign n14863 = n3939 | n11143 ;
  assign n14864 = n14862 &  n14863 ;
  assign n14866 = ( n4430 & n14865 ) | ( n4430 & n14864 ) | ( n14865 & n14864 ) ;
  assign n14867 = ( n11699 & ~n601 ) | ( n11699 & n14866 ) | ( ~n601 & n14866 ) ;
  assign n14868 = ~n11699 & n14867 ;
  assign n14869 = ( x29 & ~n14866 ) | ( x29 & n14868 ) | ( ~n14866 & n14868 ) ;
  assign n14870 = ( n14866 & ~x29 ) | ( n14866 & n14868 ) | ( ~x29 & n14868 ) ;
  assign n14871 = ( n14869 & ~n14868 ) | ( n14869 & n14870 ) | ( ~n14868 & n14870 ) ;
  assign n14893 = ~n3644 & n11572 ;
  assign n14888 = n3653 | n11149 ;
  assign n14889 = n3657 &  n11152 ;
  assign n14890 = n3652 &  n11155 ;
  assign n14891 = n14889 | n14890 ;
  assign n14892 = ( n14888 & ~n14891 ) | ( n14888 & 1'b0 ) | ( ~n14891 & 1'b0 ) ;
  assign n14894 = ( n3644 & n14893 ) | ( n3644 & n14892 ) | ( n14893 & n14892 ) ;
  assign n14872 = n2036 | n4227 ;
  assign n14873 = ( n377 & ~n3569 ) | ( n377 & n14872 ) | ( ~n3569 & n14872 ) ;
  assign n14874 = n3569 | n14873 ;
  assign n14875 = ( n3227 & ~n14874 ) | ( n3227 & n3692 ) | ( ~n14874 & n3692 ) ;
  assign n14876 = ~n3227 & n14875 ;
  assign n14877 = ( n6241 & n1982 ) | ( n6241 & n14876 ) | ( n1982 & n14876 ) ;
  assign n14878 = ~n1982 & n14877 ;
  assign n14879 = ( n1491 & ~n1650 ) | ( n1491 & n14878 ) | ( ~n1650 & n14878 ) ;
  assign n14880 = ~n1491 & n14879 ;
  assign n14881 = ( n374 & ~n527 ) | ( n374 & n14880 ) | ( ~n527 & n14880 ) ;
  assign n14882 = ~n374 & n14881 ;
  assign n14883 = ( n531 & ~n52 ) | ( n531 & n14882 ) | ( ~n52 & n14882 ) ;
  assign n14884 = ~n531 & n14883 ;
  assign n14885 = ( n459 & ~n151 ) | ( n459 & n14884 ) | ( ~n151 & n14884 ) ;
  assign n14886 = ~n459 & n14885 ;
  assign n14887 = ~n432 & n14886 ;
  assign n14966 = ( n14894 & ~n14887 ) | ( n14894 & n14965 ) | ( ~n14887 & n14965 ) ;
  assign n14967 = ( n14887 & ~n14894 ) | ( n14887 & n14965 ) | ( ~n14894 & n14965 ) ;
  assign n14968 = ( n14966 & ~n14965 ) | ( n14966 & n14967 ) | ( ~n14965 & n14967 ) ;
  assign n14996 = ( n14980 & ~n14970 ) | ( n14980 & n14995 ) | ( ~n14970 & n14995 ) ;
  assign n14997 = ( n14871 & ~n14968 ) | ( n14871 & n14996 ) | ( ~n14968 & n14996 ) ;
  assign n14998 = ( n14871 & ~n14996 ) | ( n14871 & n14968 ) | ( ~n14996 & n14968 ) ;
  assign n14999 = ( n14997 & ~n14871 ) | ( n14997 & n14998 ) | ( ~n14871 & n14998 ) ;
  assign n15028 = ( n14861 & n14999 ) | ( n14861 & n15027 ) | ( n14999 & n15027 ) ;
  assign n15029 = ( n14999 & ~n14861 ) | ( n14999 & n15027 ) | ( ~n14861 & n15027 ) ;
  assign n15030 = ( n14861 & ~n15028 ) | ( n14861 & n15029 ) | ( ~n15028 & n15029 ) ;
  assign n15034 = ~n5135 & n11122 ;
  assign n15031 = n5010 | n11128 ;
  assign n15032 = ~n5067 & n11125 ;
  assign n15033 = ( n15031 & ~n15032 ) | ( n15031 & 1'b0 ) | ( ~n15032 & 1'b0 ) ;
  assign n15035 = ( n5135 & n15034 ) | ( n5135 & n15033 ) | ( n15034 & n15033 ) ;
  assign n15036 = ~n5012 & n12100 ;
  assign n15037 = ( n15035 & ~n15036 ) | ( n15035 & 1'b0 ) | ( ~n15036 & 1'b0 ) ;
  assign n15038 = x23 &  n15037 ;
  assign n15039 = x23 | n15037 ;
  assign n15040 = ~n15038 & n15039 ;
  assign n15067 = ( n15050 & ~n15052 ) | ( n15050 & n15066 ) | ( ~n15052 & n15066 ) ;
  assign n15068 = ( n15030 & ~n15040 ) | ( n15030 & n15067 ) | ( ~n15040 & n15067 ) ;
  assign n15069 = ( n15030 & ~n15067 ) | ( n15030 & n15040 ) | ( ~n15067 & n15040 ) ;
  assign n15070 = ( n15068 & ~n15030 ) | ( n15068 & n15069 ) | ( ~n15030 & n15069 ) ;
  assign n15099 = ( n14851 & n15070 ) | ( n14851 & n15098 ) | ( n15070 & n15098 ) ;
  assign n15100 = ( n15070 & ~n14851 ) | ( n15070 & n15098 ) | ( ~n14851 & n15098 ) ;
  assign n15101 = ( n14851 & ~n15099 ) | ( n14851 & n15100 ) | ( ~n15099 & n15100 ) ;
  assign n15105 = ~n6395 & n11104 ;
  assign n15102 = n5970 | n11110 ;
  assign n15103 = ~n6170 & n11107 ;
  assign n15104 = ( n15102 & ~n15103 ) | ( n15102 & 1'b0 ) | ( ~n15103 & 1'b0 ) ;
  assign n15106 = ( n6395 & n15105 ) | ( n6395 & n15104 ) | ( n15105 & n15104 ) ;
  assign n15107 = ~n5972 & n12662 ;
  assign n15108 = ( n15106 & ~n15107 ) | ( n15106 & 1'b0 ) | ( ~n15107 & 1'b0 ) ;
  assign n15109 = x17 &  n15108 ;
  assign n15110 = x17 | n15108 ;
  assign n15111 = ~n15109 & n15110 ;
  assign n15138 = ( n15121 & ~n15123 ) | ( n15121 & n15137 ) | ( ~n15123 & n15137 ) ;
  assign n15139 = ( n15101 & ~n15111 ) | ( n15101 & n15138 ) | ( ~n15111 & n15138 ) ;
  assign n15140 = ( n15101 & ~n15138 ) | ( n15101 & n15111 ) | ( ~n15138 & n15111 ) ;
  assign n15141 = ( n15139 & ~n15101 ) | ( n15139 & n15140 ) | ( ~n15101 & n15140 ) ;
  assign n15170 = ( n14841 & n15141 ) | ( n14841 & n15169 ) | ( n15141 & n15169 ) ;
  assign n15171 = ( n15141 & ~n14841 ) | ( n15141 & n15169 ) | ( ~n14841 & n15169 ) ;
  assign n15172 = ( n14841 & ~n15170 ) | ( n14841 & n15171 ) | ( ~n15170 & n15171 ) ;
  assign n15176 = ~n7783 & n11081 ;
  assign n15173 = ( n7253 & ~n11093 ) | ( n7253 & 1'b0 ) | ( ~n11093 & 1'b0 ) ;
  assign n15174 = n7518 | n11091 ;
  assign n15175 = ~n15173 & n15174 ;
  assign n15177 = ( n7783 & n15176 ) | ( n7783 & n15175 ) | ( n15176 & n15175 ) ;
  assign n15178 = n7255 | n13775 ;
  assign n15179 = n15177 &  n15178 ;
  assign n15180 = x11 &  n15179 ;
  assign n15181 = x11 | n15179 ;
  assign n15182 = ~n15180 & n15181 ;
  assign n15209 = ( n15192 & ~n15194 ) | ( n15192 & n15208 ) | ( ~n15194 & n15208 ) ;
  assign n15210 = ( n15172 & ~n15182 ) | ( n15172 & n15209 ) | ( ~n15182 & n15209 ) ;
  assign n15211 = ( n15172 & ~n15209 ) | ( n15172 & n15182 ) | ( ~n15209 & n15182 ) ;
  assign n15212 = ( n15210 & ~n15172 ) | ( n15210 & n15211 ) | ( ~n15172 & n15211 ) ;
  assign n15241 = ( n14831 & n15212 ) | ( n14831 & n15240 ) | ( n15212 & n15240 ) ;
  assign n15242 = ( n15212 & ~n14831 ) | ( n15212 & n15240 ) | ( ~n14831 & n15240 ) ;
  assign n15243 = ( n14831 & ~n15241 ) | ( n14831 & n15242 ) | ( ~n15241 & n15242 ) ;
  assign n15247 = n14553 | n9997 ;
  assign n15244 = n9160 | n14071 ;
  assign n15245 = n9558 | n14355 ;
  assign n15246 = n15244 &  n15245 ;
  assign n15248 = ( n9997 & ~n15247 ) | ( n9997 & n15246 ) | ( ~n15247 & n15246 ) ;
  assign n15249 = ~n9155 & n14562 ;
  assign n15250 = ( n15248 & ~n15249 ) | ( n15248 & 1'b0 ) | ( ~n15249 & 1'b0 ) ;
  assign n15251 = x5 &  n15250 ;
  assign n15252 = x5 | n15250 ;
  assign n15253 = ~n15251 & n15252 ;
  assign n15280 = ( n15263 & ~n15265 ) | ( n15263 & n15279 ) | ( ~n15265 & n15279 ) ;
  assign n15281 = ( n15243 & ~n15253 ) | ( n15243 & n15280 ) | ( ~n15253 & n15280 ) ;
  assign n15282 = ( n15243 & ~n15280 ) | ( n15243 & n15253 ) | ( ~n15280 & n15253 ) ;
  assign n15283 = ( n15281 & ~n15243 ) | ( n15281 & n15282 ) | ( ~n15243 & n15282 ) ;
  assign n15318 = ( n14821 & n15283 ) | ( n14821 & n15317 ) | ( n15283 & n15317 ) ;
  assign n15319 = ( n15283 & ~n14821 ) | ( n15283 & n15317 ) | ( ~n14821 & n15317 ) ;
  assign n15320 = ( n14821 & ~n15318 ) | ( n14821 & n15319 ) | ( ~n15318 & n15319 ) ;
  assign n15328 = ~n4430 & n15320 ;
  assign n15323 = n523 | n15322 ;
  assign n15326 = n3939 | n15325 ;
  assign n15327 = n15323 &  n15326 ;
  assign n15329 = ( n4430 & n15328 ) | ( n4430 & n15327 ) | ( n15328 & n15327 ) ;
  assign n15333 = ( n15320 & n15325 ) | ( n15320 & n15331 ) | ( n15325 & n15331 ) ;
  assign n15332 = ( n15320 & ~n15325 ) | ( n15320 & n15331 ) | ( ~n15325 & n15331 ) ;
  assign n15334 = ( n15325 & ~n15333 ) | ( n15325 & n15332 ) | ( ~n15333 & n15332 ) ;
  assign n15335 = n601 | n15334 ;
  assign n15336 = n15329 &  n15335 ;
  assign n15337 = x29 &  n15336 ;
  assign n15338 = x29 | n15336 ;
  assign n15339 = ~n15337 & n15338 ;
  assign n15427 = ( n14758 & ~n15426 ) | ( n14758 & n15339 ) | ( ~n15426 & n15339 ) ;
  assign n15428 = ( n14758 & ~n15339 ) | ( n14758 & n15426 ) | ( ~n15339 & n15426 ) ;
  assign n15429 = ( n15427 & ~n14758 ) | ( n15427 & n15428 ) | ( ~n14758 & n15428 ) ;
  assign n15433 = ~n4962 & n15322 ;
  assign n15430 = n4482 | n14528 ;
  assign n15431 = ~n4495 & n14745 ;
  assign n15432 = ( n15430 & ~n15431 ) | ( n15430 & 1'b0 ) | ( ~n15431 & 1'b0 ) ;
  assign n15434 = ( n4962 & n15433 ) | ( n4962 & n15432 ) | ( n15433 & n15432 ) ;
  assign n15435 = ( n4478 & n15361 ) | ( n4478 & n15434 ) | ( n15361 & n15434 ) ;
  assign n15436 = ~n4478 & n15435 ;
  assign n15437 = ( x26 & ~n15434 ) | ( x26 & n15436 ) | ( ~n15434 & n15436 ) ;
  assign n15438 = ( n15434 & ~x26 ) | ( n15434 & n15436 ) | ( ~x26 & n15436 ) ;
  assign n15439 = ( n15437 & ~n15436 ) | ( n15437 & n15438 ) | ( ~n15436 & n15438 ) ;
  assign n15440 = ( n15391 & ~n15408 ) | ( n15391 & n15407 ) | ( ~n15408 & n15407 ) ;
  assign n15441 = ( n15409 & ~n15407 ) | ( n15409 & n15440 ) | ( ~n15407 & n15440 ) ;
  assign n15445 = n14745 | n4962 ;
  assign n15442 = n4482 | n14261 ;
  assign n15443 = n4495 | n14528 ;
  assign n15444 = n15442 &  n15443 ;
  assign n15446 = ( n4962 & ~n15445 ) | ( n4962 & n15444 ) | ( ~n15445 & n15444 ) ;
  assign n15447 = ( n4478 & n14749 ) | ( n4478 & n15446 ) | ( n14749 & n15446 ) ;
  assign n15448 = ~n4478 & n15447 ;
  assign n15449 = ( x26 & ~n15446 ) | ( x26 & n15448 ) | ( ~n15446 & n15448 ) ;
  assign n15450 = ( n15446 & ~x26 ) | ( n15446 & n15448 ) | ( ~x26 & n15448 ) ;
  assign n15451 = ( n15449 & ~n15448 ) | ( n15449 & n15450 ) | ( ~n15448 & n15450 ) ;
  assign n15452 = ( n15396 & ~x29 ) | ( n15396 & n15397 ) | ( ~x29 & n15397 ) ;
  assign n15453 = ( n15396 & ~n15452 ) | ( n15396 & 1'b0 ) | ( ~n15452 & 1'b0 ) ;
  assign n15454 = ( n15404 & ~x29 ) | ( n15404 & n15453 ) | ( ~x29 & n15453 ) ;
  assign n15455 = ( x29 & ~n15404 ) | ( x29 & n15453 ) | ( ~n15404 & n15453 ) ;
  assign n15456 = ( n15454 & ~n15453 ) | ( n15454 & n15455 ) | ( ~n15453 & n15455 ) ;
  assign n15457 = x29 &  n15397 ;
  assign n15458 = ~n15396 & n15457 ;
  assign n15459 = ( n15396 & ~n15457 ) | ( n15396 & 1'b0 ) | ( ~n15457 & 1'b0 ) ;
  assign n15460 = n15458 | n15459 ;
  assign n15490 = ~n4962 & n14261 ;
  assign n15487 = n4482 | n13785 ;
  assign n15488 = n4495 | n13998 ;
  assign n15489 = n15487 &  n15488 ;
  assign n15491 = ( n4962 & n15490 ) | ( n4962 & n15489 ) | ( n15490 & n15489 ) ;
  assign n15492 = n4478 | n14267 ;
  assign n15493 = n15491 &  n15492 ;
  assign n15494 = x26 &  n15493 ;
  assign n15495 = x26 | n15493 ;
  assign n15496 = ~n15494 & n15495 ;
  assign n15474 = n13790 | n4478 ;
  assign n15471 = n4495 | n13787 ;
  assign n15472 = n4962 | n13785 ;
  assign n15473 = n15471 &  n15472 ;
  assign n15475 = ( n4478 & ~n15474 ) | ( n4478 & n15473 ) | ( ~n15474 & n15473 ) ;
  assign n15482 = ~n4478 & n14001 ;
  assign n15480 = ~n4962 & n13998 ;
  assign n15477 = n4482 | n13787 ;
  assign n15478 = n4495 | n13785 ;
  assign n15479 = n15477 &  n15478 ;
  assign n15481 = ( n4962 & n15480 ) | ( n4962 & n15479 ) | ( n15480 & n15479 ) ;
  assign n15483 = ( n4478 & n15482 ) | ( n4478 & n15481 ) | ( n15482 & n15481 ) ;
  assign n15476 = ( n4474 & ~n13787 ) | ( n4474 & 1'b0 ) | ( ~n13787 & 1'b0 ) ;
  assign n15484 = ( n15475 & ~n15483 ) | ( n15475 & n15476 ) | ( ~n15483 & n15476 ) ;
  assign n15485 = ( x26 & ~n15475 ) | ( x26 & n15484 ) | ( ~n15475 & n15484 ) ;
  assign n15486 = ( x26 & ~n15485 ) | ( x26 & 1'b0 ) | ( ~n15485 & 1'b0 ) ;
  assign n15497 = ( n15397 & ~n15496 ) | ( n15397 & n15486 ) | ( ~n15496 & n15486 ) ;
  assign n15464 = ~n4962 & n14528 ;
  assign n15461 = n4482 | n13998 ;
  assign n15462 = n4495 | n14261 ;
  assign n15463 = n15461 &  n15462 ;
  assign n15465 = ( n4962 & n15464 ) | ( n4962 & n15463 ) | ( n15464 & n15463 ) ;
  assign n15466 = ( n4478 & ~n14532 ) | ( n4478 & n15465 ) | ( ~n14532 & n15465 ) ;
  assign n15467 = ~n4478 & n15466 ;
  assign n15468 = ( x26 & ~n15465 ) | ( x26 & n15467 ) | ( ~n15465 & n15467 ) ;
  assign n15469 = ( n15465 & ~x26 ) | ( n15465 & n15467 ) | ( ~x26 & n15467 ) ;
  assign n15470 = ( n15468 & ~n15467 ) | ( n15468 & n15469 ) | ( ~n15467 & n15469 ) ;
  assign n15498 = ( n15460 & ~n15497 ) | ( n15460 & n15470 ) | ( ~n15497 & n15470 ) ;
  assign n15499 = ( n15451 & n15456 ) | ( n15451 & n15498 ) | ( n15456 & n15498 ) ;
  assign n15500 = ( n15439 & n15441 ) | ( n15439 & n15499 ) | ( n15441 & n15499 ) ;
  assign n15501 = ( n15409 & n15412 ) | ( n15409 & n15422 ) | ( n15412 & n15422 ) ;
  assign n15502 = ( n15409 & ~n15412 ) | ( n15409 & n15422 ) | ( ~n15412 & n15422 ) ;
  assign n15503 = ( n15412 & ~n15501 ) | ( n15412 & n15502 ) | ( ~n15501 & n15502 ) ;
  assign n15509 = ~n4478 & n15346 ;
  assign n15507 = ~n4962 & n15325 ;
  assign n15504 = ~n4482 & n14745 ;
  assign n15505 = n4495 | n15322 ;
  assign n15506 = ~n15504 & n15505 ;
  assign n15508 = ( n4962 & n15507 ) | ( n4962 & n15506 ) | ( n15507 & n15506 ) ;
  assign n15510 = ( n4478 & n15509 ) | ( n4478 & n15508 ) | ( n15509 & n15508 ) ;
  assign n15512 = x26 &  n15510 ;
  assign n15511 = ~x26 & n15510 ;
  assign n15513 = ( x26 & ~n15512 ) | ( x26 & n15511 ) | ( ~n15512 & n15511 ) ;
  assign n15514 = ( n15500 & n15503 ) | ( n15500 & n15513 ) | ( n15503 & n15513 ) ;
  assign n15516 = ( n15379 & n15381 ) | ( n15379 & n15423 ) | ( n15381 & n15423 ) ;
  assign n15515 = ( n15379 & ~n15381 ) | ( n15379 & n15423 ) | ( ~n15381 & n15423 ) ;
  assign n15517 = ( n15381 & ~n15516 ) | ( n15381 & n15515 ) | ( ~n15516 & n15515 ) ;
  assign n15523 = ~n4478 & n15334 ;
  assign n15521 = ~n4962 & n15320 ;
  assign n15518 = n4482 | n15322 ;
  assign n15519 = n4495 | n15325 ;
  assign n15520 = n15518 &  n15519 ;
  assign n15522 = ( n4962 & n15521 ) | ( n4962 & n15520 ) | ( n15521 & n15520 ) ;
  assign n15524 = ( n4478 & n15523 ) | ( n4478 & n15522 ) | ( n15523 & n15522 ) ;
  assign n15526 = x26 &  n15524 ;
  assign n15525 = ~x26 & n15524 ;
  assign n15527 = ( x26 & ~n15526 ) | ( x26 & n15525 ) | ( ~n15526 & n15525 ) ;
  assign n15528 = ( n15514 & ~n15517 ) | ( n15514 & n15527 ) | ( ~n15517 & n15527 ) ;
  assign n15529 = ( n15369 & ~n15366 ) | ( n15369 & n15424 ) | ( ~n15366 & n15424 ) ;
  assign n15530 = ( n15366 & ~n15424 ) | ( n15366 & n15369 ) | ( ~n15424 & n15369 ) ;
  assign n15531 = ( n15529 & ~n15369 ) | ( n15529 & n15530 ) | ( ~n15369 & n15530 ) ;
  assign n15532 = ( n15243 & n15253 ) | ( n15243 & n15280 ) | ( n15253 & n15280 ) ;
  assign n15536 = ~n9997 & n14803 ;
  assign n15533 = n9160 | n14355 ;
  assign n15534 = ~n9558 & n14553 ;
  assign n15535 = ( n15533 & ~n15534 ) | ( n15533 & 1'b0 ) | ( ~n15534 & 1'b0 ) ;
  assign n15537 = ( n9997 & n15536 ) | ( n9997 & n15535 ) | ( n15536 & n15535 ) ;
  assign n15538 = ~n9155 & n15310 ;
  assign n15539 = ( n15537 & ~n15538 ) | ( n15537 & 1'b0 ) | ( ~n15538 & 1'b0 ) ;
  assign n15543 = ~n8764 & n14071 ;
  assign n15540 = ( n8105 & ~n11078 ) | ( n8105 & 1'b0 ) | ( ~n11078 & 1'b0 ) ;
  assign n15541 = n8429 | n13836 ;
  assign n15542 = ~n15540 & n15541 ;
  assign n15544 = ( n8764 & n15543 ) | ( n8764 & n15542 ) | ( n15543 & n15542 ) ;
  assign n15545 = ( n14079 & ~n8107 ) | ( n14079 & n15544 ) | ( ~n8107 & n15544 ) ;
  assign n15546 = ~n14079 & n15545 ;
  assign n15548 = ( x8 & n15544 ) | ( x8 & n15546 ) | ( n15544 & n15546 ) ;
  assign n15547 = ( x8 & ~n15546 ) | ( x8 & n15544 ) | ( ~n15546 & n15544 ) ;
  assign n15549 = ( n15546 & ~n15548 ) | ( n15546 & n15547 ) | ( ~n15548 & n15547 ) ;
  assign n15553 = ~n7097 & n11093 ;
  assign n15550 = n6530 | n11098 ;
  assign n15551 = n6983 | n11095 ;
  assign n15552 = n15550 &  n15551 ;
  assign n15554 = ( n7097 & n15553 ) | ( n7097 & n15552 ) | ( n15553 & n15552 ) ;
  assign n15555 = ( n12997 & ~n6532 ) | ( n12997 & n15554 ) | ( ~n6532 & n15554 ) ;
  assign n15556 = ~n12997 & n15555 ;
  assign n15557 = ( x14 & ~n15554 ) | ( x14 & n15556 ) | ( ~n15554 & n15556 ) ;
  assign n15558 = ( n15554 & ~x14 ) | ( n15554 & n15556 ) | ( ~x14 & n15556 ) ;
  assign n15559 = ( n15557 & ~n15556 ) | ( n15557 & n15558 ) | ( ~n15556 & n15558 ) ;
  assign n15563 = ~n5837 & n11110 ;
  assign n15560 = n5339 &  n11116 ;
  assign n15561 = n5761 | n11113 ;
  assign n15562 = ~n15560 & n15561 ;
  assign n15564 = ( n5837 & n15563 ) | ( n5837 & n15562 ) | ( n15563 & n15562 ) ;
  assign n15565 = ( n5341 & ~n15564 ) | ( n5341 & n12352 ) | ( ~n15564 & n12352 ) ;
  assign n15566 = ( n12352 & ~n15565 ) | ( n12352 & 1'b0 ) | ( ~n15565 & 1'b0 ) ;
  assign n15568 = ( x20 & n15564 ) | ( x20 & n15566 ) | ( n15564 & n15566 ) ;
  assign n15567 = ( x20 & ~n15566 ) | ( x20 & n15564 ) | ( ~n15566 & n15564 ) ;
  assign n15569 = ( n15566 & ~n15568 ) | ( n15566 & n15567 ) | ( ~n15568 & n15567 ) ;
  assign n15573 = ~n4962 & n11128 ;
  assign n15570 = ~n4482 & n11134 ;
  assign n15571 = n4495 | n11131 ;
  assign n15572 = ~n15570 & n15571 ;
  assign n15574 = ( n4962 & n15573 ) | ( n4962 & n15572 ) | ( n15573 & n15572 ) ;
  assign n15575 = ( n11871 & ~n4478 ) | ( n11871 & n15574 ) | ( ~n4478 & n15574 ) ;
  assign n15576 = ~n11871 & n15575 ;
  assign n15577 = ( x26 & ~n15574 ) | ( x26 & n15576 ) | ( ~n15574 & n15576 ) ;
  assign n15578 = ( n15574 & ~x26 ) | ( n15574 & n15576 ) | ( ~x26 & n15576 ) ;
  assign n15579 = ( n15577 & ~n15576 ) | ( n15577 & n15578 ) | ( ~n15576 & n15578 ) ;
  assign n15583 = ~n4430 & n11137 ;
  assign n15580 = n523 | n11143 ;
  assign n15581 = n3939 | n11140 ;
  assign n15582 = n15580 &  n15581 ;
  assign n15584 = ( n4430 & n15583 ) | ( n4430 & n15582 ) | ( n15583 & n15582 ) ;
  assign n15585 = ( n11687 & ~n601 ) | ( n11687 & n15584 ) | ( ~n601 & n15584 ) ;
  assign n15586 = ~n11687 & n15585 ;
  assign n15588 = ( x29 & n15584 ) | ( x29 & n15586 ) | ( n15584 & n15586 ) ;
  assign n15587 = ( x29 & ~n15586 ) | ( x29 & n15584 ) | ( ~n15586 & n15584 ) ;
  assign n15589 = ( n15586 & ~n15588 ) | ( n15586 & n15587 ) | ( ~n15588 & n15587 ) ;
  assign n15621 = n3644 | n11554 ;
  assign n15616 = n3653 | n11146 ;
  assign n15617 = ( n3657 & ~n11149 ) | ( n3657 & 1'b0 ) | ( ~n11149 & 1'b0 ) ;
  assign n15618 = n3652 &  n11152 ;
  assign n15619 = n15617 | n15618 ;
  assign n15620 = ( n15616 & ~n15619 ) | ( n15616 & 1'b0 ) | ( ~n15619 & 1'b0 ) ;
  assign n15622 = ( n3644 & ~n15621 ) | ( n3644 & n15620 ) | ( ~n15621 & n15620 ) ;
  assign n15590 = n243 | n4016 ;
  assign n15591 = ( n382 & n484 ) | ( n382 & n15590 ) | ( n484 & n15590 ) ;
  assign n15592 = ( n484 & ~n15591 ) | ( n484 & 1'b0 ) | ( ~n15591 & 1'b0 ) ;
  assign n15593 = ( n670 & ~n572 ) | ( n670 & n15592 ) | ( ~n572 & n15592 ) ;
  assign n15594 = ~n670 & n15593 ;
  assign n15595 = n208 | n5454 ;
  assign n15596 = ( n187 & ~n231 ) | ( n187 & n15595 ) | ( ~n231 & n15595 ) ;
  assign n15597 = n231 | n15596 ;
  assign n15598 = ( n332 & n644 ) | ( n332 & n15597 ) | ( n644 & n15597 ) ;
  assign n15599 = ( n644 & ~n15598 ) | ( n644 & 1'b0 ) | ( ~n15598 & 1'b0 ) ;
  assign n15600 = n3504 | n4342 ;
  assign n15601 = ( n3527 & ~n3091 ) | ( n3527 & n15600 ) | ( ~n3091 & n15600 ) ;
  assign n15602 = n3091 | n15601 ;
  assign n15603 = ( n463 & ~n1728 ) | ( n463 & n15602 ) | ( ~n1728 & n15602 ) ;
  assign n15604 = n1728 | n15603 ;
  assign n15605 = ( n15594 & ~n15599 ) | ( n15594 & n15604 ) | ( ~n15599 & n15604 ) ;
  assign n15606 = ( n5246 & ~n15594 ) | ( n5246 & n15605 ) | ( ~n15594 & n15605 ) ;
  assign n15607 = ( n5246 & ~n15606 ) | ( n5246 & 1'b0 ) | ( ~n15606 & 1'b0 ) ;
  assign n15608 = ( n1428 & ~n673 ) | ( n1428 & n15607 ) | ( ~n673 & n15607 ) ;
  assign n15609 = ~n1428 & n15608 ;
  assign n15610 = ( n62 & ~n122 ) | ( n62 & n15609 ) | ( ~n122 & n15609 ) ;
  assign n15611 = ~n62 & n15610 ;
  assign n15612 = ( n161 & ~n271 ) | ( n161 & n15611 ) | ( ~n271 & n15611 ) ;
  assign n15613 = ~n161 & n15612 ;
  assign n15614 = ( n151 & ~n627 ) | ( n151 & n15613 ) | ( ~n627 & n15613 ) ;
  assign n15615 = ~n151 & n15614 ;
  assign n15623 = ( n14887 & n14894 ) | ( n14887 & n14965 ) | ( n14894 & n14965 ) ;
  assign n15624 = ( n15622 & ~n15615 ) | ( n15622 & n15623 ) | ( ~n15615 & n15623 ) ;
  assign n15625 = ( n15615 & ~n15622 ) | ( n15615 & n15623 ) | ( ~n15622 & n15623 ) ;
  assign n15626 = ( n15624 & ~n15623 ) | ( n15624 & n15625 ) | ( ~n15623 & n15625 ) ;
  assign n15627 = ( n14871 & n14968 ) | ( n14871 & n14996 ) | ( n14968 & n14996 ) ;
  assign n15628 = ( n15589 & ~n15626 ) | ( n15589 & n15627 ) | ( ~n15626 & n15627 ) ;
  assign n15629 = ( n15589 & ~n15627 ) | ( n15589 & n15626 ) | ( ~n15627 & n15626 ) ;
  assign n15630 = ( n15628 & ~n15589 ) | ( n15628 & n15629 ) | ( ~n15589 & n15629 ) ;
  assign n15631 = ( n15028 & n15579 ) | ( n15028 & n15630 ) | ( n15579 & n15630 ) ;
  assign n15632 = ( n15028 & ~n15579 ) | ( n15028 & n15630 ) | ( ~n15579 & n15630 ) ;
  assign n15633 = ( n15579 & ~n15631 ) | ( n15579 & n15632 ) | ( ~n15631 & n15632 ) ;
  assign n15644 = ( n15030 & n15040 ) | ( n15030 & n15067 ) | ( n15040 & n15067 ) ;
  assign n15637 = n11119 | n5135 ;
  assign n15634 = ~n5010 & n11125 ;
  assign n15635 = n5067 | n11122 ;
  assign n15636 = ~n15634 & n15635 ;
  assign n15638 = ( n5135 & ~n15637 ) | ( n5135 & n15636 ) | ( ~n15637 & n15636 ) ;
  assign n15639 = ~n5012 & n12088 ;
  assign n15640 = ( n15638 & ~n15639 ) | ( n15638 & 1'b0 ) | ( ~n15639 & 1'b0 ) ;
  assign n15641 = x23 &  n15640 ;
  assign n15642 = x23 | n15640 ;
  assign n15643 = ~n15641 & n15642 ;
  assign n15645 = ( n15633 & ~n15644 ) | ( n15633 & n15643 ) | ( ~n15644 & n15643 ) ;
  assign n15646 = ( n15633 & ~n15643 ) | ( n15633 & n15644 ) | ( ~n15643 & n15644 ) ;
  assign n15647 = ( n15645 & ~n15633 ) | ( n15645 & n15646 ) | ( ~n15633 & n15646 ) ;
  assign n15648 = ( n15099 & n15569 ) | ( n15099 & n15647 ) | ( n15569 & n15647 ) ;
  assign n15649 = ( n15099 & ~n15569 ) | ( n15099 & n15647 ) | ( ~n15569 & n15647 ) ;
  assign n15650 = ( n15569 & ~n15648 ) | ( n15569 & n15649 ) | ( ~n15648 & n15649 ) ;
  assign n15661 = ( n15101 & n15111 ) | ( n15101 & n15138 ) | ( n15111 & n15138 ) ;
  assign n15654 = ~n6395 & n11101 ;
  assign n15651 = ~n5970 & n11107 ;
  assign n15652 = n6170 | n11104 ;
  assign n15653 = ~n15651 & n15652 ;
  assign n15655 = ( n6395 & n15654 ) | ( n6395 & n15653 ) | ( n15654 & n15653 ) ;
  assign n15656 = n5972 | n12650 ;
  assign n15657 = n15655 &  n15656 ;
  assign n15658 = x17 &  n15657 ;
  assign n15659 = x17 | n15657 ;
  assign n15660 = ~n15658 & n15659 ;
  assign n15662 = ( n15650 & ~n15661 ) | ( n15650 & n15660 ) | ( ~n15661 & n15660 ) ;
  assign n15663 = ( n15650 & ~n15660 ) | ( n15650 & n15661 ) | ( ~n15660 & n15661 ) ;
  assign n15664 = ( n15662 & ~n15650 ) | ( n15662 & n15663 ) | ( ~n15650 & n15663 ) ;
  assign n15665 = ( n15170 & n15559 ) | ( n15170 & n15664 ) | ( n15559 & n15664 ) ;
  assign n15666 = ( n15170 & ~n15559 ) | ( n15170 & n15664 ) | ( ~n15559 & n15664 ) ;
  assign n15667 = ( n15559 & ~n15665 ) | ( n15559 & n15666 ) | ( ~n15665 & n15666 ) ;
  assign n15678 = ( n15172 & n15182 ) | ( n15172 & n15209 ) | ( n15182 & n15209 ) ;
  assign n15671 = ~n7783 & n11085 ;
  assign n15668 = ( n7253 & ~n11091 ) | ( n7253 & 1'b0 ) | ( ~n11091 & 1'b0 ) ;
  assign n15669 = n7518 | n11081 ;
  assign n15670 = ~n15668 & n15669 ;
  assign n15672 = ( n7783 & n15671 ) | ( n7783 & n15670 ) | ( n15671 & n15670 ) ;
  assign n15673 = n7255 | n13377 ;
  assign n15674 = n15672 &  n15673 ;
  assign n15675 = x11 &  n15674 ;
  assign n15676 = x11 | n15674 ;
  assign n15677 = ~n15675 & n15676 ;
  assign n15679 = ( n15667 & ~n15678 ) | ( n15667 & n15677 ) | ( ~n15678 & n15677 ) ;
  assign n15680 = ( n15667 & ~n15677 ) | ( n15667 & n15678 ) | ( ~n15677 & n15678 ) ;
  assign n15681 = ( n15679 & ~n15667 ) | ( n15679 & n15680 ) | ( ~n15667 & n15680 ) ;
  assign n15682 = ( n15241 & n15549 ) | ( n15241 & n15681 ) | ( n15549 & n15681 ) ;
  assign n15683 = ( n15241 & ~n15549 ) | ( n15241 & n15681 ) | ( ~n15549 & n15681 ) ;
  assign n15684 = ( n15549 & ~n15682 ) | ( n15549 & n15683 ) | ( ~n15682 & n15683 ) ;
  assign n15685 = ( x5 & ~n15539 ) | ( x5 & n15684 ) | ( ~n15539 & n15684 ) ;
  assign n15686 = ( n15539 & ~x5 ) | ( n15539 & n15684 ) | ( ~x5 & n15684 ) ;
  assign n15687 = ( n15685 & ~n15684 ) | ( n15685 & n15686 ) | ( ~n15684 & n15686 ) ;
  assign n15688 = ( n10486 & ~n10499 ) | ( n10486 & 1'b0 ) | ( ~n10499 & 1'b0 ) ;
  assign n15689 = ( n14800 & ~n15688 ) | ( n14800 & 1'b0 ) | ( ~n15688 & 1'b0 ) ;
  assign n15690 = ~n10015 & n14807 ;
  assign n15691 = n15689 | n15690 ;
  assign n15692 = n14807 | n14814 ;
  assign n15693 = ~n10017 & n15692 ;
  assign n15694 = n15691 | n15693 ;
  assign n15695 = ( x2 & ~n15687 ) | ( x2 & n15694 ) | ( ~n15687 & n15694 ) ;
  assign n15696 = ( x2 & ~n15694 ) | ( x2 & n15687 ) | ( ~n15694 & n15687 ) ;
  assign n15697 = ( n15695 & ~x2 ) | ( n15695 & n15696 ) | ( ~x2 & n15696 ) ;
  assign n15698 = ( n15318 & n15532 ) | ( n15318 & n15697 ) | ( n15532 & n15697 ) ;
  assign n15699 = ( n15318 & ~n15532 ) | ( n15318 & n15697 ) | ( ~n15532 & n15697 ) ;
  assign n15700 = ( ~n15532 & n15698 ) | ( ~n15532 & ~n15699 ) | ( n15698 & ~n15699 ) ;
  assign n15707 = ( n15320 & n15333 ) | ( n15320 & n15700 ) | ( n15333 & n15700 ) ;
  assign n15706 = ( n15333 & ~n15320 ) | ( n15333 & n15700 ) | ( ~n15320 & n15700 ) ;
  assign n15708 = ( n15320 & ~n15707 ) | ( n15320 & n15706 ) | ( ~n15707 & n15706 ) ;
  assign n15704 = ~n4962 & n15700 ;
  assign n15701 = n4482 | n15325 ;
  assign n15702 = n4495 | n15320 ;
  assign n15703 = n15701 &  n15702 ;
  assign n15705 = ( n4962 & n15704 ) | ( n4962 & n15703 ) | ( n15704 & n15703 ) ;
  assign n15709 = ( n15705 & ~n4478 ) | ( n15705 & n15708 ) | ( ~n4478 & n15708 ) ;
  assign n15710 = ~n15708 & n15709 ;
  assign n15712 = ( x26 & n15705 ) | ( x26 & n15710 ) | ( n15705 & n15710 ) ;
  assign n15711 = ( x26 & ~n15710 ) | ( x26 & n15705 ) | ( ~n15710 & n15705 ) ;
  assign n15713 = ( n15710 & ~n15712 ) | ( n15710 & n15711 ) | ( ~n15712 & n15711 ) ;
  assign n15714 = ( n15528 & n15531 ) | ( n15528 & n15713 ) | ( n15531 & n15713 ) ;
  assign n15715 = ( n15354 & ~n15351 ) | ( n15354 & n15425 ) | ( ~n15351 & n15425 ) ;
  assign n15716 = ( n15351 & ~n15425 ) | ( n15351 & n15354 ) | ( ~n15425 & n15354 ) ;
  assign n15717 = ( n15715 & ~n15354 ) | ( n15715 & n15716 ) | ( ~n15354 & n15716 ) ;
  assign n15718 = x5 &  n15539 ;
  assign n15719 = x5 | n15539 ;
  assign n15720 = ( n15684 & ~n15718 ) | ( n15684 & n15719 ) | ( ~n15718 & n15719 ) ;
  assign n15722 = ( x2 & n15687 ) | ( x2 & n15694 ) | ( n15687 & n15694 ) ;
  assign n15721 = x2 &  n15694 ;
  assign n15723 = ( n15720 & ~n15722 ) | ( n15720 & n15721 ) | ( ~n15722 & n15721 ) ;
  assign n15724 = ( n15589 & n15626 ) | ( n15589 & n15627 ) | ( n15626 & n15627 ) ;
  assign n15725 = n4962 &  n11125 ;
  assign n15726 = n4482 | n11131 ;
  assign n15727 = n4495 | n11128 ;
  assign n15728 = n15726 &  n15727 ;
  assign n15729 = ( n15725 & ~n11125 ) | ( n15725 & n15728 ) | ( ~n11125 & n15728 ) ;
  assign n15730 = ~n4478 & n11859 ;
  assign n15731 = ( n15729 & ~n15730 ) | ( n15729 & 1'b0 ) | ( ~n15730 & 1'b0 ) ;
  assign n15732 = x26 &  n15731 ;
  assign n15733 = x26 | n15731 ;
  assign n15734 = ~n15732 & n15733 ;
  assign n15735 = ( x2 & ~n14800 ) | ( x2 & 1'b0 ) | ( ~n14800 & 1'b0 ) ;
  assign n15736 = ( x1 & ~x0 ) | ( x1 & x2 ) | ( ~x0 & x2 ) ;
  assign n15737 = x0 | n15736 ;
  assign n15738 = ~x2 & n15737 ;
  assign n15739 = ~n14547 & n14551 ;
  assign n15740 = ( n14547 & ~n14798 ) | ( n14547 & n15739 ) | ( ~n14798 & n15739 ) ;
  assign n15741 = ( n14798 & n15738 ) | ( n14798 & n15740 ) | ( n15738 & n15740 ) ;
  assign n15742 = n15735 | n15741 ;
  assign n15743 = n3644 | n11542 ;
  assign n15744 = ( n3652 & ~n11149 ) | ( n3652 & 1'b0 ) | ( ~n11149 & 1'b0 ) ;
  assign n15745 = ( n3657 & ~n11146 ) | ( n3657 & 1'b0 ) | ( ~n11146 & 1'b0 ) ;
  assign n15746 = n15744 | n15745 ;
  assign n15747 = ~n3653 & n11143 ;
  assign n15748 = ( n3653 & ~n15746 ) | ( n3653 & n15747 ) | ( ~n15746 & n15747 ) ;
  assign n15749 = n15743 &  n15748 ;
  assign n15750 = ( n1130 & ~n1357 ) | ( n1130 & n3552 ) | ( ~n1357 & n3552 ) ;
  assign n15751 = n1357 | n15750 ;
  assign n15752 = ( n2848 & ~n1796 ) | ( n2848 & n15751 ) | ( ~n1796 & n15751 ) ;
  assign n15753 = n1796 | n15752 ;
  assign n15754 = ( n2702 & ~n677 ) | ( n2702 & n15753 ) | ( ~n677 & n15753 ) ;
  assign n15755 = n677 | n15754 ;
  assign n15756 = ( n194 & ~n15755 ) | ( n194 & n344 ) | ( ~n15755 & n344 ) ;
  assign n15757 = ~n194 & n15756 ;
  assign n15758 = ( n735 & ~n274 ) | ( n735 & n15757 ) | ( ~n274 & n15757 ) ;
  assign n15759 = ~n735 & n15758 ;
  assign n15760 = ( n452 & ~n494 ) | ( n452 & n15759 ) | ( ~n494 & n15759 ) ;
  assign n15761 = ( n239 & ~n452 ) | ( n239 & n15760 ) | ( ~n452 & n15760 ) ;
  assign n15762 = ~n239 & n15761 ;
  assign n15763 = ~n236 & n15762 ;
  assign n15764 = ~n213 & n15763 ;
  assign n15765 = n1603 | n2433 ;
  assign n15766 = ( n2625 & ~n15765 ) | ( n2625 & n198 ) | ( ~n15765 & n198 ) ;
  assign n15767 = ( n15766 & ~n2625 ) | ( n15766 & 1'b0 ) | ( ~n2625 & 1'b0 ) ;
  assign n15768 = ~n11301 & n15767 ;
  assign n15769 = ( n11262 & ~n15768 ) | ( n11262 & n14918 ) | ( ~n15768 & n14918 ) ;
  assign n15770 = ( n15764 & ~n14918 ) | ( n15764 & n15769 ) | ( ~n14918 & n15769 ) ;
  assign n15771 = ( n15764 & ~n15770 ) | ( n15764 & 1'b0 ) | ( ~n15770 & 1'b0 ) ;
  assign n15772 = ( n61 & ~n70 ) | ( n61 & n15771 ) | ( ~n70 & n15771 ) ;
  assign n15773 = ~n61 & n15772 ;
  assign n15774 = ( n15773 & ~n722 ) | ( n15773 & n796 ) | ( ~n722 & n796 ) ;
  assign n15775 = ( n15774 & ~n796 ) | ( n15774 & 1'b0 ) | ( ~n796 & 1'b0 ) ;
  assign n15776 = ( n457 & ~n761 ) | ( n457 & n15775 ) | ( ~n761 & n15775 ) ;
  assign n15777 = ~n457 & n15776 ;
  assign n15778 = ( n255 & ~n603 ) | ( n255 & n15777 ) | ( ~n603 & n15777 ) ;
  assign n15779 = ~n255 & n15778 ;
  assign n15780 = ( n15742 & ~n15749 ) | ( n15742 & n15779 ) | ( ~n15749 & n15779 ) ;
  assign n15781 = ( n15749 & ~n15742 ) | ( n15749 & n15779 ) | ( ~n15742 & n15779 ) ;
  assign n15782 = ( n15780 & ~n15779 ) | ( n15780 & n15781 ) | ( ~n15779 & n15781 ) ;
  assign n15788 = n11242 | n601 ;
  assign n15786 = n11134 | n4430 ;
  assign n15783 = n523 | n11140 ;
  assign n15784 = n3939 | n11137 ;
  assign n15785 = n15783 &  n15784 ;
  assign n15787 = ( n4430 & ~n15786 ) | ( n4430 & n15785 ) | ( ~n15786 & n15785 ) ;
  assign n15789 = ( n601 & ~n15788 ) | ( n601 & n15787 ) | ( ~n15788 & n15787 ) ;
  assign n15790 = x29 &  n15789 ;
  assign n15791 = x29 | n15789 ;
  assign n15792 = ~n15790 & n15791 ;
  assign n15793 = ( n15615 & n15622 ) | ( n15615 & n15623 ) | ( n15622 & n15623 ) ;
  assign n15795 = ( n15782 & n15792 ) | ( n15782 & n15793 ) | ( n15792 & n15793 ) ;
  assign n15794 = ( n15792 & ~n15782 ) | ( n15792 & n15793 ) | ( ~n15782 & n15793 ) ;
  assign n15796 = ( n15782 & ~n15795 ) | ( n15782 & n15794 ) | ( ~n15795 & n15794 ) ;
  assign n15797 = ( n15724 & n15734 ) | ( n15724 & n15796 ) | ( n15734 & n15796 ) ;
  assign n15798 = ( n15734 & ~n15724 ) | ( n15734 & n15796 ) | ( ~n15724 & n15796 ) ;
  assign n15799 = ( n15724 & ~n15797 ) | ( n15724 & n15798 ) | ( ~n15797 & n15798 ) ;
  assign n15803 = n11116 | n5135 ;
  assign n15800 = n5010 | n11122 ;
  assign n15801 = ~n5067 & n11119 ;
  assign n15802 = ( n15800 & ~n15801 ) | ( n15800 & 1'b0 ) | ( ~n15801 & 1'b0 ) ;
  assign n15804 = ( n5135 & ~n15803 ) | ( n5135 & n15802 ) | ( ~n15803 & n15802 ) ;
  assign n15805 = n5012 | n11230 ;
  assign n15806 = n15804 &  n15805 ;
  assign n15807 = x23 &  n15806 ;
  assign n15808 = x23 | n15806 ;
  assign n15809 = ~n15807 & n15808 ;
  assign n15811 = ( n15631 & n15799 ) | ( n15631 & n15809 ) | ( n15799 & n15809 ) ;
  assign n15810 = ( n15631 & ~n15799 ) | ( n15631 & n15809 ) | ( ~n15799 & n15809 ) ;
  assign n15812 = ( n15799 & ~n15811 ) | ( n15799 & n15810 ) | ( ~n15811 & n15810 ) ;
  assign n15816 = n11107 | n5837 ;
  assign n15813 = ( n5339 & ~n11113 ) | ( n5339 & 1'b0 ) | ( ~n11113 & 1'b0 ) ;
  assign n15814 = n5761 | n11110 ;
  assign n15815 = ~n15813 & n15814 ;
  assign n15817 = ( n5837 & ~n15816 ) | ( n5837 & n15815 ) | ( ~n15816 & n15815 ) ;
  assign n15818 = ~n5341 & n12340 ;
  assign n15819 = ( n15817 & ~n15818 ) | ( n15817 & 1'b0 ) | ( ~n15818 & 1'b0 ) ;
  assign n15820 = x20 &  n15819 ;
  assign n15821 = x20 | n15819 ;
  assign n15822 = ~n15820 & n15821 ;
  assign n15823 = ( n15633 & n15643 ) | ( n15633 & n15644 ) | ( n15643 & n15644 ) ;
  assign n15825 = ( n15812 & n15822 ) | ( n15812 & n15823 ) | ( n15822 & n15823 ) ;
  assign n15824 = ( n15822 & ~n15812 ) | ( n15822 & n15823 ) | ( ~n15812 & n15823 ) ;
  assign n15826 = ( n15812 & ~n15825 ) | ( n15812 & n15824 ) | ( ~n15825 & n15824 ) ;
  assign n15830 = ~n6395 & n11098 ;
  assign n15827 = n5970 | n11104 ;
  assign n15828 = n6170 | n11101 ;
  assign n15829 = n15827 &  n15828 ;
  assign n15831 = ( n6395 & n15830 ) | ( n6395 & n15829 ) | ( n15830 & n15829 ) ;
  assign n15832 = n5972 | n11218 ;
  assign n15833 = n15831 &  n15832 ;
  assign n15834 = x17 &  n15833 ;
  assign n15835 = x17 | n15833 ;
  assign n15836 = ~n15834 & n15835 ;
  assign n15838 = ( n15648 & n15826 ) | ( n15648 & n15836 ) | ( n15826 & n15836 ) ;
  assign n15837 = ( n15648 & ~n15826 ) | ( n15648 & n15836 ) | ( ~n15826 & n15836 ) ;
  assign n15839 = ( n15826 & ~n15838 ) | ( n15826 & n15837 ) | ( ~n15838 & n15837 ) ;
  assign n15843 = ~n7097 & n11091 ;
  assign n15840 = n6530 | n11095 ;
  assign n15841 = n6983 | n11093 ;
  assign n15842 = n15840 &  n15841 ;
  assign n15844 = ( n7097 & n15843 ) | ( n7097 & n15842 ) | ( n15843 & n15842 ) ;
  assign n15845 = n6532 | n12984 ;
  assign n15846 = n15844 &  n15845 ;
  assign n15847 = x14 &  n15846 ;
  assign n15848 = x14 | n15846 ;
  assign n15849 = ~n15847 & n15848 ;
  assign n15850 = ( n15650 & n15660 ) | ( n15650 & n15661 ) | ( n15660 & n15661 ) ;
  assign n15852 = ( n15839 & n15849 ) | ( n15839 & n15850 ) | ( n15849 & n15850 ) ;
  assign n15851 = ( n15849 & ~n15839 ) | ( n15849 & n15850 ) | ( ~n15839 & n15850 ) ;
  assign n15853 = ( n15839 & ~n15852 ) | ( n15839 & n15851 ) | ( ~n15852 & n15851 ) ;
  assign n15857 = ~n7783 & n11078 ;
  assign n15854 = ( n7253 & ~n11081 ) | ( n7253 & 1'b0 ) | ( ~n11081 & 1'b0 ) ;
  assign n15855 = n7518 | n11085 ;
  assign n15856 = ~n15854 & n15855 ;
  assign n15858 = ( n7783 & n15857 ) | ( n7783 & n15856 ) | ( n15857 & n15856 ) ;
  assign n15859 = n7255 | n11206 ;
  assign n15860 = n15858 &  n15859 ;
  assign n15861 = x11 &  n15860 ;
  assign n15862 = x11 | n15860 ;
  assign n15863 = ~n15861 & n15862 ;
  assign n15865 = ( n15665 & n15853 ) | ( n15665 & n15863 ) | ( n15853 & n15863 ) ;
  assign n15864 = ( n15665 & ~n15853 ) | ( n15665 & n15863 ) | ( ~n15853 & n15863 ) ;
  assign n15866 = ( n15853 & ~n15865 ) | ( n15853 & n15864 ) | ( ~n15865 & n15864 ) ;
  assign n15867 = ( n8105 & ~n13836 ) | ( n8105 & 1'b0 ) | ( ~n13836 & 1'b0 ) ;
  assign n15868 = n8429 | n14071 ;
  assign n15869 = ~n15867 & n15868 ;
  assign n15870 = ~n8764 & n14355 ;
  assign n15871 = ( n8764 & n15869 ) | ( n8764 & n15870 ) | ( n15869 & n15870 ) ;
  assign n15872 = n8107 | n14363 ;
  assign n15873 = n15871 &  n15872 ;
  assign n15874 = x8 &  n15873 ;
  assign n15875 = x8 | n15873 ;
  assign n15876 = ~n15874 & n15875 ;
  assign n15877 = ( n15667 & n15677 ) | ( n15667 & n15678 ) | ( n15677 & n15678 ) ;
  assign n15879 = ( n15866 & n15876 ) | ( n15866 & n15877 ) | ( n15876 & n15877 ) ;
  assign n15878 = ( n15876 & ~n15866 ) | ( n15876 & n15877 ) | ( ~n15866 & n15877 ) ;
  assign n15880 = ( n15866 & ~n15879 ) | ( n15866 & n15878 ) | ( ~n15879 & n15878 ) ;
  assign n15884 = n14807 | n9997 ;
  assign n15881 = ~n9160 & n14553 ;
  assign n15882 = n9558 | n14803 ;
  assign n15883 = ~n15881 & n15882 ;
  assign n15885 = ( n9997 & ~n15884 ) | ( n9997 & n15883 ) | ( ~n15884 & n15883 ) ;
  assign n15886 = ~n9155 & n15294 ;
  assign n15887 = ( n15885 & ~n15886 ) | ( n15885 & 1'b0 ) | ( ~n15886 & 1'b0 ) ;
  assign n15888 = x5 &  n15887 ;
  assign n15889 = x5 | n15887 ;
  assign n15890 = ~n15888 & n15889 ;
  assign n15892 = ( n15682 & n15880 ) | ( n15682 & n15890 ) | ( n15880 & n15890 ) ;
  assign n15891 = ( n15682 & ~n15880 ) | ( n15682 & n15890 ) | ( ~n15880 & n15890 ) ;
  assign n15893 = ( n15880 & ~n15892 ) | ( n15880 & n15891 ) | ( ~n15892 & n15891 ) ;
  assign n15894 = ( n15318 & ~n15697 ) | ( n15318 & n15532 ) | ( ~n15697 & n15532 ) ;
  assign n15895 = ( n15723 & n15893 ) | ( n15723 & n15894 ) | ( n15893 & n15894 ) ;
  assign n15896 = ( n15893 & ~n15723 ) | ( n15893 & n15894 ) | ( ~n15723 & n15894 ) ;
  assign n15897 = ( ~n15723 & n15895 ) | ( ~n15723 & ~n15896 ) | ( n15895 & ~n15896 ) ;
  assign n15899 = ( n15700 & n15707 ) | ( n15700 & n15897 ) | ( n15707 & n15897 ) ;
  assign n15898 = ( n15707 & ~n15700 ) | ( n15707 & n15897 ) | ( ~n15700 & n15897 ) ;
  assign n15900 = ( n15700 & ~n15899 ) | ( n15700 & n15898 ) | ( ~n15899 & n15898 ) ;
  assign n15906 = ~n4478 & n15900 ;
  assign n15904 = ~n4962 & n15897 ;
  assign n15901 = n4482 | n15320 ;
  assign n15902 = n4495 | n15700 ;
  assign n15903 = n15901 &  n15902 ;
  assign n15905 = ( n4962 & n15904 ) | ( n4962 & n15903 ) | ( n15904 & n15903 ) ;
  assign n15907 = ( n4478 & n15906 ) | ( n4478 & n15905 ) | ( n15906 & n15905 ) ;
  assign n15909 = x26 &  n15907 ;
  assign n15908 = ~x26 & n15907 ;
  assign n15910 = ( x26 & ~n15909 ) | ( x26 & n15908 ) | ( ~n15909 & n15908 ) ;
  assign n15911 = ( n15714 & n15717 ) | ( n15714 & n15910 ) | ( n15717 & n15910 ) ;
  assign n15939 = n301 | n412 ;
  assign n15940 = n602 | n15939 ;
  assign n15941 = ( n14761 & ~n2610 ) | ( n14761 & n15940 ) | ( ~n2610 & n15940 ) ;
  assign n15942 = n2610 | n15941 ;
  assign n15912 = n2632 | n3889 ;
  assign n15913 = ( n1191 & ~n2035 ) | ( n1191 & n15912 ) | ( ~n2035 & n15912 ) ;
  assign n15914 = n2035 | n15913 ;
  assign n15915 = ( n1454 & ~n1585 ) | ( n1454 & n15914 ) | ( ~n1585 & n15914 ) ;
  assign n15916 = n1585 | n15915 ;
  assign n15917 = ( n372 & ~n224 ) | ( n372 & n15916 ) | ( ~n224 & n15916 ) ;
  assign n15918 = n224 | n15917 ;
  assign n15919 = ( n15918 & ~n454 ) | ( n15918 & n540 ) | ( ~n454 & n540 ) ;
  assign n15920 = n454 | n15919 ;
  assign n15921 = ( n135 & ~n643 ) | ( n135 & n15920 ) | ( ~n643 & n15920 ) ;
  assign n15922 = n643 | n15921 ;
  assign n15923 = n358 | n15922 ;
  assign n15927 = n1062 | n1808 ;
  assign n15928 = n4373 | n15927 ;
  assign n15929 = ( n15928 & ~n1549 ) | ( n15928 & n3070 ) | ( ~n1549 & n3070 ) ;
  assign n15930 = n1549 | n15929 ;
  assign n15924 = n1360 | n11262 ;
  assign n15925 = ( n374 & ~n126 ) | ( n374 & n15924 ) | ( ~n126 & n15924 ) ;
  assign n15926 = n126 | n15925 ;
  assign n15931 = ( n3984 & n15930 ) | ( n3984 & n15926 ) | ( n15930 & n15926 ) ;
  assign n15932 = ( n3984 & ~n15931 ) | ( n3984 & 1'b0 ) | ( ~n15931 & 1'b0 ) ;
  assign n15933 = ( n1512 & ~n3377 ) | ( n1512 & n15932 ) | ( ~n3377 & n15932 ) ;
  assign n15934 = ~n1512 & n15933 ;
  assign n15935 = ( n15934 & ~n2666 ) | ( n15934 & n15923 ) | ( ~n2666 & n15923 ) ;
  assign n15936 = ( n218 & ~n15923 ) | ( n218 & n15935 ) | ( ~n15923 & n15935 ) ;
  assign n15937 = ~n218 & n15936 ;
  assign n15938 = ~n191 & n15937 ;
  assign n15943 = ( n1624 & ~n15942 ) | ( n1624 & n15938 ) | ( ~n15942 & n15938 ) ;
  assign n15944 = ( n15943 & ~n1624 ) | ( n15943 & 1'b0 ) | ( ~n1624 & 1'b0 ) ;
  assign n15945 = ( n1627 & ~n2840 ) | ( n1627 & n15944 ) | ( ~n2840 & n15944 ) ;
  assign n15946 = ~n1627 & n15945 ;
  assign n15947 = ( n1511 & ~n2128 ) | ( n1511 & n15946 ) | ( ~n2128 & n15946 ) ;
  assign n15948 = ~n1511 & n15947 ;
  assign n15949 = ( n1761 & ~n715 ) | ( n1761 & n15948 ) | ( ~n715 & n15948 ) ;
  assign n15950 = ~n1761 & n15949 ;
  assign n15951 = ( n383 & ~n15950 ) | ( n383 & n624 ) | ( ~n15950 & n624 ) ;
  assign n15952 = ( n624 & ~n15951 ) | ( n624 & 1'b0 ) | ( ~n15951 & 1'b0 ) ;
  assign n15953 = ( n349 & ~n789 ) | ( n349 & n15952 ) | ( ~n789 & n15952 ) ;
  assign n15954 = ~n349 & n15953 ;
  assign n15955 = ( n524 & ~n15954 ) | ( n524 & n526 ) | ( ~n15954 & n526 ) ;
  assign n15956 = ( n524 & ~n15955 ) | ( n524 & 1'b0 ) | ( ~n15955 & 1'b0 ) ;
  assign n15957 = ( n336 & ~n229 ) | ( n336 & n15956 ) | ( ~n229 & n15956 ) ;
  assign n15958 = ~n336 & n15957 ;
  assign n15959 = ~n663 & n15958 ;
  assign n15960 = ( n15742 & ~n15781 ) | ( n15742 & n15959 ) | ( ~n15781 & n15959 ) ;
  assign n15961 = ( n15781 & ~n15742 ) | ( n15781 & n15959 ) | ( ~n15742 & n15959 ) ;
  assign n15962 = ( n15960 & ~n15959 ) | ( n15960 & n15961 ) | ( ~n15959 & n15961 ) ;
  assign n15963 = n3644 | n11699 ;
  assign n15964 = ( n3652 & ~n11146 ) | ( n3652 & 1'b0 ) | ( ~n11146 & 1'b0 ) ;
  assign n15965 = ( n3657 & ~n11143 ) | ( n3657 & 1'b0 ) | ( ~n11143 & 1'b0 ) ;
  assign n15966 = n15964 | n15965 ;
  assign n15967 = ~n3653 & n11140 ;
  assign n15968 = ( n3653 & ~n15966 ) | ( n3653 & n15967 ) | ( ~n15966 & n15967 ) ;
  assign n15969 = n15963 &  n15968 ;
  assign n15970 = ( n15794 & n15962 ) | ( n15794 & n15969 ) | ( n15962 & n15969 ) ;
  assign n15971 = ( n15962 & ~n15794 ) | ( n15962 & n15969 ) | ( ~n15794 & n15969 ) ;
  assign n15972 = ( n15794 & ~n15970 ) | ( n15794 & n15971 ) | ( ~n15970 & n15971 ) ;
  assign n15976 = ~n4430 & n11131 ;
  assign n15973 = n523 | n11137 ;
  assign n15974 = ~n3939 & n11134 ;
  assign n15975 = ( n15973 & ~n15974 ) | ( n15973 & 1'b0 ) | ( ~n15974 & 1'b0 ) ;
  assign n15977 = ( n4430 & n15976 ) | ( n4430 & n15975 ) | ( n15976 & n15975 ) ;
  assign n15978 = ~n601 & n11888 ;
  assign n15979 = ( n15977 & ~n15978 ) | ( n15977 & 1'b0 ) | ( ~n15978 & 1'b0 ) ;
  assign n15980 = x29 &  n15979 ;
  assign n15981 = x29 | n15979 ;
  assign n15982 = ~n15980 & n15981 ;
  assign n15986 = ~n4962 & n11122 ;
  assign n15983 = ~n4495 & n11125 ;
  assign n15984 = n4482 | n11128 ;
  assign n15985 = ~n15983 & n15984 ;
  assign n15987 = ( n4962 & n15986 ) | ( n4962 & n15985 ) | ( n15986 & n15985 ) ;
  assign n15988 = ~n4478 & n12100 ;
  assign n15989 = ( n15987 & ~n15988 ) | ( n15987 & 1'b0 ) | ( ~n15988 & 1'b0 ) ;
  assign n15990 = x26 &  n15989 ;
  assign n15991 = x26 | n15989 ;
  assign n15992 = ~n15990 & n15991 ;
  assign n15994 = ( n15972 & n15982 ) | ( n15972 & n15992 ) | ( n15982 & n15992 ) ;
  assign n15993 = ( n15982 & ~n15972 ) | ( n15982 & n15992 ) | ( ~n15972 & n15992 ) ;
  assign n15995 = ( n15972 & ~n15994 ) | ( n15972 & n15993 ) | ( ~n15994 & n15993 ) ;
  assign n15996 = ~n5010 & n11119 ;
  assign n15997 = ~n5067 & n11116 ;
  assign n15998 = n15996 | n15997 ;
  assign n15999 = ~n5135 & n11113 ;
  assign n16000 = ( n5135 & ~n15998 ) | ( n5135 & n15999 ) | ( ~n15998 & n15999 ) ;
  assign n16001 = n5012 | n12369 ;
  assign n16002 = n16000 &  n16001 ;
  assign n16003 = x23 &  n16002 ;
  assign n16004 = x23 | n16002 ;
  assign n16005 = ~n16003 & n16004 ;
  assign n16006 = ( n15724 & ~n15796 ) | ( n15724 & n15734 ) | ( ~n15796 & n15734 ) ;
  assign n16008 = ( n15995 & n16005 ) | ( n15995 & n16006 ) | ( n16005 & n16006 ) ;
  assign n16007 = ( n16005 & ~n15995 ) | ( n16005 & n16006 ) | ( ~n15995 & n16006 ) ;
  assign n16009 = ( n15995 & ~n16008 ) | ( n15995 & n16007 ) | ( ~n16008 & n16007 ) ;
  assign n16010 = ( n5339 & ~n11110 ) | ( n5339 & 1'b0 ) | ( ~n11110 & 1'b0 ) ;
  assign n16011 = ~n5761 & n11107 ;
  assign n16012 = n16010 | n16011 ;
  assign n16013 = ~n5837 & n11104 ;
  assign n16014 = ( n5837 & ~n16012 ) | ( n5837 & n16013 ) | ( ~n16012 & n16013 ) ;
  assign n16015 = ~n5341 & n12662 ;
  assign n16016 = ( n16014 & ~n16015 ) | ( n16014 & 1'b0 ) | ( ~n16015 & 1'b0 ) ;
  assign n16017 = x20 &  n16016 ;
  assign n16018 = x20 | n16016 ;
  assign n16019 = ~n16017 & n16018 ;
  assign n16021 = ( n15810 & n16009 ) | ( n15810 & n16019 ) | ( n16009 & n16019 ) ;
  assign n16020 = ( n15810 & ~n16009 ) | ( n15810 & n16019 ) | ( ~n16009 & n16019 ) ;
  assign n16022 = ( n16009 & ~n16021 ) | ( n16009 & n16020 ) | ( ~n16021 & n16020 ) ;
  assign n16026 = ~n6395 & n11095 ;
  assign n16023 = n5970 | n11101 ;
  assign n16024 = n6170 | n11098 ;
  assign n16025 = n16023 &  n16024 ;
  assign n16027 = ( n6395 & n16026 ) | ( n6395 & n16025 ) | ( n16026 & n16025 ) ;
  assign n16028 = n5972 | n13014 ;
  assign n16029 = n16027 &  n16028 ;
  assign n16030 = x17 &  n16029 ;
  assign n16031 = x17 | n16029 ;
  assign n16032 = ~n16030 & n16031 ;
  assign n16034 = ( n15824 & n16022 ) | ( n15824 & n16032 ) | ( n16022 & n16032 ) ;
  assign n16033 = ( n15824 & ~n16022 ) | ( n15824 & n16032 ) | ( ~n16022 & n16032 ) ;
  assign n16035 = ( n16022 & ~n16034 ) | ( n16022 & n16033 ) | ( ~n16034 & n16033 ) ;
  assign n16039 = ~n7097 & n11081 ;
  assign n16036 = n6530 | n11093 ;
  assign n16037 = n6983 | n11091 ;
  assign n16038 = n16036 &  n16037 ;
  assign n16040 = ( n7097 & n16039 ) | ( n7097 & n16038 ) | ( n16039 & n16038 ) ;
  assign n16041 = n6532 | n13775 ;
  assign n16042 = n16040 &  n16041 ;
  assign n16043 = x14 &  n16042 ;
  assign n16044 = x14 | n16042 ;
  assign n16045 = ~n16043 & n16044 ;
  assign n16047 = ( n15837 & n16035 ) | ( n15837 & n16045 ) | ( n16035 & n16045 ) ;
  assign n16046 = ( n15837 & ~n16035 ) | ( n15837 & n16045 ) | ( ~n16035 & n16045 ) ;
  assign n16048 = ( n16035 & ~n16047 ) | ( n16035 & n16046 ) | ( ~n16047 & n16046 ) ;
  assign n16052 = ~n7783 & n13836 ;
  assign n16049 = ( n7253 & ~n11085 ) | ( n7253 & 1'b0 ) | ( ~n11085 & 1'b0 ) ;
  assign n16050 = n7518 | n11078 ;
  assign n16051 = ~n16049 & n16050 ;
  assign n16053 = ( n7783 & n16052 ) | ( n7783 & n16051 ) | ( n16052 & n16051 ) ;
  assign n16054 = n7255 | n13844 ;
  assign n16055 = n16053 &  n16054 ;
  assign n16056 = x11 &  n16055 ;
  assign n16057 = x11 | n16055 ;
  assign n16058 = ~n16056 & n16057 ;
  assign n16060 = ( n15851 & n16048 ) | ( n15851 & n16058 ) | ( n16048 & n16058 ) ;
  assign n16059 = ( n15851 & ~n16048 ) | ( n15851 & n16058 ) | ( ~n16048 & n16058 ) ;
  assign n16061 = ( n16048 & ~n16060 ) | ( n16048 & n16059 ) | ( ~n16060 & n16059 ) ;
  assign n16065 = n14553 | n8764 ;
  assign n16062 = ( n8105 & ~n14071 ) | ( n8105 & 1'b0 ) | ( ~n14071 & 1'b0 ) ;
  assign n16063 = n8429 | n14355 ;
  assign n16064 = ~n16062 & n16063 ;
  assign n16066 = ( n8764 & ~n16065 ) | ( n8764 & n16064 ) | ( ~n16065 & n16064 ) ;
  assign n16067 = ~n8107 & n14562 ;
  assign n16068 = ( n16066 & ~n16067 ) | ( n16066 & 1'b0 ) | ( ~n16067 & 1'b0 ) ;
  assign n16069 = x8 &  n16068 ;
  assign n16070 = x8 | n16068 ;
  assign n16071 = ~n16069 & n16070 ;
  assign n16073 = ( n15864 & n16061 ) | ( n15864 & n16071 ) | ( n16061 & n16071 ) ;
  assign n16072 = ( n15864 & ~n16061 ) | ( n15864 & n16071 ) | ( ~n16061 & n16071 ) ;
  assign n16074 = ( n16061 & ~n16073 ) | ( n16061 & n16072 ) | ( ~n16073 & n16072 ) ;
  assign n16078 = n14800 | n9997 ;
  assign n16075 = n9160 | n14803 ;
  assign n16076 = ~n9558 & n14807 ;
  assign n16077 = ( n16075 & ~n16076 ) | ( n16075 & 1'b0 ) | ( ~n16076 & 1'b0 ) ;
  assign n16079 = ( n9997 & ~n16078 ) | ( n9997 & n16077 ) | ( ~n16078 & n16077 ) ;
  assign n16080 = n9155 | n14816 ;
  assign n16081 = n16079 &  n16080 ;
  assign n16082 = x5 &  n16081 ;
  assign n16083 = x5 | n16081 ;
  assign n16084 = ~n16082 & n16083 ;
  assign n16086 = ( n15878 & n16074 ) | ( n15878 & n16084 ) | ( n16074 & n16084 ) ;
  assign n16085 = ( n15878 & ~n16074 ) | ( n15878 & n16084 ) | ( ~n16074 & n16084 ) ;
  assign n16087 = ( n16074 & ~n16086 ) | ( n16074 & n16085 ) | ( ~n16086 & n16085 ) ;
  assign n16088 = ( n15723 & ~n15893 ) | ( n15723 & n15894 ) | ( ~n15893 & n15894 ) ;
  assign n16089 = ( n15891 & n16087 ) | ( n15891 & n16088 ) | ( n16087 & n16088 ) ;
  assign n16090 = ( n16087 & ~n15891 ) | ( n16087 & n16088 ) | ( ~n15891 & n16088 ) ;
  assign n16091 = ( ~n15891 & n16089 ) | ( ~n15891 & ~n16090 ) | ( n16089 & ~n16090 ) ;
  assign n16093 = ( n15897 & n15899 ) | ( n15897 & n16091 ) | ( n15899 & n16091 ) ;
  assign n16092 = ( n15899 & ~n15897 ) | ( n15899 & n16091 ) | ( ~n15897 & n16091 ) ;
  assign n16094 = ( n15897 & ~n16093 ) | ( n15897 & n16092 ) | ( ~n16093 & n16092 ) ;
  assign n16100 = ~n4478 & n16094 ;
  assign n16098 = ~n4962 & n16091 ;
  assign n16095 = n4482 | n15700 ;
  assign n16096 = n4495 | n15897 ;
  assign n16097 = n16095 &  n16096 ;
  assign n16099 = ( n4962 & n16098 ) | ( n4962 & n16097 ) | ( n16098 & n16097 ) ;
  assign n16101 = ( n4478 & n16100 ) | ( n4478 & n16099 ) | ( n16100 & n16099 ) ;
  assign n16103 = x26 &  n16101 ;
  assign n16102 = ~x26 & n16101 ;
  assign n16104 = ( x26 & ~n16103 ) | ( x26 & n16102 ) | ( ~n16103 & n16102 ) ;
  assign n16105 = ( n15429 & ~n15911 ) | ( n15429 & n16104 ) | ( ~n15911 & n16104 ) ;
  assign n16106 = ( n15429 & ~n16104 ) | ( n15429 & n15911 ) | ( ~n16104 & n15911 ) ;
  assign n16107 = ( n16105 & ~n15429 ) | ( n16105 & n16106 ) | ( ~n15429 & n16106 ) ;
  assign n16108 = n3644 | n11687 ;
  assign n16109 = ( n3652 & ~n11143 ) | ( n3652 & 1'b0 ) | ( ~n11143 & 1'b0 ) ;
  assign n16110 = ( n3657 & ~n11140 ) | ( n3657 & 1'b0 ) | ( ~n11140 & 1'b0 ) ;
  assign n16111 = n16109 | n16110 ;
  assign n16112 = ~n3653 & n11137 ;
  assign n16113 = ( n3653 & ~n16111 ) | ( n3653 & n16112 ) | ( ~n16111 & n16112 ) ;
  assign n16114 = n16108 &  n16113 ;
  assign n16115 = n2130 | n3159 ;
  assign n16116 = ( n973 & ~n2764 ) | ( n973 & n16115 ) | ( ~n2764 & n16115 ) ;
  assign n16117 = n2764 | n16116 ;
  assign n16118 = ( n3800 & n16117 ) | ( n3800 & n4114 ) | ( n16117 & n4114 ) ;
  assign n16119 = ( n4114 & ~n16118 ) | ( n4114 & 1'b0 ) | ( ~n16118 & 1'b0 ) ;
  assign n16120 = ( n341 & ~n3502 ) | ( n341 & n16119 ) | ( ~n3502 & n16119 ) ;
  assign n16121 = ~n341 & n16120 ;
  assign n16122 = ( n814 & ~n52 ) | ( n814 & n16121 ) | ( ~n52 & n16121 ) ;
  assign n16123 = ~n814 & n16122 ;
  assign n16124 = ( n267 & ~n188 ) | ( n267 & n16123 ) | ( ~n188 & n16123 ) ;
  assign n16125 = ~n267 & n16124 ;
  assign n16126 = ( n148 & n197 ) | ( n148 & n16125 ) | ( n197 & n16125 ) ;
  assign n16127 = ~n148 & n16126 ;
  assign n16128 = ( n603 & ~n492 ) | ( n603 & n16127 ) | ( ~n492 & n16127 ) ;
  assign n16129 = ~n603 & n16128 ;
  assign n16130 = ( n285 & ~n628 ) | ( n285 & n16129 ) | ( ~n628 & n16129 ) ;
  assign n16131 = ~n285 & n16130 ;
  assign n16133 = n15742 &  n16131 ;
  assign n16132 = ( n15742 & ~n16131 ) | ( n15742 & 1'b0 ) | ( ~n16131 & 1'b0 ) ;
  assign n16134 = ( n16131 & ~n16133 ) | ( n16131 & n16132 ) | ( ~n16133 & n16132 ) ;
  assign n16135 = ( n16114 & ~n15961 ) | ( n16114 & n16134 ) | ( ~n15961 & n16134 ) ;
  assign n16136 = ( n15961 & ~n16114 ) | ( n15961 & n16134 ) | ( ~n16114 & n16134 ) ;
  assign n16137 = ( n16135 & ~n16134 ) | ( n16135 & n16136 ) | ( ~n16134 & n16136 ) ;
  assign n16141 = ~n4430 & n11128 ;
  assign n16138 = ~n523 & n11134 ;
  assign n16139 = n3939 | n11131 ;
  assign n16140 = ~n16138 & n16139 ;
  assign n16142 = ( n4430 & n16141 ) | ( n4430 & n16140 ) | ( n16141 & n16140 ) ;
  assign n16143 = n601 | n11871 ;
  assign n16144 = n16142 &  n16143 ;
  assign n16145 = x29 &  n16144 ;
  assign n16146 = x29 | n16144 ;
  assign n16147 = ~n16145 & n16146 ;
  assign n16148 = ( n15794 & ~n15962 ) | ( n15794 & n15969 ) | ( ~n15962 & n15969 ) ;
  assign n16149 = ( n16137 & n16147 ) | ( n16137 & n16148 ) | ( n16147 & n16148 ) ;
  assign n16150 = ( n16147 & ~n16137 ) | ( n16147 & n16148 ) | ( ~n16137 & n16148 ) ;
  assign n16151 = ( n16137 & ~n16149 ) | ( n16137 & n16150 ) | ( ~n16149 & n16150 ) ;
  assign n16152 = n4962 &  n11119 ;
  assign n16153 = ~n4482 & n11125 ;
  assign n16154 = n4495 | n11122 ;
  assign n16155 = ~n16153 & n16154 ;
  assign n16156 = ( n16152 & ~n11119 ) | ( n16152 & n16155 ) | ( ~n11119 & n16155 ) ;
  assign n16157 = ~n4478 & n12088 ;
  assign n16158 = ( n16156 & ~n16157 ) | ( n16156 & 1'b0 ) | ( ~n16157 & 1'b0 ) ;
  assign n16159 = x26 &  n16158 ;
  assign n16160 = x26 | n16158 ;
  assign n16161 = ~n16159 & n16160 ;
  assign n16162 = ( n15993 & n16151 ) | ( n15993 & n16161 ) | ( n16151 & n16161 ) ;
  assign n16163 = ( n16151 & ~n15993 ) | ( n16151 & n16161 ) | ( ~n15993 & n16161 ) ;
  assign n16164 = ( n15993 & ~n16162 ) | ( n15993 & n16163 ) | ( ~n16162 & n16163 ) ;
  assign n16168 = ~n5135 & n11110 ;
  assign n16165 = ~n5010 & n11116 ;
  assign n16166 = n5067 | n11113 ;
  assign n16167 = ~n16165 & n16166 ;
  assign n16169 = ( n5135 & n16168 ) | ( n5135 & n16167 ) | ( n16168 & n16167 ) ;
  assign n16170 = ~n5012 & n12352 ;
  assign n16171 = ( n16169 & ~n16170 ) | ( n16169 & 1'b0 ) | ( ~n16170 & 1'b0 ) ;
  assign n16173 = ( x23 & n16164 ) | ( x23 & n16171 ) | ( n16164 & n16171 ) ;
  assign n16172 = ( n16164 & ~x23 ) | ( n16164 & n16171 ) | ( ~x23 & n16171 ) ;
  assign n16174 = ( x23 & ~n16173 ) | ( x23 & n16172 ) | ( ~n16173 & n16172 ) ;
  assign n16178 = ~n5837 & n11101 ;
  assign n16175 = n5339 &  n11107 ;
  assign n16176 = n5761 | n11104 ;
  assign n16177 = ~n16175 & n16176 ;
  assign n16179 = ( n5837 & n16178 ) | ( n5837 & n16177 ) | ( n16178 & n16177 ) ;
  assign n16180 = n5341 | n12650 ;
  assign n16181 = n16179 &  n16180 ;
  assign n16182 = x20 &  n16181 ;
  assign n16183 = x20 | n16181 ;
  assign n16184 = ~n16182 & n16183 ;
  assign n16186 = ( n16007 & n16174 ) | ( n16007 & n16184 ) | ( n16174 & n16184 ) ;
  assign n16185 = ( n16007 & ~n16174 ) | ( n16007 & n16184 ) | ( ~n16174 & n16184 ) ;
  assign n16187 = ( n16174 & ~n16186 ) | ( n16174 & n16185 ) | ( ~n16186 & n16185 ) ;
  assign n16191 = ~n6395 & n11093 ;
  assign n16188 = n5970 | n11098 ;
  assign n16189 = n6170 | n11095 ;
  assign n16190 = n16188 &  n16189 ;
  assign n16192 = ( n6395 & n16191 ) | ( n6395 & n16190 ) | ( n16191 & n16190 ) ;
  assign n16193 = n5972 | n12997 ;
  assign n16194 = n16192 &  n16193 ;
  assign n16195 = x17 &  n16194 ;
  assign n16196 = x17 | n16194 ;
  assign n16197 = ~n16195 & n16196 ;
  assign n16199 = ( n16020 & n16187 ) | ( n16020 & n16197 ) | ( n16187 & n16197 ) ;
  assign n16198 = ( n16020 & ~n16187 ) | ( n16020 & n16197 ) | ( ~n16187 & n16197 ) ;
  assign n16200 = ( n16187 & ~n16199 ) | ( n16187 & n16198 ) | ( ~n16199 & n16198 ) ;
  assign n16204 = ~n7097 & n11085 ;
  assign n16201 = n6530 | n11091 ;
  assign n16202 = n6983 | n11081 ;
  assign n16203 = n16201 &  n16202 ;
  assign n16205 = ( n7097 & n16204 ) | ( n7097 & n16203 ) | ( n16204 & n16203 ) ;
  assign n16206 = n6532 | n13377 ;
  assign n16207 = n16205 &  n16206 ;
  assign n16208 = x14 &  n16207 ;
  assign n16209 = x14 | n16207 ;
  assign n16210 = ~n16208 & n16209 ;
  assign n16212 = ( n16033 & n16200 ) | ( n16033 & n16210 ) | ( n16200 & n16210 ) ;
  assign n16211 = ( n16033 & ~n16200 ) | ( n16033 & n16210 ) | ( ~n16200 & n16210 ) ;
  assign n16213 = ( n16200 & ~n16212 ) | ( n16200 & n16211 ) | ( ~n16212 & n16211 ) ;
  assign n16217 = ~n7783 & n14071 ;
  assign n16214 = ( n7253 & ~n11078 ) | ( n7253 & 1'b0 ) | ( ~n11078 & 1'b0 ) ;
  assign n16215 = n7518 | n13836 ;
  assign n16216 = ~n16214 & n16215 ;
  assign n16218 = ( n7783 & n16217 ) | ( n7783 & n16216 ) | ( n16217 & n16216 ) ;
  assign n16219 = n7255 | n14079 ;
  assign n16220 = n16218 &  n16219 ;
  assign n16221 = x11 &  n16220 ;
  assign n16222 = x11 | n16220 ;
  assign n16223 = ~n16221 & n16222 ;
  assign n16224 = ( n16046 & ~n16213 ) | ( n16046 & n16223 ) | ( ~n16213 & n16223 ) ;
  assign n16334 = ( x26 & ~n16158 ) | ( x26 & n16151 ) | ( ~n16158 & n16151 ) ;
  assign n16335 = ( x26 & ~n16151 ) | ( x26 & n16158 ) | ( ~n16151 & n16158 ) ;
  assign n16336 = ( n16334 & ~x26 ) | ( n16334 & n16335 ) | ( ~x26 & n16335 ) ;
  assign n16337 = x23 &  n16171 ;
  assign n16338 = x23 | n16171 ;
  assign n16339 = ~n16337 & n16338 ;
  assign n16340 = ( n15993 & ~n16336 ) | ( n15993 & n16339 ) | ( ~n16336 & n16339 ) ;
  assign n16310 = n11116 | n4962 ;
  assign n16307 = n4482 | n11122 ;
  assign n16308 = ~n4495 & n11119 ;
  assign n16309 = ( n16307 & ~n16308 ) | ( n16307 & 1'b0 ) | ( ~n16308 & 1'b0 ) ;
  assign n16311 = ( n4962 & ~n16310 ) | ( n4962 & n16309 ) | ( ~n16310 & n16309 ) ;
  assign n16312 = n4478 | n11230 ;
  assign n16313 = n16311 &  n16312 ;
  assign n16314 = x26 &  n16313 ;
  assign n16315 = x26 | n16313 ;
  assign n16316 = ~n16314 & n16315 ;
  assign n16248 = ( n15742 & ~n15961 ) | ( n15742 & n16131 ) | ( ~n15961 & n16131 ) ;
  assign n16249 = ( n15961 & ~n15742 ) | ( n15961 & n16131 ) | ( ~n15742 & n16131 ) ;
  assign n16250 = ( n16248 & ~n16131 ) | ( n16248 & n16249 ) | ( ~n16131 & n16249 ) ;
  assign n16251 = ( n16114 & ~n16250 ) | ( n16114 & n16148 ) | ( ~n16250 & n16148 ) ;
  assign n16252 = n4430 &  n11125 ;
  assign n16253 = n523 | n11131 ;
  assign n16254 = n3939 | n11128 ;
  assign n16255 = n16253 &  n16254 ;
  assign n16256 = ( n16252 & ~n11125 ) | ( n16252 & n16255 ) | ( ~n11125 & n16255 ) ;
  assign n16257 = ~n601 & n11859 ;
  assign n16258 = ( n16256 & ~n16257 ) | ( n16256 & 1'b0 ) | ( ~n16257 & 1'b0 ) ;
  assign n16259 = x29 &  n16258 ;
  assign n16260 = x29 | n16258 ;
  assign n16261 = ~n16259 & n16260 ;
  assign n16294 = ~n3644 & n11242 ;
  assign n16298 = n11134 | n3653 ;
  assign n16295 = ( n3652 & ~n11140 ) | ( n3652 & 1'b0 ) | ( ~n11140 & 1'b0 ) ;
  assign n16296 = ( n3657 & ~n11137 ) | ( n3657 & 1'b0 ) | ( ~n11137 & 1'b0 ) ;
  assign n16297 = n16295 | n16296 ;
  assign n16299 = ( n16298 & ~n3653 ) | ( n16298 & n16297 ) | ( ~n3653 & n16297 ) ;
  assign n16300 = n16294 | n16299 ;
  assign n16288 = ~x5 & n15742 ;
  assign n16289 = x5 | n15742 ;
  assign n16290 = ( n16288 & ~n15742 ) | ( n16288 & n16289 ) | ( ~n15742 & n16289 ) ;
  assign n16262 = ( n9154 & ~n9151 ) | ( n9154 & n9158 ) | ( ~n9151 & n9158 ) ;
  assign n16263 = n9151 | n16262 ;
  assign n16264 = n14800 &  n16263 ;
  assign n16265 = n278 | n2208 ;
  assign n16266 = ( n866 & ~n124 ) | ( n866 & n16265 ) | ( ~n124 & n16265 ) ;
  assign n16267 = n124 | n16266 ;
  assign n16268 = ( n722 & ~n193 ) | ( n722 & n16267 ) | ( ~n193 & n16267 ) ;
  assign n16269 = n193 | n16268 ;
  assign n16270 = ( n188 & ~n404 ) | ( n188 & n16269 ) | ( ~n404 & n16269 ) ;
  assign n16271 = n404 | n16270 ;
  assign n16272 = ( n343 & n909 ) | ( n343 & n16271 ) | ( n909 & n16271 ) ;
  assign n16273 = ( n343 & ~n16272 ) | ( n343 & 1'b0 ) | ( ~n16272 & 1'b0 ) ;
  assign n16274 = n197 &  n16273 ;
  assign n16275 = ( n1485 & ~n4371 ) | ( n1485 & 1'b0 ) | ( ~n4371 & 1'b0 ) ;
  assign n16276 = ( n6294 & ~n6775 ) | ( n6294 & n16275 ) | ( ~n6775 & n16275 ) ;
  assign n16277 = ~n6294 & n16276 ;
  assign n16278 = ( n4173 & n16274 ) | ( n4173 & n16277 ) | ( n16274 & n16277 ) ;
  assign n16279 = ~n4173 & n16278 ;
  assign n16280 = ( n2427 & n15938 ) | ( n2427 & n16279 ) | ( n15938 & n16279 ) ;
  assign n16281 = ~n2427 & n16280 ;
  assign n16282 = ( n1046 & n4090 ) | ( n1046 & n16281 ) | ( n4090 & n16281 ) ;
  assign n16283 = ~n1046 & n16282 ;
  assign n16284 = ( n241 & ~n242 ) | ( n241 & n16283 ) | ( ~n242 & n16283 ) ;
  assign n16285 = ~n241 & n16284 ;
  assign n16286 = ( n761 & ~n256 ) | ( n761 & n16285 ) | ( ~n256 & n16285 ) ;
  assign n16287 = ~n761 & n16286 ;
  assign n16291 = ( n16264 & n16287 ) | ( n16264 & n16290 ) | ( n16287 & n16290 ) ;
  assign n16292 = ( n16264 & ~n16290 ) | ( n16264 & n16287 ) | ( ~n16290 & n16287 ) ;
  assign n16293 = ( n16290 & ~n16291 ) | ( n16290 & n16292 ) | ( ~n16291 & n16292 ) ;
  assign n16302 = ( n16249 & n16293 ) | ( n16249 & n16300 ) | ( n16293 & n16300 ) ;
  assign n16301 = ( n16249 & ~n16300 ) | ( n16249 & n16293 ) | ( ~n16300 & n16293 ) ;
  assign n16303 = ( n16300 & ~n16302 ) | ( n16300 & n16301 ) | ( ~n16302 & n16301 ) ;
  assign n16304 = ( n16251 & n16261 ) | ( n16251 & n16303 ) | ( n16261 & n16303 ) ;
  assign n16305 = ( n16261 & ~n16251 ) | ( n16261 & n16303 ) | ( ~n16251 & n16303 ) ;
  assign n16306 = ( n16251 & ~n16304 ) | ( n16251 & n16305 ) | ( ~n16304 & n16305 ) ;
  assign n16317 = ( n16114 & n16148 ) | ( n16114 & n16250 ) | ( n16148 & n16250 ) ;
  assign n16318 = ( n16114 & ~n16148 ) | ( n16114 & n16250 ) | ( ~n16148 & n16250 ) ;
  assign n16319 = ( n16148 & ~n16317 ) | ( n16148 & n16318 ) | ( ~n16317 & n16318 ) ;
  assign n16320 = ( n16147 & ~n16319 ) | ( n16147 & n16161 ) | ( ~n16319 & n16161 ) ;
  assign n16321 = ( n16316 & ~n16306 ) | ( n16316 & n16320 ) | ( ~n16306 & n16320 ) ;
  assign n16322 = ( n16306 & ~n16316 ) | ( n16306 & n16320 ) | ( ~n16316 & n16320 ) ;
  assign n16323 = ( n16321 & ~n16320 ) | ( n16321 & n16322 ) | ( ~n16320 & n16322 ) ;
  assign n16327 = n11107 | n5135 ;
  assign n16324 = n5010 | n11113 ;
  assign n16325 = n5067 | n11110 ;
  assign n16326 = n16324 &  n16325 ;
  assign n16328 = ( n5135 & ~n16327 ) | ( n5135 & n16326 ) | ( ~n16327 & n16326 ) ;
  assign n16329 = ~n5012 & n12340 ;
  assign n16330 = ( n16328 & ~n16329 ) | ( n16328 & 1'b0 ) | ( ~n16329 & 1'b0 ) ;
  assign n16331 = x23 &  n16330 ;
  assign n16332 = x23 | n16330 ;
  assign n16333 = ~n16331 & n16332 ;
  assign n16341 = ( n16323 & n16333 ) | ( n16323 & n16340 ) | ( n16333 & n16340 ) ;
  assign n16342 = ( n16323 & ~n16340 ) | ( n16323 & n16333 ) | ( ~n16340 & n16333 ) ;
  assign n16343 = ( n16340 & ~n16341 ) | ( n16340 & n16342 ) | ( ~n16341 & n16342 ) ;
  assign n16344 = ( n5339 & ~n11104 ) | ( n5339 & 1'b0 ) | ( ~n11104 & 1'b0 ) ;
  assign n16345 = n5761 | n11101 ;
  assign n16346 = ~n16344 & n16345 ;
  assign n16347 = ~n5837 & n11098 ;
  assign n16348 = ( n5837 & n16346 ) | ( n5837 & n16347 ) | ( n16346 & n16347 ) ;
  assign n16349 = n5341 | n11218 ;
  assign n16350 = n16348 &  n16349 ;
  assign n16351 = x20 &  n16350 ;
  assign n16352 = x20 | n16350 ;
  assign n16353 = ~n16351 & n16352 ;
  assign n16354 = ( n16185 & n16343 ) | ( n16185 & n16353 ) | ( n16343 & n16353 ) ;
  assign n16355 = ( n16343 & ~n16185 ) | ( n16343 & n16353 ) | ( ~n16185 & n16353 ) ;
  assign n16356 = ( n16185 & ~n16354 ) | ( n16185 & n16355 ) | ( ~n16354 & n16355 ) ;
  assign n16360 = ~n6395 & n11091 ;
  assign n16357 = n5970 | n11095 ;
  assign n16358 = n6170 | n11093 ;
  assign n16359 = n16357 &  n16358 ;
  assign n16361 = ( n6395 & n16360 ) | ( n6395 & n16359 ) | ( n16360 & n16359 ) ;
  assign n16362 = n5972 | n12984 ;
  assign n16363 = n16361 &  n16362 ;
  assign n16364 = x17 &  n16363 ;
  assign n16365 = x17 | n16363 ;
  assign n16366 = ~n16364 & n16365 ;
  assign n16367 = ( n16198 & n16356 ) | ( n16198 & n16366 ) | ( n16356 & n16366 ) ;
  assign n16368 = ( n16356 & ~n16198 ) | ( n16356 & n16366 ) | ( ~n16198 & n16366 ) ;
  assign n16369 = ( n16198 & ~n16367 ) | ( n16198 & n16368 ) | ( ~n16367 & n16368 ) ;
  assign n16373 = ~n7097 & n11078 ;
  assign n16370 = n6530 | n11081 ;
  assign n16371 = n6983 | n11085 ;
  assign n16372 = n16370 &  n16371 ;
  assign n16374 = ( n7097 & n16373 ) | ( n7097 & n16372 ) | ( n16373 & n16372 ) ;
  assign n16375 = n6532 | n11206 ;
  assign n16376 = n16374 &  n16375 ;
  assign n16377 = x14 &  n16376 ;
  assign n16378 = x14 | n16376 ;
  assign n16379 = ~n16377 & n16378 ;
  assign n16380 = ( n16211 & n16369 ) | ( n16211 & n16379 ) | ( n16369 & n16379 ) ;
  assign n16381 = ( n16369 & ~n16211 ) | ( n16369 & n16379 ) | ( ~n16211 & n16379 ) ;
  assign n16382 = ( n16211 & ~n16380 ) | ( n16211 & n16381 ) | ( ~n16380 & n16381 ) ;
  assign n16383 = ( n7253 & ~n13836 ) | ( n7253 & 1'b0 ) | ( ~n13836 & 1'b0 ) ;
  assign n16384 = n7518 | n14071 ;
  assign n16385 = ~n16383 & n16384 ;
  assign n16386 = ~n7783 & n14355 ;
  assign n16387 = ( n7783 & n16385 ) | ( n7783 & n16386 ) | ( n16385 & n16386 ) ;
  assign n16388 = n7255 | n14363 ;
  assign n16389 = n16387 &  n16388 ;
  assign n16390 = x11 &  n16389 ;
  assign n16391 = x11 | n16389 ;
  assign n16392 = ~n16390 & n16391 ;
  assign n16393 = ( n16224 & n16382 ) | ( n16224 & n16392 ) | ( n16382 & n16392 ) ;
  assign n16394 = ( n16382 & ~n16224 ) | ( n16382 & n16392 ) | ( ~n16224 & n16392 ) ;
  assign n16395 = ( n16224 & ~n16393 ) | ( n16224 & n16394 ) | ( ~n16393 & n16394 ) ;
  assign n16225 = ( n16046 & n16213 ) | ( n16046 & n16223 ) | ( n16213 & n16223 ) ;
  assign n16226 = ( n16213 & ~n16225 ) | ( n16213 & n16224 ) | ( ~n16225 & n16224 ) ;
  assign n16227 = ( n8105 & ~n14355 ) | ( n8105 & 1'b0 ) | ( ~n14355 & 1'b0 ) ;
  assign n16228 = ~n8429 & n14553 ;
  assign n16229 = n16227 | n16228 ;
  assign n16230 = ~n8764 & n14803 ;
  assign n16231 = ( n8764 & ~n16229 ) | ( n8764 & n16230 ) | ( ~n16229 & n16230 ) ;
  assign n16232 = ~n8107 & n15310 ;
  assign n16233 = ( n16231 & ~n16232 ) | ( n16231 & 1'b0 ) | ( ~n16232 & 1'b0 ) ;
  assign n16234 = x8 &  n16233 ;
  assign n16235 = x8 | n16233 ;
  assign n16236 = ~n16234 & n16235 ;
  assign n16237 = ( n16059 & ~n16226 ) | ( n16059 & n16236 ) | ( ~n16226 & n16236 ) ;
  assign n16241 = n8764 | n14807 ;
  assign n16238 = n8105 &  n14553 ;
  assign n16239 = n8429 | n14803 ;
  assign n16240 = ~n16238 & n16239 ;
  assign n16242 = ( n8764 & ~n16241 ) | ( n8764 & n16240 ) | ( ~n16241 & n16240 ) ;
  assign n16243 = ~n8107 & n15294 ;
  assign n16244 = ( n16242 & ~n16243 ) | ( n16242 & 1'b0 ) | ( ~n16243 & 1'b0 ) ;
  assign n16245 = x8 &  n16244 ;
  assign n16246 = x8 | n16244 ;
  assign n16247 = ~n16245 & n16246 ;
  assign n16576 = ( n16237 & n16247 ) | ( n16237 & n16395 ) | ( n16247 & n16395 ) ;
  assign n16396 = ( n16237 & ~n16395 ) | ( n16237 & n16247 ) | ( ~n16395 & n16247 ) ;
  assign n16577 = ( n16395 & ~n16576 ) | ( n16395 & n16396 ) | ( ~n16576 & n16396 ) ;
  assign n16564 = n9558 &  n9997 ;
  assign n16565 = ( n14800 & ~n16564 ) | ( n14800 & 1'b0 ) | ( ~n16564 & 1'b0 ) ;
  assign n16566 = ~n9160 & n14807 ;
  assign n16567 = n16565 | n16566 ;
  assign n16568 = ( n9155 & n15692 ) | ( n9155 & n16567 ) | ( n15692 & n16567 ) ;
  assign n16569 = ( n15692 & ~n16568 ) | ( n15692 & 1'b0 ) | ( ~n16568 & 1'b0 ) ;
  assign n16570 = ( n16567 & ~x5 ) | ( n16567 & n16569 ) | ( ~x5 & n16569 ) ;
  assign n16571 = ( x5 & ~n16567 ) | ( x5 & n16569 ) | ( ~n16567 & n16569 ) ;
  assign n16572 = ( n16570 & ~n16569 ) | ( n16570 & n16571 ) | ( ~n16569 & n16571 ) ;
  assign n16573 = ( n16059 & n16226 ) | ( n16059 & n16236 ) | ( n16226 & n16236 ) ;
  assign n16574 = ( n16226 & ~n16573 ) | ( n16226 & n16237 ) | ( ~n16573 & n16237 ) ;
  assign n16575 = ( n16572 & ~n16072 ) | ( n16572 & n16574 ) | ( ~n16072 & n16574 ) ;
  assign n16578 = n16072 | n16572 ;
  assign n16579 = n16072 &  n16572 ;
  assign n16580 = ( n16578 & ~n16579 ) | ( n16578 & 1'b0 ) | ( ~n16579 & 1'b0 ) ;
  assign n16581 = n16574 &  n16580 ;
  assign n16582 = n16574 | n16580 ;
  assign n16583 = ~n16581 & n16582 ;
  assign n16584 = ( n15891 & ~n16087 ) | ( n15891 & n16088 ) | ( ~n16087 & n16088 ) ;
  assign n16585 = ( n16085 & n16583 ) | ( n16085 & n16584 ) | ( n16583 & n16584 ) ;
  assign n16593 = ( n16575 & n16577 ) | ( n16575 & n16585 ) | ( n16577 & n16585 ) ;
  assign n16594 = ( n16575 & ~n16577 ) | ( n16575 & n16585 ) | ( ~n16577 & n16585 ) ;
  assign n16595 = ( n16577 & ~n16593 ) | ( n16577 & n16594 ) | ( ~n16593 & n16594 ) ;
  assign n16613 = ~n5135 & n16595 ;
  assign n16610 = n5010 | n16091 ;
  assign n16590 = ( n16583 & ~n16085 ) | ( n16583 & n16584 ) | ( ~n16085 & n16584 ) ;
  assign n16591 = ( n16085 & ~n16585 ) | ( n16085 & n16590 ) | ( ~n16585 & n16590 ) ;
  assign n16611 = n5067 | n16591 ;
  assign n16612 = n16610 &  n16611 ;
  assign n16614 = ( n5135 & n16613 ) | ( n5135 & n16612 ) | ( n16613 & n16612 ) ;
  assign n16600 = ( n16091 & n16093 ) | ( n16091 & n16591 ) | ( n16093 & n16591 ) ;
  assign n16601 = ( n16591 & n16595 ) | ( n16591 & n16600 ) | ( n16595 & n16600 ) ;
  assign n16615 = ( n16595 & ~n16591 ) | ( n16595 & n16600 ) | ( ~n16591 & n16600 ) ;
  assign n16616 = ( n16591 & ~n16601 ) | ( n16591 & n16615 ) | ( ~n16601 & n16615 ) ;
  assign n16617 = n5012 | n16616 ;
  assign n16618 = n16614 &  n16617 ;
  assign n16619 = x23 &  n16618 ;
  assign n16620 = x23 | n16618 ;
  assign n16621 = ~n16619 & n16620 ;
  assign n16622 = ( n15714 & ~n15910 ) | ( n15714 & n15717 ) | ( ~n15910 & n15717 ) ;
  assign n16623 = ( n15717 & ~n15714 ) | ( n15717 & n15910 ) | ( ~n15714 & n15910 ) ;
  assign n16624 = ( n16622 & ~n15717 ) | ( n16622 & n16623 ) | ( ~n15717 & n16623 ) ;
  assign n16628 = ~n5135 & n16591 ;
  assign n16625 = n5010 | n15897 ;
  assign n16626 = n5067 | n16091 ;
  assign n16627 = n16625 &  n16626 ;
  assign n16629 = ( n5135 & n16628 ) | ( n5135 & n16627 ) | ( n16628 & n16627 ) ;
  assign n16630 = ( n16093 & ~n16091 ) | ( n16093 & n16591 ) | ( ~n16091 & n16591 ) ;
  assign n16631 = ( n16091 & ~n16600 ) | ( n16091 & n16630 ) | ( ~n16600 & n16630 ) ;
  assign n16632 = n5012 | n16631 ;
  assign n16633 = n16629 &  n16632 ;
  assign n16634 = x23 &  n16633 ;
  assign n16635 = x23 | n16633 ;
  assign n16636 = ~n16634 & n16635 ;
  assign n16637 = ( n15528 & ~n15713 ) | ( n15528 & n15531 ) | ( ~n15713 & n15531 ) ;
  assign n16638 = ( n15531 & ~n15528 ) | ( n15531 & n15713 ) | ( ~n15528 & n15713 ) ;
  assign n16639 = ( n16637 & ~n15531 ) | ( n16637 & n16638 ) | ( ~n15531 & n16638 ) ;
  assign n16643 = ~n5135 & n16091 ;
  assign n16640 = n5010 | n15700 ;
  assign n16641 = n5067 | n15897 ;
  assign n16642 = n16640 &  n16641 ;
  assign n16644 = ( n5135 & n16643 ) | ( n5135 & n16642 ) | ( n16643 & n16642 ) ;
  assign n16645 = n5012 | n16094 ;
  assign n16646 = n16644 &  n16645 ;
  assign n16647 = x23 &  n16646 ;
  assign n16648 = x23 | n16646 ;
  assign n16649 = ~n16647 & n16648 ;
  assign n16650 = ( n15517 & ~n15514 ) | ( n15517 & n15527 ) | ( ~n15514 & n15527 ) ;
  assign n16651 = ( n15514 & ~n15527 ) | ( n15514 & n15517 ) | ( ~n15527 & n15517 ) ;
  assign n16652 = ( n16650 & ~n15517 ) | ( n16650 & n16651 ) | ( ~n15517 & n16651 ) ;
  assign n16656 = ~n5135 & n15897 ;
  assign n16653 = n5010 | n15320 ;
  assign n16654 = n5067 | n15700 ;
  assign n16655 = n16653 &  n16654 ;
  assign n16657 = ( n5135 & n16656 ) | ( n5135 & n16655 ) | ( n16656 & n16655 ) ;
  assign n16658 = ( n5012 & ~n15900 ) | ( n5012 & n16657 ) | ( ~n15900 & n16657 ) ;
  assign n16659 = ~n5012 & n16658 ;
  assign n16660 = ( x23 & ~n16657 ) | ( x23 & n16659 ) | ( ~n16657 & n16659 ) ;
  assign n16661 = ( n16657 & ~x23 ) | ( n16657 & n16659 ) | ( ~x23 & n16659 ) ;
  assign n16662 = ( n16660 & ~n16659 ) | ( n16660 & n16661 ) | ( ~n16659 & n16661 ) ;
  assign n16663 = ( n15503 & ~n15500 ) | ( n15503 & n15513 ) | ( ~n15500 & n15513 ) ;
  assign n16664 = ( n15500 & ~n15513 ) | ( n15500 & n15503 ) | ( ~n15513 & n15503 ) ;
  assign n16665 = ( n16663 & ~n15503 ) | ( n16663 & n16664 ) | ( ~n15503 & n16664 ) ;
  assign n16666 = ( n15439 & ~n15499 ) | ( n15439 & n15441 ) | ( ~n15499 & n15441 ) ;
  assign n16667 = ( n15441 & ~n15439 ) | ( n15441 & n15499 ) | ( ~n15439 & n15499 ) ;
  assign n16668 = ( n16666 & ~n15441 ) | ( n16666 & n16667 ) | ( ~n15441 & n16667 ) ;
  assign n16672 = ~n5135 & n15700 ;
  assign n16669 = n5010 | n15325 ;
  assign n16670 = n5067 | n15320 ;
  assign n16671 = n16669 &  n16670 ;
  assign n16673 = ( n5135 & n16672 ) | ( n5135 & n16671 ) | ( n16672 & n16671 ) ;
  assign n16674 = ( n5012 & ~n15708 ) | ( n5012 & n16673 ) | ( ~n15708 & n16673 ) ;
  assign n16675 = ~n5012 & n16674 ;
  assign n16677 = ( x23 & n16673 ) | ( x23 & n16675 ) | ( n16673 & n16675 ) ;
  assign n16676 = ( x23 & ~n16675 ) | ( x23 & n16673 ) | ( ~n16675 & n16673 ) ;
  assign n16678 = ( n16675 & ~n16677 ) | ( n16675 & n16676 ) | ( ~n16677 & n16676 ) ;
  assign n16679 = ( n15451 & ~n15498 ) | ( n15451 & n15456 ) | ( ~n15498 & n15456 ) ;
  assign n16680 = ( n15456 & ~n15451 ) | ( n15456 & n15498 ) | ( ~n15451 & n15498 ) ;
  assign n16681 = ( n16679 & ~n15456 ) | ( n16679 & n16680 ) | ( ~n15456 & n16680 ) ;
  assign n16685 = ~n5135 & n15320 ;
  assign n16682 = n5010 | n15322 ;
  assign n16683 = n5067 | n15325 ;
  assign n16684 = n16682 &  n16683 ;
  assign n16686 = ( n5135 & n16685 ) | ( n5135 & n16684 ) | ( n16685 & n16684 ) ;
  assign n16687 = ( n5012 & ~n15334 ) | ( n5012 & n16686 ) | ( ~n15334 & n16686 ) ;
  assign n16688 = ~n5012 & n16687 ;
  assign n16689 = ( x23 & ~n16686 ) | ( x23 & n16688 ) | ( ~n16686 & n16688 ) ;
  assign n16690 = ( n16686 & ~x23 ) | ( n16686 & n16688 ) | ( ~x23 & n16688 ) ;
  assign n16691 = ( n16689 & ~n16688 ) | ( n16689 & n16690 ) | ( ~n16688 & n16690 ) ;
  assign n16695 = ~n5135 & n15325 ;
  assign n16692 = ~n5010 & n14745 ;
  assign n16693 = n5067 | n15322 ;
  assign n16694 = ~n16692 & n16693 ;
  assign n16696 = ( n5135 & n16695 ) | ( n5135 & n16694 ) | ( n16695 & n16694 ) ;
  assign n16697 = n5012 | n15346 ;
  assign n16698 = n16696 &  n16697 ;
  assign n16699 = x23 &  n16698 ;
  assign n16700 = x23 | n16698 ;
  assign n16701 = ~n16699 & n16700 ;
  assign n16702 = ( n15470 & ~n15460 ) | ( n15470 & n15497 ) | ( ~n15460 & n15497 ) ;
  assign n16703 = ( n15498 & ~n15470 ) | ( n15498 & n16702 ) | ( ~n15470 & n16702 ) ;
  assign n16705 = ( n15397 & n15486 ) | ( n15397 & n15496 ) | ( n15486 & n15496 ) ;
  assign n16704 = ( n15397 & ~n15486 ) | ( n15397 & n15496 ) | ( ~n15486 & n15496 ) ;
  assign n16706 = ( n15486 & ~n16705 ) | ( n15486 & n16704 ) | ( ~n16705 & n16704 ) ;
  assign n16710 = ~n5135 & n15322 ;
  assign n16707 = n5010 | n14528 ;
  assign n16708 = ~n5067 & n14745 ;
  assign n16709 = ( n16707 & ~n16708 ) | ( n16707 & 1'b0 ) | ( ~n16708 & 1'b0 ) ;
  assign n16711 = ( n5135 & n16710 ) | ( n5135 & n16709 ) | ( n16710 & n16709 ) ;
  assign n16712 = ( n5012 & ~n16711 ) | ( n5012 & n15361 ) | ( ~n16711 & n15361 ) ;
  assign n16713 = ( n15361 & ~n16712 ) | ( n15361 & 1'b0 ) | ( ~n16712 & 1'b0 ) ;
  assign n16714 = ( x23 & ~n16711 ) | ( x23 & n16713 ) | ( ~n16711 & n16713 ) ;
  assign n16715 = ( n16711 & ~x23 ) | ( n16711 & n16713 ) | ( ~x23 & n16713 ) ;
  assign n16716 = ( n16714 & ~n16713 ) | ( n16714 & n16715 ) | ( ~n16713 & n16715 ) ;
  assign n16720 = n14745 | n5135 ;
  assign n16717 = n5010 | n14261 ;
  assign n16718 = n5067 | n14528 ;
  assign n16719 = n16717 &  n16718 ;
  assign n16721 = ( n5135 & ~n16720 ) | ( n5135 & n16719 ) | ( ~n16720 & n16719 ) ;
  assign n16722 = ~n5012 & n14749 ;
  assign n16723 = ( n16721 & ~n16722 ) | ( n16721 & 1'b0 ) | ( ~n16722 & 1'b0 ) ;
  assign n16724 = x23 &  n16723 ;
  assign n16725 = x23 | n16723 ;
  assign n16726 = ~n16724 & n16725 ;
  assign n16727 = ( n15475 & ~x26 ) | ( n15475 & n15476 ) | ( ~x26 & n15476 ) ;
  assign n16728 = ( n15475 & ~n16727 ) | ( n15475 & 1'b0 ) | ( ~n16727 & 1'b0 ) ;
  assign n16729 = ( n15483 & ~x26 ) | ( n15483 & n16728 ) | ( ~x26 & n16728 ) ;
  assign n16730 = ( x26 & ~n15483 ) | ( x26 & n16728 ) | ( ~n15483 & n16728 ) ;
  assign n16731 = ( n16729 & ~n16728 ) | ( n16729 & n16730 ) | ( ~n16728 & n16730 ) ;
  assign n16732 = x26 &  n15476 ;
  assign n16733 = ~n15475 & n16732 ;
  assign n16734 = ( n15475 & ~n16732 ) | ( n15475 & 1'b0 ) | ( ~n16732 & 1'b0 ) ;
  assign n16735 = n16733 | n16734 ;
  assign n16765 = ~n5135 & n14261 ;
  assign n16762 = n5010 | n13785 ;
  assign n16763 = n5067 | n13998 ;
  assign n16764 = n16762 &  n16763 ;
  assign n16766 = ( n5135 & n16765 ) | ( n5135 & n16764 ) | ( n16765 & n16764 ) ;
  assign n16767 = n5012 | n14267 ;
  assign n16768 = n16766 &  n16767 ;
  assign n16769 = x23 &  n16768 ;
  assign n16770 = x23 | n16768 ;
  assign n16771 = ~n16769 & n16770 ;
  assign n16749 = n13790 | n5012 ;
  assign n16746 = n5067 | n13787 ;
  assign n16747 = n5135 | n13785 ;
  assign n16748 = n16746 &  n16747 ;
  assign n16750 = ( n5012 & ~n16749 ) | ( n5012 & n16748 ) | ( ~n16749 & n16748 ) ;
  assign n16757 = ~n5012 & n14001 ;
  assign n16755 = ~n5135 & n13998 ;
  assign n16752 = n5010 | n13787 ;
  assign n16753 = n5067 | n13785 ;
  assign n16754 = n16752 &  n16753 ;
  assign n16756 = ( n5135 & n16755 ) | ( n5135 & n16754 ) | ( n16755 & n16754 ) ;
  assign n16758 = ( n5012 & n16757 ) | ( n5012 & n16756 ) | ( n16757 & n16756 ) ;
  assign n16751 = ( n5005 & ~n13787 ) | ( n5005 & 1'b0 ) | ( ~n13787 & 1'b0 ) ;
  assign n16759 = ( n16750 & ~n16758 ) | ( n16750 & n16751 ) | ( ~n16758 & n16751 ) ;
  assign n16760 = ( x23 & ~n16750 ) | ( x23 & n16759 ) | ( ~n16750 & n16759 ) ;
  assign n16761 = ( x23 & ~n16760 ) | ( x23 & 1'b0 ) | ( ~n16760 & 1'b0 ) ;
  assign n16772 = ( n15476 & ~n16771 ) | ( n15476 & n16761 ) | ( ~n16771 & n16761 ) ;
  assign n16739 = ~n5135 & n14528 ;
  assign n16736 = n5010 | n13998 ;
  assign n16737 = n5067 | n14261 ;
  assign n16738 = n16736 &  n16737 ;
  assign n16740 = ( n5135 & n16739 ) | ( n5135 & n16738 ) | ( n16739 & n16738 ) ;
  assign n16741 = ( n14532 & ~n5012 ) | ( n14532 & n16740 ) | ( ~n5012 & n16740 ) ;
  assign n16742 = ~n14532 & n16741 ;
  assign n16743 = ( x23 & ~n16740 ) | ( x23 & n16742 ) | ( ~n16740 & n16742 ) ;
  assign n16744 = ( n16740 & ~x23 ) | ( n16740 & n16742 ) | ( ~x23 & n16742 ) ;
  assign n16745 = ( n16743 & ~n16742 ) | ( n16743 & n16744 ) | ( ~n16742 & n16744 ) ;
  assign n16773 = ( n16735 & ~n16772 ) | ( n16735 & n16745 ) | ( ~n16772 & n16745 ) ;
  assign n16774 = ( n16726 & n16731 ) | ( n16726 & n16773 ) | ( n16731 & n16773 ) ;
  assign n16775 = ( n16706 & n16716 ) | ( n16706 & n16774 ) | ( n16716 & n16774 ) ;
  assign n16776 = ( n16701 & ~n16703 ) | ( n16701 & n16775 ) | ( ~n16703 & n16775 ) ;
  assign n16777 = ( n16681 & n16691 ) | ( n16681 & n16776 ) | ( n16691 & n16776 ) ;
  assign n16778 = ( n16668 & n16678 ) | ( n16668 & n16777 ) | ( n16678 & n16777 ) ;
  assign n16779 = ( n16662 & n16665 ) | ( n16662 & n16778 ) | ( n16665 & n16778 ) ;
  assign n16780 = ( n16649 & ~n16652 ) | ( n16649 & n16779 ) | ( ~n16652 & n16779 ) ;
  assign n16781 = ( n16636 & n16639 ) | ( n16636 & n16780 ) | ( n16639 & n16780 ) ;
  assign n16782 = ( n16621 & n16624 ) | ( n16621 & n16781 ) | ( n16624 & n16781 ) ;
  assign n16586 = ( n16575 & ~n16585 ) | ( n16575 & n16577 ) | ( ~n16585 & n16577 ) ;
  assign n16447 = x5 | n16264 ;
  assign n16448 = x5 &  n16264 ;
  assign n16449 = ( n16447 & ~n16448 ) | ( n16447 & 1'b0 ) | ( ~n16448 & 1'b0 ) ;
  assign n16450 = ( n15742 & n16287 ) | ( n15742 & n16449 ) | ( n16287 & n16449 ) ;
  assign n16397 = n713 | n911 ;
  assign n16398 = n603 | n16397 ;
  assign n16399 = n1534 | n16398 ;
  assign n16400 = ( n795 & ~n2035 ) | ( n795 & n16399 ) | ( ~n2035 & n16399 ) ;
  assign n16401 = n2035 | n16400 ;
  assign n16402 = ( n718 & ~n207 ) | ( n718 & n16401 ) | ( ~n207 & n16401 ) ;
  assign n16403 = n207 | n16402 ;
  assign n16404 = ( n384 & ~n214 ) | ( n384 & n16403 ) | ( ~n214 & n16403 ) ;
  assign n16405 = n214 | n16404 ;
  assign n16406 = ( n568 & ~n631 ) | ( n568 & n16405 ) | ( ~n631 & n16405 ) ;
  assign n16407 = n631 | n16406 ;
  assign n16408 = ( n1232 & ~n1278 ) | ( n1232 & n14619 ) | ( ~n1278 & n14619 ) ;
  assign n16409 = n1278 | n16408 ;
  assign n16410 = ( n272 & ~n722 ) | ( n272 & n16409 ) | ( ~n722 & n16409 ) ;
  assign n16411 = n722 | n16410 ;
  assign n16412 = ( n135 & ~n556 ) | ( n135 & n16411 ) | ( ~n556 & n16411 ) ;
  assign n16413 = n556 | n16412 ;
  assign n16414 = n670 | n16413 ;
  assign n16425 = n1466 | n2808 ;
  assign n16426 = n1342 | n16425 ;
  assign n16415 = n1618 | n2254 ;
  assign n16416 = ( n4697 & ~n3031 ) | ( n4697 & n16415 ) | ( ~n3031 & n16415 ) ;
  assign n16417 = n3031 | n16416 ;
  assign n16418 = ( n1581 & ~n1490 ) | ( n1581 & n16417 ) | ( ~n1490 & n16417 ) ;
  assign n16419 = n1490 | n16418 ;
  assign n16420 = ( n253 & ~n232 ) | ( n253 & n16419 ) | ( ~n232 & n16419 ) ;
  assign n16421 = n232 | n16420 ;
  assign n16422 = ( n216 & ~n572 ) | ( n216 & n16421 ) | ( ~n572 & n16421 ) ;
  assign n16423 = n572 | n16422 ;
  assign n16424 = n627 | n16423 ;
  assign n16427 = ( n4309 & ~n16426 ) | ( n4309 & n16424 ) | ( ~n16426 & n16424 ) ;
  assign n16428 = ( n3129 & ~n16427 ) | ( n3129 & n16424 ) | ( ~n16427 & n16424 ) ;
  assign n16429 = ( n3129 & ~n16428 ) | ( n3129 & 1'b0 ) | ( ~n16428 & 1'b0 ) ;
  assign n16430 = ( n16407 & ~n16414 ) | ( n16407 & n16429 ) | ( ~n16414 & n16429 ) ;
  assign n16431 = ( n887 & ~n16407 ) | ( n887 & n16430 ) | ( ~n16407 & n16430 ) ;
  assign n16432 = ~n887 & n16431 ;
  assign n16433 = ( n3245 & ~n16432 ) | ( n3245 & n645 ) | ( ~n16432 & n645 ) ;
  assign n16434 = ( n645 & ~n16433 ) | ( n645 & 1'b0 ) | ( ~n16433 & 1'b0 ) ;
  assign n16435 = ( n673 & ~n341 ) | ( n673 & n16434 ) | ( ~n341 & n16434 ) ;
  assign n16436 = ~n673 & n16435 ;
  assign n16437 = ( n16436 & ~n105 ) | ( n16436 & n376 ) | ( ~n105 & n376 ) ;
  assign n16438 = ( n16437 & ~n376 ) | ( n16437 & 1'b0 ) | ( ~n376 & 1'b0 ) ;
  assign n16439 = ~n95 & n16438 ;
  assign n16445 = n11888 | n3644 ;
  assign n16440 = n3653 | n11131 ;
  assign n16441 = n3657 &  n11134 ;
  assign n16442 = ( n3652 & ~n11137 ) | ( n3652 & 1'b0 ) | ( ~n11137 & 1'b0 ) ;
  assign n16443 = n16441 | n16442 ;
  assign n16444 = ( n16440 & ~n16443 ) | ( n16440 & 1'b0 ) | ( ~n16443 & 1'b0 ) ;
  assign n16446 = ( n3644 & ~n16445 ) | ( n3644 & n16444 ) | ( ~n16445 & n16444 ) ;
  assign n16452 = ( n16439 & n16446 ) | ( n16439 & n16450 ) | ( n16446 & n16450 ) ;
  assign n16451 = ( n16439 & ~n16450 ) | ( n16439 & n16446 ) | ( ~n16450 & n16446 ) ;
  assign n16453 = ( n16450 & ~n16452 ) | ( n16450 & n16451 ) | ( ~n16452 & n16451 ) ;
  assign n16457 = ~n4430 & n11122 ;
  assign n16454 = n523 | n11128 ;
  assign n16455 = ~n3939 & n11125 ;
  assign n16456 = ( n16454 & ~n16455 ) | ( n16454 & 1'b0 ) | ( ~n16455 & 1'b0 ) ;
  assign n16458 = ( n4430 & n16457 ) | ( n4430 & n16456 ) | ( n16457 & n16456 ) ;
  assign n16459 = ( n601 & ~n16458 ) | ( n601 & n12100 ) | ( ~n16458 & n12100 ) ;
  assign n16460 = ( n12100 & ~n16459 ) | ( n12100 & 1'b0 ) | ( ~n16459 & 1'b0 ) ;
  assign n16461 = ( x29 & ~n16458 ) | ( x29 & n16460 ) | ( ~n16458 & n16460 ) ;
  assign n16462 = ( n16458 & ~x29 ) | ( n16458 & n16460 ) | ( ~x29 & n16460 ) ;
  assign n16463 = ( n16461 & ~n16460 ) | ( n16461 & n16462 ) | ( ~n16460 & n16462 ) ;
  assign n16464 = ( n16453 & ~n16301 ) | ( n16453 & n16463 ) | ( ~n16301 & n16463 ) ;
  assign n16465 = ( n16301 & ~n16463 ) | ( n16301 & n16453 ) | ( ~n16463 & n16453 ) ;
  assign n16466 = ( n16464 & ~n16453 ) | ( n16464 & n16465 ) | ( ~n16453 & n16465 ) ;
  assign n16467 = ( n16251 & ~n16303 ) | ( n16251 & n16261 ) | ( ~n16303 & n16261 ) ;
  assign n16469 = ~n4482 & n11119 ;
  assign n16470 = ~n4495 & n11116 ;
  assign n16471 = n16469 | n16470 ;
  assign n16468 = ( n4962 & ~n11113 ) | ( n4962 & 1'b0 ) | ( ~n11113 & 1'b0 ) ;
  assign n16472 = ( n11113 & ~n16471 ) | ( n11113 & n16468 ) | ( ~n16471 & n16468 ) ;
  assign n16473 = n4478 | n12369 ;
  assign n16474 = n16472 &  n16473 ;
  assign n16475 = x26 &  n16474 ;
  assign n16476 = x26 | n16474 ;
  assign n16477 = ~n16475 & n16476 ;
  assign n16478 = ( n16466 & ~n16467 ) | ( n16466 & n16477 ) | ( ~n16467 & n16477 ) ;
  assign n16479 = ( n16466 & ~n16477 ) | ( n16466 & n16467 ) | ( ~n16477 & n16467 ) ;
  assign n16480 = ( n16478 & ~n16466 ) | ( n16478 & n16479 ) | ( ~n16466 & n16479 ) ;
  assign n16484 = ~n5135 & n11104 ;
  assign n16481 = n5010 | n11110 ;
  assign n16482 = ~n5067 & n11107 ;
  assign n16483 = ( n16481 & ~n16482 ) | ( n16481 & 1'b0 ) | ( ~n16482 & 1'b0 ) ;
  assign n16485 = ( n5135 & n16484 ) | ( n5135 & n16483 ) | ( n16484 & n16483 ) ;
  assign n16486 = ~n5012 & n12662 ;
  assign n16487 = ( n16485 & ~n16486 ) | ( n16485 & 1'b0 ) | ( ~n16486 & 1'b0 ) ;
  assign n16488 = x23 &  n16487 ;
  assign n16489 = x23 | n16487 ;
  assign n16490 = ~n16488 & n16489 ;
  assign n16492 = ( n16321 & n16480 ) | ( n16321 & n16490 ) | ( n16480 & n16490 ) ;
  assign n16491 = ( n16321 & ~n16480 ) | ( n16321 & n16490 ) | ( ~n16480 & n16490 ) ;
  assign n16493 = ( n16480 & ~n16492 ) | ( n16480 & n16491 ) | ( ~n16492 & n16491 ) ;
  assign n16497 = ~n5837 & n11095 ;
  assign n16494 = ( n5339 & ~n11101 ) | ( n5339 & 1'b0 ) | ( ~n11101 & 1'b0 ) ;
  assign n16495 = n5761 | n11098 ;
  assign n16496 = ~n16494 & n16495 ;
  assign n16498 = ( n5837 & n16497 ) | ( n5837 & n16496 ) | ( n16497 & n16496 ) ;
  assign n16499 = n5341 | n13014 ;
  assign n16500 = n16498 &  n16499 ;
  assign n16501 = x20 &  n16500 ;
  assign n16502 = x20 | n16500 ;
  assign n16503 = ~n16501 & n16502 ;
  assign n16504 = ( n16333 & ~n16323 ) | ( n16333 & n16340 ) | ( ~n16323 & n16340 ) ;
  assign n16506 = ( n16493 & n16503 ) | ( n16493 & n16504 ) | ( n16503 & n16504 ) ;
  assign n16505 = ( n16503 & ~n16493 ) | ( n16503 & n16504 ) | ( ~n16493 & n16504 ) ;
  assign n16507 = ( n16493 & ~n16506 ) | ( n16493 & n16505 ) | ( ~n16506 & n16505 ) ;
  assign n16511 = ~n6395 & n11081 ;
  assign n16508 = n5970 | n11093 ;
  assign n16509 = n6170 | n11091 ;
  assign n16510 = n16508 &  n16509 ;
  assign n16512 = ( n6395 & n16511 ) | ( n6395 & n16510 ) | ( n16511 & n16510 ) ;
  assign n16513 = n5972 | n13775 ;
  assign n16514 = n16512 &  n16513 ;
  assign n16515 = x17 &  n16514 ;
  assign n16516 = x17 | n16514 ;
  assign n16517 = ~n16515 & n16516 ;
  assign n16518 = ( n16185 & ~n16343 ) | ( n16185 & n16353 ) | ( ~n16343 & n16353 ) ;
  assign n16520 = ( n16507 & n16517 ) | ( n16507 & n16518 ) | ( n16517 & n16518 ) ;
  assign n16519 = ( n16517 & ~n16507 ) | ( n16517 & n16518 ) | ( ~n16507 & n16518 ) ;
  assign n16521 = ( n16507 & ~n16520 ) | ( n16507 & n16519 ) | ( ~n16520 & n16519 ) ;
  assign n16525 = ~n7097 & n13836 ;
  assign n16522 = n6530 | n11085 ;
  assign n16523 = n6983 | n11078 ;
  assign n16524 = n16522 &  n16523 ;
  assign n16526 = ( n7097 & n16525 ) | ( n7097 & n16524 ) | ( n16525 & n16524 ) ;
  assign n16527 = n6532 | n13844 ;
  assign n16528 = n16526 &  n16527 ;
  assign n16529 = x14 &  n16528 ;
  assign n16530 = x14 | n16528 ;
  assign n16531 = ~n16529 & n16530 ;
  assign n16532 = ( n16198 & ~n16356 ) | ( n16198 & n16366 ) | ( ~n16356 & n16366 ) ;
  assign n16534 = ( n16521 & n16531 ) | ( n16521 & n16532 ) | ( n16531 & n16532 ) ;
  assign n16533 = ( n16531 & ~n16521 ) | ( n16531 & n16532 ) | ( ~n16521 & n16532 ) ;
  assign n16535 = ( n16521 & ~n16534 ) | ( n16521 & n16533 ) | ( ~n16534 & n16533 ) ;
  assign n16539 = n14553 | n7783 ;
  assign n16536 = ( n7253 & ~n14071 ) | ( n7253 & 1'b0 ) | ( ~n14071 & 1'b0 ) ;
  assign n16537 = n7518 | n14355 ;
  assign n16538 = ~n16536 & n16537 ;
  assign n16540 = ( n7783 & ~n16539 ) | ( n7783 & n16538 ) | ( ~n16539 & n16538 ) ;
  assign n16541 = ~n7255 & n14562 ;
  assign n16542 = ( n16540 & ~n16541 ) | ( n16540 & 1'b0 ) | ( ~n16541 & 1'b0 ) ;
  assign n16543 = x11 &  n16542 ;
  assign n16544 = x11 | n16542 ;
  assign n16545 = ~n16543 & n16544 ;
  assign n16546 = ( n16211 & ~n16369 ) | ( n16211 & n16379 ) | ( ~n16369 & n16379 ) ;
  assign n16548 = ( n16535 & n16545 ) | ( n16535 & n16546 ) | ( n16545 & n16546 ) ;
  assign n16547 = ( n16545 & ~n16535 ) | ( n16545 & n16546 ) | ( ~n16535 & n16546 ) ;
  assign n16549 = ( n16535 & ~n16548 ) | ( n16535 & n16547 ) | ( ~n16548 & n16547 ) ;
  assign n16553 = n14800 | n8764 ;
  assign n16550 = ( n8105 & ~n14803 ) | ( n8105 & 1'b0 ) | ( ~n14803 & 1'b0 ) ;
  assign n16551 = ~n8429 & n14807 ;
  assign n16552 = n16550 | n16551 ;
  assign n16554 = ( n16553 & ~n8764 ) | ( n16553 & n16552 ) | ( ~n8764 & n16552 ) ;
  assign n16555 = n8107 | n14816 ;
  assign n16556 = ~n16554 & n16555 ;
  assign n16557 = x8 &  n16556 ;
  assign n16558 = x8 | n16556 ;
  assign n16559 = ~n16557 & n16558 ;
  assign n16560 = ( n16224 & ~n16382 ) | ( n16224 & n16392 ) | ( ~n16382 & n16392 ) ;
  assign n16562 = ( n16549 & n16559 ) | ( n16549 & n16560 ) | ( n16559 & n16560 ) ;
  assign n16561 = ( n16559 & ~n16549 ) | ( n16559 & n16560 ) | ( ~n16549 & n16560 ) ;
  assign n16563 = ( n16549 & ~n16562 ) | ( n16549 & n16561 ) | ( ~n16562 & n16561 ) ;
  assign n16587 = ( n16396 & ~n16586 ) | ( n16396 & n16563 ) | ( ~n16586 & n16563 ) ;
  assign n16588 = ( n16396 & ~n16563 ) | ( n16396 & n16586 ) | ( ~n16563 & n16586 ) ;
  assign n16589 = ( ~n16396 & n16587 ) | ( ~n16396 & n16588 ) | ( n16587 & n16588 ) ;
  assign n16598 = ~n5135 & n16589 ;
  assign n16592 = n5010 | n16591 ;
  assign n16596 = n5067 | n16595 ;
  assign n16597 = n16592 &  n16596 ;
  assign n16599 = ( n5135 & n16598 ) | ( n5135 & n16597 ) | ( n16598 & n16597 ) ;
  assign n16603 = ( n16589 & n16595 ) | ( n16589 & n16601 ) | ( n16595 & n16601 ) ;
  assign n16602 = ( n16589 & ~n16595 ) | ( n16589 & n16601 ) | ( ~n16595 & n16601 ) ;
  assign n16604 = ( n16595 & ~n16603 ) | ( n16595 & n16602 ) | ( ~n16603 & n16602 ) ;
  assign n16605 = n5012 | n16604 ;
  assign n16606 = n16599 &  n16605 ;
  assign n16607 = x23 &  n16606 ;
  assign n16608 = x23 | n16606 ;
  assign n16609 = ~n16607 & n16608 ;
  assign n16783 = ( n16107 & ~n16782 ) | ( n16107 & n16609 ) | ( ~n16782 & n16609 ) ;
  assign n16784 = ( n16107 & ~n16609 ) | ( n16107 & n16782 ) | ( ~n16609 & n16782 ) ;
  assign n16785 = ( n16783 & ~n16107 ) | ( n16783 & n16784 ) | ( ~n16107 & n16784 ) ;
  assign n16786 = ( n16665 & ~n16662 ) | ( n16665 & n16778 ) | ( ~n16662 & n16778 ) ;
  assign n16787 = ( n16662 & ~n16778 ) | ( n16662 & n16665 ) | ( ~n16778 & n16665 ) ;
  assign n16788 = ( n16786 & ~n16665 ) | ( n16786 & n16787 ) | ( ~n16665 & n16787 ) ;
  assign n16792 = ~n5837 & n16595 ;
  assign n16789 = ( n5339 & ~n16091 ) | ( n5339 & 1'b0 ) | ( ~n16091 & 1'b0 ) ;
  assign n16790 = n5761 | n16591 ;
  assign n16791 = ~n16789 & n16790 ;
  assign n16793 = ( n5837 & n16792 ) | ( n5837 & n16791 ) | ( n16792 & n16791 ) ;
  assign n16794 = ( n5341 & ~n16616 ) | ( n5341 & n16793 ) | ( ~n16616 & n16793 ) ;
  assign n16795 = ~n5341 & n16794 ;
  assign n16797 = ( x20 & n16793 ) | ( x20 & n16795 ) | ( n16793 & n16795 ) ;
  assign n16796 = ( x20 & ~n16795 ) | ( x20 & n16793 ) | ( ~n16795 & n16793 ) ;
  assign n16798 = ( n16795 & ~n16797 ) | ( n16795 & n16796 ) | ( ~n16797 & n16796 ) ;
  assign n16802 = ~n5837 & n16591 ;
  assign n16799 = ( n5339 & ~n15897 ) | ( n5339 & 1'b0 ) | ( ~n15897 & 1'b0 ) ;
  assign n16800 = n5761 | n16091 ;
  assign n16801 = ~n16799 & n16800 ;
  assign n16803 = ( n5837 & n16802 ) | ( n5837 & n16801 ) | ( n16802 & n16801 ) ;
  assign n16804 = ( n5341 & ~n16631 ) | ( n5341 & n16803 ) | ( ~n16631 & n16803 ) ;
  assign n16805 = ~n5341 & n16804 ;
  assign n16806 = ( x20 & ~n16803 ) | ( x20 & n16805 ) | ( ~n16803 & n16805 ) ;
  assign n16807 = ( n16803 & ~x20 ) | ( n16803 & n16805 ) | ( ~x20 & n16805 ) ;
  assign n16808 = ( n16806 & ~n16805 ) | ( n16806 & n16807 ) | ( ~n16805 & n16807 ) ;
  assign n16809 = ( n16668 & ~n16678 ) | ( n16668 & n16777 ) | ( ~n16678 & n16777 ) ;
  assign n16810 = ( n16678 & ~n16778 ) | ( n16678 & n16809 ) | ( ~n16778 & n16809 ) ;
  assign n16814 = ~n5837 & n16091 ;
  assign n16811 = ( n5339 & ~n15700 ) | ( n5339 & 1'b0 ) | ( ~n15700 & 1'b0 ) ;
  assign n16812 = n5761 | n15897 ;
  assign n16813 = ~n16811 & n16812 ;
  assign n16815 = ( n5837 & n16814 ) | ( n5837 & n16813 ) | ( n16814 & n16813 ) ;
  assign n16816 = ( n5341 & ~n16094 ) | ( n5341 & n16815 ) | ( ~n16094 & n16815 ) ;
  assign n16817 = ~n5341 & n16816 ;
  assign n16818 = ( x20 & ~n16815 ) | ( x20 & n16817 ) | ( ~n16815 & n16817 ) ;
  assign n16819 = ( n16815 & ~x20 ) | ( n16815 & n16817 ) | ( ~x20 & n16817 ) ;
  assign n16820 = ( n16818 & ~n16817 ) | ( n16818 & n16819 ) | ( ~n16817 & n16819 ) ;
  assign n16821 = ( n16681 & ~n16691 ) | ( n16681 & n16776 ) | ( ~n16691 & n16776 ) ;
  assign n16822 = ( n16691 & ~n16777 ) | ( n16691 & n16821 ) | ( ~n16777 & n16821 ) ;
  assign n16829 = ~n5837 & n15897 ;
  assign n16826 = ( n5339 & ~n15320 ) | ( n5339 & 1'b0 ) | ( ~n15320 & 1'b0 ) ;
  assign n16827 = n5761 | n15700 ;
  assign n16828 = ~n16826 & n16827 ;
  assign n16830 = ( n5837 & n16829 ) | ( n5837 & n16828 ) | ( n16829 & n16828 ) ;
  assign n16831 = ( n15900 & ~n5341 ) | ( n15900 & n16830 ) | ( ~n5341 & n16830 ) ;
  assign n16832 = ~n15900 & n16831 ;
  assign n16833 = ( x20 & ~n16830 ) | ( x20 & n16832 ) | ( ~n16830 & n16832 ) ;
  assign n16834 = ( n16830 & ~x20 ) | ( n16830 & n16832 ) | ( ~x20 & n16832 ) ;
  assign n16835 = ( n16833 & ~n16832 ) | ( n16833 & n16834 ) | ( ~n16832 & n16834 ) ;
  assign n16823 = ( n16703 & ~n16701 ) | ( n16703 & n16775 ) | ( ~n16701 & n16775 ) ;
  assign n16824 = ( n16701 & ~n16775 ) | ( n16701 & n16703 ) | ( ~n16775 & n16703 ) ;
  assign n16825 = ( n16823 & ~n16703 ) | ( n16823 & n16824 ) | ( ~n16703 & n16824 ) ;
  assign n16836 = ( n16716 & ~n16706 ) | ( n16716 & n16774 ) | ( ~n16706 & n16774 ) ;
  assign n16837 = ( n16706 & ~n16774 ) | ( n16706 & n16716 ) | ( ~n16774 & n16716 ) ;
  assign n16838 = ( n16836 & ~n16716 ) | ( n16836 & n16837 ) | ( ~n16716 & n16837 ) ;
  assign n16842 = ~n5837 & n15700 ;
  assign n16839 = ( n5339 & ~n15325 ) | ( n5339 & 1'b0 ) | ( ~n15325 & 1'b0 ) ;
  assign n16840 = n5761 | n15320 ;
  assign n16841 = ~n16839 & n16840 ;
  assign n16843 = ( n5837 & n16842 ) | ( n5837 & n16841 ) | ( n16842 & n16841 ) ;
  assign n16844 = ( n15708 & ~n5341 ) | ( n15708 & n16843 ) | ( ~n5341 & n16843 ) ;
  assign n16845 = ~n15708 & n16844 ;
  assign n16847 = ( x20 & n16843 ) | ( x20 & n16845 ) | ( n16843 & n16845 ) ;
  assign n16846 = ( x20 & ~n16845 ) | ( x20 & n16843 ) | ( ~n16845 & n16843 ) ;
  assign n16848 = ( n16845 & ~n16847 ) | ( n16845 & n16846 ) | ( ~n16847 & n16846 ) ;
  assign n16849 = ( n16726 & ~n16773 ) | ( n16726 & n16731 ) | ( ~n16773 & n16731 ) ;
  assign n16850 = ( n16731 & ~n16726 ) | ( n16731 & n16773 ) | ( ~n16726 & n16773 ) ;
  assign n16851 = ( n16849 & ~n16731 ) | ( n16849 & n16850 ) | ( ~n16731 & n16850 ) ;
  assign n16855 = ~n5837 & n15320 ;
  assign n16852 = ( n5339 & ~n15322 ) | ( n5339 & 1'b0 ) | ( ~n15322 & 1'b0 ) ;
  assign n16853 = n5761 | n15325 ;
  assign n16854 = ~n16852 & n16853 ;
  assign n16856 = ( n5837 & n16855 ) | ( n5837 & n16854 ) | ( n16855 & n16854 ) ;
  assign n16857 = ( n15334 & ~n5341 ) | ( n15334 & n16856 ) | ( ~n5341 & n16856 ) ;
  assign n16858 = ~n15334 & n16857 ;
  assign n16859 = ( x20 & ~n16856 ) | ( x20 & n16858 ) | ( ~n16856 & n16858 ) ;
  assign n16860 = ( n16856 & ~x20 ) | ( n16856 & n16858 ) | ( ~x20 & n16858 ) ;
  assign n16861 = ( n16859 & ~n16858 ) | ( n16859 & n16860 ) | ( ~n16858 & n16860 ) ;
  assign n16865 = ~n5837 & n15325 ;
  assign n16862 = n5339 &  n14745 ;
  assign n16863 = n5761 | n15322 ;
  assign n16864 = ~n16862 & n16863 ;
  assign n16866 = ( n5837 & n16865 ) | ( n5837 & n16864 ) | ( n16865 & n16864 ) ;
  assign n16867 = n5341 | n15346 ;
  assign n16868 = n16866 &  n16867 ;
  assign n16869 = x20 &  n16868 ;
  assign n16870 = x20 | n16868 ;
  assign n16871 = ~n16869 & n16870 ;
  assign n16872 = ( n16745 & ~n16735 ) | ( n16745 & n16772 ) | ( ~n16735 & n16772 ) ;
  assign n16873 = ( n16773 & ~n16745 ) | ( n16773 & n16872 ) | ( ~n16745 & n16872 ) ;
  assign n16875 = ( n15476 & n16761 ) | ( n15476 & n16771 ) | ( n16761 & n16771 ) ;
  assign n16874 = ( n15476 & ~n16761 ) | ( n15476 & n16771 ) | ( ~n16761 & n16771 ) ;
  assign n16876 = ( n16761 & ~n16875 ) | ( n16761 & n16874 ) | ( ~n16875 & n16874 ) ;
  assign n16877 = ( n5339 & ~n14528 ) | ( n5339 & 1'b0 ) | ( ~n14528 & 1'b0 ) ;
  assign n16878 = ~n5761 & n14745 ;
  assign n16879 = n16877 | n16878 ;
  assign n16880 = ~n5837 & n15322 ;
  assign n16881 = ( n5837 & ~n16879 ) | ( n5837 & n16880 ) | ( ~n16879 & n16880 ) ;
  assign n16882 = ( n5341 & ~n16881 ) | ( n5341 & n15361 ) | ( ~n16881 & n15361 ) ;
  assign n16883 = ( n15361 & ~n16882 ) | ( n15361 & 1'b0 ) | ( ~n16882 & 1'b0 ) ;
  assign n16884 = ( x20 & ~n16881 ) | ( x20 & n16883 ) | ( ~n16881 & n16883 ) ;
  assign n16885 = ( n16881 & ~x20 ) | ( n16881 & n16883 ) | ( ~x20 & n16883 ) ;
  assign n16886 = ( n16884 & ~n16883 ) | ( n16884 & n16885 ) | ( ~n16883 & n16885 ) ;
  assign n16890 = n14745 | n5837 ;
  assign n16887 = ( n5339 & ~n14261 ) | ( n5339 & 1'b0 ) | ( ~n14261 & 1'b0 ) ;
  assign n16888 = n5761 | n14528 ;
  assign n16889 = ~n16887 & n16888 ;
  assign n16891 = ( n5837 & ~n16890 ) | ( n5837 & n16889 ) | ( ~n16890 & n16889 ) ;
  assign n16892 = ~n5341 & n14749 ;
  assign n16893 = ( n16891 & ~n16892 ) | ( n16891 & 1'b0 ) | ( ~n16892 & 1'b0 ) ;
  assign n16894 = x20 &  n16893 ;
  assign n16895 = x20 | n16893 ;
  assign n16896 = ~n16894 & n16895 ;
  assign n16897 = ( n16750 & ~x23 ) | ( n16750 & n16751 ) | ( ~x23 & n16751 ) ;
  assign n16898 = ( n16750 & ~n16897 ) | ( n16750 & 1'b0 ) | ( ~n16897 & 1'b0 ) ;
  assign n16899 = ( n16758 & ~x23 ) | ( n16758 & n16898 ) | ( ~x23 & n16898 ) ;
  assign n16900 = ( x23 & ~n16758 ) | ( x23 & n16898 ) | ( ~n16758 & n16898 ) ;
  assign n16901 = ( n16899 & ~n16898 ) | ( n16899 & n16900 ) | ( ~n16898 & n16900 ) ;
  assign n16902 = x23 &  n16751 ;
  assign n16903 = ~n16750 & n16902 ;
  assign n16904 = ( n16750 & ~n16902 ) | ( n16750 & 1'b0 ) | ( ~n16902 & 1'b0 ) ;
  assign n16905 = n16903 | n16904 ;
  assign n16932 = ( n5339 & ~n13785 ) | ( n5339 & 1'b0 ) | ( ~n13785 & 1'b0 ) ;
  assign n16933 = n5761 | n13998 ;
  assign n16934 = ~n16932 & n16933 ;
  assign n16935 = ~n5837 & n14261 ;
  assign n16936 = ( n5837 & n16934 ) | ( n5837 & n16935 ) | ( n16934 & n16935 ) ;
  assign n16937 = n5341 | n14267 ;
  assign n16938 = n16936 &  n16937 ;
  assign n16939 = x20 &  n16938 ;
  assign n16940 = x20 | n16938 ;
  assign n16941 = ~n16939 & n16940 ;
  assign n16916 = ( n5337 & ~n13787 ) | ( n5337 & 1'b0 ) | ( ~n13787 & 1'b0 ) ;
  assign n16920 = n13790 | n5341 ;
  assign n16917 = n5761 | n13787 ;
  assign n16918 = n5837 | n13785 ;
  assign n16919 = n16917 &  n16918 ;
  assign n16921 = ( n5341 & ~n16920 ) | ( n5341 & n16919 ) | ( ~n16920 & n16919 ) ;
  assign n16927 = ~n5341 & n14001 ;
  assign n16925 = ~n5837 & n13998 ;
  assign n16922 = ( n5339 & ~n13787 ) | ( n5339 & 1'b0 ) | ( ~n13787 & 1'b0 ) ;
  assign n16923 = n5761 | n13785 ;
  assign n16924 = ~n16922 & n16923 ;
  assign n16926 = ( n5837 & n16925 ) | ( n5837 & n16924 ) | ( n16925 & n16924 ) ;
  assign n16928 = ( n5341 & n16927 ) | ( n5341 & n16926 ) | ( n16927 & n16926 ) ;
  assign n16929 = ( n16916 & n16921 ) | ( n16916 & n16928 ) | ( n16921 & n16928 ) ;
  assign n16930 = ( x20 & ~n16929 ) | ( x20 & n16916 ) | ( ~n16929 & n16916 ) ;
  assign n16931 = ( x20 & ~n16930 ) | ( x20 & 1'b0 ) | ( ~n16930 & 1'b0 ) ;
  assign n16942 = ( n16751 & ~n16941 ) | ( n16751 & n16931 ) | ( ~n16941 & n16931 ) ;
  assign n16909 = ~n5837 & n14528 ;
  assign n16906 = ( n5339 & ~n13998 ) | ( n5339 & 1'b0 ) | ( ~n13998 & 1'b0 ) ;
  assign n16907 = n5761 | n14261 ;
  assign n16908 = ~n16906 & n16907 ;
  assign n16910 = ( n5837 & n16909 ) | ( n5837 & n16908 ) | ( n16909 & n16908 ) ;
  assign n16911 = ( n14532 & ~n5341 ) | ( n14532 & n16910 ) | ( ~n5341 & n16910 ) ;
  assign n16912 = ~n14532 & n16911 ;
  assign n16913 = ( x20 & ~n16910 ) | ( x20 & n16912 ) | ( ~n16910 & n16912 ) ;
  assign n16914 = ( n16910 & ~x20 ) | ( n16910 & n16912 ) | ( ~x20 & n16912 ) ;
  assign n16915 = ( n16913 & ~n16912 ) | ( n16913 & n16914 ) | ( ~n16912 & n16914 ) ;
  assign n16943 = ( n16905 & ~n16942 ) | ( n16905 & n16915 ) | ( ~n16942 & n16915 ) ;
  assign n16944 = ( n16896 & n16901 ) | ( n16896 & n16943 ) | ( n16901 & n16943 ) ;
  assign n16945 = ( n16876 & n16886 ) | ( n16876 & n16944 ) | ( n16886 & n16944 ) ;
  assign n16946 = ( n16871 & ~n16873 ) | ( n16871 & n16945 ) | ( ~n16873 & n16945 ) ;
  assign n16947 = ( n16851 & n16861 ) | ( n16851 & n16946 ) | ( n16861 & n16946 ) ;
  assign n16948 = ( n16838 & n16848 ) | ( n16838 & n16947 ) | ( n16848 & n16947 ) ;
  assign n16949 = ( n16835 & ~n16825 ) | ( n16835 & n16948 ) | ( ~n16825 & n16948 ) ;
  assign n16950 = ( n16820 & n16822 ) | ( n16820 & n16949 ) | ( n16822 & n16949 ) ;
  assign n16951 = ( n16808 & n16810 ) | ( n16808 & n16950 ) | ( n16810 & n16950 ) ;
  assign n16952 = ( n16788 & n16798 ) | ( n16788 & n16951 ) | ( n16798 & n16951 ) ;
  assign n16953 = ( n16649 & ~n16779 ) | ( n16649 & n16652 ) | ( ~n16779 & n16652 ) ;
  assign n16954 = ( n16652 & ~n16649 ) | ( n16652 & n16779 ) | ( ~n16649 & n16779 ) ;
  assign n16955 = ( n16953 & ~n16652 ) | ( n16953 & n16954 ) | ( ~n16652 & n16954 ) ;
  assign n16959 = ~n5837 & n16589 ;
  assign n16956 = ( n5339 & ~n16591 ) | ( n5339 & 1'b0 ) | ( ~n16591 & 1'b0 ) ;
  assign n16957 = n5761 | n16595 ;
  assign n16958 = ~n16956 & n16957 ;
  assign n16960 = ( n5837 & n16959 ) | ( n5837 & n16958 ) | ( n16959 & n16958 ) ;
  assign n16961 = ( n5341 & ~n16604 ) | ( n5341 & n16960 ) | ( ~n16604 & n16960 ) ;
  assign n16962 = ~n5341 & n16961 ;
  assign n16964 = ( x20 & n16960 ) | ( x20 & n16962 ) | ( n16960 & n16962 ) ;
  assign n16963 = ( x20 & ~n16962 ) | ( x20 & n16960 ) | ( ~n16962 & n16960 ) ;
  assign n16965 = ( n16962 & ~n16964 ) | ( n16962 & n16963 ) | ( ~n16964 & n16963 ) ;
  assign n16966 = ( n16952 & ~n16955 ) | ( n16952 & n16965 ) | ( ~n16955 & n16965 ) ;
  assign n16967 = ( n16639 & ~n16636 ) | ( n16639 & n16780 ) | ( ~n16636 & n16780 ) ;
  assign n16968 = ( n16636 & ~n16780 ) | ( n16636 & n16639 ) | ( ~n16780 & n16639 ) ;
  assign n16969 = ( n16967 & ~n16639 ) | ( n16967 & n16968 ) | ( ~n16639 & n16968 ) ;
  assign n16970 = ( n16467 & ~n16466 ) | ( n16467 & n16477 ) | ( ~n16466 & n16477 ) ;
  assign n17000 = ( n16301 & ~n16453 ) | ( n16301 & n16463 ) | ( ~n16453 & n16463 ) ;
  assign n16972 = n235 | n2091 ;
  assign n16973 = n229 | n16972 ;
  assign n16974 = n1498 | n5552 ;
  assign n16975 = ( n16973 & ~n2960 ) | ( n16973 & n16974 ) | ( ~n2960 & n16974 ) ;
  assign n16976 = n2960 | n16975 ;
  assign n16977 = ( n128 & ~n1221 ) | ( n128 & n16976 ) | ( ~n1221 & n16976 ) ;
  assign n16978 = ( n1221 & n2878 ) | ( n1221 & n16977 ) | ( n2878 & n16977 ) ;
  assign n16979 = ( n2878 & ~n16978 ) | ( n2878 & 1'b0 ) | ( ~n16978 & 1'b0 ) ;
  assign n16980 = ( n575 & ~n16979 ) | ( n575 & n1163 ) | ( ~n16979 & n1163 ) ;
  assign n16981 = ( n1163 & ~n16980 ) | ( n1163 & 1'b0 ) | ( ~n16980 & 1'b0 ) ;
  assign n16982 = ( n604 & n2731 ) | ( n604 & n16981 ) | ( n2731 & n16981 ) ;
  assign n16983 = ~n604 & n16982 ;
  assign n16984 = ( n243 & ~n345 ) | ( n243 & n16983 ) | ( ~n345 & n16983 ) ;
  assign n16985 = ~n243 & n16984 ;
  assign n16986 = ( n678 & ~n193 ) | ( n678 & n16985 ) | ( ~n193 & n16985 ) ;
  assign n16987 = ~n678 & n16986 ;
  assign n16988 = ( n169 & ~n627 ) | ( n169 & n16987 ) | ( ~n627 & n16987 ) ;
  assign n16989 = ~n169 & n16988 ;
  assign n16971 = ( n16446 & ~n16439 ) | ( n16446 & n16450 ) | ( ~n16439 & n16450 ) ;
  assign n16991 = ( n16439 & n16971 ) | ( n16439 & n16989 ) | ( n16971 & n16989 ) ;
  assign n16990 = ( n16439 & ~n16989 ) | ( n16439 & n16971 ) | ( ~n16989 & n16971 ) ;
  assign n16992 = ( n16989 & ~n16991 ) | ( n16989 & n16990 ) | ( ~n16991 & n16990 ) ;
  assign n16993 = n3644 | n11871 ;
  assign n16994 = n3652 &  n11134 ;
  assign n16995 = ( n3657 & ~n11131 ) | ( n3657 & 1'b0 ) | ( ~n11131 & 1'b0 ) ;
  assign n16996 = n16994 | n16995 ;
  assign n16997 = ~n3653 & n11128 ;
  assign n16998 = ( n3653 & ~n16996 ) | ( n3653 & n16997 ) | ( ~n16996 & n16997 ) ;
  assign n16999 = n16993 &  n16998 ;
  assign n17001 = ( n16992 & n16999 ) | ( n16992 & n17000 ) | ( n16999 & n17000 ) ;
  assign n17002 = ( n16992 & ~n17000 ) | ( n16992 & n16999 ) | ( ~n17000 & n16999 ) ;
  assign n17003 = ( n17000 & ~n17001 ) | ( n17000 & n17002 ) | ( ~n17001 & n17002 ) ;
  assign n17004 = n4430 &  n11119 ;
  assign n17005 = ~n523 & n11125 ;
  assign n17006 = n3939 | n11122 ;
  assign n17007 = ~n17005 & n17006 ;
  assign n17008 = ( n17004 & ~n11119 ) | ( n17004 & n17007 ) | ( ~n11119 & n17007 ) ;
  assign n17009 = ~n601 & n12088 ;
  assign n17010 = ( n17008 & ~n17009 ) | ( n17008 & 1'b0 ) | ( ~n17009 & 1'b0 ) ;
  assign n17011 = x29 &  n17010 ;
  assign n17012 = x29 | n17010 ;
  assign n17013 = ~n17011 & n17012 ;
  assign n17017 = ~n4962 & n11110 ;
  assign n17014 = ~n4482 & n11116 ;
  assign n17015 = n4495 | n11113 ;
  assign n17016 = ~n17014 & n17015 ;
  assign n17018 = ( n4962 & n17017 ) | ( n4962 & n17016 ) | ( n17017 & n17016 ) ;
  assign n17019 = ~n4478 & n12352 ;
  assign n17020 = ( n17018 & ~n17019 ) | ( n17018 & 1'b0 ) | ( ~n17019 & 1'b0 ) ;
  assign n17021 = x26 &  n17020 ;
  assign n17022 = x26 | n17020 ;
  assign n17023 = ~n17021 & n17022 ;
  assign n17025 = ( n17003 & n17013 ) | ( n17003 & n17023 ) | ( n17013 & n17023 ) ;
  assign n17024 = ( n17013 & ~n17003 ) | ( n17013 & n17023 ) | ( ~n17003 & n17023 ) ;
  assign n17026 = ( n17003 & ~n17025 ) | ( n17003 & n17024 ) | ( ~n17025 & n17024 ) ;
  assign n17030 = ~n5135 & n11101 ;
  assign n17027 = ~n5010 & n11107 ;
  assign n17028 = n5067 | n11104 ;
  assign n17029 = ~n17027 & n17028 ;
  assign n17031 = ( n5135 & n17030 ) | ( n5135 & n17029 ) | ( n17030 & n17029 ) ;
  assign n17032 = n5012 | n12650 ;
  assign n17033 = n17031 &  n17032 ;
  assign n17034 = x23 &  n17033 ;
  assign n17035 = x23 | n17033 ;
  assign n17036 = ~n17034 & n17035 ;
  assign n17037 = ( n16970 & n17026 ) | ( n16970 & n17036 ) | ( n17026 & n17036 ) ;
  assign n17038 = ( n17026 & ~n16970 ) | ( n17026 & n17036 ) | ( ~n16970 & n17036 ) ;
  assign n17039 = ( n16970 & ~n17037 ) | ( n16970 & n17038 ) | ( ~n17037 & n17038 ) ;
  assign n17040 = ( n5339 & ~n11098 ) | ( n5339 & 1'b0 ) | ( ~n11098 & 1'b0 ) ;
  assign n17041 = n5761 | n11095 ;
  assign n17042 = ~n17040 & n17041 ;
  assign n17043 = ~n5837 & n11093 ;
  assign n17044 = ( n5837 & n17042 ) | ( n5837 & n17043 ) | ( n17042 & n17043 ) ;
  assign n17045 = n5341 | n12997 ;
  assign n17046 = n17044 &  n17045 ;
  assign n17047 = x20 &  n17046 ;
  assign n17048 = x20 | n17046 ;
  assign n17049 = ~n17047 & n17048 ;
  assign n17051 = ( n16491 & n17039 ) | ( n16491 & n17049 ) | ( n17039 & n17049 ) ;
  assign n17050 = ( n16491 & ~n17039 ) | ( n16491 & n17049 ) | ( ~n17039 & n17049 ) ;
  assign n17052 = ( n17039 & ~n17051 ) | ( n17039 & n17050 ) | ( ~n17051 & n17050 ) ;
  assign n17056 = ~n6395 & n11085 ;
  assign n17053 = n5970 | n11091 ;
  assign n17054 = n6170 | n11081 ;
  assign n17055 = n17053 &  n17054 ;
  assign n17057 = ( n6395 & n17056 ) | ( n6395 & n17055 ) | ( n17056 & n17055 ) ;
  assign n17058 = n5972 | n13377 ;
  assign n17059 = n17057 &  n17058 ;
  assign n17060 = x17 &  n17059 ;
  assign n17061 = x17 | n17059 ;
  assign n17062 = ~n17060 & n17061 ;
  assign n17064 = ( n16505 & n17052 ) | ( n16505 & n17062 ) | ( n17052 & n17062 ) ;
  assign n17063 = ( n16505 & ~n17052 ) | ( n16505 & n17062 ) | ( ~n17052 & n17062 ) ;
  assign n17065 = ( n17052 & ~n17064 ) | ( n17052 & n17063 ) | ( ~n17064 & n17063 ) ;
  assign n17069 = ~n7097 & n14071 ;
  assign n17066 = n6530 | n11078 ;
  assign n17067 = n6983 | n13836 ;
  assign n17068 = n17066 &  n17067 ;
  assign n17070 = ( n7097 & n17069 ) | ( n7097 & n17068 ) | ( n17069 & n17068 ) ;
  assign n17071 = n6532 | n14079 ;
  assign n17072 = n17070 &  n17071 ;
  assign n17073 = x14 &  n17072 ;
  assign n17074 = x14 | n17072 ;
  assign n17075 = ~n17073 & n17074 ;
  assign n17076 = ( n16519 & n17065 ) | ( n16519 & n17075 ) | ( n17065 & n17075 ) ;
  assign n17077 = ( n17065 & ~n16519 ) | ( n17065 & n17075 ) | ( ~n16519 & n17075 ) ;
  assign n17078 = ( n16519 & ~n17076 ) | ( n16519 & n17077 ) | ( ~n17076 & n17077 ) ;
  assign n17079 = ( n7253 & ~n14355 ) | ( n7253 & 1'b0 ) | ( ~n14355 & 1'b0 ) ;
  assign n17080 = ~n7518 & n14553 ;
  assign n17081 = n17079 | n17080 ;
  assign n17082 = ~n7783 & n14803 ;
  assign n17083 = ( n7783 & ~n17081 ) | ( n7783 & n17082 ) | ( ~n17081 & n17082 ) ;
  assign n17084 = ~n7255 & n15310 ;
  assign n17085 = ( n17083 & ~n17084 ) | ( n17083 & 1'b0 ) | ( ~n17084 & 1'b0 ) ;
  assign n17086 = x11 &  n17085 ;
  assign n17087 = x11 | n17085 ;
  assign n17088 = ~n17086 & n17087 ;
  assign n17090 = ( n16533 & n17078 ) | ( n16533 & n17088 ) | ( n17078 & n17088 ) ;
  assign n17089 = ( n16533 & ~n17078 ) | ( n16533 & n17088 ) | ( ~n17078 & n17088 ) ;
  assign n17091 = ( n17078 & ~n17090 ) | ( n17078 & n17089 ) | ( ~n17090 & n17089 ) ;
  assign n17092 = n8429 &  n8764 ;
  assign n17093 = ( n14800 & ~n17092 ) | ( n14800 & 1'b0 ) | ( ~n17092 & 1'b0 ) ;
  assign n17094 = n8105 &  n14807 ;
  assign n17095 = n17093 | n17094 ;
  assign n17096 = ( n8107 & n15692 ) | ( n8107 & n17095 ) | ( n15692 & n17095 ) ;
  assign n17097 = ( n15692 & ~n17096 ) | ( n15692 & 1'b0 ) | ( ~n17096 & 1'b0 ) ;
  assign n17098 = ( n17095 & ~x8 ) | ( n17095 & n17097 ) | ( ~x8 & n17097 ) ;
  assign n17099 = ( x8 & ~n17095 ) | ( x8 & n17097 ) | ( ~n17095 & n17097 ) ;
  assign n17100 = ( n17098 & ~n17097 ) | ( n17098 & n17099 ) | ( ~n17097 & n17099 ) ;
  assign n17101 = ( n16547 & n17091 ) | ( n16547 & n17100 ) | ( n17091 & n17100 ) ;
  assign n17102 = ( n17091 & ~n16547 ) | ( n17091 & n17100 ) | ( ~n16547 & n17100 ) ;
  assign n17103 = ( n16547 & ~n17101 ) | ( n16547 & n17102 ) | ( ~n17101 & n17102 ) ;
  assign n17104 = ( n16563 & ~n16396 ) | ( n16563 & n16586 ) | ( ~n16396 & n16586 ) ;
  assign n17105 = ( n16561 & ~n17103 ) | ( n16561 & n17104 ) | ( ~n17103 & n17104 ) ;
  assign n17106 = ( n16561 & ~n17104 ) | ( n16561 & n17103 ) | ( ~n17104 & n17103 ) ;
  assign n17107 = ( n17105 & ~n16561 ) | ( n17105 & n17106 ) | ( ~n16561 & n17106 ) ;
  assign n17111 = n17107 | n5837 ;
  assign n17108 = ( n5339 & ~n16595 ) | ( n5339 & 1'b0 ) | ( ~n16595 & 1'b0 ) ;
  assign n17109 = n5761 | n16589 ;
  assign n17110 = ~n17108 & n17109 ;
  assign n17112 = ( n5837 & ~n17111 ) | ( n5837 & n17110 ) | ( ~n17111 & n17110 ) ;
  assign n17113 = ( n16589 & ~n16603 ) | ( n16589 & n17107 ) | ( ~n16603 & n17107 ) ;
  assign n17114 = ( n16589 & ~n17107 ) | ( n16589 & n16603 ) | ( ~n17107 & n16603 ) ;
  assign n17115 = ( n17113 & ~n16589 ) | ( n17113 & n17114 ) | ( ~n16589 & n17114 ) ;
  assign n17116 = ( n5341 & ~n17112 ) | ( n5341 & n17115 ) | ( ~n17112 & n17115 ) ;
  assign n17117 = ( n17115 & ~n17116 ) | ( n17115 & 1'b0 ) | ( ~n17116 & 1'b0 ) ;
  assign n17118 = ( x20 & ~n17112 ) | ( x20 & n17117 ) | ( ~n17112 & n17117 ) ;
  assign n17119 = ( n17112 & ~x20 ) | ( n17112 & n17117 ) | ( ~x20 & n17117 ) ;
  assign n17120 = ( n17118 & ~n17117 ) | ( n17118 & n17119 ) | ( ~n17117 & n17119 ) ;
  assign n17121 = ( n16966 & n16969 ) | ( n16966 & n17120 ) | ( n16969 & n17120 ) ;
  assign n17122 = ( n16624 & ~n16621 ) | ( n16624 & n16781 ) | ( ~n16621 & n16781 ) ;
  assign n17123 = ( n16621 & ~n16781 ) | ( n16621 & n16624 ) | ( ~n16781 & n16624 ) ;
  assign n17124 = ( n17122 & ~n16624 ) | ( n17122 & n17123 ) | ( ~n16624 & n17123 ) ;
  assign n17254 = ( n16519 & ~n17065 ) | ( n16519 & n17075 ) | ( ~n17065 & n17075 ) ;
  assign n17148 = ~n5135 & n11098 ;
  assign n17145 = n5010 | n11104 ;
  assign n17146 = n5067 | n11101 ;
  assign n17147 = n17145 &  n17146 ;
  assign n17149 = ( n5135 & n17148 ) | ( n5135 & n17147 ) | ( n17148 & n17147 ) ;
  assign n17150 = n5012 | n11218 ;
  assign n17151 = n17149 &  n17150 ;
  assign n17152 = x23 &  n17151 ;
  assign n17153 = x23 | n17151 ;
  assign n17154 = ~n17152 & n17153 ;
  assign n17168 = n11116 | n4430 ;
  assign n17165 = n523 | n11122 ;
  assign n17166 = ~n3939 & n11119 ;
  assign n17167 = ( n17165 & ~n17166 ) | ( n17165 & 1'b0 ) | ( ~n17166 & 1'b0 ) ;
  assign n17169 = ( n4430 & ~n17168 ) | ( n4430 & n17167 ) | ( ~n17168 & n17167 ) ;
  assign n17170 = n601 | n11230 ;
  assign n17171 = n17169 &  n17170 ;
  assign n17172 = x29 &  n17171 ;
  assign n17173 = x29 | n17171 ;
  assign n17174 = ~n17172 & n17173 ;
  assign n17175 = ( n16971 & ~n16439 ) | ( n16971 & n16989 ) | ( ~n16439 & n16989 ) ;
  assign n17176 = ~n3644 & n11859 ;
  assign n17180 = n11125 | n3653 ;
  assign n17177 = ( n3652 & ~n11131 ) | ( n3652 & 1'b0 ) | ( ~n11131 & 1'b0 ) ;
  assign n17178 = ( n3657 & ~n11128 ) | ( n3657 & 1'b0 ) | ( ~n11128 & 1'b0 ) ;
  assign n17179 = n17177 | n17178 ;
  assign n17181 = ( n17180 & ~n3653 ) | ( n17180 & n17179 ) | ( ~n3653 & n17179 ) ;
  assign n17182 = n17176 | n17181 ;
  assign n17183 = ( n8100 & ~n8097 ) | ( n8100 & n8103 ) | ( ~n8097 & n8103 ) ;
  assign n17184 = n8097 | n17183 ;
  assign n17185 = n14800 &  n17184 ;
  assign n17186 = n272 | n531 ;
  assign n17187 = n214 | n17186 ;
  assign n17188 = ( n127 & ~n243 ) | ( n127 & n17187 ) | ( ~n243 & n17187 ) ;
  assign n17189 = n243 | n17188 ;
  assign n17190 = ( n123 & ~n169 ) | ( n123 & n17189 ) | ( ~n169 & n17189 ) ;
  assign n17191 = n169 | n17190 ;
  assign n17192 = n990 | n2766 ;
  assign n17193 = ( n5428 & ~n1731 ) | ( n5428 & n17192 ) | ( ~n1731 & n17192 ) ;
  assign n17194 = n1731 | n17193 ;
  assign n17195 = ( n2593 & ~n17194 ) | ( n2593 & n3872 ) | ( ~n17194 & n3872 ) ;
  assign n17196 = ~n2593 & n17195 ;
  assign n17197 = ( n14281 & ~n2059 ) | ( n14281 & n17196 ) | ( ~n2059 & n17196 ) ;
  assign n17198 = n2059 &  n17197 ;
  assign n17199 = ( n17191 & ~n1306 ) | ( n17191 & n17198 ) | ( ~n1306 & n17198 ) ;
  assign n17200 = ( n1484 & ~n17191 ) | ( n1484 & n17199 ) | ( ~n17191 & n17199 ) ;
  assign n17201 = ~n1484 & n17200 ;
  assign n17202 = ( n69 & ~n345 ) | ( n69 & n17201 ) | ( ~n345 & n17201 ) ;
  assign n17203 = ~n69 & n17202 ;
  assign n17204 = ( n165 & ~n91 ) | ( n165 & n17203 ) | ( ~n91 & n17203 ) ;
  assign n17205 = ~n165 & n17204 ;
  assign n17206 = ( n17205 & ~n43 ) | ( n17205 & n454 ) | ( ~n43 & n454 ) ;
  assign n17207 = ( n17206 & ~n454 ) | ( n17206 & 1'b0 ) | ( ~n454 & 1'b0 ) ;
  assign n17208 = n16439 | n17207 ;
  assign n17209 = n16439 &  n17207 ;
  assign n17210 = ( n17208 & ~n17209 ) | ( n17208 & 1'b0 ) | ( ~n17209 & 1'b0 ) ;
  assign n17211 = ( n17185 & ~x8 ) | ( n17185 & n17210 ) | ( ~x8 & n17210 ) ;
  assign n17212 = ( x8 & ~n17210 ) | ( x8 & n17185 ) | ( ~n17210 & n17185 ) ;
  assign n17213 = ( n17211 & ~n17185 ) | ( n17211 & n17212 ) | ( ~n17185 & n17212 ) ;
  assign n17215 = ( n17175 & n17182 ) | ( n17175 & n17213 ) | ( n17182 & n17213 ) ;
  assign n17214 = ( n17182 & ~n17175 ) | ( n17182 & n17213 ) | ( ~n17175 & n17213 ) ;
  assign n17216 = ( n17175 & ~n17215 ) | ( n17175 & n17214 ) | ( ~n17215 & n17214 ) ;
  assign n17217 = ( n16999 & ~n16992 ) | ( n16999 & n17000 ) | ( ~n16992 & n17000 ) ;
  assign n17218 = ( n17174 & n17216 ) | ( n17174 & n17217 ) | ( n17216 & n17217 ) ;
  assign n17219 = ( n17216 & ~n17174 ) | ( n17216 & n17217 ) | ( ~n17174 & n17217 ) ;
  assign n17220 = ( n17174 & ~n17218 ) | ( n17174 & n17219 ) | ( ~n17218 & n17219 ) ;
  assign n17158 = n11107 | n4962 ;
  assign n17155 = n4482 | n11113 ;
  assign n17156 = n4495 | n11110 ;
  assign n17157 = n17155 &  n17156 ;
  assign n17159 = ( n4962 & ~n17158 ) | ( n4962 & n17157 ) | ( ~n17158 & n17157 ) ;
  assign n17160 = ~n4478 & n12340 ;
  assign n17161 = ( n17159 & ~n17160 ) | ( n17159 & 1'b0 ) | ( ~n17160 & 1'b0 ) ;
  assign n17162 = x26 &  n17161 ;
  assign n17163 = x26 | n17161 ;
  assign n17164 = ~n17162 & n17163 ;
  assign n17221 = ( n17024 & ~n17220 ) | ( n17024 & n17164 ) | ( ~n17220 & n17164 ) ;
  assign n17222 = ( n17164 & ~n17024 ) | ( n17164 & n17220 ) | ( ~n17024 & n17220 ) ;
  assign n17223 = ( n17221 & ~n17164 ) | ( n17221 & n17222 ) | ( ~n17164 & n17222 ) ;
  assign n17224 = ( n16970 & ~n17026 ) | ( n16970 & n17036 ) | ( ~n17026 & n17036 ) ;
  assign n17225 = ( n17154 & ~n17223 ) | ( n17154 & n17224 ) | ( ~n17223 & n17224 ) ;
  assign n17226 = ( n17154 & ~n17224 ) | ( n17154 & n17223 ) | ( ~n17224 & n17223 ) ;
  assign n17227 = ( n17225 & ~n17154 ) | ( n17225 & n17226 ) | ( ~n17154 & n17226 ) ;
  assign n17138 = ~n5837 & n11091 ;
  assign n17135 = ( n5339 & ~n11095 ) | ( n5339 & 1'b0 ) | ( ~n11095 & 1'b0 ) ;
  assign n17136 = n5761 | n11093 ;
  assign n17137 = ~n17135 & n17136 ;
  assign n17139 = ( n5837 & n17138 ) | ( n5837 & n17137 ) | ( n17138 & n17137 ) ;
  assign n17140 = n5341 | n12984 ;
  assign n17141 = n17139 &  n17140 ;
  assign n17142 = x20 &  n17141 ;
  assign n17143 = x20 | n17141 ;
  assign n17144 = ~n17142 & n17143 ;
  assign n17228 = ( n17050 & ~n17227 ) | ( n17050 & n17144 ) | ( ~n17227 & n17144 ) ;
  assign n17229 = ( n17144 & ~n17050 ) | ( n17144 & n17227 ) | ( ~n17050 & n17227 ) ;
  assign n17230 = ( n17228 & ~n17144 ) | ( n17228 & n17229 ) | ( ~n17144 & n17229 ) ;
  assign n17234 = ~n6395 & n11078 ;
  assign n17231 = n5970 | n11081 ;
  assign n17232 = n6170 | n11085 ;
  assign n17233 = n17231 &  n17232 ;
  assign n17235 = ( n6395 & n17234 ) | ( n6395 & n17233 ) | ( n17234 & n17233 ) ;
  assign n17236 = n5972 | n11206 ;
  assign n17237 = n17235 &  n17236 ;
  assign n17238 = x17 &  n17237 ;
  assign n17239 = x17 | n17237 ;
  assign n17240 = ~n17238 & n17239 ;
  assign n17241 = ( n17063 & n17230 ) | ( n17063 & n17240 ) | ( n17230 & n17240 ) ;
  assign n17242 = ( n17230 & ~n17063 ) | ( n17230 & n17240 ) | ( ~n17063 & n17240 ) ;
  assign n17243 = ( n17063 & ~n17241 ) | ( n17063 & n17242 ) | ( ~n17241 & n17242 ) ;
  assign n17247 = ~n7097 & n14355 ;
  assign n17244 = n6530 | n13836 ;
  assign n17245 = n6983 | n14071 ;
  assign n17246 = n17244 &  n17245 ;
  assign n17248 = ( n7097 & n17247 ) | ( n7097 & n17246 ) | ( n17247 & n17246 ) ;
  assign n17249 = n6532 | n14363 ;
  assign n17250 = n17248 &  n17249 ;
  assign n17251 = x14 &  n17250 ;
  assign n17252 = x14 | n17250 ;
  assign n17253 = ~n17251 & n17252 ;
  assign n17255 = ( n17243 & n17253 ) | ( n17243 & n17254 ) | ( n17253 & n17254 ) ;
  assign n17256 = ( n17243 & ~n17254 ) | ( n17243 & n17253 ) | ( ~n17254 & n17253 ) ;
  assign n17257 = ( n17254 & ~n17255 ) | ( n17254 & n17256 ) | ( ~n17255 & n17256 ) ;
  assign n17128 = n7783 | n14807 ;
  assign n17125 = n7253 &  n14553 ;
  assign n17126 = n7518 | n14803 ;
  assign n17127 = ~n17125 & n17126 ;
  assign n17129 = ( n7783 & ~n17128 ) | ( n7783 & n17127 ) | ( ~n17128 & n17127 ) ;
  assign n17130 = ~n7255 & n15294 ;
  assign n17131 = ( n17129 & ~n17130 ) | ( n17129 & 1'b0 ) | ( ~n17130 & 1'b0 ) ;
  assign n17132 = x11 &  n17131 ;
  assign n17133 = x11 | n17131 ;
  assign n17134 = ~n17132 & n17133 ;
  assign n17258 = ( n17089 & n17134 ) | ( n17089 & n17257 ) | ( n17134 & n17257 ) ;
  assign n17259 = ( n17089 & ~n17257 ) | ( n17089 & n17134 ) | ( ~n17257 & n17134 ) ;
  assign n17260 = ( n17257 & ~n17258 ) | ( n17257 & n17259 ) | ( ~n17258 & n17259 ) ;
  assign n17261 = ( n17102 & n17106 ) | ( n17102 & n17260 ) | ( n17106 & n17260 ) ;
  assign n17262 = ( n17102 & ~n17260 ) | ( n17102 & n17106 ) | ( ~n17260 & n17106 ) ;
  assign n17263 = ( n17260 & ~n17261 ) | ( n17260 & n17262 ) | ( ~n17261 & n17262 ) ;
  assign n17269 = ( n17107 & n17114 ) | ( n17107 & n17263 ) | ( n17114 & n17263 ) ;
  assign n17270 = ( n17114 & ~n17107 ) | ( n17114 & n17263 ) | ( ~n17107 & n17263 ) ;
  assign n17271 = ( n17107 & ~n17269 ) | ( n17107 & n17270 ) | ( ~n17269 & n17270 ) ;
  assign n17264 = ( n5339 & ~n16589 ) | ( n5339 & 1'b0 ) | ( ~n16589 & 1'b0 ) ;
  assign n17265 = ~n5761 & n17107 ;
  assign n17266 = n17264 | n17265 ;
  assign n17267 = ~n5837 & n17263 ;
  assign n17268 = ( n5837 & ~n17266 ) | ( n5837 & n17267 ) | ( ~n17266 & n17267 ) ;
  assign n17272 = ( n5341 & ~n17268 ) | ( n5341 & n17271 ) | ( ~n17268 & n17271 ) ;
  assign n17273 = ( n17271 & ~n17272 ) | ( n17271 & 1'b0 ) | ( ~n17272 & 1'b0 ) ;
  assign n17275 = ( x20 & n17268 ) | ( x20 & n17273 ) | ( n17268 & n17273 ) ;
  assign n17274 = ( x20 & ~n17273 ) | ( x20 & n17268 ) | ( ~n17273 & n17268 ) ;
  assign n17276 = ( n17273 & ~n17275 ) | ( n17273 & n17274 ) | ( ~n17275 & n17274 ) ;
  assign n17277 = ( n17121 & n17124 ) | ( n17121 & n17276 ) | ( n17124 & n17276 ) ;
  assign n17402 = ( n17102 & ~n17106 ) | ( n17102 & n17260 ) | ( ~n17106 & n17260 ) ;
  assign n17278 = ( n17253 & ~n17243 ) | ( n17253 & n17254 ) | ( ~n17243 & n17254 ) ;
  assign n17279 = ( n17063 & ~n17230 ) | ( n17063 & n17240 ) | ( ~n17230 & n17240 ) ;
  assign n17280 = ( n17175 & ~n17182 ) | ( n17175 & n17213 ) | ( ~n17182 & n17213 ) ;
  assign n17281 = n2786 | n3729 ;
  assign n17282 = ( n1343 & n4689 ) | ( n1343 & n17281 ) | ( n4689 & n17281 ) ;
  assign n17283 = ( n1343 & ~n17282 ) | ( n1343 & 1'b0 ) | ( ~n17282 & 1'b0 ) ;
  assign n17284 = n15599 &  n17283 ;
  assign n17285 = ( n6289 & ~n17284 ) | ( n6289 & n16274 ) | ( ~n17284 & n16274 ) ;
  assign n17286 = ( n3492 & ~n16274 ) | ( n3492 & n17285 ) | ( ~n16274 & n17285 ) ;
  assign n17287 = ( n3492 & ~n17286 ) | ( n3492 & 1'b0 ) | ( ~n17286 & 1'b0 ) ;
  assign n17288 = ( n455 & ~n865 ) | ( n455 & n17287 ) | ( ~n865 & n17287 ) ;
  assign n17289 = ( n17288 & ~n455 ) | ( n17288 & 1'b0 ) | ( ~n455 & 1'b0 ) ;
  assign n17290 = ( n712 & ~n218 ) | ( n712 & n17289 ) | ( ~n218 & n17289 ) ;
  assign n17291 = ~n712 & n17290 ;
  assign n17292 = ( n678 & ~n133 ) | ( n678 & n17291 ) | ( ~n133 & n17291 ) ;
  assign n17293 = ~n678 & n17292 ;
  assign n17294 = ( n228 & ~n574 ) | ( n228 & n17293 ) | ( ~n574 & n17293 ) ;
  assign n17295 = ~n228 & n17294 ;
  assign n17296 = ( n630 & ~n353 ) | ( n630 & n17295 ) | ( ~n353 & n17295 ) ;
  assign n17297 = ~n630 & n17296 ;
  assign n17305 = ~x8 & n17185 ;
  assign n17306 = ( n17208 & ~n17211 ) | ( n17208 & n17305 ) | ( ~n17211 & n17305 ) ;
  assign n17303 = n12100 | n3644 ;
  assign n17298 = n3653 | n11122 ;
  assign n17299 = n3657 &  n11125 ;
  assign n17300 = ( n3652 & ~n11128 ) | ( n3652 & 1'b0 ) | ( ~n11128 & 1'b0 ) ;
  assign n17301 = n17299 | n17300 ;
  assign n17302 = ( n17298 & ~n17301 ) | ( n17298 & 1'b0 ) | ( ~n17301 & 1'b0 ) ;
  assign n17304 = ( n3644 & ~n17303 ) | ( n3644 & n17302 ) | ( ~n17303 & n17302 ) ;
  assign n17307 = ( n17297 & ~n17306 ) | ( n17297 & n17304 ) | ( ~n17306 & n17304 ) ;
  assign n17308 = ( n17297 & ~n17304 ) | ( n17297 & n17306 ) | ( ~n17304 & n17306 ) ;
  assign n17309 = ( n17307 & ~n17297 ) | ( n17307 & n17308 ) | ( ~n17297 & n17308 ) ;
  assign n17310 = ~n17280 & n17309 ;
  assign n17311 = ( n17280 & ~n17309 ) | ( n17280 & 1'b0 ) | ( ~n17309 & 1'b0 ) ;
  assign n17312 = n17310 | n17311 ;
  assign n17318 = ~n601 & n12369 ;
  assign n17314 = ~n523 & n11119 ;
  assign n17315 = ~n3939 & n11116 ;
  assign n17316 = n17314 | n17315 ;
  assign n17313 = ( n4430 & ~n11113 ) | ( n4430 & 1'b0 ) | ( ~n11113 & 1'b0 ) ;
  assign n17317 = ( n11113 & ~n17316 ) | ( n11113 & n17313 ) | ( ~n17316 & n17313 ) ;
  assign n17319 = ( n601 & n17318 ) | ( n601 & n17317 ) | ( n17318 & n17317 ) ;
  assign n17320 = ( n17312 & ~x29 ) | ( n17312 & n17319 ) | ( ~x29 & n17319 ) ;
  assign n17321 = ( x29 & ~n17312 ) | ( x29 & n17319 ) | ( ~n17312 & n17319 ) ;
  assign n17322 = ( n17320 & ~n17319 ) | ( n17320 & n17321 ) | ( ~n17319 & n17321 ) ;
  assign n17323 = ( n17174 & ~n17216 ) | ( n17174 & n17217 ) | ( ~n17216 & n17217 ) ;
  assign n17327 = ~n4962 & n11104 ;
  assign n17324 = n4482 | n11110 ;
  assign n17325 = ~n4495 & n11107 ;
  assign n17326 = ( n17324 & ~n17325 ) | ( n17324 & 1'b0 ) | ( ~n17325 & 1'b0 ) ;
  assign n17328 = ( n4962 & n17327 ) | ( n4962 & n17326 ) | ( n17327 & n17326 ) ;
  assign n17329 = ~n4478 & n12662 ;
  assign n17330 = ( n17328 & ~n17329 ) | ( n17328 & 1'b0 ) | ( ~n17329 & 1'b0 ) ;
  assign n17331 = x26 &  n17330 ;
  assign n17332 = x26 | n17330 ;
  assign n17333 = ~n17331 & n17332 ;
  assign n17334 = ( n17322 & ~n17323 ) | ( n17322 & n17333 ) | ( ~n17323 & n17333 ) ;
  assign n17335 = ( n17322 & ~n17333 ) | ( n17322 & n17323 ) | ( ~n17333 & n17323 ) ;
  assign n17336 = ( n17334 & ~n17322 ) | ( n17334 & n17335 ) | ( ~n17322 & n17335 ) ;
  assign n17340 = ~n5135 & n11095 ;
  assign n17337 = n5010 | n11101 ;
  assign n17338 = n5067 | n11098 ;
  assign n17339 = n17337 &  n17338 ;
  assign n17341 = ( n5135 & n17340 ) | ( n5135 & n17339 ) | ( n17340 & n17339 ) ;
  assign n17342 = n5012 | n13014 ;
  assign n17343 = n17341 &  n17342 ;
  assign n17344 = x23 &  n17343 ;
  assign n17345 = x23 | n17343 ;
  assign n17346 = ~n17344 & n17345 ;
  assign n17347 = ( n17221 & n17336 ) | ( n17221 & n17346 ) | ( n17336 & n17346 ) ;
  assign n17348 = ( n17336 & ~n17221 ) | ( n17336 & n17346 ) | ( ~n17221 & n17346 ) ;
  assign n17349 = ( n17221 & ~n17347 ) | ( n17221 & n17348 ) | ( ~n17347 & n17348 ) ;
  assign n17353 = ~n5837 & n11081 ;
  assign n17350 = ( n5339 & ~n11093 ) | ( n5339 & 1'b0 ) | ( ~n11093 & 1'b0 ) ;
  assign n17351 = n5761 | n11091 ;
  assign n17352 = ~n17350 & n17351 ;
  assign n17354 = ( n5837 & n17353 ) | ( n5837 & n17352 ) | ( n17353 & n17352 ) ;
  assign n17355 = n5341 | n13775 ;
  assign n17356 = n17354 &  n17355 ;
  assign n17357 = x20 &  n17356 ;
  assign n17358 = x20 | n17356 ;
  assign n17359 = ~n17357 & n17358 ;
  assign n17360 = ( n17225 & n17349 ) | ( n17225 & n17359 ) | ( n17349 & n17359 ) ;
  assign n17361 = ( n17349 & ~n17225 ) | ( n17349 & n17359 ) | ( ~n17225 & n17359 ) ;
  assign n17362 = ( n17225 & ~n17360 ) | ( n17225 & n17361 ) | ( ~n17360 & n17361 ) ;
  assign n17366 = ~n6395 & n13836 ;
  assign n17363 = n5970 | n11085 ;
  assign n17364 = n6170 | n11078 ;
  assign n17365 = n17363 &  n17364 ;
  assign n17367 = ( n6395 & n17366 ) | ( n6395 & n17365 ) | ( n17366 & n17365 ) ;
  assign n17368 = n5972 | n13844 ;
  assign n17369 = n17367 &  n17368 ;
  assign n17370 = x17 &  n17369 ;
  assign n17371 = x17 | n17369 ;
  assign n17372 = ~n17370 & n17371 ;
  assign n17373 = ( n17228 & n17362 ) | ( n17228 & n17372 ) | ( n17362 & n17372 ) ;
  assign n17374 = ( n17362 & ~n17228 ) | ( n17362 & n17372 ) | ( ~n17228 & n17372 ) ;
  assign n17375 = ( n17228 & ~n17373 ) | ( n17228 & n17374 ) | ( ~n17373 & n17374 ) ;
  assign n17379 = n14553 | n7097 ;
  assign n17376 = n6530 | n14071 ;
  assign n17377 = n6983 | n14355 ;
  assign n17378 = n17376 &  n17377 ;
  assign n17380 = ( n7097 & ~n17379 ) | ( n7097 & n17378 ) | ( ~n17379 & n17378 ) ;
  assign n17381 = ~n6532 & n14562 ;
  assign n17382 = ( n17380 & ~n17381 ) | ( n17380 & 1'b0 ) | ( ~n17381 & 1'b0 ) ;
  assign n17383 = x14 &  n17382 ;
  assign n17384 = x14 | n17382 ;
  assign n17385 = ~n17383 & n17384 ;
  assign n17386 = ( n17279 & n17375 ) | ( n17279 & n17385 ) | ( n17375 & n17385 ) ;
  assign n17387 = ( n17375 & ~n17279 ) | ( n17375 & n17385 ) | ( ~n17279 & n17385 ) ;
  assign n17388 = ( n17279 & ~n17386 ) | ( n17279 & n17387 ) | ( ~n17386 & n17387 ) ;
  assign n17392 = n14800 | n7783 ;
  assign n17389 = ( n7253 & ~n14803 ) | ( n7253 & 1'b0 ) | ( ~n14803 & 1'b0 ) ;
  assign n17390 = ~n7518 & n14807 ;
  assign n17391 = n17389 | n17390 ;
  assign n17393 = ( n17392 & ~n7783 ) | ( n17392 & n17391 ) | ( ~n7783 & n17391 ) ;
  assign n17394 = n7255 | n14816 ;
  assign n17395 = ~n17393 & n17394 ;
  assign n17396 = x11 &  n17395 ;
  assign n17397 = x11 | n17395 ;
  assign n17398 = ~n17396 & n17397 ;
  assign n17399 = ( n17278 & n17388 ) | ( n17278 & n17398 ) | ( n17388 & n17398 ) ;
  assign n17400 = ( n17388 & ~n17278 ) | ( n17388 & n17398 ) | ( ~n17278 & n17398 ) ;
  assign n17401 = ( n17278 & ~n17399 ) | ( n17278 & n17400 ) | ( ~n17399 & n17400 ) ;
  assign n17403 = ( n17259 & ~n17402 ) | ( n17259 & n17401 ) | ( ~n17402 & n17401 ) ;
  assign n17404 = ( n17259 & ~n17401 ) | ( n17259 & n17402 ) | ( ~n17401 & n17402 ) ;
  assign n17405 = ( ~n17259 & n17403 ) | ( ~n17259 & n17404 ) | ( n17403 & n17404 ) ;
  assign n17412 = ( n17263 & n17270 ) | ( n17263 & n17405 ) | ( n17270 & n17405 ) ;
  assign n17411 = ( n17270 & ~n17263 ) | ( n17270 & n17405 ) | ( ~n17263 & n17405 ) ;
  assign n17413 = ( n17263 & ~n17412 ) | ( n17263 & n17411 ) | ( ~n17412 & n17411 ) ;
  assign n17409 = ~n5837 & n17405 ;
  assign n17406 = n5339 &  n17107 ;
  assign n17407 = n5761 | n17263 ;
  assign n17408 = ~n17406 & n17407 ;
  assign n17410 = ( n5837 & n17409 ) | ( n5837 & n17408 ) | ( n17409 & n17408 ) ;
  assign n17414 = ( n17410 & ~n5341 ) | ( n17410 & n17413 ) | ( ~n5341 & n17413 ) ;
  assign n17415 = ~n17413 & n17414 ;
  assign n17417 = ( x20 & n17410 ) | ( x20 & n17415 ) | ( n17410 & n17415 ) ;
  assign n17416 = ( x20 & ~n17415 ) | ( x20 & n17410 ) | ( ~n17415 & n17410 ) ;
  assign n17418 = ( n17415 & ~n17417 ) | ( n17415 & n17416 ) | ( ~n17417 & n17416 ) ;
  assign n17419 = ( n16785 & ~n17277 ) | ( n16785 & n17418 ) | ( ~n17277 & n17418 ) ;
  assign n17420 = ( n16785 & ~n17418 ) | ( n16785 & n17277 ) | ( ~n17418 & n17277 ) ;
  assign n17421 = ( n17419 & ~n16785 ) | ( n17419 & n17420 ) | ( ~n16785 & n17420 ) ;
  assign n17422 = ( n17225 & ~n17349 ) | ( n17225 & n17359 ) | ( ~n17349 & n17359 ) ;
  assign n17423 = ( n17221 & ~n17336 ) | ( n17221 & n17346 ) | ( ~n17336 & n17346 ) ;
  assign n17424 = ( n17323 & ~n17322 ) | ( n17323 & n17333 ) | ( ~n17322 & n17333 ) ;
  assign n17425 = n1123 | n2550 ;
  assign n17426 = ( n738 & ~n1169 ) | ( n738 & n17425 ) | ( ~n1169 & n17425 ) ;
  assign n17427 = n1169 | n17426 ;
  assign n17428 = ( n4788 & ~n11281 ) | ( n4788 & n17427 ) | ( ~n11281 & n17427 ) ;
  assign n17429 = ( n4788 & ~n17428 ) | ( n4788 & 1'b0 ) | ( ~n17428 & 1'b0 ) ;
  assign n17430 = ( n1679 & ~n14137 ) | ( n1679 & n17429 ) | ( ~n14137 & n17429 ) ;
  assign n17431 = ~n1679 & n17430 ;
  assign n17432 = ( n842 & ~n717 ) | ( n842 & n17431 ) | ( ~n717 & n17431 ) ;
  assign n17433 = ~n842 & n17432 ;
  assign n17434 = ( n126 & ~n673 ) | ( n126 & n17433 ) | ( ~n673 & n17433 ) ;
  assign n17435 = ~n126 & n17434 ;
  assign n17436 = ( n231 & ~n242 ) | ( n231 & n17435 ) | ( ~n242 & n17435 ) ;
  assign n17437 = ~n231 & n17436 ;
  assign n17438 = ( n627 & ~n451 ) | ( n627 & n17437 ) | ( ~n451 & n17437 ) ;
  assign n17439 = ~n627 & n17438 ;
  assign n17440 = ~n140 & n17439 ;
  assign n17441 = ( n17304 & ~n17297 ) | ( n17304 & n17306 ) | ( ~n17297 & n17306 ) ;
  assign n17442 = ( n17440 & ~n17297 ) | ( n17440 & n17441 ) | ( ~n17297 & n17441 ) ;
  assign n17443 = ( n17297 & ~n17440 ) | ( n17297 & n17441 ) | ( ~n17440 & n17441 ) ;
  assign n17444 = ( n17442 & ~n17441 ) | ( n17442 & n17443 ) | ( ~n17441 & n17443 ) ;
  assign n17445 = ~n3644 & n12088 ;
  assign n17446 = n3652 &  n11125 ;
  assign n17447 = ( n3657 & ~n11122 ) | ( n3657 & 1'b0 ) | ( ~n11122 & 1'b0 ) ;
  assign n17448 = n17446 | n17447 ;
  assign n17449 = n3653 | n11119 ;
  assign n17450 = ( n17448 & ~n3653 ) | ( n17448 & n17449 ) | ( ~n3653 & n17449 ) ;
  assign n17451 = n17445 | n17450 ;
  assign n17455 = ~n4430 & n11110 ;
  assign n17452 = ~n523 & n11116 ;
  assign n17453 = n3939 | n11113 ;
  assign n17454 = ~n17452 & n17453 ;
  assign n17456 = ( n4430 & n17455 ) | ( n4430 & n17454 ) | ( n17455 & n17454 ) ;
  assign n17457 = ( n601 & ~n17456 ) | ( n601 & n12352 ) | ( ~n17456 & n12352 ) ;
  assign n17458 = ( n12352 & ~n17457 ) | ( n12352 & 1'b0 ) | ( ~n17457 & 1'b0 ) ;
  assign n17460 = ( x29 & n17456 ) | ( x29 & n17458 ) | ( n17456 & n17458 ) ;
  assign n17459 = ( x29 & ~n17458 ) | ( x29 & n17456 ) | ( ~n17458 & n17456 ) ;
  assign n17461 = ( n17458 & ~n17460 ) | ( n17458 & n17459 ) | ( ~n17460 & n17459 ) ;
  assign n17462 = ( n17444 & ~n17451 ) | ( n17444 & n17461 ) | ( ~n17451 & n17461 ) ;
  assign n17463 = ( n17451 & ~n17444 ) | ( n17451 & n17461 ) | ( ~n17444 & n17461 ) ;
  assign n17464 = ( n17462 & ~n17461 ) | ( n17462 & n17463 ) | ( ~n17461 & n17463 ) ;
  assign n17471 = ~n4962 & n11101 ;
  assign n17468 = ~n4482 & n11107 ;
  assign n17469 = n4495 | n11104 ;
  assign n17470 = ~n17468 & n17469 ;
  assign n17472 = ( n4962 & n17471 ) | ( n4962 & n17470 ) | ( n17471 & n17470 ) ;
  assign n17473 = n4478 | n12650 ;
  assign n17474 = n17472 &  n17473 ;
  assign n17475 = x26 &  n17474 ;
  assign n17476 = x26 | n17474 ;
  assign n17477 = ~n17475 & n17476 ;
  assign n17465 = ~x29 & n17319 ;
  assign n17466 = ( x29 & ~n17319 ) | ( x29 & n17311 ) | ( ~n17319 & n17311 ) ;
  assign n17467 = ( n17465 & ~n17310 ) | ( n17465 & n17466 ) | ( ~n17310 & n17466 ) ;
  assign n17478 = ( n17464 & ~n17477 ) | ( n17464 & n17467 ) | ( ~n17477 & n17467 ) ;
  assign n17479 = ( n17464 & ~n17467 ) | ( n17464 & n17477 ) | ( ~n17467 & n17477 ) ;
  assign n17480 = ( n17478 & ~n17464 ) | ( n17478 & n17479 ) | ( ~n17464 & n17479 ) ;
  assign n17484 = ~n5135 & n11093 ;
  assign n17481 = n5010 | n11098 ;
  assign n17482 = n5067 | n11095 ;
  assign n17483 = n17481 &  n17482 ;
  assign n17485 = ( n5135 & n17484 ) | ( n5135 & n17483 ) | ( n17484 & n17483 ) ;
  assign n17486 = n5012 | n12997 ;
  assign n17487 = n17485 &  n17486 ;
  assign n17488 = x23 &  n17487 ;
  assign n17489 = x23 | n17487 ;
  assign n17490 = ~n17488 & n17489 ;
  assign n17491 = ( n17424 & ~n17480 ) | ( n17424 & n17490 ) | ( ~n17480 & n17490 ) ;
  assign n17492 = ( n17424 & ~n17490 ) | ( n17424 & n17480 ) | ( ~n17490 & n17480 ) ;
  assign n17493 = ( n17491 & ~n17424 ) | ( n17491 & n17492 ) | ( ~n17424 & n17492 ) ;
  assign n17497 = ~n5837 & n11085 ;
  assign n17494 = ( n5339 & ~n11091 ) | ( n5339 & 1'b0 ) | ( ~n11091 & 1'b0 ) ;
  assign n17495 = n5761 | n11081 ;
  assign n17496 = ~n17494 & n17495 ;
  assign n17498 = ( n5837 & n17497 ) | ( n5837 & n17496 ) | ( n17497 & n17496 ) ;
  assign n17499 = n5341 | n13377 ;
  assign n17500 = n17498 &  n17499 ;
  assign n17501 = x20 &  n17500 ;
  assign n17502 = x20 | n17500 ;
  assign n17503 = ~n17501 & n17502 ;
  assign n17504 = ( n17423 & ~n17493 ) | ( n17423 & n17503 ) | ( ~n17493 & n17503 ) ;
  assign n17505 = ( n17423 & ~n17503 ) | ( n17423 & n17493 ) | ( ~n17503 & n17493 ) ;
  assign n17506 = ( n17504 & ~n17423 ) | ( n17504 & n17505 ) | ( ~n17423 & n17505 ) ;
  assign n17510 = ~n6395 & n14071 ;
  assign n17507 = n5970 | n11078 ;
  assign n17508 = n6170 | n13836 ;
  assign n17509 = n17507 &  n17508 ;
  assign n17511 = ( n6395 & n17510 ) | ( n6395 & n17509 ) | ( n17510 & n17509 ) ;
  assign n17512 = n5972 | n14079 ;
  assign n17513 = n17511 &  n17512 ;
  assign n17514 = x17 &  n17513 ;
  assign n17515 = x17 | n17513 ;
  assign n17516 = ~n17514 & n17515 ;
  assign n17517 = ( n17422 & ~n17506 ) | ( n17422 & n17516 ) | ( ~n17506 & n17516 ) ;
  assign n17518 = ( n17422 & ~n17516 ) | ( n17422 & n17506 ) | ( ~n17516 & n17506 ) ;
  assign n17519 = ( n17517 & ~n17422 ) | ( n17517 & n17518 ) | ( ~n17422 & n17518 ) ;
  assign n17520 = ( n17228 & ~n17362 ) | ( n17228 & n17372 ) | ( ~n17362 & n17372 ) ;
  assign n17524 = ~n7097 & n14803 ;
  assign n17521 = n6530 | n14355 ;
  assign n17522 = ~n6983 & n14553 ;
  assign n17523 = ( n17521 & ~n17522 ) | ( n17521 & 1'b0 ) | ( ~n17522 & 1'b0 ) ;
  assign n17525 = ( n7097 & n17524 ) | ( n7097 & n17523 ) | ( n17524 & n17523 ) ;
  assign n17526 = ~n6532 & n15310 ;
  assign n17527 = ( n17525 & ~n17526 ) | ( n17525 & 1'b0 ) | ( ~n17526 & 1'b0 ) ;
  assign n17528 = x14 &  n17527 ;
  assign n17529 = x14 | n17527 ;
  assign n17530 = ~n17528 & n17529 ;
  assign n17531 = ( n17519 & n17520 ) | ( n17519 & n17530 ) | ( n17520 & n17530 ) ;
  assign n17545 = ~n6395 & n14355 ;
  assign n17542 = n5970 | n13836 ;
  assign n17543 = n6170 | n14071 ;
  assign n17544 = n17542 &  n17543 ;
  assign n17546 = ( n6395 & n17545 ) | ( n6395 & n17544 ) | ( n17545 & n17544 ) ;
  assign n17547 = n5972 | n14363 ;
  assign n17548 = n17546 &  n17547 ;
  assign n17549 = x17 &  n17548 ;
  assign n17550 = x17 | n17548 ;
  assign n17551 = ~n17549 & n17550 ;
  assign n17555 = ~n5837 & n11078 ;
  assign n17552 = ( n5339 & ~n11081 ) | ( n5339 & 1'b0 ) | ( ~n11081 & 1'b0 ) ;
  assign n17553 = n5761 | n11085 ;
  assign n17554 = ~n17552 & n17553 ;
  assign n17556 = ( n5837 & n17555 ) | ( n5837 & n17554 ) | ( n17555 & n17554 ) ;
  assign n17557 = n5341 | n11206 ;
  assign n17558 = n17556 &  n17557 ;
  assign n17559 = x20 &  n17558 ;
  assign n17560 = x20 | n17558 ;
  assign n17561 = ~n17559 & n17560 ;
  assign n17565 = ~n5135 & n11091 ;
  assign n17562 = n5010 | n11095 ;
  assign n17563 = n5067 | n11093 ;
  assign n17564 = n17562 &  n17563 ;
  assign n17566 = ( n5135 & n17565 ) | ( n5135 & n17564 ) | ( n17565 & n17564 ) ;
  assign n17567 = n5012 | n12984 ;
  assign n17568 = n17566 &  n17567 ;
  assign n17569 = x23 &  n17568 ;
  assign n17570 = x23 | n17568 ;
  assign n17571 = ~n17569 & n17570 ;
  assign n17575 = ~n4962 & n11098 ;
  assign n17572 = n4482 | n11104 ;
  assign n17573 = n4495 | n11101 ;
  assign n17574 = n17572 &  n17573 ;
  assign n17576 = ( n4962 & n17575 ) | ( n4962 & n17574 ) | ( n17575 & n17574 ) ;
  assign n17577 = n4478 | n11218 ;
  assign n17578 = n17576 &  n17577 ;
  assign n17579 = x26 &  n17578 ;
  assign n17580 = x26 | n17578 ;
  assign n17581 = ~n17579 & n17580 ;
  assign n17589 = ( n7248 & ~n7245 ) | ( n7248 & n7251 ) | ( ~n7245 & n7251 ) ;
  assign n17590 = n7245 | n17589 ;
  assign n17591 = n14800 &  n17590 ;
  assign n17596 = n963 | n3173 ;
  assign n17597 = ( n3326 & ~n2044 ) | ( n3326 & n17596 ) | ( ~n2044 & n17596 ) ;
  assign n17598 = n2044 | n17597 ;
  assign n17599 = ( n2074 & n6057 ) | ( n2074 & n17598 ) | ( n6057 & n17598 ) ;
  assign n17600 = ( n2074 & ~n17599 ) | ( n2074 & 1'b0 ) | ( ~n17599 & 1'b0 ) ;
  assign n17601 = ( n1122 & n1510 ) | ( n1122 & n17600 ) | ( n1510 & n17600 ) ;
  assign n17602 = ~n1510 & n17601 ;
  assign n17592 = ~n2092 & n3043 ;
  assign n17593 = ( n148 & ~n274 ) | ( n148 & n17592 ) | ( ~n274 & n17592 ) ;
  assign n17594 = ~n148 & n17593 ;
  assign n17595 = ~n95 & n17594 ;
  assign n17603 = ( n1282 & ~n17602 ) | ( n1282 & n17595 ) | ( ~n17602 & n17595 ) ;
  assign n17604 = ( n81 & ~n17603 ) | ( n81 & n17595 ) | ( ~n17603 & n17595 ) ;
  assign n17605 = ~n81 & n17604 ;
  assign n17606 = ( n224 & ~n134 ) | ( n224 & n17605 ) | ( ~n134 & n17605 ) ;
  assign n17607 = ~n224 & n17606 ;
  assign n17608 = ( n165 & ~n222 ) | ( n165 & n17607 ) | ( ~n222 & n17607 ) ;
  assign n17609 = ~n165 & n17608 ;
  assign n17610 = ~n558 & n17609 ;
  assign n17611 = n17297 | n17610 ;
  assign n17612 = n17297 &  n17610 ;
  assign n17613 = ( n17611 & ~n17612 ) | ( n17611 & 1'b0 ) | ( ~n17612 & 1'b0 ) ;
  assign n17614 = ( n17591 & ~x11 ) | ( n17591 & n17613 ) | ( ~x11 & n17613 ) ;
  assign n17615 = ( x11 & ~n17613 ) | ( x11 & n17591 ) | ( ~n17613 & n17591 ) ;
  assign n17616 = ( n17614 & ~n17591 ) | ( n17614 & n17615 ) | ( ~n17591 & n17615 ) ;
  assign n17582 = n3644 | n11230 ;
  assign n17586 = n11116 | n3653 ;
  assign n17583 = ( n3652 & ~n11122 ) | ( n3652 & 1'b0 ) | ( ~n11122 & 1'b0 ) ;
  assign n17584 = n3657 &  n11119 ;
  assign n17585 = n17583 | n17584 ;
  assign n17587 = ( n17586 & ~n3653 ) | ( n17586 & n17585 ) | ( ~n3653 & n17585 ) ;
  assign n17588 = ( n17582 & ~n17587 ) | ( n17582 & 1'b0 ) | ( ~n17587 & 1'b0 ) ;
  assign n17617 = ( n17442 & n17588 ) | ( n17442 & n17616 ) | ( n17588 & n17616 ) ;
  assign n17618 = ( n17442 & ~n17616 ) | ( n17442 & n17588 ) | ( ~n17616 & n17588 ) ;
  assign n17619 = ( n17616 & ~n17617 ) | ( n17616 & n17618 ) | ( ~n17617 & n17618 ) ;
  assign n17620 = ( n17444 & ~n17461 ) | ( n17444 & n17451 ) | ( ~n17461 & n17451 ) ;
  assign n17624 = n11107 | n4430 ;
  assign n17621 = n523 | n11113 ;
  assign n17622 = n3939 | n11110 ;
  assign n17623 = n17621 &  n17622 ;
  assign n17625 = ( n4430 & ~n17624 ) | ( n4430 & n17623 ) | ( ~n17624 & n17623 ) ;
  assign n17626 = ~n601 & n12340 ;
  assign n17627 = ( n17625 & ~n17626 ) | ( n17625 & 1'b0 ) | ( ~n17626 & 1'b0 ) ;
  assign n17628 = x29 &  n17627 ;
  assign n17629 = x29 | n17627 ;
  assign n17630 = ~n17628 & n17629 ;
  assign n17631 = ( n17619 & n17620 ) | ( n17619 & n17630 ) | ( n17620 & n17630 ) ;
  assign n17632 = ( n17620 & ~n17619 ) | ( n17620 & n17630 ) | ( ~n17619 & n17630 ) ;
  assign n17633 = ( n17619 & ~n17631 ) | ( n17619 & n17632 ) | ( ~n17631 & n17632 ) ;
  assign n17634 = ( n17464 & n17467 ) | ( n17464 & n17477 ) | ( n17467 & n17477 ) ;
  assign n17635 = ( n17581 & n17633 ) | ( n17581 & n17634 ) | ( n17633 & n17634 ) ;
  assign n17636 = ( n17633 & ~n17581 ) | ( n17633 & n17634 ) | ( ~n17581 & n17634 ) ;
  assign n17637 = ( n17581 & ~n17635 ) | ( n17581 & n17636 ) | ( ~n17635 & n17636 ) ;
  assign n17638 = ( n17424 & n17480 ) | ( n17424 & n17490 ) | ( n17480 & n17490 ) ;
  assign n17639 = ( n17571 & ~n17637 ) | ( n17571 & n17638 ) | ( ~n17637 & n17638 ) ;
  assign n17640 = ( n17571 & ~n17638 ) | ( n17571 & n17637 ) | ( ~n17638 & n17637 ) ;
  assign n17641 = ( n17639 & ~n17571 ) | ( n17639 & n17640 ) | ( ~n17571 & n17640 ) ;
  assign n17642 = ( n17423 & n17493 ) | ( n17423 & n17503 ) | ( n17493 & n17503 ) ;
  assign n17643 = ( n17561 & ~n17641 ) | ( n17561 & n17642 ) | ( ~n17641 & n17642 ) ;
  assign n17644 = ( n17561 & ~n17642 ) | ( n17561 & n17641 ) | ( ~n17642 & n17641 ) ;
  assign n17645 = ( n17643 & ~n17561 ) | ( n17643 & n17644 ) | ( ~n17561 & n17644 ) ;
  assign n17646 = ( n17422 & n17506 ) | ( n17422 & n17516 ) | ( n17506 & n17516 ) ;
  assign n17647 = ( n17551 & ~n17645 ) | ( n17551 & n17646 ) | ( ~n17645 & n17646 ) ;
  assign n17648 = ( n17551 & ~n17646 ) | ( n17551 & n17645 ) | ( ~n17646 & n17645 ) ;
  assign n17649 = ( n17647 & ~n17551 ) | ( n17647 & n17648 ) | ( ~n17551 & n17648 ) ;
  assign n17535 = n14807 | n7097 ;
  assign n17532 = ~n6530 & n14553 ;
  assign n17533 = n6983 | n14803 ;
  assign n17534 = ~n17532 & n17533 ;
  assign n17536 = ( n7097 & ~n17535 ) | ( n7097 & n17534 ) | ( ~n17535 & n17534 ) ;
  assign n17537 = ~n6532 & n15294 ;
  assign n17538 = ( n17536 & ~n17537 ) | ( n17536 & 1'b0 ) | ( ~n17537 & 1'b0 ) ;
  assign n17539 = x14 &  n17538 ;
  assign n17540 = x14 | n17538 ;
  assign n17541 = ~n17539 & n17540 ;
  assign n17650 = ( n17531 & ~n17649 ) | ( n17531 & n17541 ) | ( ~n17649 & n17541 ) ;
  assign n17772 = ( n17541 & ~n17531 ) | ( n17541 & n17649 ) | ( ~n17531 & n17649 ) ;
  assign n17773 = ( n17650 & ~n17541 ) | ( n17650 & n17772 ) | ( ~n17541 & n17772 ) ;
  assign n17758 = ( n17279 & ~n17375 ) | ( n17279 & n17385 ) | ( ~n17375 & n17385 ) ;
  assign n17759 = n7518 &  n7783 ;
  assign n17760 = ( n14800 & ~n17759 ) | ( n14800 & 1'b0 ) | ( ~n17759 & 1'b0 ) ;
  assign n17761 = n7253 &  n14807 ;
  assign n17762 = n17760 | n17761 ;
  assign n17763 = ( n7255 & n15692 ) | ( n7255 & n17762 ) | ( n15692 & n17762 ) ;
  assign n17764 = ( n15692 & ~n17763 ) | ( n15692 & 1'b0 ) | ( ~n17763 & 1'b0 ) ;
  assign n17765 = ( n17762 & ~x11 ) | ( n17762 & n17764 ) | ( ~x11 & n17764 ) ;
  assign n17766 = ( x11 & ~n17762 ) | ( x11 & n17764 ) | ( ~n17762 & n17764 ) ;
  assign n17767 = ( n17765 & ~n17764 ) | ( n17765 & n17766 ) | ( ~n17764 & n17766 ) ;
  assign n17768 = ( n17520 & ~n17519 ) | ( n17520 & n17530 ) | ( ~n17519 & n17530 ) ;
  assign n17769 = ( n17519 & ~n17530 ) | ( n17519 & n17520 ) | ( ~n17530 & n17520 ) ;
  assign n17770 = ( n17768 & ~n17520 ) | ( n17768 & n17769 ) | ( ~n17520 & n17769 ) ;
  assign n17771 = ( n17758 & ~n17767 ) | ( n17758 & n17770 ) | ( ~n17767 & n17770 ) ;
  assign n17774 = ( n17758 & ~n17770 ) | ( n17758 & n17767 ) | ( ~n17770 & n17767 ) ;
  assign n17775 = ( n17767 & ~n17758 ) | ( n17767 & n17770 ) | ( ~n17758 & n17770 ) ;
  assign n17776 = ( n17774 & ~n17767 ) | ( n17774 & n17775 ) | ( ~n17767 & n17775 ) ;
  assign n17777 = ( n17278 & ~n17388 ) | ( n17278 & n17398 ) | ( ~n17388 & n17398 ) ;
  assign n17778 = ( n17401 & ~n17259 ) | ( n17401 & n17402 ) | ( ~n17259 & n17402 ) ;
  assign n17779 = ( n17776 & ~n17777 ) | ( n17776 & n17778 ) | ( ~n17777 & n17778 ) ;
  assign n17789 = ( n17771 & ~n17773 ) | ( n17771 & n17779 ) | ( ~n17773 & n17779 ) ;
  assign n17790 = ( n17771 & n17773 ) | ( n17771 & n17779 ) | ( n17773 & n17779 ) ;
  assign n17791 = ( n17773 & n17789 ) | ( n17773 & ~n17790 ) | ( n17789 & ~n17790 ) ;
  assign n17808 = ~n6395 & n17791 ;
  assign n17805 = n5970 | n17405 ;
  assign n17785 = ( n17776 & ~n17778 ) | ( n17776 & n17777 ) | ( ~n17778 & n17777 ) ;
  assign n17786 = ( n17777 & ~n17776 ) | ( n17777 & n17778 ) | ( ~n17776 & n17778 ) ;
  assign n17787 = ( n17785 & ~n17777 ) | ( n17785 & n17786 ) | ( ~n17777 & n17786 ) ;
  assign n17806 = n6170 | n17787 ;
  assign n17807 = n17805 &  n17806 ;
  assign n17809 = ( n6395 & n17808 ) | ( n6395 & n17807 ) | ( n17808 & n17807 ) ;
  assign n17795 = ( n17405 & n17412 ) | ( n17405 & n17787 ) | ( n17412 & n17787 ) ;
  assign n17796 = ( n17787 & n17791 ) | ( n17787 & n17795 ) | ( n17791 & n17795 ) ;
  assign n17810 = ( n17791 & ~n17787 ) | ( n17791 & n17795 ) | ( ~n17787 & n17795 ) ;
  assign n17811 = ( n17787 & ~n17796 ) | ( n17787 & n17810 ) | ( ~n17796 & n17810 ) ;
  assign n17812 = n5972 | n17811 ;
  assign n17813 = n17809 &  n17812 ;
  assign n17814 = x17 &  n17813 ;
  assign n17815 = x17 | n17813 ;
  assign n17816 = ~n17814 & n17815 ;
  assign n17817 = ( n17121 & ~n17276 ) | ( n17121 & n17124 ) | ( ~n17276 & n17124 ) ;
  assign n17818 = ( n17124 & ~n17121 ) | ( n17124 & n17276 ) | ( ~n17121 & n17276 ) ;
  assign n17819 = ( n17817 & ~n17124 ) | ( n17817 & n17818 ) | ( ~n17124 & n17818 ) ;
  assign n17823 = ~n6395 & n17787 ;
  assign n17820 = n5970 | n17263 ;
  assign n17821 = n6170 | n17405 ;
  assign n17822 = n17820 &  n17821 ;
  assign n17824 = ( n6395 & n17823 ) | ( n6395 & n17822 ) | ( n17823 & n17822 ) ;
  assign n17825 = ( n17412 & ~n17405 ) | ( n17412 & n17787 ) | ( ~n17405 & n17787 ) ;
  assign n17826 = ( n17405 & ~n17795 ) | ( n17405 & n17825 ) | ( ~n17795 & n17825 ) ;
  assign n17827 = n5972 | n17826 ;
  assign n17828 = n17824 &  n17827 ;
  assign n17829 = x17 &  n17828 ;
  assign n17830 = x17 | n17828 ;
  assign n17831 = ~n17829 & n17830 ;
  assign n17832 = ( n16966 & ~n17120 ) | ( n16966 & n16969 ) | ( ~n17120 & n16969 ) ;
  assign n17833 = ( n16969 & ~n16966 ) | ( n16969 & n17120 ) | ( ~n16966 & n17120 ) ;
  assign n17834 = ( n17832 & ~n16969 ) | ( n17832 & n17833 ) | ( ~n16969 & n17833 ) ;
  assign n17838 = ~n6395 & n17405 ;
  assign n17835 = ~n5970 & n17107 ;
  assign n17836 = n6170 | n17263 ;
  assign n17837 = ~n17835 & n17836 ;
  assign n17839 = ( n6395 & n17838 ) | ( n6395 & n17837 ) | ( n17838 & n17837 ) ;
  assign n17840 = ( n5972 & ~n17413 ) | ( n5972 & n17839 ) | ( ~n17413 & n17839 ) ;
  assign n17841 = ~n5972 & n17840 ;
  assign n17843 = ( x17 & n17839 ) | ( x17 & n17841 ) | ( n17839 & n17841 ) ;
  assign n17842 = ( x17 & ~n17841 ) | ( x17 & n17839 ) | ( ~n17841 & n17839 ) ;
  assign n17844 = ( n17841 & ~n17843 ) | ( n17841 & n17842 ) | ( ~n17843 & n17842 ) ;
  assign n17845 = ( n16955 & ~n16952 ) | ( n16955 & n16965 ) | ( ~n16952 & n16965 ) ;
  assign n17846 = ( n16952 & ~n16965 ) | ( n16952 & n16955 ) | ( ~n16965 & n16955 ) ;
  assign n17847 = ( n17845 & ~n16955 ) | ( n17845 & n17846 ) | ( ~n16955 & n17846 ) ;
  assign n17851 = ~n6395 & n17263 ;
  assign n17848 = n5970 | n16589 ;
  assign n17849 = ~n6170 & n17107 ;
  assign n17850 = ( n17848 & ~n17849 ) | ( n17848 & 1'b0 ) | ( ~n17849 & 1'b0 ) ;
  assign n17852 = ( n6395 & n17851 ) | ( n6395 & n17850 ) | ( n17851 & n17850 ) ;
  assign n17853 = ( n5972 & n17271 ) | ( n5972 & n17852 ) | ( n17271 & n17852 ) ;
  assign n17854 = ~n5972 & n17853 ;
  assign n17856 = ( x17 & n17852 ) | ( x17 & n17854 ) | ( n17852 & n17854 ) ;
  assign n17855 = ( x17 & ~n17854 ) | ( x17 & n17852 ) | ( ~n17854 & n17852 ) ;
  assign n17857 = ( n17854 & ~n17856 ) | ( n17854 & n17855 ) | ( ~n17856 & n17855 ) ;
  assign n17858 = ( n16788 & ~n16798 ) | ( n16788 & n16951 ) | ( ~n16798 & n16951 ) ;
  assign n17859 = ( n16798 & ~n16952 ) | ( n16798 & n17858 ) | ( ~n16952 & n17858 ) ;
  assign n17860 = ( n16808 & ~n16950 ) | ( n16808 & n16810 ) | ( ~n16950 & n16810 ) ;
  assign n17861 = ( n16810 & ~n16808 ) | ( n16810 & n16950 ) | ( ~n16808 & n16950 ) ;
  assign n17862 = ( n17860 & ~n16810 ) | ( n17860 & n17861 ) | ( ~n16810 & n17861 ) ;
  assign n17866 = n17107 | n6395 ;
  assign n17863 = n5970 | n16595 ;
  assign n17864 = n6170 | n16589 ;
  assign n17865 = n17863 &  n17864 ;
  assign n17867 = ( n6395 & ~n17866 ) | ( n6395 & n17865 ) | ( ~n17866 & n17865 ) ;
  assign n17868 = ( n5972 & n17115 ) | ( n5972 & n17867 ) | ( n17115 & n17867 ) ;
  assign n17869 = ~n5972 & n17868 ;
  assign n17870 = ( x17 & ~n17867 ) | ( x17 & n17869 ) | ( ~n17867 & n17869 ) ;
  assign n17871 = ( n17867 & ~x17 ) | ( n17867 & n17869 ) | ( ~x17 & n17869 ) ;
  assign n17872 = ( n17870 & ~n17869 ) | ( n17870 & n17871 ) | ( ~n17869 & n17871 ) ;
  assign n17873 = ( n16822 & ~n16820 ) | ( n16822 & n16949 ) | ( ~n16820 & n16949 ) ;
  assign n17874 = ( n16820 & ~n16949 ) | ( n16820 & n16822 ) | ( ~n16949 & n16822 ) ;
  assign n17875 = ( n17873 & ~n16822 ) | ( n17873 & n17874 ) | ( ~n16822 & n17874 ) ;
  assign n17879 = ~n6395 & n16589 ;
  assign n17876 = n5970 | n16591 ;
  assign n17877 = n6170 | n16595 ;
  assign n17878 = n17876 &  n17877 ;
  assign n17880 = ( n6395 & n17879 ) | ( n6395 & n17878 ) | ( n17879 & n17878 ) ;
  assign n17881 = ( n16604 & ~n5972 ) | ( n16604 & n17880 ) | ( ~n5972 & n17880 ) ;
  assign n17882 = ~n16604 & n17881 ;
  assign n17884 = ( x17 & n17880 ) | ( x17 & n17882 ) | ( n17880 & n17882 ) ;
  assign n17883 = ( x17 & ~n17882 ) | ( x17 & n17880 ) | ( ~n17882 & n17880 ) ;
  assign n17885 = ( n17882 & ~n17884 ) | ( n17882 & n17883 ) | ( ~n17884 & n17883 ) ;
  assign n17889 = ~n6395 & n16595 ;
  assign n17886 = n5970 | n16091 ;
  assign n17887 = n6170 | n16591 ;
  assign n17888 = n17886 &  n17887 ;
  assign n17890 = ( n6395 & n17889 ) | ( n6395 & n17888 ) | ( n17889 & n17888 ) ;
  assign n17891 = n5972 | n16616 ;
  assign n17892 = n17890 &  n17891 ;
  assign n17893 = x17 &  n17892 ;
  assign n17894 = x17 | n17892 ;
  assign n17895 = ~n17893 & n17894 ;
  assign n17896 = ( n16825 & ~n16948 ) | ( n16825 & n16835 ) | ( ~n16948 & n16835 ) ;
  assign n17897 = ( n16949 & ~n16835 ) | ( n16949 & n17896 ) | ( ~n16835 & n17896 ) ;
  assign n17901 = ~n6395 & n16591 ;
  assign n17898 = n5970 | n15897 ;
  assign n17899 = n6170 | n16091 ;
  assign n17900 = n17898 &  n17899 ;
  assign n17902 = ( n6395 & n17901 ) | ( n6395 & n17900 ) | ( n17901 & n17900 ) ;
  assign n17903 = n5972 | n16631 ;
  assign n17904 = n17902 &  n17903 ;
  assign n17905 = x17 &  n17904 ;
  assign n17906 = x17 | n17904 ;
  assign n17907 = ~n17905 & n17906 ;
  assign n17908 = ( n16838 & ~n16848 ) | ( n16838 & n16947 ) | ( ~n16848 & n16947 ) ;
  assign n17909 = ( n16848 & ~n16948 ) | ( n16848 & n17908 ) | ( ~n16948 & n17908 ) ;
  assign n17913 = ~n6395 & n16091 ;
  assign n17910 = n5970 | n15700 ;
  assign n17911 = n6170 | n15897 ;
  assign n17912 = n17910 &  n17911 ;
  assign n17914 = ( n6395 & n17913 ) | ( n6395 & n17912 ) | ( n17913 & n17912 ) ;
  assign n17915 = n5972 | n16094 ;
  assign n17916 = n17914 &  n17915 ;
  assign n17917 = x17 &  n17916 ;
  assign n17918 = x17 | n17916 ;
  assign n17919 = ~n17917 & n17918 ;
  assign n17920 = ( n16851 & ~n16861 ) | ( n16851 & n16946 ) | ( ~n16861 & n16946 ) ;
  assign n17921 = ( n16861 & ~n16947 ) | ( n16861 & n17920 ) | ( ~n16947 & n17920 ) ;
  assign n17928 = ~n6395 & n15897 ;
  assign n17925 = n5970 | n15320 ;
  assign n17926 = n6170 | n15700 ;
  assign n17927 = n17925 &  n17926 ;
  assign n17929 = ( n6395 & n17928 ) | ( n6395 & n17927 ) | ( n17928 & n17927 ) ;
  assign n17930 = ( n15900 & ~n5972 ) | ( n15900 & n17929 ) | ( ~n5972 & n17929 ) ;
  assign n17931 = ~n15900 & n17930 ;
  assign n17932 = ( x17 & ~n17929 ) | ( x17 & n17931 ) | ( ~n17929 & n17931 ) ;
  assign n17933 = ( n17929 & ~x17 ) | ( n17929 & n17931 ) | ( ~x17 & n17931 ) ;
  assign n17934 = ( n17932 & ~n17931 ) | ( n17932 & n17933 ) | ( ~n17931 & n17933 ) ;
  assign n17922 = ( n16873 & ~n16871 ) | ( n16873 & n16945 ) | ( ~n16871 & n16945 ) ;
  assign n17923 = ( n16871 & ~n16945 ) | ( n16871 & n16873 ) | ( ~n16945 & n16873 ) ;
  assign n17924 = ( n17922 & ~n16873 ) | ( n17922 & n17923 ) | ( ~n16873 & n17923 ) ;
  assign n17935 = ( n16886 & ~n16876 ) | ( n16886 & n16944 ) | ( ~n16876 & n16944 ) ;
  assign n17936 = ( n16876 & ~n16944 ) | ( n16876 & n16886 ) | ( ~n16944 & n16886 ) ;
  assign n17937 = ( n17935 & ~n16886 ) | ( n17935 & n17936 ) | ( ~n16886 & n17936 ) ;
  assign n17941 = ~n6395 & n15700 ;
  assign n17938 = n5970 | n15325 ;
  assign n17939 = n6170 | n15320 ;
  assign n17940 = n17938 &  n17939 ;
  assign n17942 = ( n6395 & n17941 ) | ( n6395 & n17940 ) | ( n17941 & n17940 ) ;
  assign n17943 = ( n15708 & ~n5972 ) | ( n15708 & n17942 ) | ( ~n5972 & n17942 ) ;
  assign n17944 = ~n15708 & n17943 ;
  assign n17946 = ( x17 & n17942 ) | ( x17 & n17944 ) | ( n17942 & n17944 ) ;
  assign n17945 = ( x17 & ~n17944 ) | ( x17 & n17942 ) | ( ~n17944 & n17942 ) ;
  assign n17947 = ( n17944 & ~n17946 ) | ( n17944 & n17945 ) | ( ~n17946 & n17945 ) ;
  assign n17948 = ( n16896 & ~n16943 ) | ( n16896 & n16901 ) | ( ~n16943 & n16901 ) ;
  assign n17949 = ( n16901 & ~n16896 ) | ( n16901 & n16943 ) | ( ~n16896 & n16943 ) ;
  assign n17950 = ( n17948 & ~n16901 ) | ( n17948 & n17949 ) | ( ~n16901 & n17949 ) ;
  assign n17954 = ~n6395 & n15320 ;
  assign n17951 = n5970 | n15322 ;
  assign n17952 = n6170 | n15325 ;
  assign n17953 = n17951 &  n17952 ;
  assign n17955 = ( n6395 & n17954 ) | ( n6395 & n17953 ) | ( n17954 & n17953 ) ;
  assign n17956 = ( n15334 & ~n5972 ) | ( n15334 & n17955 ) | ( ~n5972 & n17955 ) ;
  assign n17957 = ~n15334 & n17956 ;
  assign n17958 = ( x17 & ~n17955 ) | ( x17 & n17957 ) | ( ~n17955 & n17957 ) ;
  assign n17959 = ( n17955 & ~x17 ) | ( n17955 & n17957 ) | ( ~x17 & n17957 ) ;
  assign n17960 = ( n17958 & ~n17957 ) | ( n17958 & n17959 ) | ( ~n17957 & n17959 ) ;
  assign n17964 = ~n6395 & n15325 ;
  assign n17961 = ~n5970 & n14745 ;
  assign n17962 = n6170 | n15322 ;
  assign n17963 = ~n17961 & n17962 ;
  assign n17965 = ( n6395 & n17964 ) | ( n6395 & n17963 ) | ( n17964 & n17963 ) ;
  assign n17966 = n5972 | n15346 ;
  assign n17967 = n17965 &  n17966 ;
  assign n17968 = x17 &  n17967 ;
  assign n17969 = x17 | n17967 ;
  assign n17970 = ~n17968 & n17969 ;
  assign n17971 = ( n16915 & ~n16905 ) | ( n16915 & n16942 ) | ( ~n16905 & n16942 ) ;
  assign n17972 = ( n16943 & ~n16915 ) | ( n16943 & n17971 ) | ( ~n16915 & n17971 ) ;
  assign n17974 = ( n16751 & n16931 ) | ( n16751 & n16941 ) | ( n16931 & n16941 ) ;
  assign n17973 = ( n16751 & ~n16931 ) | ( n16751 & n16941 ) | ( ~n16931 & n16941 ) ;
  assign n17975 = ( n16931 & ~n17974 ) | ( n16931 & n17973 ) | ( ~n17974 & n17973 ) ;
  assign n17979 = ~n6395 & n15322 ;
  assign n17976 = n5970 | n14528 ;
  assign n17977 = ~n6170 & n14745 ;
  assign n17978 = ( n17976 & ~n17977 ) | ( n17976 & 1'b0 ) | ( ~n17977 & 1'b0 ) ;
  assign n17980 = ( n6395 & n17979 ) | ( n6395 & n17978 ) | ( n17979 & n17978 ) ;
  assign n17981 = ( n5972 & ~n17980 ) | ( n5972 & n15361 ) | ( ~n17980 & n15361 ) ;
  assign n17982 = ( n15361 & ~n17981 ) | ( n15361 & 1'b0 ) | ( ~n17981 & 1'b0 ) ;
  assign n17983 = ( x17 & ~n17980 ) | ( x17 & n17982 ) | ( ~n17980 & n17982 ) ;
  assign n17984 = ( n17980 & ~x17 ) | ( n17980 & n17982 ) | ( ~x17 & n17982 ) ;
  assign n17985 = ( n17983 & ~n17982 ) | ( n17983 & n17984 ) | ( ~n17982 & n17984 ) ;
  assign n17989 = n14745 | n6395 ;
  assign n17986 = n5970 | n14261 ;
  assign n17987 = n6170 | n14528 ;
  assign n17988 = n17986 &  n17987 ;
  assign n17990 = ( n6395 & ~n17989 ) | ( n6395 & n17988 ) | ( ~n17989 & n17988 ) ;
  assign n17991 = ~n5972 & n14749 ;
  assign n17992 = ( n17990 & ~n17991 ) | ( n17990 & 1'b0 ) | ( ~n17991 & 1'b0 ) ;
  assign n17993 = x17 &  n17992 ;
  assign n17994 = x17 | n17992 ;
  assign n17995 = ~n17993 & n17994 ;
  assign n17996 = ( x20 & n16916 ) | ( x20 & n16921 ) | ( n16916 & n16921 ) ;
  assign n17997 = ~n16916 & n17996 ;
  assign n17998 = ( n16928 & ~x20 ) | ( n16928 & n17997 ) | ( ~x20 & n17997 ) ;
  assign n17999 = ( x20 & ~n16928 ) | ( x20 & n17997 ) | ( ~n16928 & n17997 ) ;
  assign n18000 = ( n17998 & ~n17997 ) | ( n17998 & n17999 ) | ( ~n17997 & n17999 ) ;
  assign n18001 = x20 &  n16916 ;
  assign n18002 = n16921 &  n18001 ;
  assign n18003 = n16921 | n18001 ;
  assign n18004 = ~n18002 & n18003 ;
  assign n18034 = ~n6395 & n14261 ;
  assign n18031 = n5970 | n13785 ;
  assign n18032 = n6170 | n13998 ;
  assign n18033 = n18031 &  n18032 ;
  assign n18035 = ( n6395 & n18034 ) | ( n6395 & n18033 ) | ( n18034 & n18033 ) ;
  assign n18036 = n5972 | n14267 ;
  assign n18037 = n18035 &  n18036 ;
  assign n18038 = x17 &  n18037 ;
  assign n18039 = x17 | n18037 ;
  assign n18040 = ~n18038 & n18039 ;
  assign n18015 = ( n5965 & ~n13787 ) | ( n5965 & 1'b0 ) | ( ~n13787 & 1'b0 ) ;
  assign n18019 = n13790 | n5972 ;
  assign n18016 = n6170 | n13787 ;
  assign n18017 = n6395 | n13785 ;
  assign n18018 = n18016 &  n18017 ;
  assign n18020 = ( n5972 & ~n18019 ) | ( n5972 & n18018 ) | ( ~n18019 & n18018 ) ;
  assign n18026 = ~n5972 & n14001 ;
  assign n18024 = ~n6395 & n13998 ;
  assign n18021 = n5970 | n13787 ;
  assign n18022 = n6170 | n13785 ;
  assign n18023 = n18021 &  n18022 ;
  assign n18025 = ( n6395 & n18024 ) | ( n6395 & n18023 ) | ( n18024 & n18023 ) ;
  assign n18027 = ( n5972 & n18026 ) | ( n5972 & n18025 ) | ( n18026 & n18025 ) ;
  assign n18028 = ( n18015 & n18020 ) | ( n18015 & n18027 ) | ( n18020 & n18027 ) ;
  assign n18029 = ( x17 & ~n18028 ) | ( x17 & n18015 ) | ( ~n18028 & n18015 ) ;
  assign n18030 = ( x17 & ~n18029 ) | ( x17 & 1'b0 ) | ( ~n18029 & 1'b0 ) ;
  assign n18041 = ( n16916 & ~n18040 ) | ( n16916 & n18030 ) | ( ~n18040 & n18030 ) ;
  assign n18008 = ~n6395 & n14528 ;
  assign n18005 = n5970 | n13998 ;
  assign n18006 = n6170 | n14261 ;
  assign n18007 = n18005 &  n18006 ;
  assign n18009 = ( n6395 & n18008 ) | ( n6395 & n18007 ) | ( n18008 & n18007 ) ;
  assign n18010 = ( n14532 & ~n5972 ) | ( n14532 & n18009 ) | ( ~n5972 & n18009 ) ;
  assign n18011 = ~n14532 & n18010 ;
  assign n18012 = ( x17 & ~n18009 ) | ( x17 & n18011 ) | ( ~n18009 & n18011 ) ;
  assign n18013 = ( n18009 & ~x17 ) | ( n18009 & n18011 ) | ( ~x17 & n18011 ) ;
  assign n18014 = ( n18012 & ~n18011 ) | ( n18012 & n18013 ) | ( ~n18011 & n18013 ) ;
  assign n18042 = ( n18004 & ~n18041 ) | ( n18004 & n18014 ) | ( ~n18041 & n18014 ) ;
  assign n18043 = ( n17995 & n18000 ) | ( n17995 & n18042 ) | ( n18000 & n18042 ) ;
  assign n18044 = ( n17975 & n17985 ) | ( n17975 & n18043 ) | ( n17985 & n18043 ) ;
  assign n18045 = ( n17970 & ~n17972 ) | ( n17970 & n18044 ) | ( ~n17972 & n18044 ) ;
  assign n18046 = ( n17950 & n17960 ) | ( n17950 & n18045 ) | ( n17960 & n18045 ) ;
  assign n18047 = ( n17937 & n17947 ) | ( n17937 & n18046 ) | ( n17947 & n18046 ) ;
  assign n18048 = ( n17934 & ~n17924 ) | ( n17934 & n18047 ) | ( ~n17924 & n18047 ) ;
  assign n18049 = ( n17919 & n17921 ) | ( n17919 & n18048 ) | ( n17921 & n18048 ) ;
  assign n18050 = ( n17907 & n17909 ) | ( n17907 & n18049 ) | ( n17909 & n18049 ) ;
  assign n18051 = ( n17895 & ~n17897 ) | ( n17895 & n18050 ) | ( ~n17897 & n18050 ) ;
  assign n18052 = ( n17875 & n17885 ) | ( n17875 & n18051 ) | ( n17885 & n18051 ) ;
  assign n18053 = ( n17862 & n17872 ) | ( n17862 & n18052 ) | ( n17872 & n18052 ) ;
  assign n18054 = ( n17857 & n17859 ) | ( n17857 & n18053 ) | ( n17859 & n18053 ) ;
  assign n18055 = ( n17844 & ~n17847 ) | ( n17844 & n18054 ) | ( ~n17847 & n18054 ) ;
  assign n18056 = ( n17831 & n17834 ) | ( n17831 & n18055 ) | ( n17834 & n18055 ) ;
  assign n18057 = ( n17816 & n17819 ) | ( n17816 & n18056 ) | ( n17819 & n18056 ) ;
  assign n17780 = ( n17773 & ~n17771 ) | ( n17773 & n17779 ) | ( ~n17771 & n17779 ) ;
  assign n17651 = ( n17581 & ~n17633 ) | ( n17581 & n17634 ) | ( ~n17633 & n17634 ) ;
  assign n17674 = ~x11 & n17591 ;
  assign n17675 = ( n17611 & ~n17614 ) | ( n17611 & n17674 ) | ( ~n17614 & n17674 ) ;
  assign n17652 = n813 &  n5472 ;
  assign n17653 = ~n206 & n17652 ;
  assign n17654 = ( n889 & n5649 ) | ( n889 & n17653 ) | ( n5649 & n17653 ) ;
  assign n17655 = ~n889 & n17654 ;
  assign n17656 = ( n1304 & n3581 ) | ( n1304 & n17655 ) | ( n3581 & n17655 ) ;
  assign n17657 = ~n3581 & n17656 ;
  assign n17658 = ( n2043 & ~n17657 ) | ( n2043 & n3890 ) | ( ~n17657 & n3890 ) ;
  assign n17659 = ( n2043 & ~n17658 ) | ( n2043 & 1'b0 ) | ( ~n17658 & 1'b0 ) ;
  assign n17660 = ( n787 & ~n257 ) | ( n787 & n17659 ) | ( ~n257 & n17659 ) ;
  assign n17661 = ~n787 & n17660 ;
  assign n17662 = ( n745 & ~n962 ) | ( n745 & n17661 ) | ( ~n962 & n17661 ) ;
  assign n17663 = ( n17662 & ~n745 ) | ( n17662 & 1'b0 ) | ( ~n745 & 1'b0 ) ;
  assign n17664 = ( n117 & ~n568 ) | ( n117 & n17663 ) | ( ~n568 & n17663 ) ;
  assign n17665 = ~n117 & n17664 ;
  assign n17666 = ~n95 & n17665 ;
  assign n17672 = ~n3644 & n12369 ;
  assign n17667 = n3653 | n11113 ;
  assign n17668 = n3657 &  n11116 ;
  assign n17669 = n3652 &  n11119 ;
  assign n17670 = n17668 | n17669 ;
  assign n17671 = ( n17667 & ~n17670 ) | ( n17667 & 1'b0 ) | ( ~n17670 & 1'b0 ) ;
  assign n17673 = ( n3644 & n17672 ) | ( n3644 & n17671 ) | ( n17672 & n17671 ) ;
  assign n17677 = ( n17666 & n17673 ) | ( n17666 & n17675 ) | ( n17673 & n17675 ) ;
  assign n17676 = ( n17666 & ~n17675 ) | ( n17666 & n17673 ) | ( ~n17675 & n17673 ) ;
  assign n17678 = ( n17675 & ~n17677 ) | ( n17675 & n17676 ) | ( ~n17677 & n17676 ) ;
  assign n17679 = ~n17617 & n17678 ;
  assign n17680 = ( n17617 & ~n17678 ) | ( n17617 & 1'b0 ) | ( ~n17678 & 1'b0 ) ;
  assign n17681 = n17679 | n17680 ;
  assign n17687 = n12662 | n601 ;
  assign n17685 = ~n4430 & n11104 ;
  assign n17682 = n523 | n11110 ;
  assign n17683 = ~n3939 & n11107 ;
  assign n17684 = ( n17682 & ~n17683 ) | ( n17682 & 1'b0 ) | ( ~n17683 & 1'b0 ) ;
  assign n17686 = ( n4430 & n17685 ) | ( n4430 & n17684 ) | ( n17685 & n17684 ) ;
  assign n17688 = ( n601 & ~n17687 ) | ( n601 & n17686 ) | ( ~n17687 & n17686 ) ;
  assign n17689 = ( n17681 & ~x29 ) | ( n17681 & n17688 ) | ( ~x29 & n17688 ) ;
  assign n17690 = ( x29 & ~n17681 ) | ( x29 & n17688 ) | ( ~n17681 & n17688 ) ;
  assign n17691 = ( n17689 & ~n17688 ) | ( n17689 & n17690 ) | ( ~n17688 & n17690 ) ;
  assign n17692 = ( n17619 & ~n17620 ) | ( n17619 & n17630 ) | ( ~n17620 & n17630 ) ;
  assign n17696 = ~n4962 & n11095 ;
  assign n17693 = n4482 | n11101 ;
  assign n17694 = n4495 | n11098 ;
  assign n17695 = n17693 &  n17694 ;
  assign n17697 = ( n4962 & n17696 ) | ( n4962 & n17695 ) | ( n17696 & n17695 ) ;
  assign n17698 = n4478 | n13014 ;
  assign n17699 = n17697 &  n17698 ;
  assign n17700 = x26 &  n17699 ;
  assign n17701 = x26 | n17699 ;
  assign n17702 = ~n17700 & n17701 ;
  assign n17703 = ( n17691 & ~n17692 ) | ( n17691 & n17702 ) | ( ~n17692 & n17702 ) ;
  assign n17704 = ( n17691 & ~n17702 ) | ( n17691 & n17692 ) | ( ~n17702 & n17692 ) ;
  assign n17705 = ( n17703 & ~n17691 ) | ( n17703 & n17704 ) | ( ~n17691 & n17704 ) ;
  assign n17709 = ~n5135 & n11081 ;
  assign n17706 = n5010 | n11093 ;
  assign n17707 = n5067 | n11091 ;
  assign n17708 = n17706 &  n17707 ;
  assign n17710 = ( n5135 & n17709 ) | ( n5135 & n17708 ) | ( n17709 & n17708 ) ;
  assign n17711 = n5012 | n13775 ;
  assign n17712 = n17710 &  n17711 ;
  assign n17713 = x23 &  n17712 ;
  assign n17714 = x23 | n17712 ;
  assign n17715 = ~n17713 & n17714 ;
  assign n17716 = ( n17651 & n17705 ) | ( n17651 & n17715 ) | ( n17705 & n17715 ) ;
  assign n17717 = ( n17705 & ~n17651 ) | ( n17705 & n17715 ) | ( ~n17651 & n17715 ) ;
  assign n17718 = ( n17651 & ~n17716 ) | ( n17651 & n17717 ) | ( ~n17716 & n17717 ) ;
  assign n17722 = ~n5837 & n13836 ;
  assign n17719 = ( n5339 & ~n11085 ) | ( n5339 & 1'b0 ) | ( ~n11085 & 1'b0 ) ;
  assign n17720 = n5761 | n11078 ;
  assign n17721 = ~n17719 & n17720 ;
  assign n17723 = ( n5837 & n17722 ) | ( n5837 & n17721 ) | ( n17722 & n17721 ) ;
  assign n17724 = n5341 | n13844 ;
  assign n17725 = n17723 &  n17724 ;
  assign n17726 = x20 &  n17725 ;
  assign n17727 = x20 | n17725 ;
  assign n17728 = ~n17726 & n17727 ;
  assign n17729 = ( n17639 & n17718 ) | ( n17639 & n17728 ) | ( n17718 & n17728 ) ;
  assign n17730 = ( n17718 & ~n17639 ) | ( n17718 & n17728 ) | ( ~n17639 & n17728 ) ;
  assign n17731 = ( n17639 & ~n17729 ) | ( n17639 & n17730 ) | ( ~n17729 & n17730 ) ;
  assign n17735 = n14553 | n6395 ;
  assign n17732 = n5970 | n14071 ;
  assign n17733 = n6170 | n14355 ;
  assign n17734 = n17732 &  n17733 ;
  assign n17736 = ( n6395 & ~n17735 ) | ( n6395 & n17734 ) | ( ~n17735 & n17734 ) ;
  assign n17737 = ~n5972 & n14562 ;
  assign n17738 = ( n17736 & ~n17737 ) | ( n17736 & 1'b0 ) | ( ~n17737 & 1'b0 ) ;
  assign n17739 = x17 &  n17738 ;
  assign n17740 = x17 | n17738 ;
  assign n17741 = ~n17739 & n17740 ;
  assign n17742 = ( n17643 & n17731 ) | ( n17643 & n17741 ) | ( n17731 & n17741 ) ;
  assign n17743 = ( n17731 & ~n17643 ) | ( n17731 & n17741 ) | ( ~n17643 & n17741 ) ;
  assign n17744 = ( n17643 & ~n17742 ) | ( n17643 & n17743 ) | ( ~n17742 & n17743 ) ;
  assign n17748 = n14800 | n7097 ;
  assign n17745 = n6530 | n14803 ;
  assign n17746 = ~n6983 & n14807 ;
  assign n17747 = ( n17745 & ~n17746 ) | ( n17745 & 1'b0 ) | ( ~n17746 & 1'b0 ) ;
  assign n17749 = ( n7097 & ~n17748 ) | ( n7097 & n17747 ) | ( ~n17748 & n17747 ) ;
  assign n17750 = n6532 | n14816 ;
  assign n17751 = n17749 &  n17750 ;
  assign n17752 = x14 &  n17751 ;
  assign n17753 = x14 | n17751 ;
  assign n17754 = ~n17752 & n17753 ;
  assign n17755 = ( n17647 & n17744 ) | ( n17647 & n17754 ) | ( n17744 & n17754 ) ;
  assign n17756 = ( n17744 & ~n17647 ) | ( n17744 & n17754 ) | ( ~n17647 & n17754 ) ;
  assign n17757 = ( n17647 & ~n17755 ) | ( n17647 & n17756 ) | ( ~n17755 & n17756 ) ;
  assign n17781 = ( n17650 & ~n17780 ) | ( n17650 & n17757 ) | ( ~n17780 & n17757 ) ;
  assign n17782 = ( n17650 & ~n17757 ) | ( n17650 & n17780 ) | ( ~n17757 & n17780 ) ;
  assign n17783 = ( n17781 & ~n17650 ) | ( n17781 & n17782 ) | ( ~n17650 & n17782 ) ;
  assign n17784 = ( n6395 & ~n17783 ) | ( n6395 & 1'b0 ) | ( ~n17783 & 1'b0 ) ;
  assign n17788 = n5970 | n17787 ;
  assign n17792 = n6170 | n17791 ;
  assign n17793 = n17788 &  n17792 ;
  assign n17794 = ( n17783 & n17784 ) | ( n17783 & n17793 ) | ( n17784 & n17793 ) ;
  assign n17798 = ( n17783 & n17791 ) | ( n17783 & n17796 ) | ( n17791 & n17796 ) ;
  assign n17797 = ( n17783 & ~n17791 ) | ( n17783 & n17796 ) | ( ~n17791 & n17796 ) ;
  assign n17799 = ( n17791 & ~n17798 ) | ( n17791 & n17797 ) | ( ~n17798 & n17797 ) ;
  assign n17800 = n5972 | n17799 ;
  assign n17801 = n17794 &  n17800 ;
  assign n17802 = x17 &  n17801 ;
  assign n17803 = x17 | n17801 ;
  assign n17804 = ~n17802 & n17803 ;
  assign n18058 = ( n17421 & ~n18057 ) | ( n17421 & n17804 ) | ( ~n18057 & n17804 ) ;
  assign n18059 = ( n17421 & ~n17804 ) | ( n17421 & n18057 ) | ( ~n17804 & n18057 ) ;
  assign n18060 = ( n18058 & ~n17421 ) | ( n18058 & n18059 ) | ( ~n17421 & n18059 ) ;
  assign n18064 = ( n7097 & ~n17783 ) | ( n7097 & 1'b0 ) | ( ~n17783 & 1'b0 ) ;
  assign n18065 = n6530 | n17787 ;
  assign n18066 = n6983 | n17791 ;
  assign n18067 = n18065 &  n18066 ;
  assign n18068 = ( n17783 & n18064 ) | ( n17783 & n18067 ) | ( n18064 & n18067 ) ;
  assign n18069 = ( n6532 & ~n17799 ) | ( n6532 & n18068 ) | ( ~n17799 & n18068 ) ;
  assign n18070 = ~n6532 & n18069 ;
  assign n18072 = ( x14 & n18068 ) | ( x14 & n18070 ) | ( n18068 & n18070 ) ;
  assign n18071 = ( x14 & ~n18070 ) | ( x14 & n18068 ) | ( ~n18070 & n18068 ) ;
  assign n18073 = ( n18070 & ~n18072 ) | ( n18070 & n18071 ) | ( ~n18072 & n18071 ) ;
  assign n18061 = ( n17844 & ~n18054 ) | ( n17844 & n17847 ) | ( ~n18054 & n17847 ) ;
  assign n18062 = ( n17847 & ~n17844 ) | ( n17847 & n18054 ) | ( ~n17844 & n18054 ) ;
  assign n18063 = ( n18061 & ~n17847 ) | ( n18061 & n18062 ) | ( ~n17847 & n18062 ) ;
  assign n18074 = ( n17859 & ~n17857 ) | ( n17859 & n18053 ) | ( ~n17857 & n18053 ) ;
  assign n18075 = ( n17857 & ~n18053 ) | ( n17857 & n17859 ) | ( ~n18053 & n17859 ) ;
  assign n18076 = ( n18074 & ~n17859 ) | ( n18074 & n18075 ) | ( ~n17859 & n18075 ) ;
  assign n18080 = ~n7097 & n17791 ;
  assign n18077 = n6530 | n17405 ;
  assign n18078 = n6983 | n17787 ;
  assign n18079 = n18077 &  n18078 ;
  assign n18081 = ( n7097 & n18080 ) | ( n7097 & n18079 ) | ( n18080 & n18079 ) ;
  assign n18082 = ( n6532 & ~n17811 ) | ( n6532 & n18081 ) | ( ~n17811 & n18081 ) ;
  assign n18083 = ~n6532 & n18082 ;
  assign n18085 = ( x14 & n18081 ) | ( x14 & n18083 ) | ( n18081 & n18083 ) ;
  assign n18084 = ( x14 & ~n18083 ) | ( x14 & n18081 ) | ( ~n18083 & n18081 ) ;
  assign n18086 = ( n18083 & ~n18085 ) | ( n18083 & n18084 ) | ( ~n18085 & n18084 ) ;
  assign n18090 = ~n7097 & n17787 ;
  assign n18087 = n6530 | n17263 ;
  assign n18088 = n6983 | n17405 ;
  assign n18089 = n18087 &  n18088 ;
  assign n18091 = ( n7097 & n18090 ) | ( n7097 & n18089 ) | ( n18090 & n18089 ) ;
  assign n18092 = ( n6532 & ~n17826 ) | ( n6532 & n18091 ) | ( ~n17826 & n18091 ) ;
  assign n18093 = ~n6532 & n18092 ;
  assign n18094 = ( x14 & ~n18091 ) | ( x14 & n18093 ) | ( ~n18091 & n18093 ) ;
  assign n18095 = ( n18091 & ~x14 ) | ( n18091 & n18093 ) | ( ~x14 & n18093 ) ;
  assign n18096 = ( n18094 & ~n18093 ) | ( n18094 & n18095 ) | ( ~n18093 & n18095 ) ;
  assign n18097 = ( n17862 & ~n17872 ) | ( n17862 & n18052 ) | ( ~n17872 & n18052 ) ;
  assign n18098 = ( n17872 & ~n18053 ) | ( n17872 & n18097 ) | ( ~n18053 & n18097 ) ;
  assign n18102 = ~n7097 & n17405 ;
  assign n18099 = ~n6530 & n17107 ;
  assign n18100 = n6983 | n17263 ;
  assign n18101 = ~n18099 & n18100 ;
  assign n18103 = ( n7097 & n18102 ) | ( n7097 & n18101 ) | ( n18102 & n18101 ) ;
  assign n18104 = n6532 | n17413 ;
  assign n18105 = n18103 &  n18104 ;
  assign n18106 = x14 &  n18105 ;
  assign n18107 = x14 | n18105 ;
  assign n18108 = ~n18106 & n18107 ;
  assign n18109 = ( n17875 & ~n17885 ) | ( n17875 & n18051 ) | ( ~n17885 & n18051 ) ;
  assign n18110 = ( n17885 & ~n18052 ) | ( n17885 & n18109 ) | ( ~n18052 & n18109 ) ;
  assign n18117 = ~n7097 & n17263 ;
  assign n18114 = n6530 | n16589 ;
  assign n18115 = ~n6983 & n17107 ;
  assign n18116 = ( n18114 & ~n18115 ) | ( n18114 & 1'b0 ) | ( ~n18115 & 1'b0 ) ;
  assign n18118 = ( n7097 & n18117 ) | ( n7097 & n18116 ) | ( n18117 & n18116 ) ;
  assign n18119 = ( n6532 & ~n18118 ) | ( n6532 & n17271 ) | ( ~n18118 & n17271 ) ;
  assign n18120 = ( n17271 & ~n18119 ) | ( n17271 & 1'b0 ) | ( ~n18119 & 1'b0 ) ;
  assign n18122 = ( x14 & n18118 ) | ( x14 & n18120 ) | ( n18118 & n18120 ) ;
  assign n18121 = ( x14 & ~n18120 ) | ( x14 & n18118 ) | ( ~n18120 & n18118 ) ;
  assign n18123 = ( n18120 & ~n18122 ) | ( n18120 & n18121 ) | ( ~n18122 & n18121 ) ;
  assign n18111 = ( n17897 & ~n17895 ) | ( n17897 & n18050 ) | ( ~n17895 & n18050 ) ;
  assign n18112 = ( n17895 & ~n18050 ) | ( n17895 & n17897 ) | ( ~n18050 & n17897 ) ;
  assign n18113 = ( n18111 & ~n17897 ) | ( n18111 & n18112 ) | ( ~n17897 & n18112 ) ;
  assign n18124 = ( n17909 & ~n17907 ) | ( n17909 & n18049 ) | ( ~n17907 & n18049 ) ;
  assign n18125 = ( n17907 & ~n18049 ) | ( n17907 & n17909 ) | ( ~n18049 & n17909 ) ;
  assign n18126 = ( n18124 & ~n17909 ) | ( n18124 & n18125 ) | ( ~n17909 & n18125 ) ;
  assign n18130 = n17107 | n7097 ;
  assign n18127 = n6530 | n16595 ;
  assign n18128 = n6983 | n16589 ;
  assign n18129 = n18127 &  n18128 ;
  assign n18131 = ( n7097 & ~n18130 ) | ( n7097 & n18129 ) | ( ~n18130 & n18129 ) ;
  assign n18132 = ( n6532 & ~n18131 ) | ( n6532 & n17115 ) | ( ~n18131 & n17115 ) ;
  assign n18133 = ( n17115 & ~n18132 ) | ( n17115 & 1'b0 ) | ( ~n18132 & 1'b0 ) ;
  assign n18134 = ( x14 & ~n18131 ) | ( x14 & n18133 ) | ( ~n18131 & n18133 ) ;
  assign n18135 = ( n18131 & ~x14 ) | ( n18131 & n18133 ) | ( ~x14 & n18133 ) ;
  assign n18136 = ( n18134 & ~n18133 ) | ( n18134 & n18135 ) | ( ~n18133 & n18135 ) ;
  assign n18137 = ( n17921 & ~n17919 ) | ( n17921 & n18048 ) | ( ~n17919 & n18048 ) ;
  assign n18138 = ( n17919 & ~n18048 ) | ( n17919 & n17921 ) | ( ~n18048 & n17921 ) ;
  assign n18139 = ( n18137 & ~n17921 ) | ( n18137 & n18138 ) | ( ~n17921 & n18138 ) ;
  assign n18143 = ~n7097 & n16589 ;
  assign n18140 = n6530 | n16591 ;
  assign n18141 = n6983 | n16595 ;
  assign n18142 = n18140 &  n18141 ;
  assign n18144 = ( n7097 & n18143 ) | ( n7097 & n18142 ) | ( n18143 & n18142 ) ;
  assign n18145 = ( n16604 & ~n6532 ) | ( n16604 & n18144 ) | ( ~n6532 & n18144 ) ;
  assign n18146 = ~n16604 & n18145 ;
  assign n18148 = ( x14 & n18144 ) | ( x14 & n18146 ) | ( n18144 & n18146 ) ;
  assign n18147 = ( x14 & ~n18146 ) | ( x14 & n18144 ) | ( ~n18146 & n18144 ) ;
  assign n18149 = ( n18146 & ~n18148 ) | ( n18146 & n18147 ) | ( ~n18148 & n18147 ) ;
  assign n18153 = ~n7097 & n16595 ;
  assign n18150 = n6530 | n16091 ;
  assign n18151 = n6983 | n16591 ;
  assign n18152 = n18150 &  n18151 ;
  assign n18154 = ( n7097 & n18153 ) | ( n7097 & n18152 ) | ( n18153 & n18152 ) ;
  assign n18155 = n6532 | n16616 ;
  assign n18156 = n18154 &  n18155 ;
  assign n18157 = x14 &  n18156 ;
  assign n18158 = x14 | n18156 ;
  assign n18159 = ~n18157 & n18158 ;
  assign n18160 = ( n17924 & ~n18047 ) | ( n17924 & n17934 ) | ( ~n18047 & n17934 ) ;
  assign n18161 = ( n18048 & ~n17934 ) | ( n18048 & n18160 ) | ( ~n17934 & n18160 ) ;
  assign n18165 = ~n7097 & n16591 ;
  assign n18162 = n6530 | n15897 ;
  assign n18163 = n6983 | n16091 ;
  assign n18164 = n18162 &  n18163 ;
  assign n18166 = ( n7097 & n18165 ) | ( n7097 & n18164 ) | ( n18165 & n18164 ) ;
  assign n18167 = n6532 | n16631 ;
  assign n18168 = n18166 &  n18167 ;
  assign n18169 = x14 &  n18168 ;
  assign n18170 = x14 | n18168 ;
  assign n18171 = ~n18169 & n18170 ;
  assign n18172 = ( n17937 & ~n17947 ) | ( n17937 & n18046 ) | ( ~n17947 & n18046 ) ;
  assign n18173 = ( n17947 & ~n18047 ) | ( n17947 & n18172 ) | ( ~n18047 & n18172 ) ;
  assign n18177 = ~n7097 & n16091 ;
  assign n18174 = n6530 | n15700 ;
  assign n18175 = n6983 | n15897 ;
  assign n18176 = n18174 &  n18175 ;
  assign n18178 = ( n7097 & n18177 ) | ( n7097 & n18176 ) | ( n18177 & n18176 ) ;
  assign n18179 = n6532 | n16094 ;
  assign n18180 = n18178 &  n18179 ;
  assign n18181 = x14 &  n18180 ;
  assign n18182 = x14 | n18180 ;
  assign n18183 = ~n18181 & n18182 ;
  assign n18184 = ( n17950 & ~n17960 ) | ( n17950 & n18045 ) | ( ~n17960 & n18045 ) ;
  assign n18185 = ( n17960 & ~n18046 ) | ( n17960 & n18184 ) | ( ~n18046 & n18184 ) ;
  assign n18192 = ~n7097 & n15897 ;
  assign n18189 = n6530 | n15320 ;
  assign n18190 = n6983 | n15700 ;
  assign n18191 = n18189 &  n18190 ;
  assign n18193 = ( n7097 & n18192 ) | ( n7097 & n18191 ) | ( n18192 & n18191 ) ;
  assign n18194 = ( n15900 & ~n6532 ) | ( n15900 & n18193 ) | ( ~n6532 & n18193 ) ;
  assign n18195 = ~n15900 & n18194 ;
  assign n18196 = ( x14 & ~n18193 ) | ( x14 & n18195 ) | ( ~n18193 & n18195 ) ;
  assign n18197 = ( n18193 & ~x14 ) | ( n18193 & n18195 ) | ( ~x14 & n18195 ) ;
  assign n18198 = ( n18196 & ~n18195 ) | ( n18196 & n18197 ) | ( ~n18195 & n18197 ) ;
  assign n18186 = ( n17972 & ~n17970 ) | ( n17972 & n18044 ) | ( ~n17970 & n18044 ) ;
  assign n18187 = ( n17970 & ~n18044 ) | ( n17970 & n17972 ) | ( ~n18044 & n17972 ) ;
  assign n18188 = ( n18186 & ~n17972 ) | ( n18186 & n18187 ) | ( ~n17972 & n18187 ) ;
  assign n18199 = ( n17985 & ~n17975 ) | ( n17985 & n18043 ) | ( ~n17975 & n18043 ) ;
  assign n18200 = ( n17975 & ~n18043 ) | ( n17975 & n17985 ) | ( ~n18043 & n17985 ) ;
  assign n18201 = ( n18199 & ~n17985 ) | ( n18199 & n18200 ) | ( ~n17985 & n18200 ) ;
  assign n18205 = ~n7097 & n15700 ;
  assign n18202 = n6530 | n15325 ;
  assign n18203 = n6983 | n15320 ;
  assign n18204 = n18202 &  n18203 ;
  assign n18206 = ( n7097 & n18205 ) | ( n7097 & n18204 ) | ( n18205 & n18204 ) ;
  assign n18207 = ( n15708 & ~n6532 ) | ( n15708 & n18206 ) | ( ~n6532 & n18206 ) ;
  assign n18208 = ~n15708 & n18207 ;
  assign n18210 = ( x14 & n18206 ) | ( x14 & n18208 ) | ( n18206 & n18208 ) ;
  assign n18209 = ( x14 & ~n18208 ) | ( x14 & n18206 ) | ( ~n18208 & n18206 ) ;
  assign n18211 = ( n18208 & ~n18210 ) | ( n18208 & n18209 ) | ( ~n18210 & n18209 ) ;
  assign n18212 = ( n17995 & ~n18042 ) | ( n17995 & n18000 ) | ( ~n18042 & n18000 ) ;
  assign n18213 = ( n18000 & ~n17995 ) | ( n18000 & n18042 ) | ( ~n17995 & n18042 ) ;
  assign n18214 = ( n18212 & ~n18000 ) | ( n18212 & n18213 ) | ( ~n18000 & n18213 ) ;
  assign n18218 = ~n7097 & n15320 ;
  assign n18215 = n6530 | n15322 ;
  assign n18216 = n6983 | n15325 ;
  assign n18217 = n18215 &  n18216 ;
  assign n18219 = ( n7097 & n18218 ) | ( n7097 & n18217 ) | ( n18218 & n18217 ) ;
  assign n18220 = ( n15334 & ~n6532 ) | ( n15334 & n18219 ) | ( ~n6532 & n18219 ) ;
  assign n18221 = ~n15334 & n18220 ;
  assign n18222 = ( x14 & ~n18219 ) | ( x14 & n18221 ) | ( ~n18219 & n18221 ) ;
  assign n18223 = ( n18219 & ~x14 ) | ( n18219 & n18221 ) | ( ~x14 & n18221 ) ;
  assign n18224 = ( n18222 & ~n18221 ) | ( n18222 & n18223 ) | ( ~n18221 & n18223 ) ;
  assign n18228 = ~n7097 & n15325 ;
  assign n18225 = ~n6530 & n14745 ;
  assign n18226 = n6983 | n15322 ;
  assign n18227 = ~n18225 & n18226 ;
  assign n18229 = ( n7097 & n18228 ) | ( n7097 & n18227 ) | ( n18228 & n18227 ) ;
  assign n18230 = n6532 | n15346 ;
  assign n18231 = n18229 &  n18230 ;
  assign n18232 = x14 &  n18231 ;
  assign n18233 = x14 | n18231 ;
  assign n18234 = ~n18232 & n18233 ;
  assign n18235 = ( n18014 & ~n18004 ) | ( n18014 & n18041 ) | ( ~n18004 & n18041 ) ;
  assign n18236 = ( n18042 & ~n18014 ) | ( n18042 & n18235 ) | ( ~n18014 & n18235 ) ;
  assign n18238 = ( n16916 & n18030 ) | ( n16916 & n18040 ) | ( n18030 & n18040 ) ;
  assign n18237 = ( n16916 & ~n18030 ) | ( n16916 & n18040 ) | ( ~n18030 & n18040 ) ;
  assign n18239 = ( n18030 & ~n18238 ) | ( n18030 & n18237 ) | ( ~n18238 & n18237 ) ;
  assign n18243 = ~n7097 & n15322 ;
  assign n18240 = n6530 | n14528 ;
  assign n18241 = ~n6983 & n14745 ;
  assign n18242 = ( n18240 & ~n18241 ) | ( n18240 & 1'b0 ) | ( ~n18241 & 1'b0 ) ;
  assign n18244 = ( n7097 & n18243 ) | ( n7097 & n18242 ) | ( n18243 & n18242 ) ;
  assign n18245 = ( n6532 & ~n18244 ) | ( n6532 & n15361 ) | ( ~n18244 & n15361 ) ;
  assign n18246 = ( n15361 & ~n18245 ) | ( n15361 & 1'b0 ) | ( ~n18245 & 1'b0 ) ;
  assign n18247 = ( x14 & ~n18244 ) | ( x14 & n18246 ) | ( ~n18244 & n18246 ) ;
  assign n18248 = ( n18244 & ~x14 ) | ( n18244 & n18246 ) | ( ~x14 & n18246 ) ;
  assign n18249 = ( n18247 & ~n18246 ) | ( n18247 & n18248 ) | ( ~n18246 & n18248 ) ;
  assign n18253 = n14745 | n7097 ;
  assign n18250 = n6530 | n14261 ;
  assign n18251 = n6983 | n14528 ;
  assign n18252 = n18250 &  n18251 ;
  assign n18254 = ( n7097 & ~n18253 ) | ( n7097 & n18252 ) | ( ~n18253 & n18252 ) ;
  assign n18255 = ~n6532 & n14749 ;
  assign n18256 = ( n18254 & ~n18255 ) | ( n18254 & 1'b0 ) | ( ~n18255 & 1'b0 ) ;
  assign n18257 = x14 &  n18256 ;
  assign n18258 = x14 | n18256 ;
  assign n18259 = ~n18257 & n18258 ;
  assign n18260 = ( x17 & n18015 ) | ( x17 & n18020 ) | ( n18015 & n18020 ) ;
  assign n18261 = ~n18015 & n18260 ;
  assign n18262 = ( n18027 & ~x17 ) | ( n18027 & n18261 ) | ( ~x17 & n18261 ) ;
  assign n18263 = ( x17 & ~n18027 ) | ( x17 & n18261 ) | ( ~n18027 & n18261 ) ;
  assign n18264 = ( n18262 & ~n18261 ) | ( n18262 & n18263 ) | ( ~n18261 & n18263 ) ;
  assign n18265 = x17 &  n18015 ;
  assign n18266 = n18020 &  n18265 ;
  assign n18267 = n18020 | n18265 ;
  assign n18268 = ~n18266 & n18267 ;
  assign n18298 = ~n7097 & n14261 ;
  assign n18295 = n6530 | n13785 ;
  assign n18296 = n6983 | n13998 ;
  assign n18297 = n18295 &  n18296 ;
  assign n18299 = ( n7097 & n18298 ) | ( n7097 & n18297 ) | ( n18298 & n18297 ) ;
  assign n18300 = n6532 | n14267 ;
  assign n18301 = n18299 &  n18300 ;
  assign n18302 = x14 &  n18301 ;
  assign n18303 = x14 | n18301 ;
  assign n18304 = ~n18302 & n18303 ;
  assign n18279 = ( n6525 & ~n13787 ) | ( n6525 & 1'b0 ) | ( ~n13787 & 1'b0 ) ;
  assign n18283 = n13790 | n6532 ;
  assign n18280 = n6983 | n13787 ;
  assign n18281 = n7097 | n13785 ;
  assign n18282 = n18280 &  n18281 ;
  assign n18284 = ( n6532 & ~n18283 ) | ( n6532 & n18282 ) | ( ~n18283 & n18282 ) ;
  assign n18290 = ~n6532 & n14001 ;
  assign n18288 = ~n7097 & n13998 ;
  assign n18285 = n6530 | n13787 ;
  assign n18286 = n6983 | n13785 ;
  assign n18287 = n18285 &  n18286 ;
  assign n18289 = ( n7097 & n18288 ) | ( n7097 & n18287 ) | ( n18288 & n18287 ) ;
  assign n18291 = ( n6532 & n18290 ) | ( n6532 & n18289 ) | ( n18290 & n18289 ) ;
  assign n18292 = ( n18279 & n18284 ) | ( n18279 & n18291 ) | ( n18284 & n18291 ) ;
  assign n18293 = ( x14 & ~n18292 ) | ( x14 & n18279 ) | ( ~n18292 & n18279 ) ;
  assign n18294 = ( x14 & ~n18293 ) | ( x14 & 1'b0 ) | ( ~n18293 & 1'b0 ) ;
  assign n18305 = ( n18015 & ~n18304 ) | ( n18015 & n18294 ) | ( ~n18304 & n18294 ) ;
  assign n18272 = ~n7097 & n14528 ;
  assign n18269 = n6530 | n13998 ;
  assign n18270 = n6983 | n14261 ;
  assign n18271 = n18269 &  n18270 ;
  assign n18273 = ( n7097 & n18272 ) | ( n7097 & n18271 ) | ( n18272 & n18271 ) ;
  assign n18274 = ( n14532 & ~n6532 ) | ( n14532 & n18273 ) | ( ~n6532 & n18273 ) ;
  assign n18275 = ~n14532 & n18274 ;
  assign n18276 = ( x14 & ~n18273 ) | ( x14 & n18275 ) | ( ~n18273 & n18275 ) ;
  assign n18277 = ( n18273 & ~x14 ) | ( n18273 & n18275 ) | ( ~x14 & n18275 ) ;
  assign n18278 = ( n18276 & ~n18275 ) | ( n18276 & n18277 ) | ( ~n18275 & n18277 ) ;
  assign n18306 = ( n18268 & ~n18305 ) | ( n18268 & n18278 ) | ( ~n18305 & n18278 ) ;
  assign n18307 = ( n18259 & n18264 ) | ( n18259 & n18306 ) | ( n18264 & n18306 ) ;
  assign n18308 = ( n18239 & n18249 ) | ( n18239 & n18307 ) | ( n18249 & n18307 ) ;
  assign n18309 = ( n18234 & ~n18236 ) | ( n18234 & n18308 ) | ( ~n18236 & n18308 ) ;
  assign n18310 = ( n18214 & n18224 ) | ( n18214 & n18309 ) | ( n18224 & n18309 ) ;
  assign n18311 = ( n18201 & n18211 ) | ( n18201 & n18310 ) | ( n18211 & n18310 ) ;
  assign n18312 = ( n18198 & ~n18188 ) | ( n18198 & n18311 ) | ( ~n18188 & n18311 ) ;
  assign n18313 = ( n18183 & n18185 ) | ( n18183 & n18312 ) | ( n18185 & n18312 ) ;
  assign n18314 = ( n18171 & n18173 ) | ( n18171 & n18313 ) | ( n18173 & n18313 ) ;
  assign n18315 = ( n18159 & ~n18161 ) | ( n18159 & n18314 ) | ( ~n18161 & n18314 ) ;
  assign n18316 = ( n18139 & n18149 ) | ( n18139 & n18315 ) | ( n18149 & n18315 ) ;
  assign n18317 = ( n18126 & n18136 ) | ( n18126 & n18316 ) | ( n18136 & n18316 ) ;
  assign n18318 = ( n18123 & ~n18113 ) | ( n18123 & n18317 ) | ( ~n18113 & n18317 ) ;
  assign n18319 = ( n18108 & n18110 ) | ( n18108 & n18318 ) | ( n18110 & n18318 ) ;
  assign n18320 = ( n18096 & n18098 ) | ( n18096 & n18319 ) | ( n18098 & n18319 ) ;
  assign n18321 = ( n18076 & n18086 ) | ( n18076 & n18320 ) | ( n18086 & n18320 ) ;
  assign n18322 = ( n18073 & ~n18063 ) | ( n18073 & n18321 ) | ( ~n18063 & n18321 ) ;
  assign n18323 = ( n17834 & ~n17831 ) | ( n17834 & n18055 ) | ( ~n17831 & n18055 ) ;
  assign n18324 = ( n17831 & ~n18055 ) | ( n17831 & n17834 ) | ( ~n18055 & n17834 ) ;
  assign n18325 = ( n18323 & ~n17834 ) | ( n18323 & n18324 ) | ( ~n17834 & n18324 ) ;
  assign n18326 = ( n17647 & ~n17744 ) | ( n17647 & n17754 ) | ( ~n17744 & n17754 ) ;
  assign n18327 = n6983 &  n7097 ;
  assign n18328 = ( n14800 & ~n18327 ) | ( n14800 & 1'b0 ) | ( ~n18327 & 1'b0 ) ;
  assign n18329 = ~n6530 & n14807 ;
  assign n18330 = n18328 | n18329 ;
  assign n18331 = ( n6532 & n15692 ) | ( n6532 & n18330 ) | ( n15692 & n18330 ) ;
  assign n18332 = ( n15692 & ~n18331 ) | ( n15692 & 1'b0 ) | ( ~n18331 & 1'b0 ) ;
  assign n18333 = ( n18330 & ~x14 ) | ( n18330 & n18332 ) | ( ~x14 & n18332 ) ;
  assign n18334 = ( x14 & ~n18330 ) | ( x14 & n18332 ) | ( ~n18330 & n18332 ) ;
  assign n18335 = ( n18333 & ~n18332 ) | ( n18333 & n18334 ) | ( ~n18332 & n18334 ) ;
  assign n18336 = ( n17643 & ~n17731 ) | ( n17643 & n17741 ) | ( ~n17731 & n17741 ) ;
  assign n18337 = ( n17651 & ~n17705 ) | ( n17651 & n17715 ) | ( ~n17705 & n17715 ) ;
  assign n18338 = ( n17692 & ~n17691 ) | ( n17692 & n17702 ) | ( ~n17691 & n17702 ) ;
  assign n18342 = ~n4430 & n11101 ;
  assign n18339 = ~n523 & n11107 ;
  assign n18340 = n3939 | n11104 ;
  assign n18341 = ~n18339 & n18340 ;
  assign n18343 = ( n4430 & n18342 ) | ( n4430 & n18341 ) | ( n18342 & n18341 ) ;
  assign n18344 = n601 | n12650 ;
  assign n18345 = n18343 &  n18344 ;
  assign n18346 = x29 &  n18345 ;
  assign n18347 = x29 | n18345 ;
  assign n18348 = ~n18346 & n18347 ;
  assign n18349 = ( n17673 & ~n17666 ) | ( n17673 & n17675 ) | ( ~n17666 & n17675 ) ;
  assign n18363 = ( n1633 & ~n4074 ) | ( n1633 & n14640 ) | ( ~n4074 & n14640 ) ;
  assign n18364 = ~n1633 & n18363 ;
  assign n18350 = n1359 | n2064 ;
  assign n18351 = ( n1343 & ~n18350 ) | ( n1343 & n3792 ) | ( ~n18350 & n3792 ) ;
  assign n18352 = ( n423 & ~n3792 ) | ( n423 & n18351 ) | ( ~n3792 & n18351 ) ;
  assign n18353 = ~n423 & n18352 ;
  assign n18354 = ( n1679 & ~n1883 ) | ( n1679 & n18353 ) | ( ~n1883 & n18353 ) ;
  assign n18355 = ~n1679 & n18354 ;
  assign n18356 = ( n1807 & ~n1001 ) | ( n1807 & n18355 ) | ( ~n1001 & n18355 ) ;
  assign n18357 = ~n1807 & n18356 ;
  assign n18358 = ( n673 & ~n260 ) | ( n673 & n18357 ) | ( ~n260 & n18357 ) ;
  assign n18359 = ~n673 & n18358 ;
  assign n18360 = ( n276 & ~n187 ) | ( n276 & n18359 ) | ( ~n187 & n18359 ) ;
  assign n18361 = ~n276 & n18360 ;
  assign n18362 = ~n666 & n18361 ;
  assign n18365 = ( n3113 & ~n18364 ) | ( n3113 & n18362 ) | ( ~n18364 & n18362 ) ;
  assign n18366 = ( n163 & ~n18365 ) | ( n163 & n18362 ) | ( ~n18365 & n18362 ) ;
  assign n18367 = ~n163 & n18366 ;
  assign n18368 = ( n1581 & ~n947 ) | ( n1581 & n18367 ) | ( ~n947 & n18367 ) ;
  assign n18369 = ~n1581 & n18368 ;
  assign n18370 = ( n18369 & ~n383 ) | ( n18369 & n2936 ) | ( ~n383 & n2936 ) ;
  assign n18371 = ( n18370 & ~n2936 ) | ( n18370 & 1'b0 ) | ( ~n2936 & 1'b0 ) ;
  assign n18372 = ( n352 & ~n18371 ) | ( n352 & n813 ) | ( ~n18371 & n813 ) ;
  assign n18373 = ( n813 & ~n18372 ) | ( n813 & 1'b0 ) | ( ~n18372 & 1'b0 ) ;
  assign n18374 = ( n909 & ~n718 ) | ( n909 & n18373 ) | ( ~n718 & n18373 ) ;
  assign n18375 = ~n909 & n18374 ;
  assign n18376 = ( n338 & ~n18375 ) | ( n338 & n524 ) | ( ~n18375 & n524 ) ;
  assign n18377 = ( n524 & ~n18376 ) | ( n524 & 1'b0 ) | ( ~n18376 & 1'b0 ) ;
  assign n18378 = ( n169 & ~n340 ) | ( n169 & n18377 ) | ( ~n340 & n18377 ) ;
  assign n18379 = ~n169 & n18378 ;
  assign n18380 = ~n617 & n18379 ;
  assign n18381 = ~n3644 & n12352 ;
  assign n18382 = n3652 &  n11116 ;
  assign n18383 = ( n3657 & ~n11113 ) | ( n3657 & 1'b0 ) | ( ~n11113 & 1'b0 ) ;
  assign n18384 = n18382 | n18383 ;
  assign n18385 = ~n3653 & n11110 ;
  assign n18386 = ( n3653 & ~n18384 ) | ( n3653 & n18385 ) | ( ~n18384 & n18385 ) ;
  assign n18387 = ~n18381 & n18386 ;
  assign n18388 = ( n18380 & ~n17666 ) | ( n18380 & n18387 ) | ( ~n17666 & n18387 ) ;
  assign n18389 = ( n17666 & ~n18380 ) | ( n17666 & n18387 ) | ( ~n18380 & n18387 ) ;
  assign n18390 = ( n18388 & ~n18387 ) | ( n18388 & n18389 ) | ( ~n18387 & n18389 ) ;
  assign n18391 = ~x29 & n17688 ;
  assign n18392 = ( x29 & ~n17688 ) | ( x29 & n17680 ) | ( ~n17688 & n17680 ) ;
  assign n18393 = ( n18391 & ~n17679 ) | ( n18391 & n18392 ) | ( ~n17679 & n18392 ) ;
  assign n18394 = ( n18349 & n18390 ) | ( n18349 & n18393 ) | ( n18390 & n18393 ) ;
  assign n18395 = ( n18390 & ~n18349 ) | ( n18390 & n18393 ) | ( ~n18349 & n18393 ) ;
  assign n18396 = ( n18349 & ~n18394 ) | ( n18349 & n18395 ) | ( ~n18394 & n18395 ) ;
  assign n18400 = ~n4962 & n11093 ;
  assign n18397 = n4482 | n11098 ;
  assign n18398 = n4495 | n11095 ;
  assign n18399 = n18397 &  n18398 ;
  assign n18401 = ( n4962 & n18400 ) | ( n4962 & n18399 ) | ( n18400 & n18399 ) ;
  assign n18402 = n4478 | n12997 ;
  assign n18403 = n18401 &  n18402 ;
  assign n18404 = x26 &  n18403 ;
  assign n18405 = x26 | n18403 ;
  assign n18406 = ~n18404 & n18405 ;
  assign n18407 = ( n18348 & ~n18396 ) | ( n18348 & n18406 ) | ( ~n18396 & n18406 ) ;
  assign n18408 = ( n18348 & ~n18406 ) | ( n18348 & n18396 ) | ( ~n18406 & n18396 ) ;
  assign n18409 = ( n18407 & ~n18348 ) | ( n18407 & n18408 ) | ( ~n18348 & n18408 ) ;
  assign n18413 = ~n5135 & n11085 ;
  assign n18410 = n5010 | n11091 ;
  assign n18411 = n5067 | n11081 ;
  assign n18412 = n18410 &  n18411 ;
  assign n18414 = ( n5135 & n18413 ) | ( n5135 & n18412 ) | ( n18413 & n18412 ) ;
  assign n18415 = n5012 | n13377 ;
  assign n18416 = n18414 &  n18415 ;
  assign n18417 = x23 &  n18416 ;
  assign n18418 = x23 | n18416 ;
  assign n18419 = ~n18417 & n18418 ;
  assign n18420 = ( n18338 & n18409 ) | ( n18338 & n18419 ) | ( n18409 & n18419 ) ;
  assign n18421 = ( n18409 & ~n18338 ) | ( n18409 & n18419 ) | ( ~n18338 & n18419 ) ;
  assign n18422 = ( n18338 & ~n18420 ) | ( n18338 & n18421 ) | ( ~n18420 & n18421 ) ;
  assign n18426 = ~n5837 & n14071 ;
  assign n18423 = ( n5339 & ~n11078 ) | ( n5339 & 1'b0 ) | ( ~n11078 & 1'b0 ) ;
  assign n18424 = n5761 | n13836 ;
  assign n18425 = ~n18423 & n18424 ;
  assign n18427 = ( n5837 & n18426 ) | ( n5837 & n18425 ) | ( n18426 & n18425 ) ;
  assign n18428 = n5341 | n14079 ;
  assign n18429 = n18427 &  n18428 ;
  assign n18430 = x20 &  n18429 ;
  assign n18431 = x20 | n18429 ;
  assign n18432 = ~n18430 & n18431 ;
  assign n18433 = ( n18337 & n18422 ) | ( n18337 & n18432 ) | ( n18422 & n18432 ) ;
  assign n18434 = ( n18422 & ~n18337 ) | ( n18422 & n18432 ) | ( ~n18337 & n18432 ) ;
  assign n18435 = ( n18337 & ~n18433 ) | ( n18337 & n18434 ) | ( ~n18433 & n18434 ) ;
  assign n18436 = ( n17639 & ~n17718 ) | ( n17639 & n17728 ) | ( ~n17718 & n17728 ) ;
  assign n18437 = ( n18435 & ~n18436 ) | ( n18435 & 1'b0 ) | ( ~n18436 & 1'b0 ) ;
  assign n18438 = ~n18435 & n18436 ;
  assign n18439 = n18437 | n18438 ;
  assign n18443 = ~n6395 & n14803 ;
  assign n18440 = n5970 | n14355 ;
  assign n18441 = ~n6170 & n14553 ;
  assign n18442 = ( n18440 & ~n18441 ) | ( n18440 & 1'b0 ) | ( ~n18441 & 1'b0 ) ;
  assign n18444 = ( n6395 & n18443 ) | ( n6395 & n18442 ) | ( n18443 & n18442 ) ;
  assign n18445 = ~n5972 & n15310 ;
  assign n18446 = ( n18444 & ~n18445 ) | ( n18444 & 1'b0 ) | ( ~n18445 & 1'b0 ) ;
  assign n18447 = ( x17 & ~n18439 ) | ( x17 & n18446 ) | ( ~n18439 & n18446 ) ;
  assign n18448 = ( n18439 & ~x17 ) | ( n18439 & n18446 ) | ( ~x17 & n18446 ) ;
  assign n18449 = ( n18447 & ~n18446 ) | ( n18447 & n18448 ) | ( ~n18446 & n18448 ) ;
  assign n18450 = ( n18335 & n18336 ) | ( n18335 & n18449 ) | ( n18336 & n18449 ) ;
  assign n18451 = ( n18336 & ~n18335 ) | ( n18336 & n18449 ) | ( ~n18335 & n18449 ) ;
  assign n18452 = ( n18335 & ~n18450 ) | ( n18335 & n18451 ) | ( ~n18450 & n18451 ) ;
  assign n18453 = ( n17757 & ~n17650 ) | ( n17757 & n17780 ) | ( ~n17650 & n17780 ) ;
  assign n18454 = ( n18452 & ~n18326 ) | ( n18452 & n18453 ) | ( ~n18326 & n18453 ) ;
  assign n18455 = ( n18326 & n18452 ) | ( n18326 & n18453 ) | ( n18452 & n18453 ) ;
  assign n18456 = ( ~n18326 & ~n18454 ) | ( ~n18326 & n18455 ) | ( ~n18454 & n18455 ) ;
  assign n18460 = ~n7097 & n18456 ;
  assign n18457 = n6530 | n17791 ;
  assign n18458 = n6983 | n17783 ;
  assign n18459 = n18457 &  n18458 ;
  assign n18461 = ( n7097 & n18460 ) | ( n7097 & n18459 ) | ( n18460 & n18459 ) ;
  assign n18463 = ( n17783 & n17798 ) | ( n17783 & n18456 ) | ( n17798 & n18456 ) ;
  assign n18462 = ( n17798 & ~n17783 ) | ( n17798 & n18456 ) | ( ~n17783 & n18456 ) ;
  assign n18464 = ( n17783 & ~n18463 ) | ( n17783 & n18462 ) | ( ~n18463 & n18462 ) ;
  assign n18465 = ( n6532 & ~n18464 ) | ( n6532 & n18461 ) | ( ~n18464 & n18461 ) ;
  assign n18466 = ~n6532 & n18465 ;
  assign n18467 = ( x14 & ~n18461 ) | ( x14 & n18466 ) | ( ~n18461 & n18466 ) ;
  assign n18468 = ( n18461 & ~x14 ) | ( n18461 & n18466 ) | ( ~x14 & n18466 ) ;
  assign n18469 = ( n18467 & ~n18466 ) | ( n18467 & n18468 ) | ( ~n18466 & n18468 ) ;
  assign n18470 = ( n18322 & n18325 ) | ( n18322 & n18469 ) | ( n18325 & n18469 ) ;
  assign n18471 = ( n17819 & ~n17816 ) | ( n17819 & n18056 ) | ( ~n17816 & n18056 ) ;
  assign n18472 = ( n17816 & ~n18056 ) | ( n17816 & n17819 ) | ( ~n18056 & n17819 ) ;
  assign n18473 = ( n18471 & ~n17819 ) | ( n18471 & n18472 ) | ( ~n17819 & n18472 ) ;
  assign n18477 = n14807 | n6395 ;
  assign n18474 = ~n5970 & n14553 ;
  assign n18475 = n6170 | n14803 ;
  assign n18476 = ~n18474 & n18475 ;
  assign n18478 = ( n6395 & ~n18477 ) | ( n6395 & n18476 ) | ( ~n18477 & n18476 ) ;
  assign n18479 = ~n5972 & n15294 ;
  assign n18480 = ( n18478 & ~n18479 ) | ( n18478 & 1'b0 ) | ( ~n18479 & 1'b0 ) ;
  assign n18481 = x17 &  n18480 ;
  assign n18482 = x17 | n18480 ;
  assign n18483 = ~n18481 & n18482 ;
  assign n18484 = ( x17 & ~n18446 ) | ( x17 & 1'b0 ) | ( ~n18446 & 1'b0 ) ;
  assign n18485 = ( n18438 & ~x17 ) | ( n18438 & n18446 ) | ( ~x17 & n18446 ) ;
  assign n18486 = ( n18484 & ~n18437 ) | ( n18484 & n18485 ) | ( ~n18437 & n18485 ) ;
  assign n18487 = ( n5339 & ~n13836 ) | ( n5339 & 1'b0 ) | ( ~n13836 & 1'b0 ) ;
  assign n18488 = n5761 | n14071 ;
  assign n18489 = ~n18487 & n18488 ;
  assign n18490 = ~n5837 & n14355 ;
  assign n18491 = ( n5837 & n18489 ) | ( n5837 & n18490 ) | ( n18489 & n18490 ) ;
  assign n18492 = n5341 | n14363 ;
  assign n18493 = n18491 &  n18492 ;
  assign n18494 = x20 &  n18493 ;
  assign n18495 = x20 | n18493 ;
  assign n18496 = ~n18494 & n18495 ;
  assign n18500 = ~n5135 & n11078 ;
  assign n18497 = n5010 | n11081 ;
  assign n18498 = n5067 | n11085 ;
  assign n18499 = n18497 &  n18498 ;
  assign n18501 = ( n5135 & n18500 ) | ( n5135 & n18499 ) | ( n18500 & n18499 ) ;
  assign n18502 = n5012 | n11206 ;
  assign n18503 = n18501 &  n18502 ;
  assign n18504 = x23 &  n18503 ;
  assign n18505 = x23 | n18503 ;
  assign n18506 = ~n18504 & n18505 ;
  assign n18520 = ~n4430 & n11098 ;
  assign n18517 = n523 | n11104 ;
  assign n18518 = n3939 | n11101 ;
  assign n18519 = n18517 &  n18518 ;
  assign n18521 = ( n4430 & n18520 ) | ( n4430 & n18519 ) | ( n18520 & n18519 ) ;
  assign n18522 = n601 | n11218 ;
  assign n18523 = n18521 &  n18522 ;
  assign n18524 = x29 &  n18523 ;
  assign n18525 = x29 | n18523 ;
  assign n18526 = ~n18524 & n18525 ;
  assign n18527 = ~n3644 & n12340 ;
  assign n18531 = n11107 | n3653 ;
  assign n18528 = ( n3652 & ~n11113 ) | ( n3652 & 1'b0 ) | ( ~n11113 & 1'b0 ) ;
  assign n18529 = ( n3657 & ~n11110 ) | ( n3657 & 1'b0 ) | ( ~n11110 & 1'b0 ) ;
  assign n18530 = n18528 | n18529 ;
  assign n18532 = ( n18531 & ~n3653 ) | ( n18531 & n18530 ) | ( ~n3653 & n18530 ) ;
  assign n18533 = n18527 | n18532 ;
  assign n18534 = ( n6522 & ~n6525 ) | ( n6522 & n6528 ) | ( ~n6525 & n6528 ) ;
  assign n18535 = n6525 | n18534 ;
  assign n18536 = n14800 &  n18535 ;
  assign n18537 = n238 | n1580 ;
  assign n18538 = ( n405 & n18537 ) | ( n405 & n786 ) | ( n18537 & n786 ) ;
  assign n18539 = ( n786 & ~n18538 ) | ( n786 & 1'b0 ) | ( ~n18538 & 1'b0 ) ;
  assign n18540 = ( n225 & ~n571 ) | ( n225 & n18539 ) | ( ~n571 & n18539 ) ;
  assign n18541 = ~n225 & n18540 ;
  assign n18542 = ( n154 & ~n2279 ) | ( n154 & n15927 ) | ( ~n2279 & n15927 ) ;
  assign n18543 = n2279 | n18542 ;
  assign n18544 = ( n4253 & ~n1584 ) | ( n4253 & n18543 ) | ( ~n1584 & n18543 ) ;
  assign n18545 = n1584 | n18544 ;
  assign n18546 = ( n2686 & ~n18541 ) | ( n2686 & n18545 ) | ( ~n18541 & n18545 ) ;
  assign n18547 = ( n2686 & ~n18546 ) | ( n2686 & 1'b0 ) | ( ~n18546 & 1'b0 ) ;
  assign n18548 = ( n1807 & ~n6627 ) | ( n1807 & n18547 ) | ( ~n6627 & n18547 ) ;
  assign n18549 = ~n1807 & n18548 ;
  assign n18550 = ( n234 & ~n2713 ) | ( n234 & n18549 ) | ( ~n2713 & n18549 ) ;
  assign n18551 = ~n234 & n18550 ;
  assign n18552 = ( n453 & ~n494 ) | ( n453 & n18551 ) | ( ~n494 & n18551 ) ;
  assign n18553 = ~n453 & n18552 ;
  assign n18554 = ( n267 & ~n909 ) | ( n267 & n18553 ) | ( ~n909 & n18553 ) ;
  assign n18555 = ~n267 & n18554 ;
  assign n18556 = ( n93 & ~n285 ) | ( n93 & n18555 ) | ( ~n285 & n18555 ) ;
  assign n18557 = ~n93 & n18556 ;
  assign n18558 = n17666 | n18557 ;
  assign n18559 = n17666 &  n18557 ;
  assign n18560 = ( n18558 & ~n18559 ) | ( n18558 & 1'b0 ) | ( ~n18559 & 1'b0 ) ;
  assign n18561 = ( n18536 & ~x14 ) | ( n18536 & n18560 ) | ( ~x14 & n18560 ) ;
  assign n18562 = ( x14 & ~n18560 ) | ( x14 & n18536 ) | ( ~n18560 & n18536 ) ;
  assign n18563 = ( n18561 & ~n18536 ) | ( n18561 & n18562 ) | ( ~n18536 & n18562 ) ;
  assign n18565 = ( n18388 & n18533 ) | ( n18388 & n18563 ) | ( n18533 & n18563 ) ;
  assign n18564 = ( n18533 & ~n18388 ) | ( n18533 & n18563 ) | ( ~n18388 & n18563 ) ;
  assign n18566 = ( n18388 & ~n18565 ) | ( n18388 & n18564 ) | ( ~n18565 & n18564 ) ;
  assign n18567 = ( n18349 & ~n18390 ) | ( n18349 & n18393 ) | ( ~n18390 & n18393 ) ;
  assign n18568 = ( n18526 & n18566 ) | ( n18526 & n18567 ) | ( n18566 & n18567 ) ;
  assign n18569 = ( n18566 & ~n18526 ) | ( n18566 & n18567 ) | ( ~n18526 & n18567 ) ;
  assign n18570 = ( n18526 & ~n18568 ) | ( n18526 & n18569 ) | ( ~n18568 & n18569 ) ;
  assign n18510 = ~n4962 & n11091 ;
  assign n18507 = n4482 | n11095 ;
  assign n18508 = n4495 | n11093 ;
  assign n18509 = n18507 &  n18508 ;
  assign n18511 = ( n4962 & n18510 ) | ( n4962 & n18509 ) | ( n18510 & n18509 ) ;
  assign n18512 = n4478 | n12984 ;
  assign n18513 = n18511 &  n18512 ;
  assign n18514 = x26 &  n18513 ;
  assign n18515 = x26 | n18513 ;
  assign n18516 = ~n18514 & n18515 ;
  assign n18571 = ( n18407 & ~n18570 ) | ( n18407 & n18516 ) | ( ~n18570 & n18516 ) ;
  assign n18572 = ( n18516 & ~n18407 ) | ( n18516 & n18570 ) | ( ~n18407 & n18570 ) ;
  assign n18573 = ( n18571 & ~n18516 ) | ( n18571 & n18572 ) | ( ~n18516 & n18572 ) ;
  assign n18574 = ( n18338 & ~n18409 ) | ( n18338 & n18419 ) | ( ~n18409 & n18419 ) ;
  assign n18575 = ( n18506 & ~n18573 ) | ( n18506 & n18574 ) | ( ~n18573 & n18574 ) ;
  assign n18576 = ( n18506 & ~n18574 ) | ( n18506 & n18573 ) | ( ~n18574 & n18573 ) ;
  assign n18577 = ( n18575 & ~n18506 ) | ( n18575 & n18576 ) | ( ~n18506 & n18576 ) ;
  assign n18578 = ( n18337 & ~n18422 ) | ( n18337 & n18432 ) | ( ~n18422 & n18432 ) ;
  assign n18579 = ( n18496 & ~n18577 ) | ( n18496 & n18578 ) | ( ~n18577 & n18578 ) ;
  assign n18580 = ( n18496 & ~n18578 ) | ( n18496 & n18577 ) | ( ~n18578 & n18577 ) ;
  assign n18581 = ( n18579 & ~n18496 ) | ( n18579 & n18580 ) | ( ~n18496 & n18580 ) ;
  assign n18582 = ( n18483 & ~n18486 ) | ( n18483 & n18581 ) | ( ~n18486 & n18581 ) ;
  assign n18583 = ( n18483 & ~n18581 ) | ( n18483 & n18486 ) | ( ~n18581 & n18486 ) ;
  assign n18584 = ( n18582 & ~n18483 ) | ( n18582 & n18583 ) | ( ~n18483 & n18583 ) ;
  assign n18585 = ( n18335 & ~n18336 ) | ( n18335 & n18449 ) | ( ~n18336 & n18449 ) ;
  assign n18586 = ( n18326 & ~n18453 ) | ( n18326 & n18452 ) | ( ~n18453 & n18452 ) ;
  assign n18587 = ( n18584 & n18585 ) | ( n18584 & n18586 ) | ( n18585 & n18586 ) ;
  assign n18588 = ( n18585 & ~n18584 ) | ( n18585 & n18586 ) | ( ~n18584 & n18586 ) ;
  assign n18589 = ( n18584 & ~n18587 ) | ( n18584 & n18588 ) | ( ~n18587 & n18588 ) ;
  assign n18596 = ( n18456 & n18463 ) | ( n18456 & n18589 ) | ( n18463 & n18589 ) ;
  assign n18595 = ( n18463 & ~n18456 ) | ( n18463 & n18589 ) | ( ~n18456 & n18589 ) ;
  assign n18597 = ( n18456 & ~n18596 ) | ( n18456 & n18595 ) | ( ~n18596 & n18595 ) ;
  assign n18593 = ~n7097 & n18589 ;
  assign n18590 = n6530 | n17783 ;
  assign n18591 = n6983 | n18456 ;
  assign n18592 = n18590 &  n18591 ;
  assign n18594 = ( n7097 & n18593 ) | ( n7097 & n18592 ) | ( n18593 & n18592 ) ;
  assign n18598 = ( n18594 & ~n6532 ) | ( n18594 & n18597 ) | ( ~n6532 & n18597 ) ;
  assign n18599 = ~n18597 & n18598 ;
  assign n18601 = ( x14 & n18594 ) | ( x14 & n18599 ) | ( n18594 & n18599 ) ;
  assign n18600 = ( x14 & ~n18599 ) | ( x14 & n18594 ) | ( ~n18599 & n18594 ) ;
  assign n18602 = ( n18599 & ~n18601 ) | ( n18599 & n18600 ) | ( ~n18601 & n18600 ) ;
  assign n18603 = ( n18470 & n18473 ) | ( n18470 & n18602 ) | ( n18473 & n18602 ) ;
  assign n18709 = ( n18584 & ~n18586 ) | ( n18584 & n18585 ) | ( ~n18586 & n18585 ) ;
  assign n18604 = ( n18388 & ~n18533 ) | ( n18388 & n18563 ) | ( ~n18533 & n18563 ) ;
  assign n18650 = ~x29 & n18604 ;
  assign n18651 = x29 | n18604 ;
  assign n18652 = ( n18650 & ~n18604 ) | ( n18650 & n18651 ) | ( ~n18604 & n18651 ) ;
  assign n18605 = n717 | n2192 ;
  assign n18606 = ( n1385 & ~n1494 ) | ( n1385 & n18605 ) | ( ~n1494 & n18605 ) ;
  assign n18607 = n1494 | n18606 ;
  assign n18608 = ( n345 & ~n359 ) | ( n345 & n18607 ) | ( ~n359 & n18607 ) ;
  assign n18609 = n359 | n18608 ;
  assign n18610 = ( n18609 & ~n349 ) | ( n18609 & n800 ) | ( ~n349 & n800 ) ;
  assign n18611 = n349 | n18610 ;
  assign n18612 = ( n340 & ~n373 ) | ( n340 & n18611 ) | ( ~n373 & n18611 ) ;
  assign n18613 = n373 | n18612 ;
  assign n18614 = n459 | n18613 ;
  assign n18615 = ( n316 & ~n2242 ) | ( n316 & n2850 ) | ( ~n2242 & n2850 ) ;
  assign n18616 = n2242 | n18615 ;
  assign n18617 = ( n3516 & ~n3788 ) | ( n3516 & n18616 ) | ( ~n3788 & n18616 ) ;
  assign n18618 = ( n3516 & ~n18617 ) | ( n3516 & 1'b0 ) | ( ~n18617 & 1'b0 ) ;
  assign n18619 = ( n2484 & ~n18614 ) | ( n2484 & n18618 ) | ( ~n18614 & n18618 ) ;
  assign n18620 = ~n2484 & n18619 ;
  assign n18621 = ( n842 & ~n3281 ) | ( n842 & n18620 ) | ( ~n3281 & n18620 ) ;
  assign n18622 = ~n842 & n18621 ;
  assign n18623 = ( n126 & n344 ) | ( n126 & n18622 ) | ( n344 & n18622 ) ;
  assign n18624 = ~n126 & n18623 ;
  assign n18625 = ( n429 & ~n674 ) | ( n429 & n18624 ) | ( ~n674 & n18624 ) ;
  assign n18626 = ~n429 & n18625 ;
  assign n18627 = ( n529 & ~n911 ) | ( n529 & n18626 ) | ( ~n911 & n18626 ) ;
  assign n18628 = ~n529 & n18627 ;
  assign n18629 = ( n478 & ~n137 ) | ( n478 & n18628 ) | ( ~n137 & n18628 ) ;
  assign n18630 = ~n478 & n18629 ;
  assign n18638 = ~x14 & n18536 ;
  assign n18639 = ( n18558 & ~n18561 ) | ( n18558 & n18638 ) | ( ~n18561 & n18638 ) ;
  assign n18636 = n12662 | n3644 ;
  assign n18631 = n3653 | n11104 ;
  assign n18632 = n3657 &  n11107 ;
  assign n18633 = ( n3652 & ~n11110 ) | ( n3652 & 1'b0 ) | ( ~n11110 & 1'b0 ) ;
  assign n18634 = n18632 | n18633 ;
  assign n18635 = ( n18631 & ~n18634 ) | ( n18631 & 1'b0 ) | ( ~n18634 & 1'b0 ) ;
  assign n18637 = ( n3644 & ~n18636 ) | ( n3644 & n18635 ) | ( ~n18636 & n18635 ) ;
  assign n18640 = ( n18630 & ~n18639 ) | ( n18630 & n18637 ) | ( ~n18639 & n18637 ) ;
  assign n18641 = ( n18630 & ~n18637 ) | ( n18630 & n18639 ) | ( ~n18637 & n18639 ) ;
  assign n18642 = ( n18640 & ~n18630 ) | ( n18640 & n18641 ) | ( ~n18630 & n18641 ) ;
  assign n18648 = ~n601 & n13014 ;
  assign n18646 = ~n4430 & n11095 ;
  assign n18643 = n523 | n11101 ;
  assign n18644 = n3939 | n11098 ;
  assign n18645 = n18643 &  n18644 ;
  assign n18647 = ( n4430 & n18646 ) | ( n4430 & n18645 ) | ( n18646 & n18645 ) ;
  assign n18649 = ( n601 & n18648 ) | ( n601 & n18647 ) | ( n18648 & n18647 ) ;
  assign n18653 = ( n18642 & n18649 ) | ( n18642 & n18652 ) | ( n18649 & n18652 ) ;
  assign n18654 = ( n18642 & ~n18652 ) | ( n18642 & n18649 ) | ( ~n18652 & n18649 ) ;
  assign n18655 = ( n18652 & ~n18653 ) | ( n18652 & n18654 ) | ( ~n18653 & n18654 ) ;
  assign n18656 = ( n18526 & ~n18566 ) | ( n18526 & n18567 ) | ( ~n18566 & n18567 ) ;
  assign n18660 = ~n4962 & n11081 ;
  assign n18657 = n4482 | n11093 ;
  assign n18658 = n4495 | n11091 ;
  assign n18659 = n18657 &  n18658 ;
  assign n18661 = ( n4962 & n18660 ) | ( n4962 & n18659 ) | ( n18660 & n18659 ) ;
  assign n18662 = n4478 | n13775 ;
  assign n18663 = n18661 &  n18662 ;
  assign n18664 = x26 &  n18663 ;
  assign n18665 = x26 | n18663 ;
  assign n18666 = ~n18664 & n18665 ;
  assign n18667 = ( n18655 & ~n18656 ) | ( n18655 & n18666 ) | ( ~n18656 & n18666 ) ;
  assign n18668 = ( n18655 & ~n18666 ) | ( n18655 & n18656 ) | ( ~n18666 & n18656 ) ;
  assign n18669 = ( n18667 & ~n18655 ) | ( n18667 & n18668 ) | ( ~n18655 & n18668 ) ;
  assign n18673 = ~n5135 & n13836 ;
  assign n18670 = n5010 | n11085 ;
  assign n18671 = n5067 | n11078 ;
  assign n18672 = n18670 &  n18671 ;
  assign n18674 = ( n5135 & n18673 ) | ( n5135 & n18672 ) | ( n18673 & n18672 ) ;
  assign n18675 = n5012 | n13844 ;
  assign n18676 = n18674 &  n18675 ;
  assign n18677 = x23 &  n18676 ;
  assign n18678 = x23 | n18676 ;
  assign n18679 = ~n18677 & n18678 ;
  assign n18680 = ( n18571 & n18669 ) | ( n18571 & n18679 ) | ( n18669 & n18679 ) ;
  assign n18681 = ( n18669 & ~n18571 ) | ( n18669 & n18679 ) | ( ~n18571 & n18679 ) ;
  assign n18682 = ( n18571 & ~n18680 ) | ( n18571 & n18681 ) | ( ~n18680 & n18681 ) ;
  assign n18686 = n14553 | n5837 ;
  assign n18683 = ( n5339 & ~n14071 ) | ( n5339 & 1'b0 ) | ( ~n14071 & 1'b0 ) ;
  assign n18684 = n5761 | n14355 ;
  assign n18685 = ~n18683 & n18684 ;
  assign n18687 = ( n5837 & ~n18686 ) | ( n5837 & n18685 ) | ( ~n18686 & n18685 ) ;
  assign n18688 = ~n5341 & n14562 ;
  assign n18689 = ( n18687 & ~n18688 ) | ( n18687 & 1'b0 ) | ( ~n18688 & 1'b0 ) ;
  assign n18690 = x20 &  n18689 ;
  assign n18691 = x20 | n18689 ;
  assign n18692 = ~n18690 & n18691 ;
  assign n18693 = ( n18575 & n18682 ) | ( n18575 & n18692 ) | ( n18682 & n18692 ) ;
  assign n18694 = ( n18682 & ~n18575 ) | ( n18682 & n18692 ) | ( ~n18575 & n18692 ) ;
  assign n18695 = ( n18575 & ~n18693 ) | ( n18575 & n18694 ) | ( ~n18693 & n18694 ) ;
  assign n18699 = n14800 | n6395 ;
  assign n18696 = n5970 | n14803 ;
  assign n18697 = ~n6170 & n14807 ;
  assign n18698 = ( n18696 & ~n18697 ) | ( n18696 & 1'b0 ) | ( ~n18697 & 1'b0 ) ;
  assign n18700 = ( n6395 & ~n18699 ) | ( n6395 & n18698 ) | ( ~n18699 & n18698 ) ;
  assign n18701 = n5972 | n14816 ;
  assign n18702 = n18700 &  n18701 ;
  assign n18703 = x17 &  n18702 ;
  assign n18704 = x17 | n18702 ;
  assign n18705 = ~n18703 & n18704 ;
  assign n18706 = ( n18579 & n18695 ) | ( n18579 & n18705 ) | ( n18695 & n18705 ) ;
  assign n18707 = ( n18695 & ~n18579 ) | ( n18695 & n18705 ) | ( ~n18579 & n18705 ) ;
  assign n18708 = ( n18579 & ~n18706 ) | ( n18579 & n18707 ) | ( ~n18706 & n18707 ) ;
  assign n18710 = ( n18583 & ~n18709 ) | ( n18583 & n18708 ) | ( ~n18709 & n18708 ) ;
  assign n18711 = ( n18583 & ~n18708 ) | ( n18583 & n18709 ) | ( ~n18708 & n18709 ) ;
  assign n18712 = ( ~n18583 & n18710 ) | ( ~n18583 & n18711 ) | ( n18710 & n18711 ) ;
  assign n18719 = ( n18589 & n18596 ) | ( n18589 & n18712 ) | ( n18596 & n18712 ) ;
  assign n18718 = ( n18596 & ~n18589 ) | ( n18596 & n18712 ) | ( ~n18589 & n18712 ) ;
  assign n18720 = ( n18589 & ~n18719 ) | ( n18589 & n18718 ) | ( ~n18719 & n18718 ) ;
  assign n18716 = ~n7097 & n18712 ;
  assign n18713 = n6530 | n18456 ;
  assign n18714 = n6983 | n18589 ;
  assign n18715 = n18713 &  n18714 ;
  assign n18717 = ( n7097 & n18716 ) | ( n7097 & n18715 ) | ( n18716 & n18715 ) ;
  assign n18721 = ( n18717 & ~n6532 ) | ( n18717 & n18720 ) | ( ~n6532 & n18720 ) ;
  assign n18722 = ~n18720 & n18721 ;
  assign n18724 = ( x14 & n18717 ) | ( x14 & n18722 ) | ( n18717 & n18722 ) ;
  assign n18723 = ( x14 & ~n18722 ) | ( x14 & n18717 ) | ( ~n18722 & n18717 ) ;
  assign n18725 = ( n18722 & ~n18724 ) | ( n18722 & n18723 ) | ( ~n18724 & n18723 ) ;
  assign n18726 = ( n18060 & ~n18603 ) | ( n18060 & n18725 ) | ( ~n18603 & n18725 ) ;
  assign n18727 = ( n18060 & ~n18725 ) | ( n18060 & n18603 ) | ( ~n18725 & n18603 ) ;
  assign n18728 = ( n18726 & ~n18060 ) | ( n18726 & n18727 ) | ( ~n18060 & n18727 ) ;
  assign n18817 = n5837 | n14807 ;
  assign n18814 = n5339 &  n14553 ;
  assign n18815 = n5761 | n14803 ;
  assign n18816 = ~n18814 & n18815 ;
  assign n18818 = ( n5837 & ~n18817 ) | ( n5837 & n18816 ) | ( ~n18817 & n18816 ) ;
  assign n18819 = ~n5341 & n15294 ;
  assign n18820 = ( n18818 & ~n18819 ) | ( n18818 & 1'b0 ) | ( ~n18819 & 1'b0 ) ;
  assign n18821 = x20 &  n18820 ;
  assign n18822 = x20 | n18820 ;
  assign n18823 = ~n18821 & n18822 ;
  assign n18802 = ( n18571 & ~n18669 ) | ( n18571 & n18679 ) | ( ~n18669 & n18679 ) ;
  assign n18729 = ( n18656 & ~n18655 ) | ( n18656 & n18666 ) | ( ~n18655 & n18666 ) ;
  assign n18730 = x29 | n18649 ;
  assign n18731 = x29 &  n18649 ;
  assign n18732 = ( n18730 & ~n18731 ) | ( n18730 & 1'b0 ) | ( ~n18731 & 1'b0 ) ;
  assign n18733 = ( n18604 & ~n18642 ) | ( n18604 & n18732 ) | ( ~n18642 & n18732 ) ;
  assign n18783 = x26 | n18733 ;
  assign n18784 = ~x26 & n18733 ;
  assign n18785 = ( n18783 & ~n18733 ) | ( n18783 & n18784 ) | ( ~n18733 & n18784 ) ;
  assign n18766 = ~n4430 & n11093 ;
  assign n18763 = n523 | n11098 ;
  assign n18764 = n3939 | n11095 ;
  assign n18765 = n18763 &  n18764 ;
  assign n18767 = ( n4430 & n18766 ) | ( n4430 & n18765 ) | ( n18766 & n18765 ) ;
  assign n18768 = ( n12997 & ~n601 ) | ( n12997 & n18767 ) | ( ~n601 & n18767 ) ;
  assign n18769 = ~n12997 & n18768 ;
  assign n18770 = ( x29 & ~n18767 ) | ( x29 & n18769 ) | ( ~n18767 & n18769 ) ;
  assign n18771 = ( n18767 & ~x29 ) | ( n18767 & n18769 ) | ( ~x29 & n18769 ) ;
  assign n18772 = ( n18770 & ~n18769 ) | ( n18770 & n18771 ) | ( ~n18769 & n18771 ) ;
  assign n18734 = n1326 | n2360 ;
  assign n18735 = ( n3157 & n3290 ) | ( n3157 & n18734 ) | ( n3290 & n18734 ) ;
  assign n18736 = ( n3157 & ~n18735 ) | ( n3157 & 1'b0 ) | ( ~n18735 & 1'b0 ) ;
  assign n18737 = ( n204 & n606 ) | ( n204 & n18736 ) | ( n606 & n18736 ) ;
  assign n18738 = ~n606 & n18737 ;
  assign n18739 = ( n3777 & ~n18738 ) | ( n3777 & n5647 ) | ( ~n18738 & n5647 ) ;
  assign n18740 = ( n4304 & ~n5647 ) | ( n4304 & n18739 ) | ( ~n5647 & n18739 ) ;
  assign n18741 = ( n4304 & ~n18740 ) | ( n4304 & 1'b0 ) | ( ~n18740 & 1'b0 ) ;
  assign n18742 = ( n885 & ~n865 ) | ( n885 & n18741 ) | ( ~n865 & n18741 ) ;
  assign n18743 = ~n885 & n18742 ;
  assign n18744 = ( n333 & ~n1426 ) | ( n333 & n18743 ) | ( ~n1426 & n18743 ) ;
  assign n18745 = ~n333 & n18744 ;
  assign n18746 = ( n490 & ~n486 ) | ( n490 & n18745 ) | ( ~n486 & n18745 ) ;
  assign n18747 = ~n490 & n18746 ;
  assign n18748 = ( n169 & ~n549 ) | ( n169 & n18747 ) | ( ~n549 & n18747 ) ;
  assign n18749 = ~n169 & n18748 ;
  assign n18750 = ( n459 & ~n149 ) | ( n459 & n18749 ) | ( ~n149 & n18749 ) ;
  assign n18751 = ~n459 & n18750 ;
  assign n18752 = ( n18637 & ~n18630 ) | ( n18637 & n18639 ) | ( ~n18630 & n18639 ) ;
  assign n18753 = ( n18630 & ~n18751 ) | ( n18630 & n18752 ) | ( ~n18751 & n18752 ) ;
  assign n18754 = ( n18630 & ~n18752 ) | ( n18630 & n18751 ) | ( ~n18752 & n18751 ) ;
  assign n18755 = ( n18753 & ~n18630 ) | ( n18753 & n18754 ) | ( ~n18630 & n18754 ) ;
  assign n18756 = n3644 | n12650 ;
  assign n18757 = n3652 &  n11107 ;
  assign n18758 = ( n3657 & ~n11104 ) | ( n3657 & 1'b0 ) | ( ~n11104 & 1'b0 ) ;
  assign n18759 = n18757 | n18758 ;
  assign n18760 = ~n3653 & n11101 ;
  assign n18761 = ( n3653 & ~n18759 ) | ( n3653 & n18760 ) | ( ~n18759 & n18760 ) ;
  assign n18762 = n18756 &  n18761 ;
  assign n18773 = ( n18755 & n18762 ) | ( n18755 & n18772 ) | ( n18762 & n18772 ) ;
  assign n18774 = ( n18755 & ~n18772 ) | ( n18755 & n18762 ) | ( ~n18772 & n18762 ) ;
  assign n18775 = ( n18772 & ~n18773 ) | ( n18772 & n18774 ) | ( ~n18773 & n18774 ) ;
  assign n18779 = ~n4962 & n11085 ;
  assign n18776 = n4482 | n11091 ;
  assign n18777 = n4495 | n11081 ;
  assign n18778 = n18776 &  n18777 ;
  assign n18780 = ( n4962 & n18779 ) | ( n4962 & n18778 ) | ( n18779 & n18778 ) ;
  assign n18781 = n4478 | n13377 ;
  assign n18782 = n18780 &  n18781 ;
  assign n18787 = ( n18775 & n18782 ) | ( n18775 & n18785 ) | ( n18782 & n18785 ) ;
  assign n18786 = ( n18775 & ~n18785 ) | ( n18775 & n18782 ) | ( ~n18785 & n18782 ) ;
  assign n18788 = ( n18785 & ~n18787 ) | ( n18785 & n18786 ) | ( ~n18787 & n18786 ) ;
  assign n18792 = ~n5135 & n14071 ;
  assign n18789 = n5010 | n11078 ;
  assign n18790 = n5067 | n13836 ;
  assign n18791 = n18789 &  n18790 ;
  assign n18793 = ( n5135 & n18792 ) | ( n5135 & n18791 ) | ( n18792 & n18791 ) ;
  assign n18794 = n5012 | n14079 ;
  assign n18795 = n18793 &  n18794 ;
  assign n18796 = x23 &  n18795 ;
  assign n18797 = x23 | n18795 ;
  assign n18798 = ~n18796 & n18797 ;
  assign n18799 = ( n18729 & n18788 ) | ( n18729 & n18798 ) | ( n18788 & n18798 ) ;
  assign n18800 = ( n18788 & ~n18729 ) | ( n18788 & n18798 ) | ( ~n18729 & n18798 ) ;
  assign n18801 = ( n18729 & ~n18799 ) | ( n18729 & n18800 ) | ( ~n18799 & n18800 ) ;
  assign n18803 = ( n5339 & ~n14355 ) | ( n5339 & 1'b0 ) | ( ~n14355 & 1'b0 ) ;
  assign n18804 = ~n5761 & n14553 ;
  assign n18805 = n18803 | n18804 ;
  assign n18806 = ~n5837 & n14803 ;
  assign n18807 = ( n5837 & ~n18805 ) | ( n5837 & n18806 ) | ( ~n18805 & n18806 ) ;
  assign n18808 = ~n5341 & n15310 ;
  assign n18809 = ( n18807 & ~n18808 ) | ( n18807 & 1'b0 ) | ( ~n18808 & 1'b0 ) ;
  assign n18810 = x20 &  n18809 ;
  assign n18811 = x20 | n18809 ;
  assign n18812 = ~n18810 & n18811 ;
  assign n18813 = ( n18802 & ~n18801 ) | ( n18802 & n18812 ) | ( ~n18801 & n18812 ) ;
  assign n18827 = ~n5135 & n14355 ;
  assign n18824 = n5010 | n13836 ;
  assign n18825 = n5067 | n14071 ;
  assign n18826 = n18824 &  n18825 ;
  assign n18828 = ( n5135 & n18827 ) | ( n5135 & n18826 ) | ( n18827 & n18826 ) ;
  assign n18829 = n5012 | n14363 ;
  assign n18830 = n18828 &  n18829 ;
  assign n18831 = x23 &  n18830 ;
  assign n18832 = x23 | n18830 ;
  assign n18833 = ~n18831 & n18832 ;
  assign n18837 = ~n4962 & n11078 ;
  assign n18834 = n4482 | n11081 ;
  assign n18835 = n4495 | n11085 ;
  assign n18836 = n18834 &  n18835 ;
  assign n18838 = ( n4962 & n18837 ) | ( n4962 & n18836 ) | ( n18837 & n18836 ) ;
  assign n18839 = n4478 | n11206 ;
  assign n18840 = n18838 &  n18839 ;
  assign n18841 = x26 &  n18840 ;
  assign n18842 = x26 | n18840 ;
  assign n18843 = ~n18841 & n18842 ;
  assign n18851 = ( n5965 & ~n5962 ) | ( n5965 & n5968 ) | ( ~n5962 & n5968 ) ;
  assign n18852 = n5962 | n18851 ;
  assign n18853 = n14800 &  n18852 ;
  assign n18868 = ( n16398 & ~n3474 ) | ( n16398 & n6777 ) | ( ~n3474 & n6777 ) ;
  assign n18869 = n3474 | n18868 ;
  assign n18865 = n207 | n490 ;
  assign n18866 = ( n18865 & ~n558 ) | ( n18865 & n643 ) | ( ~n558 & n643 ) ;
  assign n18867 = n558 | n18866 ;
  assign n18854 = n66 | x23 ;
  assign n18855 = ( x23 & ~n18854 ) | ( x23 & n38 ) | ( ~n18854 & n38 ) ;
  assign n18856 = ( n228 & ~n1491 ) | ( n228 & n572 ) | ( ~n1491 & n572 ) ;
  assign n18857 = n1491 | n18856 ;
  assign n18858 = ( n4834 & ~n2515 ) | ( n4834 & n18857 ) | ( ~n2515 & n18857 ) ;
  assign n18859 = n2515 | n18858 ;
  assign n18860 = ( n372 & ~n735 ) | ( n372 & n18859 ) | ( ~n735 & n18859 ) ;
  assign n18861 = n735 | n18860 ;
  assign n18862 = ( n492 & ~n336 ) | ( n492 & n18861 ) | ( ~n336 & n18861 ) ;
  assign n18863 = n336 | n18862 ;
  assign n18864 = ( n38 & ~n18855 ) | ( n38 & n18863 ) | ( ~n18855 & n18863 ) ;
  assign n18870 = ( n18869 & ~n18867 ) | ( n18869 & n18864 ) | ( ~n18867 & n18864 ) ;
  assign n18871 = ( n3756 & n18870 ) | ( n3756 & n18867 ) | ( n18870 & n18867 ) ;
  assign n18872 = ( n3756 & ~n18871 ) | ( n3756 & 1'b0 ) | ( ~n18871 & 1'b0 ) ;
  assign n18873 = ( n5246 & ~n3392 ) | ( n5246 & n18872 ) | ( ~n3392 & n18872 ) ;
  assign n18874 = n3392 &  n18873 ;
  assign n18875 = ( n2484 & ~n3213 ) | ( n2484 & n18874 ) | ( ~n3213 & n18874 ) ;
  assign n18876 = ( n18875 & ~n2484 ) | ( n18875 & 1'b0 ) | ( ~n2484 & 1'b0 ) ;
  assign n18877 = ( n624 & ~n18876 ) | ( n624 & n2309 ) | ( ~n18876 & n2309 ) ;
  assign n18878 = ( n624 & ~n18877 ) | ( n624 & 1'b0 ) | ( ~n18877 & 1'b0 ) ;
  assign n18879 = ( n775 & ~n18878 ) | ( n775 & n813 ) | ( ~n18878 & n813 ) ;
  assign n18880 = ( n813 & ~n18879 ) | ( n813 & 1'b0 ) | ( ~n18879 & 1'b0 ) ;
  assign n18881 = ( n670 & ~n574 ) | ( n670 & n18880 ) | ( ~n574 & n18880 ) ;
  assign n18882 = ~n670 & n18881 ;
  assign n18883 = n18751 | n18882 ;
  assign n18884 = n18751 &  n18882 ;
  assign n18885 = ( n18883 & ~n18884 ) | ( n18883 & 1'b0 ) | ( ~n18884 & 1'b0 ) ;
  assign n18886 = ( n18853 & ~x17 ) | ( n18853 & n18885 ) | ( ~x17 & n18885 ) ;
  assign n18887 = ( x17 & ~n18885 ) | ( x17 & n18853 ) | ( ~n18885 & n18853 ) ;
  assign n18888 = ( n18886 & ~n18853 ) | ( n18886 & n18887 ) | ( ~n18853 & n18887 ) ;
  assign n18844 = n3644 | n11218 ;
  assign n18845 = ( n3652 & ~n11104 ) | ( n3652 & 1'b0 ) | ( ~n11104 & 1'b0 ) ;
  assign n18846 = ( n3657 & ~n11101 ) | ( n3657 & 1'b0 ) | ( ~n11101 & 1'b0 ) ;
  assign n18847 = n18845 | n18846 ;
  assign n18848 = ~n3653 & n11098 ;
  assign n18849 = ( n3653 & ~n18847 ) | ( n3653 & n18848 ) | ( ~n18847 & n18848 ) ;
  assign n18850 = n18844 &  n18849 ;
  assign n18889 = ( n18753 & n18850 ) | ( n18753 & n18888 ) | ( n18850 & n18888 ) ;
  assign n18890 = ( n18753 & ~n18888 ) | ( n18753 & n18850 ) | ( ~n18888 & n18850 ) ;
  assign n18891 = ( n18888 & ~n18889 ) | ( n18888 & n18890 ) | ( ~n18889 & n18890 ) ;
  assign n18892 = ( n18762 & ~n18755 ) | ( n18762 & n18772 ) | ( ~n18755 & n18772 ) ;
  assign n18896 = ~n4430 & n11091 ;
  assign n18893 = n523 | n11095 ;
  assign n18894 = n3939 | n11093 ;
  assign n18895 = n18893 &  n18894 ;
  assign n18897 = ( n4430 & n18896 ) | ( n4430 & n18895 ) | ( n18896 & n18895 ) ;
  assign n18898 = n601 | n12984 ;
  assign n18899 = n18897 &  n18898 ;
  assign n18900 = x29 &  n18899 ;
  assign n18901 = x29 | n18899 ;
  assign n18902 = ~n18900 & n18901 ;
  assign n18903 = ( n18891 & ~n18892 ) | ( n18891 & n18902 ) | ( ~n18892 & n18902 ) ;
  assign n18904 = ( n18891 & ~n18902 ) | ( n18891 & n18892 ) | ( ~n18902 & n18892 ) ;
  assign n18905 = ( n18903 & ~n18891 ) | ( n18903 & n18904 ) | ( ~n18891 & n18904 ) ;
  assign n18906 = x26 | n18782 ;
  assign n18907 = x26 &  n18782 ;
  assign n18908 = ( n18906 & ~n18907 ) | ( n18906 & 1'b0 ) | ( ~n18907 & 1'b0 ) ;
  assign n18909 = ( n18733 & ~n18775 ) | ( n18733 & n18908 ) | ( ~n18775 & n18908 ) ;
  assign n18910 = ( n18843 & ~n18905 ) | ( n18843 & n18909 ) | ( ~n18905 & n18909 ) ;
  assign n18911 = ( n18843 & ~n18909 ) | ( n18843 & n18905 ) | ( ~n18909 & n18905 ) ;
  assign n18912 = ( n18910 & ~n18843 ) | ( n18910 & n18911 ) | ( ~n18843 & n18911 ) ;
  assign n18913 = ( n18729 & ~n18788 ) | ( n18729 & n18798 ) | ( ~n18788 & n18798 ) ;
  assign n18914 = ( n18833 & n18912 ) | ( n18833 & n18913 ) | ( n18912 & n18913 ) ;
  assign n18915 = ( n18912 & ~n18833 ) | ( n18912 & n18913 ) | ( ~n18833 & n18913 ) ;
  assign n18916 = ( n18833 & ~n18914 ) | ( n18833 & n18915 ) | ( ~n18914 & n18915 ) ;
  assign n18917 = ( n18813 & n18823 ) | ( n18813 & n18916 ) | ( n18823 & n18916 ) ;
  assign n19029 = ( n18813 & ~n18823 ) | ( n18813 & n18916 ) | ( ~n18823 & n18916 ) ;
  assign n19030 = ( n18823 & ~n18917 ) | ( n18823 & n19029 ) | ( ~n18917 & n19029 ) ;
  assign n19016 = n6170 &  n6395 ;
  assign n19017 = ( n14800 & ~n19016 ) | ( n14800 & 1'b0 ) | ( ~n19016 & 1'b0 ) ;
  assign n19018 = ~n5970 & n14807 ;
  assign n19019 = n19017 | n19018 ;
  assign n19020 = ( n5972 & n15692 ) | ( n5972 & n19019 ) | ( n15692 & n19019 ) ;
  assign n19021 = ( n15692 & ~n19020 ) | ( n15692 & 1'b0 ) | ( ~n19020 & 1'b0 ) ;
  assign n19022 = ( n19019 & ~x17 ) | ( n19019 & n19021 ) | ( ~x17 & n19021 ) ;
  assign n19023 = ( x17 & ~n19019 ) | ( x17 & n19021 ) | ( ~n19019 & n19021 ) ;
  assign n19024 = ( n19022 & ~n19021 ) | ( n19022 & n19023 ) | ( ~n19021 & n19023 ) ;
  assign n19015 = ( n18575 & ~n18682 ) | ( n18575 & n18692 ) | ( ~n18682 & n18692 ) ;
  assign n19025 = ( n18801 & n18802 ) | ( n18801 & n18812 ) | ( n18802 & n18812 ) ;
  assign n19026 = ( n18801 & ~n18802 ) | ( n18801 & n18812 ) | ( ~n18802 & n18812 ) ;
  assign n19027 = ( n18802 & ~n19025 ) | ( n18802 & n19026 ) | ( ~n19025 & n19026 ) ;
  assign n19028 = ( n19024 & ~n19015 ) | ( n19024 & n19027 ) | ( ~n19015 & n19027 ) ;
  assign n19031 = ( n19015 & n19024 ) | ( n19015 & n19027 ) | ( n19024 & n19027 ) ;
  assign n19032 = ( n19015 & ~n19024 ) | ( n19015 & n19027 ) | ( ~n19024 & n19027 ) ;
  assign n19033 = ( n19024 & ~n19031 ) | ( n19024 & n19032 ) | ( ~n19031 & n19032 ) ;
  assign n19035 = ( n18708 & ~n18583 ) | ( n18708 & n18709 ) | ( ~n18583 & n18709 ) ;
  assign n19034 = ( n18579 & ~n18695 ) | ( n18579 & n18705 ) | ( ~n18695 & n18705 ) ;
  assign n19036 = ( n19033 & ~n19035 ) | ( n19033 & n19034 ) | ( ~n19035 & n19034 ) ;
  assign n19046 = ( n19028 & n19030 ) | ( n19028 & n19036 ) | ( n19030 & n19036 ) ;
  assign n19045 = ( n19028 & ~n19030 ) | ( n19028 & n19036 ) | ( ~n19030 & n19036 ) ;
  assign n19047 = ( n19030 & ~n19046 ) | ( n19030 & n19045 ) | ( ~n19046 & n19045 ) ;
  assign n19065 = n19047 | n7783 ;
  assign n19062 = ( n7253 & ~n18712 ) | ( n7253 & 1'b0 ) | ( ~n18712 & 1'b0 ) ;
  assign n19041 = ( n19033 & ~n19034 ) | ( n19033 & n19035 ) | ( ~n19034 & n19035 ) ;
  assign n19042 = ( n19033 & n19034 ) | ( n19033 & n19035 ) | ( n19034 & n19035 ) ;
  assign n19043 = ( ~n19034 & ~n19041 ) | ( ~n19034 & n19042 ) | ( ~n19041 & n19042 ) ;
  assign n19063 = n7518 | n19043 ;
  assign n19064 = ~n19062 & n19063 ;
  assign n19066 = ( n7783 & ~n19065 ) | ( n7783 & n19064 ) | ( ~n19065 & n19064 ) ;
  assign n19052 = ( n18712 & n18719 ) | ( n18712 & n19043 ) | ( n18719 & n19043 ) ;
  assign n19053 = ( n19043 & ~n19047 ) | ( n19043 & n19052 ) | ( ~n19047 & n19052 ) ;
  assign n19067 = ( n19043 & ~n19052 ) | ( n19043 & n19047 ) | ( ~n19052 & n19047 ) ;
  assign n19068 = ( n19053 & ~n19043 ) | ( n19053 & n19067 ) | ( ~n19043 & n19067 ) ;
  assign n19069 = ~n7255 & n19068 ;
  assign n19070 = ( n19066 & ~n19069 ) | ( n19066 & 1'b0 ) | ( ~n19069 & 1'b0 ) ;
  assign n19071 = x11 &  n19070 ;
  assign n19072 = x11 | n19070 ;
  assign n19073 = ~n19071 & n19072 ;
  assign n19074 = ( n18470 & ~n18602 ) | ( n18470 & n18473 ) | ( ~n18602 & n18473 ) ;
  assign n19075 = ( n18473 & ~n18470 ) | ( n18473 & n18602 ) | ( ~n18470 & n18602 ) ;
  assign n19076 = ( n19074 & ~n18473 ) | ( n19074 & n19075 ) | ( ~n18473 & n19075 ) ;
  assign n19080 = ~n7783 & n19043 ;
  assign n19077 = ( n7253 & ~n18589 ) | ( n7253 & 1'b0 ) | ( ~n18589 & 1'b0 ) ;
  assign n19078 = n7518 | n18712 ;
  assign n19079 = ~n19077 & n19078 ;
  assign n19081 = ( n7783 & n19080 ) | ( n7783 & n19079 ) | ( n19080 & n19079 ) ;
  assign n19082 = ( n18719 & ~n18712 ) | ( n18719 & n19043 ) | ( ~n18712 & n19043 ) ;
  assign n19083 = ( n18712 & ~n19052 ) | ( n18712 & n19082 ) | ( ~n19052 & n19082 ) ;
  assign n19084 = ( n7255 & ~n19083 ) | ( n7255 & n19081 ) | ( ~n19083 & n19081 ) ;
  assign n19085 = ~n7255 & n19084 ;
  assign n19086 = ( x11 & ~n19081 ) | ( x11 & n19085 ) | ( ~n19081 & n19085 ) ;
  assign n19087 = ( n19081 & ~x11 ) | ( n19081 & n19085 ) | ( ~x11 & n19085 ) ;
  assign n19088 = ( n19086 & ~n19085 ) | ( n19086 & n19087 ) | ( ~n19085 & n19087 ) ;
  assign n19089 = ( n18322 & ~n18469 ) | ( n18322 & n18325 ) | ( ~n18469 & n18325 ) ;
  assign n19090 = ( n18325 & ~n18322 ) | ( n18325 & n18469 ) | ( ~n18322 & n18469 ) ;
  assign n19091 = ( n19089 & ~n18325 ) | ( n19089 & n19090 ) | ( ~n18325 & n19090 ) ;
  assign n19095 = ~n7783 & n18712 ;
  assign n19092 = ( n7253 & ~n18456 ) | ( n7253 & 1'b0 ) | ( ~n18456 & 1'b0 ) ;
  assign n19093 = n7518 | n18589 ;
  assign n19094 = ~n19092 & n19093 ;
  assign n19096 = ( n7783 & n19095 ) | ( n7783 & n19094 ) | ( n19095 & n19094 ) ;
  assign n19097 = ( n7255 & ~n18720 ) | ( n7255 & n19096 ) | ( ~n18720 & n19096 ) ;
  assign n19098 = ~n7255 & n19097 ;
  assign n19100 = ( x11 & n19096 ) | ( x11 & n19098 ) | ( n19096 & n19098 ) ;
  assign n19099 = ( x11 & ~n19098 ) | ( x11 & n19096 ) | ( ~n19098 & n19096 ) ;
  assign n19101 = ( n19098 & ~n19100 ) | ( n19098 & n19099 ) | ( ~n19100 & n19099 ) ;
  assign n19102 = ( n18063 & ~n18321 ) | ( n18063 & n18073 ) | ( ~n18321 & n18073 ) ;
  assign n19103 = ( n18322 & ~n18073 ) | ( n18322 & n19102 ) | ( ~n18073 & n19102 ) ;
  assign n19107 = ~n7783 & n18589 ;
  assign n19104 = ( n7253 & ~n17783 ) | ( n7253 & 1'b0 ) | ( ~n17783 & 1'b0 ) ;
  assign n19105 = n7518 | n18456 ;
  assign n19106 = ~n19104 & n19105 ;
  assign n19108 = ( n7783 & n19107 ) | ( n7783 & n19106 ) | ( n19107 & n19106 ) ;
  assign n19109 = ( n7255 & ~n18597 ) | ( n7255 & n19108 ) | ( ~n18597 & n19108 ) ;
  assign n19110 = ~n7255 & n19109 ;
  assign n19112 = ( x11 & n19108 ) | ( x11 & n19110 ) | ( n19108 & n19110 ) ;
  assign n19111 = ( x11 & ~n19110 ) | ( x11 & n19108 ) | ( ~n19110 & n19108 ) ;
  assign n19113 = ( n19110 & ~n19112 ) | ( n19110 & n19111 ) | ( ~n19112 & n19111 ) ;
  assign n19114 = ( n18076 & ~n18086 ) | ( n18076 & n18320 ) | ( ~n18086 & n18320 ) ;
  assign n19115 = ( n18086 & ~n18321 ) | ( n18086 & n19114 ) | ( ~n18321 & n19114 ) ;
  assign n19116 = ( n18096 & ~n18319 ) | ( n18096 & n18098 ) | ( ~n18319 & n18098 ) ;
  assign n19117 = ( n18098 & ~n18096 ) | ( n18098 & n18319 ) | ( ~n18096 & n18319 ) ;
  assign n19118 = ( n19116 & ~n18098 ) | ( n19116 & n19117 ) | ( ~n18098 & n19117 ) ;
  assign n19122 = ~n7783 & n18456 ;
  assign n19119 = ( n7253 & ~n17791 ) | ( n7253 & 1'b0 ) | ( ~n17791 & 1'b0 ) ;
  assign n19120 = n7518 | n17783 ;
  assign n19121 = ~n19119 & n19120 ;
  assign n19123 = ( n7783 & n19122 ) | ( n7783 & n19121 ) | ( n19122 & n19121 ) ;
  assign n19124 = ( n18464 & ~n7255 ) | ( n18464 & n19123 ) | ( ~n7255 & n19123 ) ;
  assign n19125 = ~n18464 & n19124 ;
  assign n19126 = ( x11 & ~n19123 ) | ( x11 & n19125 ) | ( ~n19123 & n19125 ) ;
  assign n19127 = ( n19123 & ~x11 ) | ( n19123 & n19125 ) | ( ~x11 & n19125 ) ;
  assign n19128 = ( n19126 & ~n19125 ) | ( n19126 & n19127 ) | ( ~n19125 & n19127 ) ;
  assign n19129 = ( n18110 & ~n18108 ) | ( n18110 & n18318 ) | ( ~n18108 & n18318 ) ;
  assign n19130 = ( n18108 & ~n18318 ) | ( n18108 & n18110 ) | ( ~n18318 & n18110 ) ;
  assign n19131 = ( n19129 & ~n18110 ) | ( n19129 & n19130 ) | ( ~n18110 & n19130 ) ;
  assign n19135 = ~n7783 & n17783 ;
  assign n19132 = ( n7253 & ~n17787 ) | ( n7253 & 1'b0 ) | ( ~n17787 & 1'b0 ) ;
  assign n19133 = n7518 | n17791 ;
  assign n19134 = ~n19132 & n19133 ;
  assign n19136 = ( n7783 & n19135 ) | ( n7783 & n19134 ) | ( n19135 & n19134 ) ;
  assign n19137 = ( n17799 & ~n7255 ) | ( n17799 & n19136 ) | ( ~n7255 & n19136 ) ;
  assign n19138 = ~n17799 & n19137 ;
  assign n19140 = ( x11 & n19136 ) | ( x11 & n19138 ) | ( n19136 & n19138 ) ;
  assign n19139 = ( x11 & ~n19138 ) | ( x11 & n19136 ) | ( ~n19138 & n19136 ) ;
  assign n19141 = ( n19138 & ~n19140 ) | ( n19138 & n19139 ) | ( ~n19140 & n19139 ) ;
  assign n19145 = ~n7783 & n17791 ;
  assign n19142 = ( n7253 & ~n17405 ) | ( n7253 & 1'b0 ) | ( ~n17405 & 1'b0 ) ;
  assign n19143 = n7518 | n17787 ;
  assign n19144 = ~n19142 & n19143 ;
  assign n19146 = ( n7783 & n19145 ) | ( n7783 & n19144 ) | ( n19145 & n19144 ) ;
  assign n19147 = n7255 | n17811 ;
  assign n19148 = n19146 &  n19147 ;
  assign n19149 = x11 &  n19148 ;
  assign n19150 = x11 | n19148 ;
  assign n19151 = ~n19149 & n19150 ;
  assign n19152 = ( n18113 & ~n18317 ) | ( n18113 & n18123 ) | ( ~n18317 & n18123 ) ;
  assign n19153 = ( n18318 & ~n18123 ) | ( n18318 & n19152 ) | ( ~n18123 & n19152 ) ;
  assign n19154 = ( n7253 & ~n17263 ) | ( n7253 & 1'b0 ) | ( ~n17263 & 1'b0 ) ;
  assign n19155 = n7518 | n17405 ;
  assign n19156 = ~n19154 & n19155 ;
  assign n19157 = ~n7783 & n17787 ;
  assign n19158 = ( n7783 & n19156 ) | ( n7783 & n19157 ) | ( n19156 & n19157 ) ;
  assign n19159 = n7255 | n17826 ;
  assign n19160 = n19158 &  n19159 ;
  assign n19161 = x11 &  n19160 ;
  assign n19162 = x11 | n19160 ;
  assign n19163 = ~n19161 & n19162 ;
  assign n19164 = ( n18126 & ~n18136 ) | ( n18126 & n18316 ) | ( ~n18136 & n18316 ) ;
  assign n19165 = ( n18136 & ~n18317 ) | ( n18136 & n19164 ) | ( ~n18317 & n19164 ) ;
  assign n19169 = ~n7783 & n17405 ;
  assign n19166 = n7253 &  n17107 ;
  assign n19167 = n7518 | n17263 ;
  assign n19168 = ~n19166 & n19167 ;
  assign n19170 = ( n7783 & n19169 ) | ( n7783 & n19168 ) | ( n19169 & n19168 ) ;
  assign n19171 = n7255 | n17413 ;
  assign n19172 = n19170 &  n19171 ;
  assign n19173 = x11 &  n19172 ;
  assign n19174 = x11 | n19172 ;
  assign n19175 = ~n19173 & n19174 ;
  assign n19176 = ( n18139 & ~n18149 ) | ( n18139 & n18315 ) | ( ~n18149 & n18315 ) ;
  assign n19177 = ( n18149 & ~n18316 ) | ( n18149 & n19176 ) | ( ~n18316 & n19176 ) ;
  assign n19181 = ( n7253 & ~n16589 ) | ( n7253 & 1'b0 ) | ( ~n16589 & 1'b0 ) ;
  assign n19182 = ~n7518 & n17107 ;
  assign n19183 = n19181 | n19182 ;
  assign n19184 = ~n7783 & n17263 ;
  assign n19185 = ( n7783 & ~n19183 ) | ( n7783 & n19184 ) | ( ~n19183 & n19184 ) ;
  assign n19186 = ( n7255 & ~n19185 ) | ( n7255 & n17271 ) | ( ~n19185 & n17271 ) ;
  assign n19187 = ( n17271 & ~n19186 ) | ( n17271 & 1'b0 ) | ( ~n19186 & 1'b0 ) ;
  assign n19189 = ( x11 & n19185 ) | ( x11 & n19187 ) | ( n19185 & n19187 ) ;
  assign n19188 = ( x11 & ~n19187 ) | ( x11 & n19185 ) | ( ~n19187 & n19185 ) ;
  assign n19190 = ( n19187 & ~n19189 ) | ( n19187 & n19188 ) | ( ~n19189 & n19188 ) ;
  assign n19178 = ( n18161 & ~n18159 ) | ( n18161 & n18314 ) | ( ~n18159 & n18314 ) ;
  assign n19179 = ( n18159 & ~n18314 ) | ( n18159 & n18161 ) | ( ~n18314 & n18161 ) ;
  assign n19180 = ( n19178 & ~n18161 ) | ( n19178 & n19179 ) | ( ~n18161 & n19179 ) ;
  assign n19191 = ( n18173 & ~n18171 ) | ( n18173 & n18313 ) | ( ~n18171 & n18313 ) ;
  assign n19192 = ( n18171 & ~n18313 ) | ( n18171 & n18173 ) | ( ~n18313 & n18173 ) ;
  assign n19193 = ( n19191 & ~n18173 ) | ( n19191 & n19192 ) | ( ~n18173 & n19192 ) ;
  assign n19197 = n17107 | n7783 ;
  assign n19194 = ( n7253 & ~n16595 ) | ( n7253 & 1'b0 ) | ( ~n16595 & 1'b0 ) ;
  assign n19195 = n7518 | n16589 ;
  assign n19196 = ~n19194 & n19195 ;
  assign n19198 = ( n7783 & ~n19197 ) | ( n7783 & n19196 ) | ( ~n19197 & n19196 ) ;
  assign n19199 = ( n7255 & ~n19198 ) | ( n7255 & n17115 ) | ( ~n19198 & n17115 ) ;
  assign n19200 = ( n17115 & ~n19199 ) | ( n17115 & 1'b0 ) | ( ~n19199 & 1'b0 ) ;
  assign n19201 = ( x11 & ~n19198 ) | ( x11 & n19200 ) | ( ~n19198 & n19200 ) ;
  assign n19202 = ( n19198 & ~x11 ) | ( n19198 & n19200 ) | ( ~x11 & n19200 ) ;
  assign n19203 = ( n19201 & ~n19200 ) | ( n19201 & n19202 ) | ( ~n19200 & n19202 ) ;
  assign n19204 = ( n18185 & ~n18183 ) | ( n18185 & n18312 ) | ( ~n18183 & n18312 ) ;
  assign n19205 = ( n18183 & ~n18312 ) | ( n18183 & n18185 ) | ( ~n18312 & n18185 ) ;
  assign n19206 = ( n19204 & ~n18185 ) | ( n19204 & n19205 ) | ( ~n18185 & n19205 ) ;
  assign n19210 = ~n7783 & n16589 ;
  assign n19207 = ( n7253 & ~n16591 ) | ( n7253 & 1'b0 ) | ( ~n16591 & 1'b0 ) ;
  assign n19208 = n7518 | n16595 ;
  assign n19209 = ~n19207 & n19208 ;
  assign n19211 = ( n7783 & n19210 ) | ( n7783 & n19209 ) | ( n19210 & n19209 ) ;
  assign n19212 = ( n16604 & ~n7255 ) | ( n16604 & n19211 ) | ( ~n7255 & n19211 ) ;
  assign n19213 = ~n16604 & n19212 ;
  assign n19215 = ( x11 & n19211 ) | ( x11 & n19213 ) | ( n19211 & n19213 ) ;
  assign n19214 = ( x11 & ~n19213 ) | ( x11 & n19211 ) | ( ~n19213 & n19211 ) ;
  assign n19216 = ( n19213 & ~n19215 ) | ( n19213 & n19214 ) | ( ~n19215 & n19214 ) ;
  assign n19220 = ~n7783 & n16595 ;
  assign n19217 = ( n7253 & ~n16091 ) | ( n7253 & 1'b0 ) | ( ~n16091 & 1'b0 ) ;
  assign n19218 = n7518 | n16591 ;
  assign n19219 = ~n19217 & n19218 ;
  assign n19221 = ( n7783 & n19220 ) | ( n7783 & n19219 ) | ( n19220 & n19219 ) ;
  assign n19222 = n7255 | n16616 ;
  assign n19223 = n19221 &  n19222 ;
  assign n19224 = x11 &  n19223 ;
  assign n19225 = x11 | n19223 ;
  assign n19226 = ~n19224 & n19225 ;
  assign n19227 = ( n18188 & ~n18311 ) | ( n18188 & n18198 ) | ( ~n18311 & n18198 ) ;
  assign n19228 = ( n18312 & ~n18198 ) | ( n18312 & n19227 ) | ( ~n18198 & n19227 ) ;
  assign n19232 = ~n7783 & n16591 ;
  assign n19229 = ( n7253 & ~n15897 ) | ( n7253 & 1'b0 ) | ( ~n15897 & 1'b0 ) ;
  assign n19230 = n7518 | n16091 ;
  assign n19231 = ~n19229 & n19230 ;
  assign n19233 = ( n7783 & n19232 ) | ( n7783 & n19231 ) | ( n19232 & n19231 ) ;
  assign n19234 = n7255 | n16631 ;
  assign n19235 = n19233 &  n19234 ;
  assign n19236 = x11 &  n19235 ;
  assign n19237 = x11 | n19235 ;
  assign n19238 = ~n19236 & n19237 ;
  assign n19239 = ( n18201 & ~n18211 ) | ( n18201 & n18310 ) | ( ~n18211 & n18310 ) ;
  assign n19240 = ( n18211 & ~n18311 ) | ( n18211 & n19239 ) | ( ~n18311 & n19239 ) ;
  assign n19244 = ~n7783 & n16091 ;
  assign n19241 = ( n7253 & ~n15700 ) | ( n7253 & 1'b0 ) | ( ~n15700 & 1'b0 ) ;
  assign n19242 = n7518 | n15897 ;
  assign n19243 = ~n19241 & n19242 ;
  assign n19245 = ( n7783 & n19244 ) | ( n7783 & n19243 ) | ( n19244 & n19243 ) ;
  assign n19246 = n7255 | n16094 ;
  assign n19247 = n19245 &  n19246 ;
  assign n19248 = x11 &  n19247 ;
  assign n19249 = x11 | n19247 ;
  assign n19250 = ~n19248 & n19249 ;
  assign n19251 = ( n18214 & ~n18224 ) | ( n18214 & n18309 ) | ( ~n18224 & n18309 ) ;
  assign n19252 = ( n18224 & ~n18310 ) | ( n18224 & n19251 ) | ( ~n18310 & n19251 ) ;
  assign n19259 = ~n7783 & n15897 ;
  assign n19256 = ( n7253 & ~n15320 ) | ( n7253 & 1'b0 ) | ( ~n15320 & 1'b0 ) ;
  assign n19257 = n7518 | n15700 ;
  assign n19258 = ~n19256 & n19257 ;
  assign n19260 = ( n7783 & n19259 ) | ( n7783 & n19258 ) | ( n19259 & n19258 ) ;
  assign n19261 = ( n15900 & ~n7255 ) | ( n15900 & n19260 ) | ( ~n7255 & n19260 ) ;
  assign n19262 = ~n15900 & n19261 ;
  assign n19263 = ( x11 & ~n19260 ) | ( x11 & n19262 ) | ( ~n19260 & n19262 ) ;
  assign n19264 = ( n19260 & ~x11 ) | ( n19260 & n19262 ) | ( ~x11 & n19262 ) ;
  assign n19265 = ( n19263 & ~n19262 ) | ( n19263 & n19264 ) | ( ~n19262 & n19264 ) ;
  assign n19253 = ( n18236 & ~n18234 ) | ( n18236 & n18308 ) | ( ~n18234 & n18308 ) ;
  assign n19254 = ( n18234 & ~n18308 ) | ( n18234 & n18236 ) | ( ~n18308 & n18236 ) ;
  assign n19255 = ( n19253 & ~n18236 ) | ( n19253 & n19254 ) | ( ~n18236 & n19254 ) ;
  assign n19266 = ( n18249 & ~n18239 ) | ( n18249 & n18307 ) | ( ~n18239 & n18307 ) ;
  assign n19267 = ( n18239 & ~n18307 ) | ( n18239 & n18249 ) | ( ~n18307 & n18249 ) ;
  assign n19268 = ( n19266 & ~n18249 ) | ( n19266 & n19267 ) | ( ~n18249 & n19267 ) ;
  assign n19272 = ~n7783 & n15700 ;
  assign n19269 = ( n7253 & ~n15325 ) | ( n7253 & 1'b0 ) | ( ~n15325 & 1'b0 ) ;
  assign n19270 = n7518 | n15320 ;
  assign n19271 = ~n19269 & n19270 ;
  assign n19273 = ( n7783 & n19272 ) | ( n7783 & n19271 ) | ( n19272 & n19271 ) ;
  assign n19274 = ( n15708 & ~n7255 ) | ( n15708 & n19273 ) | ( ~n7255 & n19273 ) ;
  assign n19275 = ~n15708 & n19274 ;
  assign n19277 = ( x11 & n19273 ) | ( x11 & n19275 ) | ( n19273 & n19275 ) ;
  assign n19276 = ( x11 & ~n19275 ) | ( x11 & n19273 ) | ( ~n19275 & n19273 ) ;
  assign n19278 = ( n19275 & ~n19277 ) | ( n19275 & n19276 ) | ( ~n19277 & n19276 ) ;
  assign n19279 = ( n18259 & ~n18306 ) | ( n18259 & n18264 ) | ( ~n18306 & n18264 ) ;
  assign n19280 = ( n18264 & ~n18259 ) | ( n18264 & n18306 ) | ( ~n18259 & n18306 ) ;
  assign n19281 = ( n19279 & ~n18264 ) | ( n19279 & n19280 ) | ( ~n18264 & n19280 ) ;
  assign n19285 = ~n7783 & n15320 ;
  assign n19282 = ( n7253 & ~n15322 ) | ( n7253 & 1'b0 ) | ( ~n15322 & 1'b0 ) ;
  assign n19283 = n7518 | n15325 ;
  assign n19284 = ~n19282 & n19283 ;
  assign n19286 = ( n7783 & n19285 ) | ( n7783 & n19284 ) | ( n19285 & n19284 ) ;
  assign n19287 = ( n15334 & ~n7255 ) | ( n15334 & n19286 ) | ( ~n7255 & n19286 ) ;
  assign n19288 = ~n15334 & n19287 ;
  assign n19289 = ( x11 & ~n19286 ) | ( x11 & n19288 ) | ( ~n19286 & n19288 ) ;
  assign n19290 = ( n19286 & ~x11 ) | ( n19286 & n19288 ) | ( ~x11 & n19288 ) ;
  assign n19291 = ( n19289 & ~n19288 ) | ( n19289 & n19290 ) | ( ~n19288 & n19290 ) ;
  assign n19295 = ~n7783 & n15325 ;
  assign n19292 = n7253 &  n14745 ;
  assign n19293 = n7518 | n15322 ;
  assign n19294 = ~n19292 & n19293 ;
  assign n19296 = ( n7783 & n19295 ) | ( n7783 & n19294 ) | ( n19295 & n19294 ) ;
  assign n19297 = n7255 | n15346 ;
  assign n19298 = n19296 &  n19297 ;
  assign n19299 = x11 &  n19298 ;
  assign n19300 = x11 | n19298 ;
  assign n19301 = ~n19299 & n19300 ;
  assign n19302 = ( n18278 & ~n18268 ) | ( n18278 & n18305 ) | ( ~n18268 & n18305 ) ;
  assign n19303 = ( n18306 & ~n18278 ) | ( n18306 & n19302 ) | ( ~n18278 & n19302 ) ;
  assign n19305 = ( n18015 & n18294 ) | ( n18015 & n18304 ) | ( n18294 & n18304 ) ;
  assign n19304 = ( n18015 & ~n18294 ) | ( n18015 & n18304 ) | ( ~n18294 & n18304 ) ;
  assign n19306 = ( n18294 & ~n19305 ) | ( n18294 & n19304 ) | ( ~n19305 & n19304 ) ;
  assign n19307 = ( n7253 & ~n14528 ) | ( n7253 & 1'b0 ) | ( ~n14528 & 1'b0 ) ;
  assign n19308 = ~n7518 & n14745 ;
  assign n19309 = n19307 | n19308 ;
  assign n19310 = ~n7783 & n15322 ;
  assign n19311 = ( n7783 & ~n19309 ) | ( n7783 & n19310 ) | ( ~n19309 & n19310 ) ;
  assign n19312 = ( n7255 & ~n19311 ) | ( n7255 & n15361 ) | ( ~n19311 & n15361 ) ;
  assign n19313 = ( n15361 & ~n19312 ) | ( n15361 & 1'b0 ) | ( ~n19312 & 1'b0 ) ;
  assign n19314 = ( x11 & ~n19311 ) | ( x11 & n19313 ) | ( ~n19311 & n19313 ) ;
  assign n19315 = ( n19311 & ~x11 ) | ( n19311 & n19313 ) | ( ~x11 & n19313 ) ;
  assign n19316 = ( n19314 & ~n19313 ) | ( n19314 & n19315 ) | ( ~n19313 & n19315 ) ;
  assign n19320 = n14745 | n7783 ;
  assign n19317 = ( n7253 & ~n14261 ) | ( n7253 & 1'b0 ) | ( ~n14261 & 1'b0 ) ;
  assign n19318 = n7518 | n14528 ;
  assign n19319 = ~n19317 & n19318 ;
  assign n19321 = ( n7783 & ~n19320 ) | ( n7783 & n19319 ) | ( ~n19320 & n19319 ) ;
  assign n19322 = ~n7255 & n14749 ;
  assign n19323 = ( n19321 & ~n19322 ) | ( n19321 & 1'b0 ) | ( ~n19322 & 1'b0 ) ;
  assign n19324 = x11 &  n19323 ;
  assign n19325 = x11 | n19323 ;
  assign n19326 = ~n19324 & n19325 ;
  assign n19327 = ( x14 & n18279 ) | ( x14 & n18284 ) | ( n18279 & n18284 ) ;
  assign n19328 = ~n18279 & n19327 ;
  assign n19329 = ( n18291 & ~x14 ) | ( n18291 & n19328 ) | ( ~x14 & n19328 ) ;
  assign n19330 = ( x14 & ~n18291 ) | ( x14 & n19328 ) | ( ~n18291 & n19328 ) ;
  assign n19331 = ( n19329 & ~n19328 ) | ( n19329 & n19330 ) | ( ~n19328 & n19330 ) ;
  assign n19332 = x14 &  n18279 ;
  assign n19333 = n18284 &  n19332 ;
  assign n19334 = n18284 | n19332 ;
  assign n19335 = ~n19333 & n19334 ;
  assign n19362 = ( n7253 & ~n13785 ) | ( n7253 & 1'b0 ) | ( ~n13785 & 1'b0 ) ;
  assign n19363 = n7518 | n13998 ;
  assign n19364 = ~n19362 & n19363 ;
  assign n19365 = ~n7783 & n14261 ;
  assign n19366 = ( n7783 & n19364 ) | ( n7783 & n19365 ) | ( n19364 & n19365 ) ;
  assign n19367 = n7255 | n14267 ;
  assign n19368 = n19366 &  n19367 ;
  assign n19369 = x11 &  n19368 ;
  assign n19370 = x11 | n19368 ;
  assign n19371 = ~n19369 & n19370 ;
  assign n19346 = ( n7251 & ~n13787 ) | ( n7251 & 1'b0 ) | ( ~n13787 & 1'b0 ) ;
  assign n19350 = n13790 | n7255 ;
  assign n19347 = n7518 | n13787 ;
  assign n19348 = n7783 | n13785 ;
  assign n19349 = n19347 &  n19348 ;
  assign n19351 = ( n7255 & ~n19350 ) | ( n7255 & n19349 ) | ( ~n19350 & n19349 ) ;
  assign n19357 = ~n7255 & n14001 ;
  assign n19355 = ~n7783 & n13998 ;
  assign n19352 = ( n7253 & ~n13787 ) | ( n7253 & 1'b0 ) | ( ~n13787 & 1'b0 ) ;
  assign n19353 = n7518 | n13785 ;
  assign n19354 = ~n19352 & n19353 ;
  assign n19356 = ( n7783 & n19355 ) | ( n7783 & n19354 ) | ( n19355 & n19354 ) ;
  assign n19358 = ( n7255 & n19357 ) | ( n7255 & n19356 ) | ( n19357 & n19356 ) ;
  assign n19359 = ( n19346 & n19351 ) | ( n19346 & n19358 ) | ( n19351 & n19358 ) ;
  assign n19360 = ( x11 & ~n19359 ) | ( x11 & n19346 ) | ( ~n19359 & n19346 ) ;
  assign n19361 = ( x11 & ~n19360 ) | ( x11 & 1'b0 ) | ( ~n19360 & 1'b0 ) ;
  assign n19372 = ( n18279 & ~n19371 ) | ( n18279 & n19361 ) | ( ~n19371 & n19361 ) ;
  assign n19339 = ~n7783 & n14528 ;
  assign n19336 = ( n7253 & ~n13998 ) | ( n7253 & 1'b0 ) | ( ~n13998 & 1'b0 ) ;
  assign n19337 = n7518 | n14261 ;
  assign n19338 = ~n19336 & n19337 ;
  assign n19340 = ( n7783 & n19339 ) | ( n7783 & n19338 ) | ( n19339 & n19338 ) ;
  assign n19341 = ( n14532 & ~n7255 ) | ( n14532 & n19340 ) | ( ~n7255 & n19340 ) ;
  assign n19342 = ~n14532 & n19341 ;
  assign n19343 = ( x11 & ~n19340 ) | ( x11 & n19342 ) | ( ~n19340 & n19342 ) ;
  assign n19344 = ( n19340 & ~x11 ) | ( n19340 & n19342 ) | ( ~x11 & n19342 ) ;
  assign n19345 = ( n19343 & ~n19342 ) | ( n19343 & n19344 ) | ( ~n19342 & n19344 ) ;
  assign n19373 = ( n19335 & ~n19372 ) | ( n19335 & n19345 ) | ( ~n19372 & n19345 ) ;
  assign n19374 = ( n19326 & n19331 ) | ( n19326 & n19373 ) | ( n19331 & n19373 ) ;
  assign n19375 = ( n19306 & n19316 ) | ( n19306 & n19374 ) | ( n19316 & n19374 ) ;
  assign n19376 = ( n19301 & ~n19303 ) | ( n19301 & n19375 ) | ( ~n19303 & n19375 ) ;
  assign n19377 = ( n19281 & n19291 ) | ( n19281 & n19376 ) | ( n19291 & n19376 ) ;
  assign n19378 = ( n19268 & n19278 ) | ( n19268 & n19377 ) | ( n19278 & n19377 ) ;
  assign n19379 = ( n19265 & ~n19255 ) | ( n19265 & n19378 ) | ( ~n19255 & n19378 ) ;
  assign n19380 = ( n19250 & n19252 ) | ( n19250 & n19379 ) | ( n19252 & n19379 ) ;
  assign n19381 = ( n19238 & n19240 ) | ( n19238 & n19380 ) | ( n19240 & n19380 ) ;
  assign n19382 = ( n19226 & ~n19228 ) | ( n19226 & n19381 ) | ( ~n19228 & n19381 ) ;
  assign n19383 = ( n19206 & n19216 ) | ( n19206 & n19382 ) | ( n19216 & n19382 ) ;
  assign n19384 = ( n19193 & n19203 ) | ( n19193 & n19383 ) | ( n19203 & n19383 ) ;
  assign n19385 = ( n19190 & ~n19180 ) | ( n19190 & n19384 ) | ( ~n19180 & n19384 ) ;
  assign n19386 = ( n19175 & n19177 ) | ( n19175 & n19385 ) | ( n19177 & n19385 ) ;
  assign n19387 = ( n19163 & n19165 ) | ( n19163 & n19386 ) | ( n19165 & n19386 ) ;
  assign n19388 = ( n19151 & ~n19153 ) | ( n19151 & n19387 ) | ( ~n19153 & n19387 ) ;
  assign n19389 = ( n19131 & n19141 ) | ( n19131 & n19388 ) | ( n19141 & n19388 ) ;
  assign n19390 = ( n19118 & n19128 ) | ( n19118 & n19389 ) | ( n19128 & n19389 ) ;
  assign n19391 = ( n19113 & n19115 ) | ( n19113 & n19390 ) | ( n19115 & n19390 ) ;
  assign n19392 = ( n19101 & ~n19103 ) | ( n19101 & n19391 ) | ( ~n19103 & n19391 ) ;
  assign n19393 = ( n19088 & n19091 ) | ( n19088 & n19392 ) | ( n19091 & n19392 ) ;
  assign n19394 = ( n19073 & n19076 ) | ( n19073 & n19393 ) | ( n19076 & n19393 ) ;
  assign n18918 = ( n18843 & n18905 ) | ( n18843 & n18909 ) | ( n18905 & n18909 ) ;
  assign n18919 = ( n485 & ~n349 ) | ( n485 & n2959 ) | ( ~n349 & n2959 ) ;
  assign n18920 = n349 | n18919 ;
  assign n18921 = ( n237 & ~n529 ) | ( n237 & n18920 ) | ( ~n529 & n18920 ) ;
  assign n18922 = n529 | n18921 ;
  assign n18923 = n196 | n18922 ;
  assign n18924 = ( n5430 & ~n960 ) | ( n5430 & n14311 ) | ( ~n960 & n14311 ) ;
  assign n18925 = n960 | n18924 ;
  assign n18926 = ( n18923 & ~n3245 ) | ( n18923 & n18925 ) | ( ~n3245 & n18925 ) ;
  assign n18927 = n3245 | n18926 ;
  assign n18928 = ( n229 & n18927 ) | ( n229 & n813 ) | ( n18927 & n813 ) ;
  assign n18929 = ( n813 & ~n18928 ) | ( n813 & 1'b0 ) | ( ~n18928 & 1'b0 ) ;
  assign n18930 = ~n166 & n18929 ;
  assign n18931 = ( n425 & ~n475 ) | ( n425 & n672 ) | ( ~n475 & n672 ) ;
  assign n18932 = n475 | n18931 ;
  assign n18933 = ( n70 & n1547 ) | ( n70 & n18932 ) | ( n1547 & n18932 ) ;
  assign n18934 = ( n1547 & ~n18933 ) | ( n1547 & 1'b0 ) | ( ~n18933 & 1'b0 ) ;
  assign n18935 = ~n117 & n18934 ;
  assign n18936 = ( n1690 & ~n1434 ) | ( n1690 & n2188 ) | ( ~n1434 & n2188 ) ;
  assign n18937 = ~n1690 & n18936 ;
  assign n18938 = ( n3267 & n18935 ) | ( n3267 & n18937 ) | ( n18935 & n18937 ) ;
  assign n18939 = ~n3267 & n18938 ;
  assign n18940 = n18930 &  n18939 ;
  assign n18941 = ( n18864 & ~n14303 ) | ( n18864 & n18940 ) | ( ~n14303 & n18940 ) ;
  assign n18942 = ( n3409 & ~n18941 ) | ( n3409 & n18864 ) | ( ~n18941 & n18864 ) ;
  assign n18943 = ( n3409 & ~n18942 ) | ( n3409 & 1'b0 ) | ( ~n18942 & 1'b0 ) ;
  assign n18944 = ( n2082 & ~n134 ) | ( n2082 & n18943 ) | ( ~n134 & n18943 ) ;
  assign n18945 = ~n2082 & n18944 ;
  assign n18946 = ( n138 & ~n150 ) | ( n138 & n18945 ) | ( ~n150 & n18945 ) ;
  assign n18947 = ~n138 & n18946 ;
  assign n18948 = ( n230 & ~n734 ) | ( n230 & n18947 ) | ( ~n734 & n18947 ) ;
  assign n18949 = ~n230 & n18948 ;
  assign n18957 = ~x17 & n18853 ;
  assign n18958 = ( n18883 & ~n18886 ) | ( n18883 & n18957 ) | ( ~n18886 & n18957 ) ;
  assign n18955 = ~n3644 & n13014 ;
  assign n18950 = n3653 | n11095 ;
  assign n18951 = ( n3657 & ~n11098 ) | ( n3657 & 1'b0 ) | ( ~n11098 & 1'b0 ) ;
  assign n18952 = ( n3652 & ~n11101 ) | ( n3652 & 1'b0 ) | ( ~n11101 & 1'b0 ) ;
  assign n18953 = n18951 | n18952 ;
  assign n18954 = ( n18950 & ~n18953 ) | ( n18950 & 1'b0 ) | ( ~n18953 & 1'b0 ) ;
  assign n18956 = ( n3644 & n18955 ) | ( n3644 & n18954 ) | ( n18955 & n18954 ) ;
  assign n18959 = ( n18949 & ~n18958 ) | ( n18949 & n18956 ) | ( ~n18958 & n18956 ) ;
  assign n18960 = ( n18949 & ~n18956 ) | ( n18949 & n18958 ) | ( ~n18956 & n18958 ) ;
  assign n18961 = ( n18959 & ~n18949 ) | ( n18959 & n18960 ) | ( ~n18949 & n18960 ) ;
  assign n18962 = ~n18889 & n18961 ;
  assign n18963 = ( n18889 & ~n18961 ) | ( n18889 & 1'b0 ) | ( ~n18961 & 1'b0 ) ;
  assign n18964 = n18962 | n18963 ;
  assign n18970 = ~n601 & n13775 ;
  assign n18968 = ~n4430 & n11081 ;
  assign n18965 = n523 | n11093 ;
  assign n18966 = n3939 | n11091 ;
  assign n18967 = n18965 &  n18966 ;
  assign n18969 = ( n4430 & n18968 ) | ( n4430 & n18967 ) | ( n18968 & n18967 ) ;
  assign n18971 = ( n601 & n18970 ) | ( n601 & n18969 ) | ( n18970 & n18969 ) ;
  assign n18972 = ( n18964 & ~x29 ) | ( n18964 & n18971 ) | ( ~x29 & n18971 ) ;
  assign n18973 = ( x29 & ~n18964 ) | ( x29 & n18971 ) | ( ~n18964 & n18971 ) ;
  assign n18974 = ( n18972 & ~n18971 ) | ( n18972 & n18973 ) | ( ~n18971 & n18973 ) ;
  assign n18975 = ( n18891 & n18892 ) | ( n18891 & n18902 ) | ( n18892 & n18902 ) ;
  assign n18979 = ~n4962 & n13836 ;
  assign n18976 = n4482 | n11085 ;
  assign n18977 = n4495 | n11078 ;
  assign n18978 = n18976 &  n18977 ;
  assign n18980 = ( n4962 & n18979 ) | ( n4962 & n18978 ) | ( n18979 & n18978 ) ;
  assign n18981 = n4478 | n13844 ;
  assign n18982 = n18980 &  n18981 ;
  assign n18983 = x26 &  n18982 ;
  assign n18984 = x26 | n18982 ;
  assign n18985 = ~n18983 & n18984 ;
  assign n18986 = ( n18974 & ~n18975 ) | ( n18974 & n18985 ) | ( ~n18975 & n18985 ) ;
  assign n18987 = ( n18974 & ~n18985 ) | ( n18974 & n18975 ) | ( ~n18985 & n18975 ) ;
  assign n18988 = ( n18986 & ~n18974 ) | ( n18986 & n18987 ) | ( ~n18974 & n18987 ) ;
  assign n18992 = n14553 | n5135 ;
  assign n18989 = n5010 | n14071 ;
  assign n18990 = n5067 | n14355 ;
  assign n18991 = n18989 &  n18990 ;
  assign n18993 = ( n5135 & ~n18992 ) | ( n5135 & n18991 ) | ( ~n18992 & n18991 ) ;
  assign n18994 = ~n5012 & n14562 ;
  assign n18995 = ( n18993 & ~n18994 ) | ( n18993 & 1'b0 ) | ( ~n18994 & 1'b0 ) ;
  assign n18996 = x23 &  n18995 ;
  assign n18997 = x23 | n18995 ;
  assign n18998 = ~n18996 & n18997 ;
  assign n18999 = ( n18918 & n18988 ) | ( n18918 & n18998 ) | ( n18988 & n18998 ) ;
  assign n19000 = ( n18988 & ~n18918 ) | ( n18988 & n18998 ) | ( ~n18918 & n18998 ) ;
  assign n19001 = ( n18918 & ~n18999 ) | ( n18918 & n19000 ) | ( ~n18999 & n19000 ) ;
  assign n19005 = n14800 | n5837 ;
  assign n19002 = ( n5339 & ~n14803 ) | ( n5339 & 1'b0 ) | ( ~n14803 & 1'b0 ) ;
  assign n19003 = ~n5761 & n14807 ;
  assign n19004 = n19002 | n19003 ;
  assign n19006 = ( n19005 & ~n5837 ) | ( n19005 & n19004 ) | ( ~n5837 & n19004 ) ;
  assign n19007 = n5341 | n14816 ;
  assign n19008 = ~n19006 & n19007 ;
  assign n19009 = x20 &  n19008 ;
  assign n19010 = x20 | n19008 ;
  assign n19011 = ~n19009 & n19010 ;
  assign n19012 = ( n18914 & n19001 ) | ( n18914 & n19011 ) | ( n19001 & n19011 ) ;
  assign n19013 = ( n19001 & ~n18914 ) | ( n19001 & n19011 ) | ( ~n18914 & n19011 ) ;
  assign n19014 = ( n18914 & ~n19012 ) | ( n18914 & n19013 ) | ( ~n19012 & n19013 ) ;
  assign n19037 = ( n19030 & ~n19028 ) | ( n19030 & n19036 ) | ( ~n19028 & n19036 ) ;
  assign n19038 = ( n18917 & n19014 ) | ( n18917 & n19037 ) | ( n19014 & n19037 ) ;
  assign n19039 = ( n19014 & ~n18917 ) | ( n19014 & n19037 ) | ( ~n18917 & n19037 ) ;
  assign n19040 = ( n18917 & ~n19038 ) | ( n18917 & n19039 ) | ( ~n19038 & n19039 ) ;
  assign n19050 = n19040 | n7783 ;
  assign n19044 = ( n7253 & ~n19043 ) | ( n7253 & 1'b0 ) | ( ~n19043 & 1'b0 ) ;
  assign n19048 = ~n7518 & n19047 ;
  assign n19049 = n19044 | n19048 ;
  assign n19051 = ( n19050 & ~n7783 ) | ( n19050 & n19049 ) | ( ~n7783 & n19049 ) ;
  assign n19054 = ( n19047 & ~n19040 ) | ( n19047 & n19053 ) | ( ~n19040 & n19053 ) ;
  assign n19055 = ( n19040 & ~n19053 ) | ( n19040 & n19047 ) | ( ~n19053 & n19047 ) ;
  assign n19056 = ( n19054 & ~n19047 ) | ( n19054 & n19055 ) | ( ~n19047 & n19055 ) ;
  assign n19057 = n7255 | n19056 ;
  assign n19058 = ~n19051 & n19057 ;
  assign n19059 = x11 &  n19058 ;
  assign n19060 = x11 | n19058 ;
  assign n19061 = ~n19059 & n19060 ;
  assign n19395 = ( n18728 & ~n19394 ) | ( n18728 & n19061 ) | ( ~n19394 & n19061 ) ;
  assign n19396 = ( n18728 & ~n19061 ) | ( n18728 & n19394 ) | ( ~n19061 & n19394 ) ;
  assign n19397 = ( n19395 & ~n18728 ) | ( n19395 & n19396 ) | ( ~n18728 & n19396 ) ;
  assign n19398 = ( n19091 & ~n19088 ) | ( n19091 & n19392 ) | ( ~n19088 & n19392 ) ;
  assign n19399 = ( n19088 & ~n19392 ) | ( n19088 & n19091 ) | ( ~n19392 & n19091 ) ;
  assign n19400 = ( n19398 & ~n19091 ) | ( n19398 & n19399 ) | ( ~n19091 & n19399 ) ;
  assign n19495 = n8105 &  n19047 ;
  assign n19496 = ~n8429 & n19040 ;
  assign n19497 = n19495 | n19496 ;
  assign n19401 = ( n18914 & ~n19001 ) | ( n18914 & n19011 ) | ( ~n19001 & n19011 ) ;
  assign n19402 = n5761 &  n5837 ;
  assign n19403 = ( n14800 & ~n19402 ) | ( n14800 & 1'b0 ) | ( ~n19402 & 1'b0 ) ;
  assign n19404 = n5339 &  n14807 ;
  assign n19405 = n19403 | n19404 ;
  assign n19406 = ( n5341 & n15692 ) | ( n5341 & n19405 ) | ( n15692 & n19405 ) ;
  assign n19407 = ( n15692 & ~n19406 ) | ( n15692 & 1'b0 ) | ( ~n19406 & 1'b0 ) ;
  assign n19408 = ( n19405 & ~x20 ) | ( n19405 & n19407 ) | ( ~x20 & n19407 ) ;
  assign n19409 = ( x20 & ~n19405 ) | ( x20 & n19407 ) | ( ~n19405 & n19407 ) ;
  assign n19410 = ( n19408 & ~n19407 ) | ( n19408 & n19409 ) | ( ~n19407 & n19409 ) ;
  assign n19411 = ( n18918 & ~n18988 ) | ( n18918 & n18998 ) | ( ~n18988 & n18998 ) ;
  assign n19415 = ~n4430 & n11085 ;
  assign n19412 = n523 | n11091 ;
  assign n19413 = n3939 | n11081 ;
  assign n19414 = n19412 &  n19413 ;
  assign n19416 = ( n4430 & n19415 ) | ( n4430 & n19414 ) | ( n19415 & n19414 ) ;
  assign n19417 = n601 | n13377 ;
  assign n19418 = n19416 &  n19417 ;
  assign n19419 = x29 &  n19418 ;
  assign n19420 = x29 | n19418 ;
  assign n19421 = ~n19419 & n19420 ;
  assign n19422 = ( n18956 & ~n18949 ) | ( n18956 & n18958 ) | ( ~n18949 & n18958 ) ;
  assign n19430 = ( n678 & ~n333 ) | ( n678 & n792 ) | ( ~n333 & n792 ) ;
  assign n19431 = n333 | n19430 ;
  assign n19432 = n216 | n19431 ;
  assign n19433 = n431 | n19432 ;
  assign n19434 = ( n738 & ~n19433 ) | ( n738 & n4841 ) | ( ~n19433 & n4841 ) ;
  assign n19435 = ( n19434 & ~n738 ) | ( n19434 & 1'b0 ) | ( ~n738 & 1'b0 ) ;
  assign n19436 = ( n2162 & n5597 ) | ( n2162 & n19435 ) | ( n5597 & n19435 ) ;
  assign n19437 = ~n2162 & n19436 ;
  assign n19438 = ( n15764 & n2887 ) | ( n15764 & n19437 ) | ( n2887 & n19437 ) ;
  assign n19439 = ~n2887 & n19438 ;
  assign n19440 = ( n2427 & ~n887 ) | ( n2427 & n19439 ) | ( ~n887 & n19439 ) ;
  assign n19441 = ~n2427 & n19440 ;
  assign n19442 = ( n1427 & ~n2191 ) | ( n1427 & n19441 ) | ( ~n2191 & n19441 ) ;
  assign n19443 = ( n72 & ~n1427 ) | ( n72 & n19442 ) | ( ~n1427 & n19442 ) ;
  assign n19444 = ~n72 & n19443 ;
  assign n19445 = ( n233 & ~n672 ) | ( n233 & n19444 ) | ( ~n672 & n19444 ) ;
  assign n19446 = ( n162 & ~n233 ) | ( n162 & n19445 ) | ( ~n233 & n19445 ) ;
  assign n19447 = ~n162 & n19446 ;
  assign n19448 = ( n571 & n3680 ) | ( n571 & n19447 ) | ( n3680 & n19447 ) ;
  assign n19449 = ~n571 & n19448 ;
  assign n19450 = ( n627 & ~n117 ) | ( n627 & n19449 ) | ( ~n117 & n19449 ) ;
  assign n19451 = ~n627 & n19450 ;
  assign n19423 = n3644 | n12997 ;
  assign n19424 = ( n3652 & ~n11098 ) | ( n3652 & 1'b0 ) | ( ~n11098 & 1'b0 ) ;
  assign n19425 = ( n3657 & ~n11095 ) | ( n3657 & 1'b0 ) | ( ~n11095 & 1'b0 ) ;
  assign n19426 = n19424 | n19425 ;
  assign n19427 = ~n3653 & n11093 ;
  assign n19428 = ( n3653 & ~n19426 ) | ( n3653 & n19427 ) | ( ~n19426 & n19427 ) ;
  assign n19429 = n19423 &  n19428 ;
  assign n19452 = ( n18949 & ~n19451 ) | ( n18949 & n19429 ) | ( ~n19451 & n19429 ) ;
  assign n19453 = ( n18949 & ~n19429 ) | ( n18949 & n19451 ) | ( ~n19429 & n19451 ) ;
  assign n19454 = ( n19452 & ~n18949 ) | ( n19452 & n19453 ) | ( ~n18949 & n19453 ) ;
  assign n19455 = ~x29 & n18971 ;
  assign n19456 = ( x29 & ~n18971 ) | ( x29 & n18963 ) | ( ~n18971 & n18963 ) ;
  assign n19457 = ( n19455 & ~n18962 ) | ( n19455 & n19456 ) | ( ~n18962 & n19456 ) ;
  assign n19458 = ( n19422 & n19454 ) | ( n19422 & n19457 ) | ( n19454 & n19457 ) ;
  assign n19459 = ( n19454 & ~n19422 ) | ( n19454 & n19457 ) | ( ~n19422 & n19457 ) ;
  assign n19460 = ( n19422 & ~n19458 ) | ( n19422 & n19459 ) | ( ~n19458 & n19459 ) ;
  assign n19464 = ~n4962 & n14071 ;
  assign n19461 = n4482 | n11078 ;
  assign n19462 = n4495 | n13836 ;
  assign n19463 = n19461 &  n19462 ;
  assign n19465 = ( n4962 & n19464 ) | ( n4962 & n19463 ) | ( n19464 & n19463 ) ;
  assign n19466 = n4478 | n14079 ;
  assign n19467 = n19465 &  n19466 ;
  assign n19468 = x26 &  n19467 ;
  assign n19469 = x26 | n19467 ;
  assign n19470 = ~n19468 & n19469 ;
  assign n19471 = ( n19421 & ~n19460 ) | ( n19421 & n19470 ) | ( ~n19460 & n19470 ) ;
  assign n19472 = ( n19421 & ~n19470 ) | ( n19421 & n19460 ) | ( ~n19470 & n19460 ) ;
  assign n19473 = ( n19471 & ~n19421 ) | ( n19471 & n19472 ) | ( ~n19421 & n19472 ) ;
  assign n19474 = ( n18975 & ~n18974 ) | ( n18975 & n18985 ) | ( ~n18974 & n18985 ) ;
  assign n19475 = ( n19473 & ~n19474 ) | ( n19473 & 1'b0 ) | ( ~n19474 & 1'b0 ) ;
  assign n19476 = ~n19473 & n19474 ;
  assign n19477 = n19475 | n19476 ;
  assign n19481 = ~n5135 & n14803 ;
  assign n19478 = n5010 | n14355 ;
  assign n19479 = ~n5067 & n14553 ;
  assign n19480 = ( n19478 & ~n19479 ) | ( n19478 & 1'b0 ) | ( ~n19479 & 1'b0 ) ;
  assign n19482 = ( n5135 & n19481 ) | ( n5135 & n19480 ) | ( n19481 & n19480 ) ;
  assign n19483 = ~n5012 & n15310 ;
  assign n19484 = ( n19482 & ~n19483 ) | ( n19482 & 1'b0 ) | ( ~n19483 & 1'b0 ) ;
  assign n19485 = ( x23 & ~n19477 ) | ( x23 & n19484 ) | ( ~n19477 & n19484 ) ;
  assign n19486 = ( n19477 & ~x23 ) | ( n19477 & n19484 ) | ( ~x23 & n19484 ) ;
  assign n19487 = ( n19485 & ~n19484 ) | ( n19485 & n19486 ) | ( ~n19484 & n19486 ) ;
  assign n19488 = ( n19410 & n19411 ) | ( n19410 & n19487 ) | ( n19411 & n19487 ) ;
  assign n19489 = ( n19411 & ~n19410 ) | ( n19411 & n19487 ) | ( ~n19410 & n19487 ) ;
  assign n19490 = ( n19410 & ~n19488 ) | ( n19410 & n19489 ) | ( ~n19488 & n19489 ) ;
  assign n19491 = ( n18917 & ~n19014 ) | ( n18917 & n19037 ) | ( ~n19014 & n19037 ) ;
  assign n19492 = ( n19401 & ~n19490 ) | ( n19401 & n19491 ) | ( ~n19490 & n19491 ) ;
  assign n19493 = ( n19401 & ~n19491 ) | ( n19401 & n19490 ) | ( ~n19491 & n19490 ) ;
  assign n19494 = ( ~n19401 & n19492 ) | ( ~n19401 & n19493 ) | ( n19492 & n19493 ) ;
  assign n19498 = ~n8764 & n19494 ;
  assign n19499 = ( n8764 & ~n19497 ) | ( n8764 & n19498 ) | ( ~n19497 & n19498 ) ;
  assign n19500 = ( n19040 & ~n19055 ) | ( n19040 & n19494 ) | ( ~n19055 & n19494 ) ;
  assign n19501 = ( n19040 & ~n19494 ) | ( n19040 & n19055 ) | ( ~n19494 & n19055 ) ;
  assign n19502 = ( n19500 & ~n19040 ) | ( n19500 & n19501 ) | ( ~n19040 & n19501 ) ;
  assign n19503 = ( n8107 & ~n19502 ) | ( n8107 & n19499 ) | ( ~n19502 & n19499 ) ;
  assign n19504 = ~n8107 & n19503 ;
  assign n19505 = ( x8 & ~n19499 ) | ( x8 & n19504 ) | ( ~n19499 & n19504 ) ;
  assign n19506 = ( n19499 & ~x8 ) | ( n19499 & n19504 ) | ( ~x8 & n19504 ) ;
  assign n19507 = ( n19505 & ~n19504 ) | ( n19505 & n19506 ) | ( ~n19504 & n19506 ) ;
  assign n19514 = n19040 | n8764 ;
  assign n19511 = ( n8105 & ~n19043 ) | ( n8105 & 1'b0 ) | ( ~n19043 & 1'b0 ) ;
  assign n19512 = ~n8429 & n19047 ;
  assign n19513 = n19511 | n19512 ;
  assign n19515 = ( n19514 & ~n8764 ) | ( n19514 & n19513 ) | ( ~n8764 & n19513 ) ;
  assign n19516 = ( n19056 & ~n8107 ) | ( n19056 & n19515 ) | ( ~n8107 & n19515 ) ;
  assign n19517 = n8107 | n19516 ;
  assign n19518 = ( x8 & ~n19515 ) | ( x8 & n19517 ) | ( ~n19515 & n19517 ) ;
  assign n19519 = ( n19515 & ~x8 ) | ( n19515 & n19517 ) | ( ~x8 & n19517 ) ;
  assign n19520 = ( n19518 & ~n19517 ) | ( n19518 & n19519 ) | ( ~n19517 & n19519 ) ;
  assign n19508 = ( n19101 & ~n19391 ) | ( n19101 & n19103 ) | ( ~n19391 & n19103 ) ;
  assign n19509 = ( n19103 & ~n19101 ) | ( n19103 & n19391 ) | ( ~n19101 & n19391 ) ;
  assign n19510 = ( n19508 & ~n19103 ) | ( n19508 & n19509 ) | ( ~n19103 & n19509 ) ;
  assign n19521 = ( n19115 & ~n19113 ) | ( n19115 & n19390 ) | ( ~n19113 & n19390 ) ;
  assign n19522 = ( n19113 & ~n19390 ) | ( n19113 & n19115 ) | ( ~n19390 & n19115 ) ;
  assign n19523 = ( n19521 & ~n19115 ) | ( n19521 & n19522 ) | ( ~n19115 & n19522 ) ;
  assign n19527 = n19047 | n8764 ;
  assign n19524 = ( n8105 & ~n18712 ) | ( n8105 & 1'b0 ) | ( ~n18712 & 1'b0 ) ;
  assign n19525 = n8429 | n19043 ;
  assign n19526 = ~n19524 & n19525 ;
  assign n19528 = ( n8764 & ~n19527 ) | ( n8764 & n19526 ) | ( ~n19527 & n19526 ) ;
  assign n19529 = ( n8107 & n19068 ) | ( n8107 & n19528 ) | ( n19068 & n19528 ) ;
  assign n19530 = ~n8107 & n19529 ;
  assign n19532 = ( x8 & n19528 ) | ( x8 & n19530 ) | ( n19528 & n19530 ) ;
  assign n19531 = ( x8 & ~n19530 ) | ( x8 & n19528 ) | ( ~n19530 & n19528 ) ;
  assign n19533 = ( n19530 & ~n19532 ) | ( n19530 & n19531 ) | ( ~n19532 & n19531 ) ;
  assign n19537 = ~n8764 & n19043 ;
  assign n19534 = ( n8105 & ~n18589 ) | ( n8105 & 1'b0 ) | ( ~n18589 & 1'b0 ) ;
  assign n19535 = n8429 | n18712 ;
  assign n19536 = ~n19534 & n19535 ;
  assign n19538 = ( n8764 & n19537 ) | ( n8764 & n19536 ) | ( n19537 & n19536 ) ;
  assign n19539 = n8107 | n19083 ;
  assign n19540 = n19538 &  n19539 ;
  assign n19541 = x8 &  n19540 ;
  assign n19542 = x8 | n19540 ;
  assign n19543 = ~n19541 & n19542 ;
  assign n19544 = ( n19118 & ~n19128 ) | ( n19118 & n19389 ) | ( ~n19128 & n19389 ) ;
  assign n19545 = ( n19128 & ~n19390 ) | ( n19128 & n19544 ) | ( ~n19390 & n19544 ) ;
  assign n19549 = ~n8764 & n18712 ;
  assign n19546 = ( n8105 & ~n18456 ) | ( n8105 & 1'b0 ) | ( ~n18456 & 1'b0 ) ;
  assign n19547 = n8429 | n18589 ;
  assign n19548 = ~n19546 & n19547 ;
  assign n19550 = ( n8764 & n19549 ) | ( n8764 & n19548 ) | ( n19549 & n19548 ) ;
  assign n19551 = n8107 | n18720 ;
  assign n19552 = n19550 &  n19551 ;
  assign n19553 = x8 &  n19552 ;
  assign n19554 = x8 | n19552 ;
  assign n19555 = ~n19553 & n19554 ;
  assign n19556 = ( n19131 & ~n19141 ) | ( n19131 & n19388 ) | ( ~n19141 & n19388 ) ;
  assign n19557 = ( n19141 & ~n19389 ) | ( n19141 & n19556 ) | ( ~n19389 & n19556 ) ;
  assign n19564 = ~n8764 & n18589 ;
  assign n19561 = ( n8105 & ~n17783 ) | ( n8105 & 1'b0 ) | ( ~n17783 & 1'b0 ) ;
  assign n19562 = n8429 | n18456 ;
  assign n19563 = ~n19561 & n19562 ;
  assign n19565 = ( n8764 & n19564 ) | ( n8764 & n19563 ) | ( n19564 & n19563 ) ;
  assign n19566 = ( n18597 & ~n8107 ) | ( n18597 & n19565 ) | ( ~n8107 & n19565 ) ;
  assign n19567 = ~n18597 & n19566 ;
  assign n19569 = ( x8 & n19565 ) | ( x8 & n19567 ) | ( n19565 & n19567 ) ;
  assign n19568 = ( x8 & ~n19567 ) | ( x8 & n19565 ) | ( ~n19567 & n19565 ) ;
  assign n19570 = ( n19567 & ~n19569 ) | ( n19567 & n19568 ) | ( ~n19569 & n19568 ) ;
  assign n19558 = ( n19153 & ~n19151 ) | ( n19153 & n19387 ) | ( ~n19151 & n19387 ) ;
  assign n19559 = ( n19151 & ~n19387 ) | ( n19151 & n19153 ) | ( ~n19387 & n19153 ) ;
  assign n19560 = ( n19558 & ~n19153 ) | ( n19558 & n19559 ) | ( ~n19153 & n19559 ) ;
  assign n19571 = ( n19165 & ~n19163 ) | ( n19165 & n19386 ) | ( ~n19163 & n19386 ) ;
  assign n19572 = ( n19163 & ~n19386 ) | ( n19163 & n19165 ) | ( ~n19386 & n19165 ) ;
  assign n19573 = ( n19571 & ~n19165 ) | ( n19571 & n19572 ) | ( ~n19165 & n19572 ) ;
  assign n19577 = ~n8764 & n18456 ;
  assign n19574 = ( n8105 & ~n17791 ) | ( n8105 & 1'b0 ) | ( ~n17791 & 1'b0 ) ;
  assign n19575 = n8429 | n17783 ;
  assign n19576 = ~n19574 & n19575 ;
  assign n19578 = ( n8764 & n19577 ) | ( n8764 & n19576 ) | ( n19577 & n19576 ) ;
  assign n19579 = ( n18464 & ~n8107 ) | ( n18464 & n19578 ) | ( ~n8107 & n19578 ) ;
  assign n19580 = ~n18464 & n19579 ;
  assign n19581 = ( x8 & ~n19578 ) | ( x8 & n19580 ) | ( ~n19578 & n19580 ) ;
  assign n19582 = ( n19578 & ~x8 ) | ( n19578 & n19580 ) | ( ~x8 & n19580 ) ;
  assign n19583 = ( n19581 & ~n19580 ) | ( n19581 & n19582 ) | ( ~n19580 & n19582 ) ;
  assign n19584 = ( n19177 & ~n19175 ) | ( n19177 & n19385 ) | ( ~n19175 & n19385 ) ;
  assign n19585 = ( n19175 & ~n19385 ) | ( n19175 & n19177 ) | ( ~n19385 & n19177 ) ;
  assign n19586 = ( n19584 & ~n19177 ) | ( n19584 & n19585 ) | ( ~n19177 & n19585 ) ;
  assign n19590 = ~n8764 & n17783 ;
  assign n19587 = ( n8105 & ~n17787 ) | ( n8105 & 1'b0 ) | ( ~n17787 & 1'b0 ) ;
  assign n19588 = n8429 | n17791 ;
  assign n19589 = ~n19587 & n19588 ;
  assign n19591 = ( n8764 & n19590 ) | ( n8764 & n19589 ) | ( n19590 & n19589 ) ;
  assign n19592 = ( n17799 & ~n8107 ) | ( n17799 & n19591 ) | ( ~n8107 & n19591 ) ;
  assign n19593 = ~n17799 & n19592 ;
  assign n19595 = ( x8 & n19591 ) | ( x8 & n19593 ) | ( n19591 & n19593 ) ;
  assign n19594 = ( x8 & ~n19593 ) | ( x8 & n19591 ) | ( ~n19593 & n19591 ) ;
  assign n19596 = ( n19593 & ~n19595 ) | ( n19593 & n19594 ) | ( ~n19595 & n19594 ) ;
  assign n19600 = ~n8764 & n17791 ;
  assign n19597 = ( n8105 & ~n17405 ) | ( n8105 & 1'b0 ) | ( ~n17405 & 1'b0 ) ;
  assign n19598 = n8429 | n17787 ;
  assign n19599 = ~n19597 & n19598 ;
  assign n19601 = ( n8764 & n19600 ) | ( n8764 & n19599 ) | ( n19600 & n19599 ) ;
  assign n19602 = n8107 | n17811 ;
  assign n19603 = n19601 &  n19602 ;
  assign n19604 = x8 &  n19603 ;
  assign n19605 = x8 | n19603 ;
  assign n19606 = ~n19604 & n19605 ;
  assign n19607 = ( n19180 & ~n19384 ) | ( n19180 & n19190 ) | ( ~n19384 & n19190 ) ;
  assign n19608 = ( n19385 & ~n19190 ) | ( n19385 & n19607 ) | ( ~n19190 & n19607 ) ;
  assign n19609 = ( n8105 & ~n17263 ) | ( n8105 & 1'b0 ) | ( ~n17263 & 1'b0 ) ;
  assign n19610 = n8429 | n17405 ;
  assign n19611 = ~n19609 & n19610 ;
  assign n19612 = ~n8764 & n17787 ;
  assign n19613 = ( n8764 & n19611 ) | ( n8764 & n19612 ) | ( n19611 & n19612 ) ;
  assign n19614 = n8107 | n17826 ;
  assign n19615 = n19613 &  n19614 ;
  assign n19616 = x8 &  n19615 ;
  assign n19617 = x8 | n19615 ;
  assign n19618 = ~n19616 & n19617 ;
  assign n19619 = ( n19193 & ~n19203 ) | ( n19193 & n19383 ) | ( ~n19203 & n19383 ) ;
  assign n19620 = ( n19203 & ~n19384 ) | ( n19203 & n19619 ) | ( ~n19384 & n19619 ) ;
  assign n19624 = ~n8764 & n17405 ;
  assign n19621 = n8105 &  n17107 ;
  assign n19622 = n8429 | n17263 ;
  assign n19623 = ~n19621 & n19622 ;
  assign n19625 = ( n8764 & n19624 ) | ( n8764 & n19623 ) | ( n19624 & n19623 ) ;
  assign n19626 = n8107 | n17413 ;
  assign n19627 = n19625 &  n19626 ;
  assign n19628 = x8 &  n19627 ;
  assign n19629 = x8 | n19627 ;
  assign n19630 = ~n19628 & n19629 ;
  assign n19631 = ( n19206 & ~n19216 ) | ( n19206 & n19382 ) | ( ~n19216 & n19382 ) ;
  assign n19632 = ( n19216 & ~n19383 ) | ( n19216 & n19631 ) | ( ~n19383 & n19631 ) ;
  assign n19636 = ( n8105 & ~n16589 ) | ( n8105 & 1'b0 ) | ( ~n16589 & 1'b0 ) ;
  assign n19637 = ~n8429 & n17107 ;
  assign n19638 = n19636 | n19637 ;
  assign n19639 = ~n8764 & n17263 ;
  assign n19640 = ( n8764 & ~n19638 ) | ( n8764 & n19639 ) | ( ~n19638 & n19639 ) ;
  assign n19641 = ( n8107 & ~n19640 ) | ( n8107 & n17271 ) | ( ~n19640 & n17271 ) ;
  assign n19642 = ( n17271 & ~n19641 ) | ( n17271 & 1'b0 ) | ( ~n19641 & 1'b0 ) ;
  assign n19644 = ( x8 & n19640 ) | ( x8 & n19642 ) | ( n19640 & n19642 ) ;
  assign n19643 = ( x8 & ~n19642 ) | ( x8 & n19640 ) | ( ~n19642 & n19640 ) ;
  assign n19645 = ( n19642 & ~n19644 ) | ( n19642 & n19643 ) | ( ~n19644 & n19643 ) ;
  assign n19633 = ( n19228 & ~n19226 ) | ( n19228 & n19381 ) | ( ~n19226 & n19381 ) ;
  assign n19634 = ( n19226 & ~n19381 ) | ( n19226 & n19228 ) | ( ~n19381 & n19228 ) ;
  assign n19635 = ( n19633 & ~n19228 ) | ( n19633 & n19634 ) | ( ~n19228 & n19634 ) ;
  assign n19646 = ( n19240 & ~n19238 ) | ( n19240 & n19380 ) | ( ~n19238 & n19380 ) ;
  assign n19647 = ( n19238 & ~n19380 ) | ( n19238 & n19240 ) | ( ~n19380 & n19240 ) ;
  assign n19648 = ( n19646 & ~n19240 ) | ( n19646 & n19647 ) | ( ~n19240 & n19647 ) ;
  assign n19652 = n17107 | n8764 ;
  assign n19649 = ( n8105 & ~n16595 ) | ( n8105 & 1'b0 ) | ( ~n16595 & 1'b0 ) ;
  assign n19650 = n8429 | n16589 ;
  assign n19651 = ~n19649 & n19650 ;
  assign n19653 = ( n8764 & ~n19652 ) | ( n8764 & n19651 ) | ( ~n19652 & n19651 ) ;
  assign n19654 = ( n8107 & ~n19653 ) | ( n8107 & n17115 ) | ( ~n19653 & n17115 ) ;
  assign n19655 = ( n17115 & ~n19654 ) | ( n17115 & 1'b0 ) | ( ~n19654 & 1'b0 ) ;
  assign n19656 = ( x8 & ~n19653 ) | ( x8 & n19655 ) | ( ~n19653 & n19655 ) ;
  assign n19657 = ( n19653 & ~x8 ) | ( n19653 & n19655 ) | ( ~x8 & n19655 ) ;
  assign n19658 = ( n19656 & ~n19655 ) | ( n19656 & n19657 ) | ( ~n19655 & n19657 ) ;
  assign n19659 = ( n19252 & ~n19250 ) | ( n19252 & n19379 ) | ( ~n19250 & n19379 ) ;
  assign n19660 = ( n19250 & ~n19379 ) | ( n19250 & n19252 ) | ( ~n19379 & n19252 ) ;
  assign n19661 = ( n19659 & ~n19252 ) | ( n19659 & n19660 ) | ( ~n19252 & n19660 ) ;
  assign n19665 = ~n8764 & n16589 ;
  assign n19662 = ( n8105 & ~n16591 ) | ( n8105 & 1'b0 ) | ( ~n16591 & 1'b0 ) ;
  assign n19663 = n8429 | n16595 ;
  assign n19664 = ~n19662 & n19663 ;
  assign n19666 = ( n8764 & n19665 ) | ( n8764 & n19664 ) | ( n19665 & n19664 ) ;
  assign n19667 = ( n16604 & ~n8107 ) | ( n16604 & n19666 ) | ( ~n8107 & n19666 ) ;
  assign n19668 = ~n16604 & n19667 ;
  assign n19670 = ( x8 & n19666 ) | ( x8 & n19668 ) | ( n19666 & n19668 ) ;
  assign n19669 = ( x8 & ~n19668 ) | ( x8 & n19666 ) | ( ~n19668 & n19666 ) ;
  assign n19671 = ( n19668 & ~n19670 ) | ( n19668 & n19669 ) | ( ~n19670 & n19669 ) ;
  assign n19675 = ~n8764 & n16595 ;
  assign n19672 = ( n8105 & ~n16091 ) | ( n8105 & 1'b0 ) | ( ~n16091 & 1'b0 ) ;
  assign n19673 = n8429 | n16591 ;
  assign n19674 = ~n19672 & n19673 ;
  assign n19676 = ( n8764 & n19675 ) | ( n8764 & n19674 ) | ( n19675 & n19674 ) ;
  assign n19677 = n8107 | n16616 ;
  assign n19678 = n19676 &  n19677 ;
  assign n19679 = x8 &  n19678 ;
  assign n19680 = x8 | n19678 ;
  assign n19681 = ~n19679 & n19680 ;
  assign n19682 = ( n19255 & ~n19378 ) | ( n19255 & n19265 ) | ( ~n19378 & n19265 ) ;
  assign n19683 = ( n19379 & ~n19265 ) | ( n19379 & n19682 ) | ( ~n19265 & n19682 ) ;
  assign n19687 = ~n8764 & n16591 ;
  assign n19684 = ( n8105 & ~n15897 ) | ( n8105 & 1'b0 ) | ( ~n15897 & 1'b0 ) ;
  assign n19685 = n8429 | n16091 ;
  assign n19686 = ~n19684 & n19685 ;
  assign n19688 = ( n8764 & n19687 ) | ( n8764 & n19686 ) | ( n19687 & n19686 ) ;
  assign n19689 = n8107 | n16631 ;
  assign n19690 = n19688 &  n19689 ;
  assign n19691 = x8 &  n19690 ;
  assign n19692 = x8 | n19690 ;
  assign n19693 = ~n19691 & n19692 ;
  assign n19694 = ( n19268 & ~n19278 ) | ( n19268 & n19377 ) | ( ~n19278 & n19377 ) ;
  assign n19695 = ( n19278 & ~n19378 ) | ( n19278 & n19694 ) | ( ~n19378 & n19694 ) ;
  assign n19699 = ~n8764 & n16091 ;
  assign n19696 = ( n8105 & ~n15700 ) | ( n8105 & 1'b0 ) | ( ~n15700 & 1'b0 ) ;
  assign n19697 = n8429 | n15897 ;
  assign n19698 = ~n19696 & n19697 ;
  assign n19700 = ( n8764 & n19699 ) | ( n8764 & n19698 ) | ( n19699 & n19698 ) ;
  assign n19701 = n8107 | n16094 ;
  assign n19702 = n19700 &  n19701 ;
  assign n19703 = x8 &  n19702 ;
  assign n19704 = x8 | n19702 ;
  assign n19705 = ~n19703 & n19704 ;
  assign n19706 = ( n19281 & ~n19291 ) | ( n19281 & n19376 ) | ( ~n19291 & n19376 ) ;
  assign n19707 = ( n19291 & ~n19377 ) | ( n19291 & n19706 ) | ( ~n19377 & n19706 ) ;
  assign n19714 = ~n8764 & n15897 ;
  assign n19711 = ( n8105 & ~n15320 ) | ( n8105 & 1'b0 ) | ( ~n15320 & 1'b0 ) ;
  assign n19712 = n8429 | n15700 ;
  assign n19713 = ~n19711 & n19712 ;
  assign n19715 = ( n8764 & n19714 ) | ( n8764 & n19713 ) | ( n19714 & n19713 ) ;
  assign n19716 = ( n15900 & ~n8107 ) | ( n15900 & n19715 ) | ( ~n8107 & n19715 ) ;
  assign n19717 = ~n15900 & n19716 ;
  assign n19718 = ( x8 & ~n19715 ) | ( x8 & n19717 ) | ( ~n19715 & n19717 ) ;
  assign n19719 = ( n19715 & ~x8 ) | ( n19715 & n19717 ) | ( ~x8 & n19717 ) ;
  assign n19720 = ( n19718 & ~n19717 ) | ( n19718 & n19719 ) | ( ~n19717 & n19719 ) ;
  assign n19708 = ( n19303 & ~n19301 ) | ( n19303 & n19375 ) | ( ~n19301 & n19375 ) ;
  assign n19709 = ( n19301 & ~n19375 ) | ( n19301 & n19303 ) | ( ~n19375 & n19303 ) ;
  assign n19710 = ( n19708 & ~n19303 ) | ( n19708 & n19709 ) | ( ~n19303 & n19709 ) ;
  assign n19721 = ( n19316 & ~n19306 ) | ( n19316 & n19374 ) | ( ~n19306 & n19374 ) ;
  assign n19722 = ( n19306 & ~n19374 ) | ( n19306 & n19316 ) | ( ~n19374 & n19316 ) ;
  assign n19723 = ( n19721 & ~n19316 ) | ( n19721 & n19722 ) | ( ~n19316 & n19722 ) ;
  assign n19727 = ~n8764 & n15700 ;
  assign n19724 = ( n8105 & ~n15325 ) | ( n8105 & 1'b0 ) | ( ~n15325 & 1'b0 ) ;
  assign n19725 = n8429 | n15320 ;
  assign n19726 = ~n19724 & n19725 ;
  assign n19728 = ( n8764 & n19727 ) | ( n8764 & n19726 ) | ( n19727 & n19726 ) ;
  assign n19729 = ( n15708 & ~n8107 ) | ( n15708 & n19728 ) | ( ~n8107 & n19728 ) ;
  assign n19730 = ~n15708 & n19729 ;
  assign n19732 = ( x8 & n19728 ) | ( x8 & n19730 ) | ( n19728 & n19730 ) ;
  assign n19731 = ( x8 & ~n19730 ) | ( x8 & n19728 ) | ( ~n19730 & n19728 ) ;
  assign n19733 = ( n19730 & ~n19732 ) | ( n19730 & n19731 ) | ( ~n19732 & n19731 ) ;
  assign n19734 = ( n19326 & ~n19373 ) | ( n19326 & n19331 ) | ( ~n19373 & n19331 ) ;
  assign n19735 = ( n19331 & ~n19326 ) | ( n19331 & n19373 ) | ( ~n19326 & n19373 ) ;
  assign n19736 = ( n19734 & ~n19331 ) | ( n19734 & n19735 ) | ( ~n19331 & n19735 ) ;
  assign n19740 = ~n8764 & n15320 ;
  assign n19737 = ( n8105 & ~n15322 ) | ( n8105 & 1'b0 ) | ( ~n15322 & 1'b0 ) ;
  assign n19738 = n8429 | n15325 ;
  assign n19739 = ~n19737 & n19738 ;
  assign n19741 = ( n8764 & n19740 ) | ( n8764 & n19739 ) | ( n19740 & n19739 ) ;
  assign n19742 = ( n15334 & ~n8107 ) | ( n15334 & n19741 ) | ( ~n8107 & n19741 ) ;
  assign n19743 = ~n15334 & n19742 ;
  assign n19744 = ( x8 & ~n19741 ) | ( x8 & n19743 ) | ( ~n19741 & n19743 ) ;
  assign n19745 = ( n19741 & ~x8 ) | ( n19741 & n19743 ) | ( ~x8 & n19743 ) ;
  assign n19746 = ( n19744 & ~n19743 ) | ( n19744 & n19745 ) | ( ~n19743 & n19745 ) ;
  assign n19750 = ~n8764 & n15325 ;
  assign n19747 = n8105 &  n14745 ;
  assign n19748 = n8429 | n15322 ;
  assign n19749 = ~n19747 & n19748 ;
  assign n19751 = ( n8764 & n19750 ) | ( n8764 & n19749 ) | ( n19750 & n19749 ) ;
  assign n19752 = n8107 | n15346 ;
  assign n19753 = n19751 &  n19752 ;
  assign n19754 = x8 &  n19753 ;
  assign n19755 = x8 | n19753 ;
  assign n19756 = ~n19754 & n19755 ;
  assign n19757 = ( n19345 & ~n19335 ) | ( n19345 & n19372 ) | ( ~n19335 & n19372 ) ;
  assign n19758 = ( n19373 & ~n19345 ) | ( n19373 & n19757 ) | ( ~n19345 & n19757 ) ;
  assign n19760 = ( n18279 & n19361 ) | ( n18279 & n19371 ) | ( n19361 & n19371 ) ;
  assign n19759 = ( n18279 & ~n19361 ) | ( n18279 & n19371 ) | ( ~n19361 & n19371 ) ;
  assign n19761 = ( n19361 & ~n19760 ) | ( n19361 & n19759 ) | ( ~n19760 & n19759 ) ;
  assign n19762 = ( n8105 & ~n14528 ) | ( n8105 & 1'b0 ) | ( ~n14528 & 1'b0 ) ;
  assign n19763 = ~n8429 & n14745 ;
  assign n19764 = n19762 | n19763 ;
  assign n19765 = ~n8764 & n15322 ;
  assign n19766 = ( n8764 & ~n19764 ) | ( n8764 & n19765 ) | ( ~n19764 & n19765 ) ;
  assign n19767 = ( n8107 & ~n19766 ) | ( n8107 & n15361 ) | ( ~n19766 & n15361 ) ;
  assign n19768 = ( n15361 & ~n19767 ) | ( n15361 & 1'b0 ) | ( ~n19767 & 1'b0 ) ;
  assign n19769 = ( x8 & ~n19766 ) | ( x8 & n19768 ) | ( ~n19766 & n19768 ) ;
  assign n19770 = ( n19766 & ~x8 ) | ( n19766 & n19768 ) | ( ~x8 & n19768 ) ;
  assign n19771 = ( n19769 & ~n19768 ) | ( n19769 & n19770 ) | ( ~n19768 & n19770 ) ;
  assign n19775 = n14745 | n8764 ;
  assign n19772 = ( n8105 & ~n14261 ) | ( n8105 & 1'b0 ) | ( ~n14261 & 1'b0 ) ;
  assign n19773 = n8429 | n14528 ;
  assign n19774 = ~n19772 & n19773 ;
  assign n19776 = ( n8764 & ~n19775 ) | ( n8764 & n19774 ) | ( ~n19775 & n19774 ) ;
  assign n19777 = ~n8107 & n14749 ;
  assign n19778 = ( n19776 & ~n19777 ) | ( n19776 & 1'b0 ) | ( ~n19777 & 1'b0 ) ;
  assign n19779 = x8 &  n19778 ;
  assign n19780 = x8 | n19778 ;
  assign n19781 = ~n19779 & n19780 ;
  assign n19782 = ( x11 & n19346 ) | ( x11 & n19351 ) | ( n19346 & n19351 ) ;
  assign n19783 = ~n19346 & n19782 ;
  assign n19784 = ( n19358 & ~x11 ) | ( n19358 & n19783 ) | ( ~x11 & n19783 ) ;
  assign n19785 = ( x11 & ~n19358 ) | ( x11 & n19783 ) | ( ~n19358 & n19783 ) ;
  assign n19786 = ( n19784 & ~n19783 ) | ( n19784 & n19785 ) | ( ~n19783 & n19785 ) ;
  assign n19787 = x11 &  n19346 ;
  assign n19788 = n19351 &  n19787 ;
  assign n19789 = n19351 | n19787 ;
  assign n19790 = ~n19788 & n19789 ;
  assign n19817 = ( n8105 & ~n13785 ) | ( n8105 & 1'b0 ) | ( ~n13785 & 1'b0 ) ;
  assign n19818 = n8429 | n13998 ;
  assign n19819 = ~n19817 & n19818 ;
  assign n19820 = ~n8764 & n14261 ;
  assign n19821 = ( n8764 & n19819 ) | ( n8764 & n19820 ) | ( n19819 & n19820 ) ;
  assign n19822 = n8107 | n14267 ;
  assign n19823 = n19821 &  n19822 ;
  assign n19824 = x8 &  n19823 ;
  assign n19825 = x8 | n19823 ;
  assign n19826 = ~n19824 & n19825 ;
  assign n19801 = ( n8103 & ~n13787 ) | ( n8103 & 1'b0 ) | ( ~n13787 & 1'b0 ) ;
  assign n19805 = n13790 | n8107 ;
  assign n19802 = n8429 | n13787 ;
  assign n19803 = n8764 | n13785 ;
  assign n19804 = n19802 &  n19803 ;
  assign n19806 = ( n8107 & ~n19805 ) | ( n8107 & n19804 ) | ( ~n19805 & n19804 ) ;
  assign n19812 = ~n8107 & n14001 ;
  assign n19810 = ~n8764 & n13998 ;
  assign n19807 = ( n8105 & ~n13787 ) | ( n8105 & 1'b0 ) | ( ~n13787 & 1'b0 ) ;
  assign n19808 = n8429 | n13785 ;
  assign n19809 = ~n19807 & n19808 ;
  assign n19811 = ( n8764 & n19810 ) | ( n8764 & n19809 ) | ( n19810 & n19809 ) ;
  assign n19813 = ( n8107 & n19812 ) | ( n8107 & n19811 ) | ( n19812 & n19811 ) ;
  assign n19814 = ( n19801 & n19806 ) | ( n19801 & n19813 ) | ( n19806 & n19813 ) ;
  assign n19815 = ( x8 & ~n19814 ) | ( x8 & n19801 ) | ( ~n19814 & n19801 ) ;
  assign n19816 = ( x8 & ~n19815 ) | ( x8 & 1'b0 ) | ( ~n19815 & 1'b0 ) ;
  assign n19827 = ( n19346 & ~n19826 ) | ( n19346 & n19816 ) | ( ~n19826 & n19816 ) ;
  assign n19794 = ~n8764 & n14528 ;
  assign n19791 = ( n8105 & ~n13998 ) | ( n8105 & 1'b0 ) | ( ~n13998 & 1'b0 ) ;
  assign n19792 = n8429 | n14261 ;
  assign n19793 = ~n19791 & n19792 ;
  assign n19795 = ( n8764 & n19794 ) | ( n8764 & n19793 ) | ( n19794 & n19793 ) ;
  assign n19796 = ( n14532 & ~n8107 ) | ( n14532 & n19795 ) | ( ~n8107 & n19795 ) ;
  assign n19797 = ~n14532 & n19796 ;
  assign n19798 = ( x8 & ~n19795 ) | ( x8 & n19797 ) | ( ~n19795 & n19797 ) ;
  assign n19799 = ( n19795 & ~x8 ) | ( n19795 & n19797 ) | ( ~x8 & n19797 ) ;
  assign n19800 = ( n19798 & ~n19797 ) | ( n19798 & n19799 ) | ( ~n19797 & n19799 ) ;
  assign n19828 = ( n19790 & ~n19827 ) | ( n19790 & n19800 ) | ( ~n19827 & n19800 ) ;
  assign n19829 = ( n19781 & n19786 ) | ( n19781 & n19828 ) | ( n19786 & n19828 ) ;
  assign n19830 = ( n19761 & n19771 ) | ( n19761 & n19829 ) | ( n19771 & n19829 ) ;
  assign n19831 = ( n19756 & ~n19758 ) | ( n19756 & n19830 ) | ( ~n19758 & n19830 ) ;
  assign n19832 = ( n19736 & n19746 ) | ( n19736 & n19831 ) | ( n19746 & n19831 ) ;
  assign n19833 = ( n19723 & n19733 ) | ( n19723 & n19832 ) | ( n19733 & n19832 ) ;
  assign n19834 = ( n19720 & ~n19710 ) | ( n19720 & n19833 ) | ( ~n19710 & n19833 ) ;
  assign n19835 = ( n19705 & n19707 ) | ( n19705 & n19834 ) | ( n19707 & n19834 ) ;
  assign n19836 = ( n19693 & n19695 ) | ( n19693 & n19835 ) | ( n19695 & n19835 ) ;
  assign n19837 = ( n19681 & ~n19683 ) | ( n19681 & n19836 ) | ( ~n19683 & n19836 ) ;
  assign n19838 = ( n19661 & n19671 ) | ( n19661 & n19837 ) | ( n19671 & n19837 ) ;
  assign n19839 = ( n19648 & n19658 ) | ( n19648 & n19838 ) | ( n19658 & n19838 ) ;
  assign n19840 = ( n19645 & ~n19635 ) | ( n19645 & n19839 ) | ( ~n19635 & n19839 ) ;
  assign n19841 = ( n19630 & n19632 ) | ( n19630 & n19840 ) | ( n19632 & n19840 ) ;
  assign n19842 = ( n19618 & n19620 ) | ( n19618 & n19841 ) | ( n19620 & n19841 ) ;
  assign n19843 = ( n19606 & ~n19608 ) | ( n19606 & n19842 ) | ( ~n19608 & n19842 ) ;
  assign n19844 = ( n19586 & n19596 ) | ( n19586 & n19843 ) | ( n19596 & n19843 ) ;
  assign n19845 = ( n19573 & n19583 ) | ( n19573 & n19844 ) | ( n19583 & n19844 ) ;
  assign n19846 = ( n19570 & ~n19560 ) | ( n19570 & n19845 ) | ( ~n19560 & n19845 ) ;
  assign n19847 = ( n19555 & n19557 ) | ( n19555 & n19846 ) | ( n19557 & n19846 ) ;
  assign n19848 = ( n19543 & n19545 ) | ( n19543 & n19847 ) | ( n19545 & n19847 ) ;
  assign n19849 = ( n19523 & n19533 ) | ( n19523 & n19848 ) | ( n19533 & n19848 ) ;
  assign n19850 = ( n19520 & ~n19510 ) | ( n19520 & n19849 ) | ( ~n19510 & n19849 ) ;
  assign n19851 = ( n19400 & n19507 ) | ( n19400 & n19850 ) | ( n19507 & n19850 ) ;
  assign n19852 = ( n19076 & ~n19073 ) | ( n19076 & n19393 ) | ( ~n19073 & n19393 ) ;
  assign n19853 = ( n19073 & ~n19393 ) | ( n19073 & n19076 ) | ( ~n19393 & n19076 ) ;
  assign n19854 = ( n19852 & ~n19076 ) | ( n19852 & n19853 ) | ( ~n19076 & n19853 ) ;
  assign n19858 = n14807 | n5135 ;
  assign n19855 = ~n5010 & n14553 ;
  assign n19856 = n5067 | n14803 ;
  assign n19857 = ~n19855 & n19856 ;
  assign n19859 = ( n5135 & ~n19858 ) | ( n5135 & n19857 ) | ( ~n19858 & n19857 ) ;
  assign n19860 = ( n5012 & n15294 ) | ( n5012 & n19859 ) | ( n15294 & n19859 ) ;
  assign n19861 = ~n5012 & n19860 ;
  assign n19862 = ( x23 & ~n19859 ) | ( x23 & n19861 ) | ( ~n19859 & n19861 ) ;
  assign n19863 = ( n19859 & ~x23 ) | ( n19859 & n19861 ) | ( ~x23 & n19861 ) ;
  assign n19864 = ( n19862 & ~n19861 ) | ( n19862 & n19863 ) | ( ~n19861 & n19863 ) ;
  assign n19865 = ( x23 & ~n19484 ) | ( x23 & 1'b0 ) | ( ~n19484 & 1'b0 ) ;
  assign n19866 = ( n19476 & ~x23 ) | ( n19476 & n19484 ) | ( ~x23 & n19484 ) ;
  assign n19867 = ( n19865 & ~n19475 ) | ( n19865 & n19866 ) | ( ~n19475 & n19866 ) ;
  assign n19927 = ( n19422 & ~n19454 ) | ( n19422 & n19457 ) | ( ~n19454 & n19457 ) ;
  assign n19931 = ~n4430 & n11078 ;
  assign n19928 = n523 | n11081 ;
  assign n19929 = n3939 | n11085 ;
  assign n19930 = n19928 &  n19929 ;
  assign n19932 = ( n4430 & n19931 ) | ( n4430 & n19930 ) | ( n19931 & n19930 ) ;
  assign n19933 = n601 | n11206 ;
  assign n19934 = n19932 &  n19933 ;
  assign n19878 = ( n19429 & ~n18949 ) | ( n19429 & n19451 ) | ( ~n18949 & n19451 ) ;
  assign n19886 = n1532 | n5413 ;
  assign n19887 = ( n1133 & n3383 ) | ( n1133 & n19886 ) | ( n3383 & n19886 ) ;
  assign n19888 = ( n3383 & ~n19887 ) | ( n3383 & 1'b0 ) | ( ~n19887 & 1'b0 ) ;
  assign n19889 = ( n2186 & ~n2764 ) | ( n2186 & n19888 ) | ( ~n2764 & n19888 ) ;
  assign n19890 = ~n2186 & n19889 ;
  assign n19891 = ( n1495 & ~n1512 ) | ( n1495 & n19890 ) | ( ~n1512 & n19890 ) ;
  assign n19892 = ~n1495 & n19891 ;
  assign n19893 = ( n126 & ~n2191 ) | ( n126 & n19892 ) | ( ~n2191 & n19892 ) ;
  assign n19894 = ~n126 & n19893 ;
  assign n19895 = ( n234 & ~n671 ) | ( n234 & n19894 ) | ( ~n671 & n19894 ) ;
  assign n19896 = ~n234 & n19895 ;
  assign n19897 = ( n351 & ~n137 ) | ( n351 & n19896 ) | ( ~n137 & n19896 ) ;
  assign n19898 = ~n351 & n19897 ;
  assign n19899 = n1732 | n4371 ;
  assign n19900 = ( n1990 & n3526 ) | ( n1990 & n19899 ) | ( n3526 & n19899 ) ;
  assign n19901 = ( n1990 & ~n19900 ) | ( n1990 & 1'b0 ) | ( ~n19900 & 1'b0 ) ;
  assign n19902 = ( n2609 & ~n19898 ) | ( n2609 & n19901 ) | ( ~n19898 & n19901 ) ;
  assign n19903 = ( n1820 & n19898 ) | ( n1820 & n19902 ) | ( n19898 & n19902 ) ;
  assign n19904 = ~n1820 & n19903 ;
  assign n19905 = ( n1581 & ~n1678 ) | ( n1581 & n19904 ) | ( ~n1678 & n19904 ) ;
  assign n19906 = ~n1581 & n19905 ;
  assign n19907 = ( n193 & ~n1876 ) | ( n193 & n19906 ) | ( ~n1876 & n19906 ) ;
  assign n19908 = ~n193 & n19907 ;
  assign n19909 = ( n167 & ~n676 ) | ( n167 & n19908 ) | ( ~n676 & n19908 ) ;
  assign n19910 = ~n167 & n19909 ;
  assign n19911 = ( n476 & ~n336 ) | ( n476 & n19910 ) | ( ~n336 & n19910 ) ;
  assign n19912 = ~n476 & n19911 ;
  assign n19913 = ( n358 & ~n155 ) | ( n358 & n19912 ) | ( ~n155 & n19912 ) ;
  assign n19914 = ~n358 & n19913 ;
  assign n19915 = n18949 &  n19914 ;
  assign n19916 = n18949 | n19914 ;
  assign n19917 = ~n19915 & n19916 ;
  assign n19918 = ( n5334 & ~n5331 ) | ( n5334 & n5337 ) | ( ~n5331 & n5337 ) ;
  assign n19919 = n5331 | n19918 ;
  assign n19920 = n14800 &  n19919 ;
  assign n19921 = ( x20 & n19917 ) | ( x20 & n19920 ) | ( n19917 & n19920 ) ;
  assign n19922 = ( n19917 & ~x20 ) | ( n19917 & n19920 ) | ( ~x20 & n19920 ) ;
  assign n19923 = ( x20 & ~n19921 ) | ( x20 & n19922 ) | ( ~n19921 & n19922 ) ;
  assign n19879 = n3644 | n12984 ;
  assign n19880 = ( n3652 & ~n11095 ) | ( n3652 & 1'b0 ) | ( ~n11095 & 1'b0 ) ;
  assign n19881 = ( n3657 & ~n11093 ) | ( n3657 & 1'b0 ) | ( ~n11093 & 1'b0 ) ;
  assign n19882 = n19880 | n19881 ;
  assign n19883 = ~n3653 & n11091 ;
  assign n19884 = ( n3653 & ~n19882 ) | ( n3653 & n19883 ) | ( ~n19882 & n19883 ) ;
  assign n19885 = n19879 &  n19884 ;
  assign n19924 = ( n19878 & ~n19923 ) | ( n19878 & n19885 ) | ( ~n19923 & n19885 ) ;
  assign n19925 = ( n19878 & ~n19885 ) | ( n19878 & n19923 ) | ( ~n19885 & n19923 ) ;
  assign n19926 = ( n19924 & ~n19878 ) | ( n19924 & n19925 ) | ( ~n19878 & n19925 ) ;
  assign n19935 = x29 | n19926 ;
  assign n19936 = ~x29 & n19926 ;
  assign n19937 = ( n19935 & ~n19926 ) | ( n19935 & n19936 ) | ( ~n19926 & n19936 ) ;
  assign n19938 = ( n19927 & ~n19934 ) | ( n19927 & n19937 ) | ( ~n19934 & n19937 ) ;
  assign n19939 = ( n19934 & ~n19927 ) | ( n19934 & n19937 ) | ( ~n19927 & n19937 ) ;
  assign n19940 = ( n19938 & ~n19937 ) | ( n19938 & n19939 ) | ( ~n19937 & n19939 ) ;
  assign n19871 = ~n4962 & n14355 ;
  assign n19868 = n4482 | n13836 ;
  assign n19869 = n4495 | n14071 ;
  assign n19870 = n19868 &  n19869 ;
  assign n19872 = ( n4962 & n19871 ) | ( n4962 & n19870 ) | ( n19871 & n19870 ) ;
  assign n19873 = ( n4478 & ~n14363 ) | ( n4478 & n19872 ) | ( ~n14363 & n19872 ) ;
  assign n19874 = ~n4478 & n19873 ;
  assign n19875 = ( x26 & ~n19872 ) | ( x26 & n19874 ) | ( ~n19872 & n19874 ) ;
  assign n19876 = ( n19872 & ~x26 ) | ( n19872 & n19874 ) | ( ~x26 & n19874 ) ;
  assign n19877 = ( n19875 & ~n19874 ) | ( n19875 & n19876 ) | ( ~n19874 & n19876 ) ;
  assign n19941 = ( n19471 & ~n19940 ) | ( n19471 & n19877 ) | ( ~n19940 & n19877 ) ;
  assign n19942 = ( n19877 & ~n19471 ) | ( n19877 & n19940 ) | ( ~n19471 & n19940 ) ;
  assign n19943 = ( n19941 & ~n19877 ) | ( n19941 & n19942 ) | ( ~n19877 & n19942 ) ;
  assign n19945 = ( n19864 & n19867 ) | ( n19864 & n19943 ) | ( n19867 & n19943 ) ;
  assign n19944 = ( n19867 & ~n19864 ) | ( n19867 & n19943 ) | ( ~n19864 & n19943 ) ;
  assign n19946 = ( n19864 & ~n19945 ) | ( n19864 & n19944 ) | ( ~n19945 & n19944 ) ;
  assign n19947 = ( n19410 & ~n19411 ) | ( n19410 & n19487 ) | ( ~n19411 & n19487 ) ;
  assign n19948 = ( n19401 & n19490 ) | ( n19401 & n19491 ) | ( n19490 & n19491 ) ;
  assign n19949 = ( n19947 & ~n19946 ) | ( n19947 & n19948 ) | ( ~n19946 & n19948 ) ;
  assign n19950 = ( n19946 & n19947 ) | ( n19946 & n19948 ) | ( n19947 & n19948 ) ;
  assign n19951 = ( ~n19946 & ~n19949 ) | ( ~n19946 & n19950 ) | ( ~n19949 & n19950 ) ;
  assign n19955 = ~n8764 & n19951 ;
  assign n19952 = n8105 &  n19040 ;
  assign n19953 = n8429 | n19494 ;
  assign n19954 = ~n19952 & n19953 ;
  assign n19956 = ( n8764 & n19955 ) | ( n8764 & n19954 ) | ( n19955 & n19954 ) ;
  assign n19957 = ( n19494 & ~n19951 ) | ( n19494 & n19501 ) | ( ~n19951 & n19501 ) ;
  assign n19958 = ( n19494 & ~n19501 ) | ( n19494 & n19951 ) | ( ~n19501 & n19951 ) ;
  assign n19959 = ( n19957 & ~n19494 ) | ( n19957 & n19958 ) | ( ~n19494 & n19958 ) ;
  assign n19960 = ( n8107 & n19956 ) | ( n8107 & n19959 ) | ( n19956 & n19959 ) ;
  assign n19961 = ~n8107 & n19960 ;
  assign n19963 = ( x8 & n19956 ) | ( x8 & n19961 ) | ( n19956 & n19961 ) ;
  assign n19962 = ( x8 & ~n19961 ) | ( x8 & n19956 ) | ( ~n19961 & n19956 ) ;
  assign n19964 = ( n19961 & ~n19963 ) | ( n19961 & n19962 ) | ( ~n19963 & n19962 ) ;
  assign n19965 = ( n19851 & n19854 ) | ( n19851 & n19964 ) | ( n19854 & n19964 ) ;
  assign n19966 = ( n19471 & n19877 ) | ( n19471 & n19940 ) | ( n19877 & n19940 ) ;
  assign n19967 = ( x20 & ~n19920 ) | ( x20 & 1'b0 ) | ( ~n19920 & 1'b0 ) ;
  assign n19968 = ( n19915 & ~x20 ) | ( n19915 & n19920 ) | ( ~x20 & n19920 ) ;
  assign n19969 = ( n19916 & n19967 ) | ( n19916 & n19968 ) | ( n19967 & n19968 ) ;
  assign n19975 = ~n3644 & n13775 ;
  assign n19970 = n3653 | n11081 ;
  assign n19971 = ( n3657 & ~n11091 ) | ( n3657 & 1'b0 ) | ( ~n11091 & 1'b0 ) ;
  assign n19972 = ( n3652 & ~n11093 ) | ( n3652 & 1'b0 ) | ( ~n11093 & 1'b0 ) ;
  assign n19973 = n19971 | n19972 ;
  assign n19974 = ( n19970 & ~n19973 ) | ( n19970 & 1'b0 ) | ( ~n19973 & 1'b0 ) ;
  assign n19976 = ( n3644 & n19975 ) | ( n3644 & n19974 ) | ( n19975 & n19974 ) ;
  assign n19977 = ( n19969 & ~n14780 ) | ( n19969 & n19976 ) | ( ~n14780 & n19976 ) ;
  assign n19978 = ( n14780 & ~n19976 ) | ( n14780 & n19969 ) | ( ~n19976 & n19969 ) ;
  assign n19979 = ( n19977 & ~n19969 ) | ( n19977 & n19978 ) | ( ~n19969 & n19978 ) ;
  assign n19980 = ( n19878 & n19885 ) | ( n19878 & n19923 ) | ( n19885 & n19923 ) ;
  assign n19986 = ~n601 & n13844 ;
  assign n19981 = n4430 | n13836 ;
  assign n19982 = n523 | n11085 ;
  assign n19983 = n3939 | n11078 ;
  assign n19984 = n19982 &  n19983 ;
  assign n19985 = n19981 &  n19984 ;
  assign n19987 = ( n601 & n19986 ) | ( n601 & n19985 ) | ( n19986 & n19985 ) ;
  assign n19989 = x29 &  n19987 ;
  assign n19988 = ~x29 & n19987 ;
  assign n19990 = ( x29 & ~n19989 ) | ( x29 & n19988 ) | ( ~n19989 & n19988 ) ;
  assign n19991 = ( n19979 & ~n19980 ) | ( n19979 & n19990 ) | ( ~n19980 & n19990 ) ;
  assign n19992 = ( n19979 & ~n19990 ) | ( n19979 & n19980 ) | ( ~n19990 & n19980 ) ;
  assign n19993 = ( n19991 & ~n19979 ) | ( n19991 & n19992 ) | ( ~n19979 & n19992 ) ;
  assign n19994 = x29 | n19934 ;
  assign n19995 = x29 &  n19934 ;
  assign n19996 = ( n19994 & ~n19995 ) | ( n19994 & 1'b0 ) | ( ~n19995 & 1'b0 ) ;
  assign n19997 = ( n19926 & n19927 ) | ( n19926 & n19996 ) | ( n19927 & n19996 ) ;
  assign n20001 = n14553 | n4962 ;
  assign n19998 = n4482 | n14071 ;
  assign n19999 = n4495 | n14355 ;
  assign n20000 = n19998 &  n19999 ;
  assign n20002 = ( n4962 & ~n20001 ) | ( n4962 & n20000 ) | ( ~n20001 & n20000 ) ;
  assign n20003 = ( n4478 & n14562 ) | ( n4478 & n20002 ) | ( n14562 & n20002 ) ;
  assign n20004 = ~n4478 & n20003 ;
  assign n20005 = ( x26 & ~n20002 ) | ( x26 & n20004 ) | ( ~n20002 & n20004 ) ;
  assign n20006 = ( n20002 & ~x26 ) | ( n20002 & n20004 ) | ( ~x26 & n20004 ) ;
  assign n20007 = ( n20005 & ~n20004 ) | ( n20005 & n20006 ) | ( ~n20004 & n20006 ) ;
  assign n20008 = ( n19993 & ~n19997 ) | ( n19993 & n20007 ) | ( ~n19997 & n20007 ) ;
  assign n20009 = ( n19993 & ~n20007 ) | ( n19993 & n19997 ) | ( ~n20007 & n19997 ) ;
  assign n20010 = ( n20008 & ~n19993 ) | ( n20008 & n20009 ) | ( ~n19993 & n20009 ) ;
  assign n20014 = n14800 | n5135 ;
  assign n20011 = n5010 | n14803 ;
  assign n20012 = ~n5067 & n14807 ;
  assign n20013 = ( n20011 & ~n20012 ) | ( n20011 & 1'b0 ) | ( ~n20012 & 1'b0 ) ;
  assign n20015 = ( n5135 & ~n20014 ) | ( n5135 & n20013 ) | ( ~n20014 & n20013 ) ;
  assign n20016 = ( n5012 & ~n14816 ) | ( n5012 & n20015 ) | ( ~n14816 & n20015 ) ;
  assign n20017 = ~n5012 & n20016 ;
  assign n20018 = ( x23 & ~n20015 ) | ( x23 & n20017 ) | ( ~n20015 & n20017 ) ;
  assign n20019 = ( n20015 & ~x23 ) | ( n20015 & n20017 ) | ( ~x23 & n20017 ) ;
  assign n20020 = ( n20018 & ~n20017 ) | ( n20018 & n20019 ) | ( ~n20017 & n20019 ) ;
  assign n20021 = ( n19966 & n20010 ) | ( n19966 & n20020 ) | ( n20010 & n20020 ) ;
  assign n20022 = ( n20010 & ~n19966 ) | ( n20010 & n20020 ) | ( ~n19966 & n20020 ) ;
  assign n20023 = ( n19966 & ~n20021 ) | ( n19966 & n20022 ) | ( ~n20021 & n20022 ) ;
  assign n20024 = ( n19946 & ~n19947 ) | ( n19946 & n19948 ) | ( ~n19947 & n19948 ) ;
  assign n20025 = ( n19945 & n20023 ) | ( n19945 & n20024 ) | ( n20023 & n20024 ) ;
  assign n20026 = ( n20023 & ~n19945 ) | ( n20023 & n20024 ) | ( ~n19945 & n20024 ) ;
  assign n20027 = ( ~n19945 & n20025 ) | ( ~n19945 & ~n20026 ) | ( n20025 & ~n20026 ) ;
  assign n20034 = ( n19951 & n19958 ) | ( n19951 & n20027 ) | ( n19958 & n20027 ) ;
  assign n20033 = ( n19958 & ~n19951 ) | ( n19958 & n20027 ) | ( ~n19951 & n20027 ) ;
  assign n20035 = ( n19951 & ~n20034 ) | ( n19951 & n20033 ) | ( ~n20034 & n20033 ) ;
  assign n20031 = ~n8764 & n20027 ;
  assign n20028 = ( n8105 & ~n19494 ) | ( n8105 & 1'b0 ) | ( ~n19494 & 1'b0 ) ;
  assign n20029 = n8429 | n19951 ;
  assign n20030 = ~n20028 & n20029 ;
  assign n20032 = ( n8764 & n20031 ) | ( n8764 & n20030 ) | ( n20031 & n20030 ) ;
  assign n20036 = ( n20032 & ~n8107 ) | ( n20032 & n20035 ) | ( ~n8107 & n20035 ) ;
  assign n20037 = ~n20035 & n20036 ;
  assign n20039 = ( x8 & n20032 ) | ( x8 & n20037 ) | ( n20032 & n20037 ) ;
  assign n20038 = ( x8 & ~n20037 ) | ( x8 & n20032 ) | ( ~n20037 & n20032 ) ;
  assign n20040 = ( n20037 & ~n20039 ) | ( n20037 & n20038 ) | ( ~n20039 & n20038 ) ;
  assign n20041 = ( n19397 & ~n19965 ) | ( n19397 & n20040 ) | ( ~n19965 & n20040 ) ;
  assign n20042 = ( n19397 & ~n20040 ) | ( n19397 & n19965 ) | ( ~n20040 & n19965 ) ;
  assign n20043 = ( n20041 & ~n19397 ) | ( n20041 & n20042 ) | ( ~n19397 & n20042 ) ;
  assign n20227 = ( n19966 & ~n20010 ) | ( n19966 & n20020 ) | ( ~n20010 & n20020 ) ;
  assign n20211 = ( n19997 & ~n19993 ) | ( n19997 & n20007 ) | ( ~n19993 & n20007 ) ;
  assign n20215 = n5067 &  n5135 ;
  assign n20216 = ( n14800 & ~n20215 ) | ( n14800 & 1'b0 ) | ( ~n20215 & 1'b0 ) ;
  assign n20217 = ~n5010 & n14807 ;
  assign n20218 = n20216 | n20217 ;
  assign n20219 = ( n5012 & ~n20218 ) | ( n5012 & n15692 ) | ( ~n20218 & n15692 ) ;
  assign n20220 = ~n5012 & n20219 ;
  assign n20221 = ( n20218 & ~x23 ) | ( n20218 & n20220 ) | ( ~x23 & n20220 ) ;
  assign n20222 = ( x23 & ~n20218 ) | ( x23 & n20220 ) | ( ~n20218 & n20220 ) ;
  assign n20223 = ( n20221 & ~n20220 ) | ( n20221 & n20222 ) | ( ~n20220 & n20222 ) ;
  assign n20045 = n3644 | n13377 ;
  assign n20046 = ( n3652 & ~n11091 ) | ( n3652 & 1'b0 ) | ( ~n11091 & 1'b0 ) ;
  assign n20047 = ( n3657 & ~n11081 ) | ( n3657 & 1'b0 ) | ( ~n11081 & 1'b0 ) ;
  assign n20048 = n20046 | n20047 ;
  assign n20049 = ~n3653 & n11085 ;
  assign n20050 = ( n3653 & ~n20048 ) | ( n3653 & n20049 ) | ( ~n20048 & n20049 ) ;
  assign n20051 = n20045 &  n20050 ;
  assign n20052 = n1196 | n6045 ;
  assign n20053 = ( n4141 & ~n1096 ) | ( n4141 & n20052 ) | ( ~n1096 & n20052 ) ;
  assign n20054 = n1096 | n20053 ;
  assign n20055 = ( n14322 & ~n18930 ) | ( n14322 & n20054 ) | ( ~n18930 & n20054 ) ;
  assign n20056 = ( n4832 & ~n14322 ) | ( n4832 & n20055 ) | ( ~n14322 & n20055 ) ;
  assign n20057 = ( n4832 & ~n20056 ) | ( n4832 & 1'b0 ) | ( ~n20056 & 1'b0 ) ;
  assign n20058 = ( n20057 & ~n1325 ) | ( n20057 & n1884 ) | ( ~n1325 & n1884 ) ;
  assign n20059 = ( n20058 & ~n1884 ) | ( n20058 & 1'b0 ) | ( ~n1884 & 1'b0 ) ;
  assign n20060 = ( n194 & ~n884 ) | ( n194 & n20059 ) | ( ~n884 & n20059 ) ;
  assign n20061 = ~n194 & n20060 ;
  assign n20062 = ( n778 & ~n255 ) | ( n778 & n20061 ) | ( ~n255 & n20061 ) ;
  assign n20063 = ~n778 & n20062 ;
  assign n20064 = ( n406 & ~n569 ) | ( n406 & n20063 ) | ( ~n569 & n20063 ) ;
  assign n20065 = ~n406 & n20064 ;
  assign n20066 = ( n19977 & ~n14780 ) | ( n19977 & n20065 ) | ( ~n14780 & n20065 ) ;
  assign n20067 = ( n14780 & ~n20065 ) | ( n14780 & n19977 ) | ( ~n20065 & n19977 ) ;
  assign n20068 = ( n20066 & ~n19977 ) | ( n20066 & n20067 ) | ( ~n19977 & n20067 ) ;
  assign n20072 = ~n4430 & n14071 ;
  assign n20069 = n523 | n11078 ;
  assign n20070 = n3939 | n13836 ;
  assign n20071 = n20069 &  n20070 ;
  assign n20073 = ( n4430 & n20072 ) | ( n4430 & n20071 ) | ( n20072 & n20071 ) ;
  assign n20074 = ( n601 & ~n14079 ) | ( n601 & n20073 ) | ( ~n14079 & n20073 ) ;
  assign n20075 = ~n601 & n20074 ;
  assign n20077 = ( x29 & n20073 ) | ( x29 & n20075 ) | ( n20073 & n20075 ) ;
  assign n20076 = ( x29 & ~n20075 ) | ( x29 & n20073 ) | ( ~n20075 & n20073 ) ;
  assign n20078 = ( n20075 & ~n20077 ) | ( n20075 & n20076 ) | ( ~n20077 & n20076 ) ;
  assign n20079 = ( n20051 & n20068 ) | ( n20051 & n20078 ) | ( n20068 & n20078 ) ;
  assign n20080 = ( n20068 & ~n20051 ) | ( n20068 & n20078 ) | ( ~n20051 & n20078 ) ;
  assign n20081 = ( n20051 & ~n20079 ) | ( n20051 & n20080 ) | ( ~n20079 & n20080 ) ;
  assign n20044 = ( n19980 & ~n19979 ) | ( n19980 & n19990 ) | ( ~n19979 & n19990 ) ;
  assign n20087 = n15310 | n4478 ;
  assign n20082 = n4962 | n14803 ;
  assign n20083 = n4482 | n14355 ;
  assign n20084 = ~n4495 & n14553 ;
  assign n20085 = ( n20083 & ~n20084 ) | ( n20083 & 1'b0 ) | ( ~n20084 & 1'b0 ) ;
  assign n20086 = n20082 &  n20085 ;
  assign n20088 = ( n4478 & ~n20087 ) | ( n4478 & n20086 ) | ( ~n20087 & n20086 ) ;
  assign n20089 = x26 | n20088 ;
  assign n20090 = ( x26 & ~n20088 ) | ( x26 & 1'b0 ) | ( ~n20088 & 1'b0 ) ;
  assign n20091 = ( n20089 & ~x26 ) | ( n20089 & n20090 ) | ( ~x26 & n20090 ) ;
  assign n20212 = ( n20081 & ~n20044 ) | ( n20081 & n20091 ) | ( ~n20044 & n20091 ) ;
  assign n20213 = ( n20044 & ~n20091 ) | ( n20044 & n20081 ) | ( ~n20091 & n20081 ) ;
  assign n20214 = ( n20212 & ~n20081 ) | ( n20212 & n20213 ) | ( ~n20081 & n20213 ) ;
  assign n20224 = ( n20211 & ~n20223 ) | ( n20211 & n20214 ) | ( ~n20223 & n20214 ) ;
  assign n20225 = ( n20211 & ~n20214 ) | ( n20211 & n20223 ) | ( ~n20214 & n20223 ) ;
  assign n20226 = ( n20224 & ~n20211 ) | ( n20224 & n20225 ) | ( ~n20211 & n20225 ) ;
  assign n20228 = ( n19945 & ~n20023 ) | ( n19945 & n20024 ) | ( ~n20023 & n20024 ) ;
  assign n20239 = ( n20227 & ~n20226 ) | ( n20227 & n20228 ) | ( ~n20226 & n20228 ) ;
  assign n20240 = ( n20226 & ~n20228 ) | ( n20226 & n20227 ) | ( ~n20228 & n20227 ) ;
  assign n20241 = ( ~n20227 & n20239 ) | ( ~n20227 & n20240 ) | ( n20239 & n20240 ) ;
  assign n20229 = ( n20226 & n20227 ) | ( n20226 & n20228 ) | ( n20227 & n20228 ) ;
  assign n20096 = n14807 | n4962 ;
  assign n20093 = ~n4482 & n14553 ;
  assign n20094 = n4495 | n14803 ;
  assign n20095 = ~n20093 & n20094 ;
  assign n20097 = ( n4962 & ~n20096 ) | ( n4962 & n20095 ) | ( ~n20096 & n20095 ) ;
  assign n20098 = ~n4478 & n15294 ;
  assign n20099 = ( n20097 & ~n20098 ) | ( n20097 & 1'b0 ) | ( ~n20098 & 1'b0 ) ;
  assign n20100 = x26 &  n20099 ;
  assign n20101 = x26 | n20099 ;
  assign n20102 = ~n20100 & n20101 ;
  assign n20092 = ( n20044 & ~n20081 ) | ( n20044 & n20091 ) | ( ~n20081 & n20091 ) ;
  assign n20103 = ( n20051 & ~n20068 ) | ( n20051 & n20078 ) | ( ~n20068 & n20078 ) ;
  assign n20129 = n3644 | n11206 ;
  assign n20130 = ( n3652 & ~n11081 ) | ( n3652 & 1'b0 ) | ( ~n11081 & 1'b0 ) ;
  assign n20131 = ( n3657 & ~n11085 ) | ( n3657 & 1'b0 ) | ( ~n11085 & 1'b0 ) ;
  assign n20132 = n20130 | n20131 ;
  assign n20133 = ~n3653 & n11078 ;
  assign n20134 = ( n3653 & ~n20132 ) | ( n3653 & n20133 ) | ( ~n20132 & n20133 ) ;
  assign n20135 = n20129 &  n20134 ;
  assign n20104 = n1207 | n4227 ;
  assign n20105 = ( n5228 & n6681 ) | ( n5228 & n20104 ) | ( n6681 & n20104 ) ;
  assign n20106 = ( n5228 & ~n20105 ) | ( n5228 & 1'b0 ) | ( ~n20105 & 1'b0 ) ;
  assign n20107 = ( n11294 & ~n16407 ) | ( n11294 & n20106 ) | ( ~n16407 & n20106 ) ;
  assign n20108 = ( n314 & ~n11294 ) | ( n314 & n20107 ) | ( ~n11294 & n20107 ) ;
  assign n20109 = ~n314 & n20108 ;
  assign n20110 = ( n604 & ~n1807 ) | ( n604 & n20109 ) | ( ~n1807 & n20109 ) ;
  assign n20111 = ~n604 & n20110 ;
  assign n20112 = ( n346 & ~n952 ) | ( n346 & n20111 ) | ( ~n952 & n20111 ) ;
  assign n20113 = ~n346 & n20112 ;
  assign n20114 = ( n424 & ~n194 ) | ( n424 & n20113 ) | ( ~n194 & n20113 ) ;
  assign n20115 = ~n424 & n20114 ;
  assign n20116 = ( n744 & ~n572 ) | ( n744 & n20115 ) | ( ~n572 & n20115 ) ;
  assign n20117 = ~n744 & n20116 ;
  assign n20118 = ( n617 & ~n670 ) | ( n617 & n20117 ) | ( ~n670 & n20117 ) ;
  assign n20119 = ~n617 & n20118 ;
  assign n20120 = n20065 &  n20119 ;
  assign n20121 = n20065 | n20119 ;
  assign n20122 = ~n20120 & n20121 ;
  assign n20123 = ( n5005 & ~n5002 ) | ( n5005 & n5008 ) | ( ~n5002 & n5008 ) ;
  assign n20124 = n5002 | n20123 ;
  assign n20125 = n14800 &  n20124 ;
  assign n20126 = ( x23 & n20122 ) | ( x23 & n20125 ) | ( n20122 & n20125 ) ;
  assign n20127 = ( n20122 & ~x23 ) | ( n20122 & n20125 ) | ( ~x23 & n20125 ) ;
  assign n20128 = ( x23 & ~n20126 ) | ( x23 & n20127 ) | ( ~n20126 & n20127 ) ;
  assign n20137 = ( n20067 & n20128 ) | ( n20067 & n20135 ) | ( n20128 & n20135 ) ;
  assign n20136 = ( n20067 & ~n20135 ) | ( n20067 & n20128 ) | ( ~n20135 & n20128 ) ;
  assign n20138 = ( n20135 & ~n20137 ) | ( n20135 & n20136 ) | ( ~n20137 & n20136 ) ;
  assign n20142 = ~n4430 & n14355 ;
  assign n20139 = n523 | n13836 ;
  assign n20140 = n3939 | n14071 ;
  assign n20141 = n20139 &  n20140 ;
  assign n20143 = ( n4430 & n20142 ) | ( n4430 & n20141 ) | ( n20142 & n20141 ) ;
  assign n20144 = n601 | n14363 ;
  assign n20145 = n20143 &  n20144 ;
  assign n20146 = x29 &  n20145 ;
  assign n20147 = x29 | n20145 ;
  assign n20148 = ~n20146 & n20147 ;
  assign n20149 = ( n20103 & ~n20138 ) | ( n20103 & n20148 ) | ( ~n20138 & n20148 ) ;
  assign n20150 = ( n20103 & ~n20148 ) | ( n20103 & n20138 ) | ( ~n20148 & n20138 ) ;
  assign n20151 = ( n20149 & ~n20103 ) | ( n20149 & n20150 ) | ( ~n20103 & n20150 ) ;
  assign n20231 = ( n20102 & ~n20092 ) | ( n20102 & n20151 ) | ( ~n20092 & n20151 ) ;
  assign n20232 = ( n20092 & ~n20151 ) | ( n20092 & n20102 ) | ( ~n20151 & n20102 ) ;
  assign n20233 = ( n20231 & ~n20102 ) | ( n20231 & n20232 ) | ( ~n20102 & n20232 ) ;
  assign n20230 = ( n20214 & ~n20211 ) | ( n20214 & n20223 ) | ( ~n20211 & n20223 ) ;
  assign n20243 = ( n20229 & ~n20233 ) | ( n20229 & n20230 ) | ( ~n20233 & n20230 ) ;
  assign n20244 = ( n20230 & ~n20229 ) | ( n20230 & n20233 ) | ( ~n20229 & n20233 ) ;
  assign n20245 = ( n20243 & ~n20230 ) | ( n20243 & n20244 ) | ( ~n20230 & n20244 ) ;
  assign n20249 = ( n20027 & n20034 ) | ( n20027 & n20241 ) | ( n20034 & n20241 ) ;
  assign n20250 = ( n20241 & ~n20245 ) | ( n20241 & n20249 ) | ( ~n20245 & n20249 ) ;
  assign n20264 = ( n20241 & ~n20249 ) | ( n20241 & n20245 ) | ( ~n20249 & n20245 ) ;
  assign n20265 = ( n20250 & ~n20241 ) | ( n20250 & n20264 ) | ( ~n20241 & n20264 ) ;
  assign n20266 = n20265 | n9155 ;
  assign n20259 = ~n9997 & n20245 ;
  assign n20260 = n9160 | n20027 ;
  assign n20261 = n9558 | n20241 ;
  assign n20262 = n20260 &  n20261 ;
  assign n20263 = ~n20259 & n20262 ;
  assign n20267 = ( n9155 & ~n20266 ) | ( n9155 & n20263 ) | ( ~n20266 & n20263 ) ;
  assign n20268 = x5 | n20267 ;
  assign n20269 = ( x5 & ~n20267 ) | ( x5 & 1'b0 ) | ( ~n20267 & 1'b0 ) ;
  assign n20270 = ( n20268 & ~x5 ) | ( n20268 & n20269 ) | ( ~x5 & n20269 ) ;
  assign n20271 = ( n19851 & ~n19964 ) | ( n19851 & n19854 ) | ( ~n19964 & n19854 ) ;
  assign n20272 = ( n19854 & ~n19851 ) | ( n19854 & n19964 ) | ( ~n19851 & n19964 ) ;
  assign n20273 = ( n20271 & ~n19854 ) | ( n20271 & n20272 ) | ( ~n19854 & n20272 ) ;
  assign n20277 = ~n9997 & n20241 ;
  assign n20274 = n9160 | n19951 ;
  assign n20275 = n9558 | n20027 ;
  assign n20276 = n20274 &  n20275 ;
  assign n20278 = ( n9997 & n20277 ) | ( n9997 & n20276 ) | ( n20277 & n20276 ) ;
  assign n20279 = ( n20027 & ~n20241 ) | ( n20027 & n20034 ) | ( ~n20241 & n20034 ) ;
  assign n20280 = ( n20241 & ~n20249 ) | ( n20241 & n20279 ) | ( ~n20249 & n20279 ) ;
  assign n20281 = ( n9155 & ~n20280 ) | ( n9155 & n20278 ) | ( ~n20280 & n20278 ) ;
  assign n20282 = ~n9155 & n20281 ;
  assign n20283 = ( x5 & ~n20278 ) | ( x5 & n20282 ) | ( ~n20278 & n20282 ) ;
  assign n20284 = ( n20278 & ~x5 ) | ( n20278 & n20282 ) | ( ~x5 & n20282 ) ;
  assign n20285 = ( n20283 & ~n20282 ) | ( n20283 & n20284 ) | ( ~n20282 & n20284 ) ;
  assign n20286 = ( n19400 & ~n19507 ) | ( n19400 & n19850 ) | ( ~n19507 & n19850 ) ;
  assign n20287 = ( n19507 & ~n19851 ) | ( n19507 & n20286 ) | ( ~n19851 & n20286 ) ;
  assign n20291 = ~n9997 & n20027 ;
  assign n20288 = n9160 | n19494 ;
  assign n20289 = n9558 | n19951 ;
  assign n20290 = n20288 &  n20289 ;
  assign n20292 = ( n9997 & n20291 ) | ( n9997 & n20290 ) | ( n20291 & n20290 ) ;
  assign n20293 = ( n9155 & ~n20035 ) | ( n9155 & n20292 ) | ( ~n20035 & n20292 ) ;
  assign n20294 = ~n9155 & n20293 ;
  assign n20296 = ( x5 & n20292 ) | ( x5 & n20294 ) | ( n20292 & n20294 ) ;
  assign n20295 = ( x5 & ~n20294 ) | ( x5 & n20292 ) | ( ~n20294 & n20292 ) ;
  assign n20297 = ( n20294 & ~n20296 ) | ( n20294 & n20295 ) | ( ~n20296 & n20295 ) ;
  assign n20298 = ( n19510 & ~n19849 ) | ( n19510 & n19520 ) | ( ~n19849 & n19520 ) ;
  assign n20299 = ( n19850 & ~n19520 ) | ( n19850 & n20298 ) | ( ~n19520 & n20298 ) ;
  assign n20303 = ~n9997 & n19951 ;
  assign n20300 = ~n9160 & n19040 ;
  assign n20301 = n9558 | n19494 ;
  assign n20302 = ~n20300 & n20301 ;
  assign n20304 = ( n9997 & n20303 ) | ( n9997 & n20302 ) | ( n20303 & n20302 ) ;
  assign n20305 = ~n9155 & n19959 ;
  assign n20306 = ( n20304 & ~n20305 ) | ( n20304 & 1'b0 ) | ( ~n20305 & 1'b0 ) ;
  assign n20307 = x5 &  n20306 ;
  assign n20308 = x5 | n20306 ;
  assign n20309 = ~n20307 & n20308 ;
  assign n20310 = ( n19523 & ~n19533 ) | ( n19523 & n19848 ) | ( ~n19533 & n19848 ) ;
  assign n20311 = ( n19533 & ~n19849 ) | ( n19533 & n20310 ) | ( ~n19849 & n20310 ) ;
  assign n20312 = ( n19543 & ~n19847 ) | ( n19543 & n19545 ) | ( ~n19847 & n19545 ) ;
  assign n20313 = ( n19545 & ~n19543 ) | ( n19545 & n19847 ) | ( ~n19543 & n19847 ) ;
  assign n20314 = ( n20312 & ~n19545 ) | ( n20312 & n20313 ) | ( ~n19545 & n20313 ) ;
  assign n20315 = ~n9160 & n19047 ;
  assign n20316 = ~n9558 & n19040 ;
  assign n20317 = n20315 | n20316 ;
  assign n20318 = ~n9997 & n19494 ;
  assign n20319 = ( n9997 & ~n20317 ) | ( n9997 & n20318 ) | ( ~n20317 & n20318 ) ;
  assign n20320 = ( n19502 & ~n9155 ) | ( n19502 & n20319 ) | ( ~n9155 & n20319 ) ;
  assign n20321 = ~n19502 & n20320 ;
  assign n20322 = ( x5 & ~n20319 ) | ( x5 & n20321 ) | ( ~n20319 & n20321 ) ;
  assign n20323 = ( n20319 & ~x5 ) | ( n20319 & n20321 ) | ( ~x5 & n20321 ) ;
  assign n20324 = ( n20322 & ~n20321 ) | ( n20322 & n20323 ) | ( ~n20321 & n20323 ) ;
  assign n20325 = ( n19557 & ~n19555 ) | ( n19557 & n19846 ) | ( ~n19555 & n19846 ) ;
  assign n20326 = ( n19555 & ~n19846 ) | ( n19555 & n19557 ) | ( ~n19846 & n19557 ) ;
  assign n20327 = ( n20325 & ~n19557 ) | ( n20325 & n20326 ) | ( ~n19557 & n20326 ) ;
  assign n20331 = n19040 | n9997 ;
  assign n20328 = n9160 | n19043 ;
  assign n20329 = ~n9558 & n19047 ;
  assign n20330 = ( n20328 & ~n20329 ) | ( n20328 & 1'b0 ) | ( ~n20329 & 1'b0 ) ;
  assign n20332 = ( n9997 & ~n20331 ) | ( n9997 & n20330 ) | ( ~n20331 & n20330 ) ;
  assign n20333 = ( n19056 & ~n9155 ) | ( n19056 & n20332 ) | ( ~n9155 & n20332 ) ;
  assign n20334 = ~n19056 & n20333 ;
  assign n20336 = ( x5 & n20332 ) | ( x5 & n20334 ) | ( n20332 & n20334 ) ;
  assign n20335 = ( x5 & ~n20334 ) | ( x5 & n20332 ) | ( ~n20334 & n20332 ) ;
  assign n20337 = ( n20334 & ~n20336 ) | ( n20334 & n20335 ) | ( ~n20336 & n20335 ) ;
  assign n20341 = n19047 | n9997 ;
  assign n20338 = n9160 | n18712 ;
  assign n20339 = n9558 | n19043 ;
  assign n20340 = n20338 &  n20339 ;
  assign n20342 = ( n9997 & ~n20341 ) | ( n9997 & n20340 ) | ( ~n20341 & n20340 ) ;
  assign n20343 = ~n9155 & n19068 ;
  assign n20344 = ( n20342 & ~n20343 ) | ( n20342 & 1'b0 ) | ( ~n20343 & 1'b0 ) ;
  assign n20345 = x5 &  n20344 ;
  assign n20346 = x5 | n20344 ;
  assign n20347 = ~n20345 & n20346 ;
  assign n20348 = ( n19560 & ~n19845 ) | ( n19560 & n19570 ) | ( ~n19845 & n19570 ) ;
  assign n20349 = ( n19846 & ~n19570 ) | ( n19846 & n20348 ) | ( ~n19570 & n20348 ) ;
  assign n20353 = ~n9997 & n19043 ;
  assign n20350 = n9160 | n18589 ;
  assign n20351 = n9558 | n18712 ;
  assign n20352 = n20350 &  n20351 ;
  assign n20354 = ( n9997 & n20353 ) | ( n9997 & n20352 ) | ( n20353 & n20352 ) ;
  assign n20355 = n9155 | n19083 ;
  assign n20356 = n20354 &  n20355 ;
  assign n20357 = x5 &  n20356 ;
  assign n20358 = x5 | n20356 ;
  assign n20359 = ~n20357 & n20358 ;
  assign n20360 = ( n19573 & ~n19583 ) | ( n19573 & n19844 ) | ( ~n19583 & n19844 ) ;
  assign n20361 = ( n19583 & ~n19845 ) | ( n19583 & n20360 ) | ( ~n19845 & n20360 ) ;
  assign n20365 = ~n9997 & n18712 ;
  assign n20362 = n9160 | n18456 ;
  assign n20363 = n9558 | n18589 ;
  assign n20364 = n20362 &  n20363 ;
  assign n20366 = ( n9997 & n20365 ) | ( n9997 & n20364 ) | ( n20365 & n20364 ) ;
  assign n20367 = n9155 | n18720 ;
  assign n20368 = n20366 &  n20367 ;
  assign n20369 = x5 &  n20368 ;
  assign n20370 = x5 | n20368 ;
  assign n20371 = ~n20369 & n20370 ;
  assign n20372 = ( n19586 & ~n19596 ) | ( n19586 & n19843 ) | ( ~n19596 & n19843 ) ;
  assign n20373 = ( n19596 & ~n19844 ) | ( n19596 & n20372 ) | ( ~n19844 & n20372 ) ;
  assign n20380 = ~n9997 & n18589 ;
  assign n20377 = n9160 | n17783 ;
  assign n20378 = n9558 | n18456 ;
  assign n20379 = n20377 &  n20378 ;
  assign n20381 = ( n9997 & n20380 ) | ( n9997 & n20379 ) | ( n20380 & n20379 ) ;
  assign n20382 = ( n18597 & ~n9155 ) | ( n18597 & n20381 ) | ( ~n9155 & n20381 ) ;
  assign n20383 = ~n18597 & n20382 ;
  assign n20385 = ( x5 & n20381 ) | ( x5 & n20383 ) | ( n20381 & n20383 ) ;
  assign n20384 = ( x5 & ~n20383 ) | ( x5 & n20381 ) | ( ~n20383 & n20381 ) ;
  assign n20386 = ( n20383 & ~n20385 ) | ( n20383 & n20384 ) | ( ~n20385 & n20384 ) ;
  assign n20374 = ( n19608 & ~n19606 ) | ( n19608 & n19842 ) | ( ~n19606 & n19842 ) ;
  assign n20375 = ( n19606 & ~n19842 ) | ( n19606 & n19608 ) | ( ~n19842 & n19608 ) ;
  assign n20376 = ( n20374 & ~n19608 ) | ( n20374 & n20375 ) | ( ~n19608 & n20375 ) ;
  assign n20387 = ( n19620 & ~n19618 ) | ( n19620 & n19841 ) | ( ~n19618 & n19841 ) ;
  assign n20388 = ( n19618 & ~n19841 ) | ( n19618 & n19620 ) | ( ~n19841 & n19620 ) ;
  assign n20389 = ( n20387 & ~n19620 ) | ( n20387 & n20388 ) | ( ~n19620 & n20388 ) ;
  assign n20393 = ~n9997 & n18456 ;
  assign n20390 = n9160 | n17791 ;
  assign n20391 = n9558 | n17783 ;
  assign n20392 = n20390 &  n20391 ;
  assign n20394 = ( n9997 & n20393 ) | ( n9997 & n20392 ) | ( n20393 & n20392 ) ;
  assign n20395 = ( n18464 & ~n9155 ) | ( n18464 & n20394 ) | ( ~n9155 & n20394 ) ;
  assign n20396 = ~n18464 & n20395 ;
  assign n20397 = ( x5 & ~n20394 ) | ( x5 & n20396 ) | ( ~n20394 & n20396 ) ;
  assign n20398 = ( n20394 & ~x5 ) | ( n20394 & n20396 ) | ( ~x5 & n20396 ) ;
  assign n20399 = ( n20397 & ~n20396 ) | ( n20397 & n20398 ) | ( ~n20396 & n20398 ) ;
  assign n20400 = ( n19632 & ~n19630 ) | ( n19632 & n19840 ) | ( ~n19630 & n19840 ) ;
  assign n20401 = ( n19630 & ~n19840 ) | ( n19630 & n19632 ) | ( ~n19840 & n19632 ) ;
  assign n20402 = ( n20400 & ~n19632 ) | ( n20400 & n20401 ) | ( ~n19632 & n20401 ) ;
  assign n20403 = ( n9997 & ~n17783 ) | ( n9997 & 1'b0 ) | ( ~n17783 & 1'b0 ) ;
  assign n20404 = n9160 | n17787 ;
  assign n20405 = n9558 | n17791 ;
  assign n20406 = n20404 &  n20405 ;
  assign n20407 = ( n17783 & n20403 ) | ( n17783 & n20406 ) | ( n20403 & n20406 ) ;
  assign n20408 = ( n17799 & ~n9155 ) | ( n17799 & n20407 ) | ( ~n9155 & n20407 ) ;
  assign n20409 = ~n17799 & n20408 ;
  assign n20411 = ( x5 & n20407 ) | ( x5 & n20409 ) | ( n20407 & n20409 ) ;
  assign n20410 = ( x5 & ~n20409 ) | ( x5 & n20407 ) | ( ~n20409 & n20407 ) ;
  assign n20412 = ( n20409 & ~n20411 ) | ( n20409 & n20410 ) | ( ~n20411 & n20410 ) ;
  assign n20416 = ~n9997 & n17791 ;
  assign n20413 = n9160 | n17405 ;
  assign n20414 = n9558 | n17787 ;
  assign n20415 = n20413 &  n20414 ;
  assign n20417 = ( n9997 & n20416 ) | ( n9997 & n20415 ) | ( n20416 & n20415 ) ;
  assign n20418 = n9155 | n17811 ;
  assign n20419 = n20417 &  n20418 ;
  assign n20420 = x5 &  n20419 ;
  assign n20421 = x5 | n20419 ;
  assign n20422 = ~n20420 & n20421 ;
  assign n20423 = ( n19635 & ~n19839 ) | ( n19635 & n19645 ) | ( ~n19839 & n19645 ) ;
  assign n20424 = ( n19840 & ~n19645 ) | ( n19840 & n20423 ) | ( ~n19645 & n20423 ) ;
  assign n20428 = ~n9997 & n17787 ;
  assign n20425 = n9160 | n17263 ;
  assign n20426 = n9558 | n17405 ;
  assign n20427 = n20425 &  n20426 ;
  assign n20429 = ( n9997 & n20428 ) | ( n9997 & n20427 ) | ( n20428 & n20427 ) ;
  assign n20430 = n9155 | n17826 ;
  assign n20431 = n20429 &  n20430 ;
  assign n20432 = x5 &  n20431 ;
  assign n20433 = x5 | n20431 ;
  assign n20434 = ~n20432 & n20433 ;
  assign n20435 = ( n19648 & ~n19658 ) | ( n19648 & n19838 ) | ( ~n19658 & n19838 ) ;
  assign n20436 = ( n19658 & ~n19839 ) | ( n19658 & n20435 ) | ( ~n19839 & n20435 ) ;
  assign n20440 = ~n9997 & n17405 ;
  assign n20437 = ~n9160 & n17107 ;
  assign n20438 = n9558 | n17263 ;
  assign n20439 = ~n20437 & n20438 ;
  assign n20441 = ( n9997 & n20440 ) | ( n9997 & n20439 ) | ( n20440 & n20439 ) ;
  assign n20442 = n9155 | n17413 ;
  assign n20443 = n20441 &  n20442 ;
  assign n20444 = x5 &  n20443 ;
  assign n20445 = x5 | n20443 ;
  assign n20446 = ~n20444 & n20445 ;
  assign n20447 = ( n19661 & ~n19671 ) | ( n19661 & n19837 ) | ( ~n19671 & n19837 ) ;
  assign n20448 = ( n19671 & ~n19838 ) | ( n19671 & n20447 ) | ( ~n19838 & n20447 ) ;
  assign n20455 = ~n9997 & n17263 ;
  assign n20452 = n9160 | n16589 ;
  assign n20453 = ~n9558 & n17107 ;
  assign n20454 = ( n20452 & ~n20453 ) | ( n20452 & 1'b0 ) | ( ~n20453 & 1'b0 ) ;
  assign n20456 = ( n9997 & n20455 ) | ( n9997 & n20454 ) | ( n20455 & n20454 ) ;
  assign n20457 = ( n9155 & ~n20456 ) | ( n9155 & n17271 ) | ( ~n20456 & n17271 ) ;
  assign n20458 = ( n17271 & ~n20457 ) | ( n17271 & 1'b0 ) | ( ~n20457 & 1'b0 ) ;
  assign n20460 = ( x5 & n20456 ) | ( x5 & n20458 ) | ( n20456 & n20458 ) ;
  assign n20459 = ( x5 & ~n20458 ) | ( x5 & n20456 ) | ( ~n20458 & n20456 ) ;
  assign n20461 = ( n20458 & ~n20460 ) | ( n20458 & n20459 ) | ( ~n20460 & n20459 ) ;
  assign n20449 = ( n19683 & ~n19681 ) | ( n19683 & n19836 ) | ( ~n19681 & n19836 ) ;
  assign n20450 = ( n19681 & ~n19836 ) | ( n19681 & n19683 ) | ( ~n19836 & n19683 ) ;
  assign n20451 = ( n20449 & ~n19683 ) | ( n20449 & n20450 ) | ( ~n19683 & n20450 ) ;
  assign n20462 = ( n19695 & ~n19693 ) | ( n19695 & n19835 ) | ( ~n19693 & n19835 ) ;
  assign n20463 = ( n19693 & ~n19835 ) | ( n19693 & n19695 ) | ( ~n19835 & n19695 ) ;
  assign n20464 = ( n20462 & ~n19695 ) | ( n20462 & n20463 ) | ( ~n19695 & n20463 ) ;
  assign n20468 = n17107 | n9997 ;
  assign n20465 = n9160 | n16595 ;
  assign n20466 = n9558 | n16589 ;
  assign n20467 = n20465 &  n20466 ;
  assign n20469 = ( n9997 & ~n20468 ) | ( n9997 & n20467 ) | ( ~n20468 & n20467 ) ;
  assign n20470 = ( n9155 & ~n20469 ) | ( n9155 & n17115 ) | ( ~n20469 & n17115 ) ;
  assign n20471 = ( n17115 & ~n20470 ) | ( n17115 & 1'b0 ) | ( ~n20470 & 1'b0 ) ;
  assign n20472 = ( x5 & ~n20469 ) | ( x5 & n20471 ) | ( ~n20469 & n20471 ) ;
  assign n20473 = ( n20469 & ~x5 ) | ( n20469 & n20471 ) | ( ~x5 & n20471 ) ;
  assign n20474 = ( n20472 & ~n20471 ) | ( n20472 & n20473 ) | ( ~n20471 & n20473 ) ;
  assign n20475 = ( n19707 & ~n19705 ) | ( n19707 & n19834 ) | ( ~n19705 & n19834 ) ;
  assign n20476 = ( n19705 & ~n19834 ) | ( n19705 & n19707 ) | ( ~n19834 & n19707 ) ;
  assign n20477 = ( n20475 & ~n19707 ) | ( n20475 & n20476 ) | ( ~n19707 & n20476 ) ;
  assign n20481 = ~n9997 & n16589 ;
  assign n20478 = n9160 | n16591 ;
  assign n20479 = n9558 | n16595 ;
  assign n20480 = n20478 &  n20479 ;
  assign n20482 = ( n9997 & n20481 ) | ( n9997 & n20480 ) | ( n20481 & n20480 ) ;
  assign n20483 = ( n16604 & ~n9155 ) | ( n16604 & n20482 ) | ( ~n9155 & n20482 ) ;
  assign n20484 = ~n16604 & n20483 ;
  assign n20486 = ( x5 & n20482 ) | ( x5 & n20484 ) | ( n20482 & n20484 ) ;
  assign n20485 = ( x5 & ~n20484 ) | ( x5 & n20482 ) | ( ~n20484 & n20482 ) ;
  assign n20487 = ( n20484 & ~n20486 ) | ( n20484 & n20485 ) | ( ~n20486 & n20485 ) ;
  assign n20491 = ~n9997 & n16595 ;
  assign n20488 = n9160 | n16091 ;
  assign n20489 = n9558 | n16591 ;
  assign n20490 = n20488 &  n20489 ;
  assign n20492 = ( n9997 & n20491 ) | ( n9997 & n20490 ) | ( n20491 & n20490 ) ;
  assign n20493 = n9155 | n16616 ;
  assign n20494 = n20492 &  n20493 ;
  assign n20495 = x5 &  n20494 ;
  assign n20496 = x5 | n20494 ;
  assign n20497 = ~n20495 & n20496 ;
  assign n20498 = ( n19710 & ~n19833 ) | ( n19710 & n19720 ) | ( ~n19833 & n19720 ) ;
  assign n20499 = ( n19834 & ~n19720 ) | ( n19834 & n20498 ) | ( ~n19720 & n20498 ) ;
  assign n20503 = ~n9997 & n16591 ;
  assign n20500 = n9160 | n15897 ;
  assign n20501 = n9558 | n16091 ;
  assign n20502 = n20500 &  n20501 ;
  assign n20504 = ( n9997 & n20503 ) | ( n9997 & n20502 ) | ( n20503 & n20502 ) ;
  assign n20505 = n9155 | n16631 ;
  assign n20506 = n20504 &  n20505 ;
  assign n20507 = x5 &  n20506 ;
  assign n20508 = x5 | n20506 ;
  assign n20509 = ~n20507 & n20508 ;
  assign n20510 = ( n19723 & ~n19733 ) | ( n19723 & n19832 ) | ( ~n19733 & n19832 ) ;
  assign n20511 = ( n19733 & ~n19833 ) | ( n19733 & n20510 ) | ( ~n19833 & n20510 ) ;
  assign n20515 = ~n9997 & n16091 ;
  assign n20512 = n9160 | n15700 ;
  assign n20513 = n9558 | n15897 ;
  assign n20514 = n20512 &  n20513 ;
  assign n20516 = ( n9997 & n20515 ) | ( n9997 & n20514 ) | ( n20515 & n20514 ) ;
  assign n20517 = n9155 | n16094 ;
  assign n20518 = n20516 &  n20517 ;
  assign n20519 = x5 &  n20518 ;
  assign n20520 = x5 | n20518 ;
  assign n20521 = ~n20519 & n20520 ;
  assign n20522 = ( n19736 & ~n19746 ) | ( n19736 & n19831 ) | ( ~n19746 & n19831 ) ;
  assign n20523 = ( n19746 & ~n19832 ) | ( n19746 & n20522 ) | ( ~n19832 & n20522 ) ;
  assign n20530 = ~n9997 & n15897 ;
  assign n20527 = n9160 | n15320 ;
  assign n20528 = n9558 | n15700 ;
  assign n20529 = n20527 &  n20528 ;
  assign n20531 = ( n9997 & n20530 ) | ( n9997 & n20529 ) | ( n20530 & n20529 ) ;
  assign n20532 = ( n15900 & ~n9155 ) | ( n15900 & n20531 ) | ( ~n9155 & n20531 ) ;
  assign n20533 = ~n15900 & n20532 ;
  assign n20534 = ( x5 & ~n20531 ) | ( x5 & n20533 ) | ( ~n20531 & n20533 ) ;
  assign n20535 = ( n20531 & ~x5 ) | ( n20531 & n20533 ) | ( ~x5 & n20533 ) ;
  assign n20536 = ( n20534 & ~n20533 ) | ( n20534 & n20535 ) | ( ~n20533 & n20535 ) ;
  assign n20524 = ( n19758 & ~n19756 ) | ( n19758 & n19830 ) | ( ~n19756 & n19830 ) ;
  assign n20525 = ( n19756 & ~n19830 ) | ( n19756 & n19758 ) | ( ~n19830 & n19758 ) ;
  assign n20526 = ( n20524 & ~n19758 ) | ( n20524 & n20525 ) | ( ~n19758 & n20525 ) ;
  assign n20537 = ( n19771 & ~n19761 ) | ( n19771 & n19829 ) | ( ~n19761 & n19829 ) ;
  assign n20538 = ( n19761 & ~n19829 ) | ( n19761 & n19771 ) | ( ~n19829 & n19771 ) ;
  assign n20539 = ( n20537 & ~n19771 ) | ( n20537 & n20538 ) | ( ~n19771 & n20538 ) ;
  assign n20543 = ~n9997 & n15700 ;
  assign n20540 = n9160 | n15325 ;
  assign n20541 = n9558 | n15320 ;
  assign n20542 = n20540 &  n20541 ;
  assign n20544 = ( n9997 & n20543 ) | ( n9997 & n20542 ) | ( n20543 & n20542 ) ;
  assign n20545 = ( n15708 & ~n9155 ) | ( n15708 & n20544 ) | ( ~n9155 & n20544 ) ;
  assign n20546 = ~n15708 & n20545 ;
  assign n20548 = ( x5 & n20544 ) | ( x5 & n20546 ) | ( n20544 & n20546 ) ;
  assign n20547 = ( x5 & ~n20546 ) | ( x5 & n20544 ) | ( ~n20546 & n20544 ) ;
  assign n20549 = ( n20546 & ~n20548 ) | ( n20546 & n20547 ) | ( ~n20548 & n20547 ) ;
  assign n20550 = ( n19781 & ~n19828 ) | ( n19781 & n19786 ) | ( ~n19828 & n19786 ) ;
  assign n20551 = ( n19786 & ~n19781 ) | ( n19786 & n19828 ) | ( ~n19781 & n19828 ) ;
  assign n20552 = ( n20550 & ~n19786 ) | ( n20550 & n20551 ) | ( ~n19786 & n20551 ) ;
  assign n20556 = ~n9997 & n15320 ;
  assign n20553 = n9160 | n15322 ;
  assign n20554 = n9558 | n15325 ;
  assign n20555 = n20553 &  n20554 ;
  assign n20557 = ( n9997 & n20556 ) | ( n9997 & n20555 ) | ( n20556 & n20555 ) ;
  assign n20558 = ( n15334 & ~n9155 ) | ( n15334 & n20557 ) | ( ~n9155 & n20557 ) ;
  assign n20559 = ~n15334 & n20558 ;
  assign n20560 = ( x5 & ~n20557 ) | ( x5 & n20559 ) | ( ~n20557 & n20559 ) ;
  assign n20561 = ( n20557 & ~x5 ) | ( n20557 & n20559 ) | ( ~x5 & n20559 ) ;
  assign n20562 = ( n20560 & ~n20559 ) | ( n20560 & n20561 ) | ( ~n20559 & n20561 ) ;
  assign n20566 = ~n9997 & n15325 ;
  assign n20563 = ~n9160 & n14745 ;
  assign n20564 = n9558 | n15322 ;
  assign n20565 = ~n20563 & n20564 ;
  assign n20567 = ( n9997 & n20566 ) | ( n9997 & n20565 ) | ( n20566 & n20565 ) ;
  assign n20568 = n9155 | n15346 ;
  assign n20569 = n20567 &  n20568 ;
  assign n20570 = x5 &  n20569 ;
  assign n20571 = x5 | n20569 ;
  assign n20572 = ~n20570 & n20571 ;
  assign n20573 = ( n19800 & ~n19790 ) | ( n19800 & n19827 ) | ( ~n19790 & n19827 ) ;
  assign n20574 = ( n19828 & ~n19800 ) | ( n19828 & n20573 ) | ( ~n19800 & n20573 ) ;
  assign n20576 = ( n19346 & n19816 ) | ( n19346 & n19826 ) | ( n19816 & n19826 ) ;
  assign n20575 = ( n19346 & ~n19816 ) | ( n19346 & n19826 ) | ( ~n19816 & n19826 ) ;
  assign n20577 = ( n19816 & ~n20576 ) | ( n19816 & n20575 ) | ( ~n20576 & n20575 ) ;
  assign n20581 = ~n9997 & n15322 ;
  assign n20578 = n9160 | n14528 ;
  assign n20579 = ~n9558 & n14745 ;
  assign n20580 = ( n20578 & ~n20579 ) | ( n20578 & 1'b0 ) | ( ~n20579 & 1'b0 ) ;
  assign n20582 = ( n9997 & n20581 ) | ( n9997 & n20580 ) | ( n20581 & n20580 ) ;
  assign n20583 = ( n9155 & ~n20582 ) | ( n9155 & n15361 ) | ( ~n20582 & n15361 ) ;
  assign n20584 = ( n15361 & ~n20583 ) | ( n15361 & 1'b0 ) | ( ~n20583 & 1'b0 ) ;
  assign n20585 = ( x5 & ~n20582 ) | ( x5 & n20584 ) | ( ~n20582 & n20584 ) ;
  assign n20586 = ( n20582 & ~x5 ) | ( n20582 & n20584 ) | ( ~x5 & n20584 ) ;
  assign n20587 = ( n20585 & ~n20584 ) | ( n20585 & n20586 ) | ( ~n20584 & n20586 ) ;
  assign n20591 = n14745 | n9997 ;
  assign n20588 = n9160 | n14261 ;
  assign n20589 = n9558 | n14528 ;
  assign n20590 = n20588 &  n20589 ;
  assign n20592 = ( n9997 & ~n20591 ) | ( n9997 & n20590 ) | ( ~n20591 & n20590 ) ;
  assign n20593 = ~n9155 & n14749 ;
  assign n20594 = ( n20592 & ~n20593 ) | ( n20592 & 1'b0 ) | ( ~n20593 & 1'b0 ) ;
  assign n20595 = x5 &  n20594 ;
  assign n20596 = x5 | n20594 ;
  assign n20597 = ~n20595 & n20596 ;
  assign n20598 = ( x8 & n19801 ) | ( x8 & n19806 ) | ( n19801 & n19806 ) ;
  assign n20599 = ~n19801 & n20598 ;
  assign n20600 = ( n19813 & ~x8 ) | ( n19813 & n20599 ) | ( ~x8 & n20599 ) ;
  assign n20601 = ( x8 & ~n19813 ) | ( x8 & n20599 ) | ( ~n19813 & n20599 ) ;
  assign n20602 = ( n20600 & ~n20599 ) | ( n20600 & n20601 ) | ( ~n20599 & n20601 ) ;
  assign n20603 = x8 &  n19801 ;
  assign n20604 = n19806 &  n20603 ;
  assign n20605 = n19806 | n20603 ;
  assign n20606 = ~n20604 & n20605 ;
  assign n20636 = ~n9997 & n14261 ;
  assign n20633 = n9160 | n13785 ;
  assign n20634 = n9558 | n13998 ;
  assign n20635 = n20633 &  n20634 ;
  assign n20637 = ( n9997 & n20636 ) | ( n9997 & n20635 ) | ( n20636 & n20635 ) ;
  assign n20638 = n9155 | n14267 ;
  assign n20639 = n20637 &  n20638 ;
  assign n20640 = x5 &  n20639 ;
  assign n20641 = x5 | n20639 ;
  assign n20642 = ~n20640 & n20641 ;
  assign n20617 = ( n9154 & ~n13787 ) | ( n9154 & 1'b0 ) | ( ~n13787 & 1'b0 ) ;
  assign n20621 = n13790 | n9155 ;
  assign n20618 = n9558 | n13787 ;
  assign n20619 = n9997 | n13785 ;
  assign n20620 = n20618 &  n20619 ;
  assign n20622 = ( n9155 & ~n20621 ) | ( n9155 & n20620 ) | ( ~n20621 & n20620 ) ;
  assign n20628 = ~n9155 & n14001 ;
  assign n20626 = ~n9997 & n13998 ;
  assign n20623 = n9160 | n13787 ;
  assign n20624 = n9558 | n13785 ;
  assign n20625 = n20623 &  n20624 ;
  assign n20627 = ( n9997 & n20626 ) | ( n9997 & n20625 ) | ( n20626 & n20625 ) ;
  assign n20629 = ( n9155 & n20628 ) | ( n9155 & n20627 ) | ( n20628 & n20627 ) ;
  assign n20630 = ( n20617 & n20622 ) | ( n20617 & n20629 ) | ( n20622 & n20629 ) ;
  assign n20631 = ( x5 & ~n20630 ) | ( x5 & n20617 ) | ( ~n20630 & n20617 ) ;
  assign n20632 = ( x5 & ~n20631 ) | ( x5 & 1'b0 ) | ( ~n20631 & 1'b0 ) ;
  assign n20643 = ( n19801 & ~n20642 ) | ( n19801 & n20632 ) | ( ~n20642 & n20632 ) ;
  assign n20610 = ~n9997 & n14528 ;
  assign n20607 = n9160 | n13998 ;
  assign n20608 = n9558 | n14261 ;
  assign n20609 = n20607 &  n20608 ;
  assign n20611 = ( n9997 & n20610 ) | ( n9997 & n20609 ) | ( n20610 & n20609 ) ;
  assign n20612 = ( n14532 & ~n9155 ) | ( n14532 & n20611 ) | ( ~n9155 & n20611 ) ;
  assign n20613 = ~n14532 & n20612 ;
  assign n20614 = ( x5 & ~n20611 ) | ( x5 & n20613 ) | ( ~n20611 & n20613 ) ;
  assign n20615 = ( n20611 & ~x5 ) | ( n20611 & n20613 ) | ( ~x5 & n20613 ) ;
  assign n20616 = ( n20614 & ~n20613 ) | ( n20614 & n20615 ) | ( ~n20613 & n20615 ) ;
  assign n20644 = ( n20606 & ~n20643 ) | ( n20606 & n20616 ) | ( ~n20643 & n20616 ) ;
  assign n20645 = ( n20597 & n20602 ) | ( n20597 & n20644 ) | ( n20602 & n20644 ) ;
  assign n20646 = ( n20577 & n20587 ) | ( n20577 & n20645 ) | ( n20587 & n20645 ) ;
  assign n20647 = ( n20572 & ~n20574 ) | ( n20572 & n20646 ) | ( ~n20574 & n20646 ) ;
  assign n20648 = ( n20552 & n20562 ) | ( n20552 & n20647 ) | ( n20562 & n20647 ) ;
  assign n20649 = ( n20539 & n20549 ) | ( n20539 & n20648 ) | ( n20549 & n20648 ) ;
  assign n20650 = ( n20536 & ~n20526 ) | ( n20536 & n20649 ) | ( ~n20526 & n20649 ) ;
  assign n20651 = ( n20521 & n20523 ) | ( n20521 & n20650 ) | ( n20523 & n20650 ) ;
  assign n20652 = ( n20509 & n20511 ) | ( n20509 & n20651 ) | ( n20511 & n20651 ) ;
  assign n20653 = ( n20497 & ~n20499 ) | ( n20497 & n20652 ) | ( ~n20499 & n20652 ) ;
  assign n20654 = ( n20477 & n20487 ) | ( n20477 & n20653 ) | ( n20487 & n20653 ) ;
  assign n20655 = ( n20464 & n20474 ) | ( n20464 & n20654 ) | ( n20474 & n20654 ) ;
  assign n20656 = ( n20461 & ~n20451 ) | ( n20461 & n20655 ) | ( ~n20451 & n20655 ) ;
  assign n20657 = ( n20446 & n20448 ) | ( n20446 & n20656 ) | ( n20448 & n20656 ) ;
  assign n20658 = ( n20434 & n20436 ) | ( n20434 & n20657 ) | ( n20436 & n20657 ) ;
  assign n20659 = ( n20422 & ~n20424 ) | ( n20422 & n20658 ) | ( ~n20424 & n20658 ) ;
  assign n20660 = ( n20402 & n20412 ) | ( n20402 & n20659 ) | ( n20412 & n20659 ) ;
  assign n20661 = ( n20389 & n20399 ) | ( n20389 & n20660 ) | ( n20399 & n20660 ) ;
  assign n20662 = ( n20386 & ~n20376 ) | ( n20386 & n20661 ) | ( ~n20376 & n20661 ) ;
  assign n20663 = ( n20371 & n20373 ) | ( n20371 & n20662 ) | ( n20373 & n20662 ) ;
  assign n20664 = ( n20359 & n20361 ) | ( n20359 & n20663 ) | ( n20361 & n20663 ) ;
  assign n20665 = ( n20347 & ~n20349 ) | ( n20347 & n20664 ) | ( ~n20349 & n20664 ) ;
  assign n20666 = ( n20327 & n20337 ) | ( n20327 & n20665 ) | ( n20337 & n20665 ) ;
  assign n20667 = ( n20314 & n20324 ) | ( n20314 & n20666 ) | ( n20324 & n20666 ) ;
  assign n20668 = ( n20309 & n20311 ) | ( n20309 & n20667 ) | ( n20311 & n20667 ) ;
  assign n20669 = ( n20297 & ~n20299 ) | ( n20297 & n20668 ) | ( ~n20299 & n20668 ) ;
  assign n20670 = ( n20285 & n20287 ) | ( n20285 & n20669 ) | ( n20287 & n20669 ) ;
  assign n20671 = ( n20270 & n20273 ) | ( n20270 & n20670 ) | ( n20273 & n20670 ) ;
  assign n20152 = ( n20092 & n20102 ) | ( n20092 & n20151 ) | ( n20102 & n20151 ) ;
  assign n20153 = n1807 | n6820 ;
  assign n20154 = ( n884 & ~n885 ) | ( n884 & n20153 ) | ( ~n885 & n20153 ) ;
  assign n20155 = n885 | n20154 ;
  assign n20156 = ( n274 & ~n281 ) | ( n274 & n20155 ) | ( ~n281 & n20155 ) ;
  assign n20157 = n281 | n20156 ;
  assign n20158 = ( n221 & ~n627 ) | ( n221 & n20157 ) | ( ~n627 & n20157 ) ;
  assign n20159 = n627 | n20158 ;
  assign n20160 = n1271 | n13800 ;
  assign n20161 = ( n997 & n20160 ) | ( n997 & n1092 ) | ( n20160 & n1092 ) ;
  assign n20162 = ( n1092 & ~n20161 ) | ( n1092 & 1'b0 ) | ( ~n20161 & 1'b0 ) ;
  assign n20163 = ( n1122 & n1283 ) | ( n1122 & n20162 ) | ( n1283 & n20162 ) ;
  assign n20164 = ~n1283 & n20163 ;
  assign n20165 = ( n413 & ~n20159 ) | ( n413 & n20164 ) | ( ~n20159 & n20164 ) ;
  assign n20166 = ~n413 & n20165 ;
  assign n20167 = ( n408 & ~n455 ) | ( n408 & n20166 ) | ( ~n455 & n20166 ) ;
  assign n20168 = ~n408 & n20167 ;
  assign n20169 = ( n460 & ~n233 ) | ( n460 & n20168 ) | ( ~n233 & n20168 ) ;
  assign n20170 = ~n460 & n20169 ;
  assign n20171 = ( x23 & ~n20125 ) | ( x23 & 1'b0 ) | ( ~n20125 & 1'b0 ) ;
  assign n20172 = ( n20120 & ~x23 ) | ( n20120 & n20125 ) | ( ~x23 & n20125 ) ;
  assign n20173 = ( n20121 & n20171 ) | ( n20121 & n20172 ) | ( n20171 & n20172 ) ;
  assign n20179 = ~n3644 & n13844 ;
  assign n20174 = n3653 | n13836 ;
  assign n20175 = ( n3657 & ~n11078 ) | ( n3657 & 1'b0 ) | ( ~n11078 & 1'b0 ) ;
  assign n20176 = ( n3652 & ~n11085 ) | ( n3652 & 1'b0 ) | ( ~n11085 & 1'b0 ) ;
  assign n20177 = n20175 | n20176 ;
  assign n20178 = ( n20174 & ~n20177 ) | ( n20174 & 1'b0 ) | ( ~n20177 & 1'b0 ) ;
  assign n20180 = ( n3644 & n20179 ) | ( n3644 & n20178 ) | ( n20179 & n20178 ) ;
  assign n20181 = ( n20170 & ~n20173 ) | ( n20170 & n20180 ) | ( ~n20173 & n20180 ) ;
  assign n20182 = ( n20170 & ~n20180 ) | ( n20170 & n20173 ) | ( ~n20180 & n20173 ) ;
  assign n20183 = ( n20181 & ~n20170 ) | ( n20181 & n20182 ) | ( ~n20170 & n20182 ) ;
  assign n20187 = n14553 | n4430 ;
  assign n20184 = n523 | n14071 ;
  assign n20185 = n3939 | n14355 ;
  assign n20186 = n20184 &  n20185 ;
  assign n20188 = ( n4430 & ~n20187 ) | ( n4430 & n20186 ) | ( ~n20187 & n20186 ) ;
  assign n20189 = ( n601 & ~n20188 ) | ( n601 & n14562 ) | ( ~n20188 & n14562 ) ;
  assign n20190 = ( n14562 & ~n20189 ) | ( n14562 & 1'b0 ) | ( ~n20189 & 1'b0 ) ;
  assign n20191 = ( x29 & ~n20188 ) | ( x29 & n20190 ) | ( ~n20188 & n20190 ) ;
  assign n20192 = ( n20188 & ~x29 ) | ( n20188 & n20190 ) | ( ~x29 & n20190 ) ;
  assign n20193 = ( n20191 & ~n20190 ) | ( n20191 & n20192 ) | ( ~n20190 & n20192 ) ;
  assign n20194 = ( n20183 & ~n20137 ) | ( n20183 & n20193 ) | ( ~n20137 & n20193 ) ;
  assign n20195 = ( n20137 & ~n20193 ) | ( n20137 & n20183 ) | ( ~n20193 & n20183 ) ;
  assign n20196 = ( n20194 & ~n20183 ) | ( n20194 & n20195 ) | ( ~n20183 & n20195 ) ;
  assign n20197 = ( n20103 & n20138 ) | ( n20103 & n20148 ) | ( n20138 & n20148 ) ;
  assign n20201 = n14800 | n4962 ;
  assign n20198 = n4482 | n14803 ;
  assign n20199 = ~n4495 & n14807 ;
  assign n20200 = ( n20198 & ~n20199 ) | ( n20198 & 1'b0 ) | ( ~n20199 & 1'b0 ) ;
  assign n20202 = ( n4962 & ~n20201 ) | ( n4962 & n20200 ) | ( ~n20201 & n20200 ) ;
  assign n20203 = n4478 | n14816 ;
  assign n20204 = n20202 &  n20203 ;
  assign n20205 = x26 &  n20204 ;
  assign n20206 = x26 | n20204 ;
  assign n20207 = ~n20205 & n20206 ;
  assign n20208 = ( n20196 & ~n20197 ) | ( n20196 & n20207 ) | ( ~n20197 & n20207 ) ;
  assign n20209 = ( n20196 & ~n20207 ) | ( n20196 & n20197 ) | ( ~n20207 & n20197 ) ;
  assign n20210 = ( n20208 & ~n20196 ) | ( n20208 & n20209 ) | ( ~n20196 & n20209 ) ;
  assign n20234 = ( n20229 & ~n20230 ) | ( n20229 & n20233 ) | ( ~n20230 & n20233 ) ;
  assign n20235 = ( n20152 & n20210 ) | ( n20152 & n20234 ) | ( n20210 & n20234 ) ;
  assign n20236 = ( n20210 & ~n20152 ) | ( n20210 & n20234 ) | ( ~n20152 & n20234 ) ;
  assign n20237 = ( n20152 & ~n20235 ) | ( n20152 & n20236 ) | ( ~n20235 & n20236 ) ;
  assign n20238 = n9997 &  n20237 ;
  assign n20242 = n9160 | n20241 ;
  assign n20246 = ~n9558 & n20245 ;
  assign n20247 = ( n20242 & ~n20246 ) | ( n20242 & 1'b0 ) | ( ~n20246 & 1'b0 ) ;
  assign n20248 = ( n20238 & ~n20237 ) | ( n20238 & n20247 ) | ( ~n20237 & n20247 ) ;
  assign n20251 = ( n20237 & ~n20245 ) | ( n20237 & n20250 ) | ( ~n20245 & n20250 ) ;
  assign n20252 = ( n20245 & ~n20237 ) | ( n20245 & n20250 ) | ( ~n20237 & n20250 ) ;
  assign n20253 = ( n20251 & ~n20250 ) | ( n20251 & n20252 ) | ( ~n20250 & n20252 ) ;
  assign n20254 = n9155 | n20253 ;
  assign n20255 = n20248 &  n20254 ;
  assign n20256 = x5 &  n20255 ;
  assign n20257 = x5 | n20255 ;
  assign n20258 = ~n20256 & n20257 ;
  assign n20672 = ( n20043 & ~n20671 ) | ( n20043 & n20258 ) | ( ~n20671 & n20258 ) ;
  assign n20673 = ( n20043 & ~n20258 ) | ( n20043 & n20671 ) | ( ~n20258 & n20671 ) ;
  assign n20674 = ( n20672 & ~n20043 ) | ( n20672 & n20673 ) | ( ~n20043 & n20673 ) ;
  assign n20675 = ( n20273 & ~n20270 ) | ( n20273 & n20670 ) | ( ~n20270 & n20670 ) ;
  assign n20676 = ( n20270 & ~n20670 ) | ( n20270 & n20273 ) | ( ~n20670 & n20273 ) ;
  assign n20677 = ( n20675 & ~n20273 ) | ( n20675 & n20676 ) | ( ~n20273 & n20676 ) ;
  assign n20737 = ( n20173 & ~n20170 ) | ( n20173 & n20180 ) | ( ~n20170 & n20180 ) ;
  assign n20704 = n3644 | n14079 ;
  assign n20705 = ( n3652 & ~n11078 ) | ( n3652 & 1'b0 ) | ( ~n11078 & 1'b0 ) ;
  assign n20706 = ( n3657 & ~n13836 ) | ( n3657 & 1'b0 ) | ( ~n13836 & 1'b0 ) ;
  assign n20707 = n20705 | n20706 ;
  assign n20708 = ~n3653 & n14071 ;
  assign n20709 = ( n3653 & ~n20707 ) | ( n3653 & n20708 ) | ( ~n20707 & n20708 ) ;
  assign n20710 = n20704 &  n20709 ;
  assign n20711 = n164 | n1602 ;
  assign n20712 = ( n710 & ~n20711 ) | ( n710 & n13800 ) | ( ~n20711 & n13800 ) ;
  assign n20713 = ( n1028 & ~n13800 ) | ( n1028 & n20712 ) | ( ~n13800 & n20712 ) ;
  assign n20714 = ( n20713 & ~n1028 ) | ( n20713 & 1'b0 ) | ( ~n1028 & 1'b0 ) ;
  assign n20715 = ( n575 & ~n20714 ) | ( n575 & n879 ) | ( ~n20714 & n879 ) ;
  assign n20716 = ( n879 & ~n20715 ) | ( n879 & 1'b0 ) | ( ~n20715 & 1'b0 ) ;
  assign n20717 = ( n789 & n989 ) | ( n789 & n20716 ) | ( n989 & n20716 ) ;
  assign n20718 = ~n789 & n20717 ;
  assign n20719 = ( n460 & ~n20718 ) | ( n460 & n484 ) | ( ~n20718 & n484 ) ;
  assign n20720 = ( n484 & ~n20719 ) | ( n484 & 1'b0 ) | ( ~n20719 & 1'b0 ) ;
  assign n20721 = ( n205 & ~n237 ) | ( n205 & n20720 ) | ( ~n237 & n20720 ) ;
  assign n20722 = ~n205 & n20721 ;
  assign n20723 = ~n417 & n20722 ;
  assign n20724 = ( n20710 & ~n20170 ) | ( n20710 & n20723 ) | ( ~n20170 & n20723 ) ;
  assign n20735 = ( n20170 & ~n20710 ) | ( n20170 & n20723 ) | ( ~n20710 & n20723 ) ;
  assign n20736 = ( n20724 & ~n20723 ) | ( n20724 & n20735 ) | ( ~n20723 & n20735 ) ;
  assign n20738 = ( n20137 & ~n20183 ) | ( n20137 & n20193 ) | ( ~n20183 & n20193 ) ;
  assign n20744 = ( n20736 & n20737 ) | ( n20736 & n20738 ) | ( n20737 & n20738 ) ;
  assign n20745 = ( n20736 & ~n20737 ) | ( n20736 & n20738 ) | ( ~n20737 & n20738 ) ;
  assign n20746 = ( n20737 & ~n20744 ) | ( n20737 & n20745 ) | ( ~n20744 & n20745 ) ;
  assign n20756 = ~n4430 & n14803 ;
  assign n20753 = n523 | n14355 ;
  assign n20754 = ~n3939 & n14553 ;
  assign n20755 = ( n20753 & ~n20754 ) | ( n20753 & 1'b0 ) | ( ~n20754 & 1'b0 ) ;
  assign n20757 = ( n4430 & n20756 ) | ( n4430 & n20755 ) | ( n20756 & n20755 ) ;
  assign n20758 = ~n601 & n15310 ;
  assign n20759 = ( n20757 & ~n20758 ) | ( n20757 & 1'b0 ) | ( ~n20758 & 1'b0 ) ;
  assign n20760 = x29 &  n20759 ;
  assign n20761 = x29 | n20759 ;
  assign n20762 = ~n20760 & n20761 ;
  assign n20747 = n4495 &  n4962 ;
  assign n20748 = ( n14800 & ~n20747 ) | ( n14800 & 1'b0 ) | ( ~n20747 & 1'b0 ) ;
  assign n20749 = ~n4482 & n14807 ;
  assign n20750 = n20748 | n20749 ;
  assign n20751 = ~n4478 & n15692 ;
  assign n20752 = n20750 | n20751 ;
  assign n20763 = ( x26 & ~n20762 ) | ( x26 & n20752 ) | ( ~n20762 & n20752 ) ;
  assign n20764 = ( n20752 & ~x26 ) | ( n20752 & n20762 ) | ( ~x26 & n20762 ) ;
  assign n20765 = ( n20763 & ~n20752 ) | ( n20763 & n20764 ) | ( ~n20752 & n20764 ) ;
  assign n20766 = n20746 | n20765 ;
  assign n20767 = ( n20746 & ~n20765 ) | ( n20746 & 1'b0 ) | ( ~n20765 & 1'b0 ) ;
  assign n20768 = ( n20766 & ~n20746 ) | ( n20766 & n20767 ) | ( ~n20746 & n20767 ) ;
  assign n20743 = ( n20197 & ~n20196 ) | ( n20197 & n20207 ) | ( ~n20196 & n20207 ) ;
  assign n20769 = ( n20152 & ~n20210 ) | ( n20152 & n20234 ) | ( ~n20210 & n20234 ) ;
  assign n20780 = ( n20743 & ~n20769 ) | ( n20743 & n20768 ) | ( ~n20769 & n20768 ) ;
  assign n20781 = ( n20768 & ~n20743 ) | ( n20768 & n20769 ) | ( ~n20743 & n20769 ) ;
  assign n20782 = ( ~n20768 & n20780 ) | ( ~n20768 & n20781 ) | ( n20780 & n20781 ) ;
  assign n20681 = n14807 | n4430 ;
  assign n20678 = ~n523 & n14553 ;
  assign n20679 = n3939 | n14803 ;
  assign n20680 = ~n20678 & n20679 ;
  assign n20682 = ( n4430 & ~n20681 ) | ( n4430 & n20680 ) | ( ~n20681 & n20680 ) ;
  assign n20683 = ~n601 & n15294 ;
  assign n20684 = ( n20682 & ~n20683 ) | ( n20682 & 1'b0 ) | ( ~n20683 & 1'b0 ) ;
  assign n20685 = x29 &  n20684 ;
  assign n20686 = x29 | n20684 ;
  assign n20687 = ~n20685 & n20686 ;
  assign n20725 = n3644 | n14363 ;
  assign n20726 = ( n3652 & ~n13836 ) | ( n3652 & 1'b0 ) | ( ~n13836 & 1'b0 ) ;
  assign n20727 = ( n3657 & ~n14071 ) | ( n3657 & 1'b0 ) | ( ~n14071 & 1'b0 ) ;
  assign n20728 = n20726 | n20727 ;
  assign n20729 = ~n3653 & n14355 ;
  assign n20730 = ( n3653 & ~n20728 ) | ( n3653 & n20729 ) | ( ~n20728 & n20729 ) ;
  assign n20731 = n20725 &  n20730 ;
  assign n20688 = n553 | n698 ;
  assign n20689 = n460 | n20688 ;
  assign n20690 = n774 &  n858 ;
  assign n20691 = ( n929 & n20689 ) | ( n929 & n20690 ) | ( n20689 & n20690 ) ;
  assign n20692 = ( n602 & ~n20689 ) | ( n602 & n20691 ) | ( ~n20689 & n20691 ) ;
  assign n20693 = ~n602 & n20692 ;
  assign n20694 = ~n237 & n20693 ;
  assign n20695 = n20170 &  n20694 ;
  assign n20696 = n20170 | n20694 ;
  assign n20697 = ~n20695 & n20696 ;
  assign n20698 = ( n4477 & ~n4474 ) | ( n4477 & n4480 ) | ( ~n4474 & n4480 ) ;
  assign n20699 = n4474 | n20698 ;
  assign n20700 = n14800 &  n20699 ;
  assign n20701 = ( x26 & n20697 ) | ( x26 & n20700 ) | ( n20697 & n20700 ) ;
  assign n20702 = ( n20697 & ~x26 ) | ( n20697 & n20700 ) | ( ~x26 & n20700 ) ;
  assign n20703 = ( x26 & ~n20701 ) | ( x26 & n20702 ) | ( ~n20701 & n20702 ) ;
  assign n20733 = ( n20703 & n20724 ) | ( n20703 & n20731 ) | ( n20724 & n20731 ) ;
  assign n20732 = ( n20703 & ~n20731 ) | ( n20703 & n20724 ) | ( ~n20731 & n20724 ) ;
  assign n20734 = ( n20731 & ~n20733 ) | ( n20731 & n20732 ) | ( ~n20733 & n20732 ) ;
  assign n20739 = ( n20737 & ~n20736 ) | ( n20737 & n20738 ) | ( ~n20736 & n20738 ) ;
  assign n20740 = ( n20687 & ~n20734 ) | ( n20687 & n20739 ) | ( ~n20734 & n20739 ) ;
  assign n20741 = ( n20687 & ~n20739 ) | ( n20687 & n20734 ) | ( ~n20739 & n20734 ) ;
  assign n20742 = ( n20740 & ~n20687 ) | ( n20740 & n20741 ) | ( ~n20687 & n20741 ) ;
  assign n20770 = ( n20743 & n20768 ) | ( n20743 & n20769 ) | ( n20768 & n20769 ) ;
  assign n20771 = ~x26 & n20752 ;
  assign n20772 = ( x26 & ~n20752 ) | ( x26 & 1'b0 ) | ( ~n20752 & 1'b0 ) ;
  assign n20773 = n20771 | n20772 ;
  assign n20774 = ( n20746 & ~n20762 ) | ( n20746 & n20773 ) | ( ~n20762 & n20773 ) ;
  assign n20775 = ( n20742 & n20770 ) | ( n20742 & n20774 ) | ( n20770 & n20774 ) ;
  assign n20776 = ( n20770 & ~n20742 ) | ( n20770 & n20774 ) | ( ~n20742 & n20774 ) ;
  assign n20777 = ( n20742 & ~n20775 ) | ( n20742 & n20776 ) | ( ~n20775 & n20776 ) ;
  assign n20786 = ( n20237 & ~n20250 ) | ( n20237 & n20245 ) | ( ~n20250 & n20245 ) ;
  assign n20787 = ( n20237 & ~n20782 ) | ( n20237 & n20786 ) | ( ~n20782 & n20786 ) ;
  assign n20788 = ( n20777 & n20782 ) | ( n20777 & n20787 ) | ( n20782 & n20787 ) ;
  assign n20789 = ( n20777 & ~n20782 ) | ( n20777 & n20787 ) | ( ~n20782 & n20787 ) ;
  assign n20790 = ( n20782 & ~n20788 ) | ( n20782 & n20789 ) | ( ~n20788 & n20789 ) ;
  assign n20791 = ~n10017 & n20790 ;
  assign n20778 = n10499 &  n20777 ;
  assign n20779 = ~n10015 & n20237 ;
  assign n20783 = n10486 | n20782 ;
  assign n20784 = ~n20779 & n20783 ;
  assign n20785 = ~n20778 & n20784 ;
  assign n20792 = ( n10017 & n20791 ) | ( n10017 & n20785 ) | ( n20791 & n20785 ) ;
  assign n20794 = x2 &  n20792 ;
  assign n20793 = ~x2 & n20792 ;
  assign n20795 = ( x2 & ~n20794 ) | ( x2 & n20793 ) | ( ~n20794 & n20793 ) ;
  assign n20796 = ( n20314 & ~n20324 ) | ( n20314 & n20666 ) | ( ~n20324 & n20666 ) ;
  assign n20797 = ( n20324 & ~n20667 ) | ( n20324 & n20796 ) | ( ~n20667 & n20796 ) ;
  assign n20806 = ( x5 & n20617 ) | ( x5 & n20622 ) | ( n20617 & n20622 ) ;
  assign n20807 = ~n20617 & n20806 ;
  assign n20808 = ( n20629 & ~x5 ) | ( n20629 & n20807 ) | ( ~x5 & n20807 ) ;
  assign n20809 = ( x5 & ~n20629 ) | ( x5 & n20807 ) | ( ~n20629 & n20807 ) ;
  assign n20810 = ( n20808 & ~n20807 ) | ( n20808 & n20809 ) | ( ~n20807 & n20809 ) ;
  assign n20839 = n10015 | n13998 ;
  assign n20840 = n10486 | n14261 ;
  assign n20841 = n20839 &  n20840 ;
  assign n20842 = n10499 &  n14528 ;
  assign n20843 = ( n20841 & ~n10499 ) | ( n20841 & n20842 ) | ( ~n10499 & n20842 ) ;
  assign n20844 = ( n14532 & ~n10017 ) | ( n14532 & n20843 ) | ( ~n10017 & n20843 ) ;
  assign n20845 = ~n14532 & n20844 ;
  assign n20846 = ( x2 & ~n20843 ) | ( x2 & n20845 ) | ( ~n20843 & n20845 ) ;
  assign n20847 = ( n20843 & ~x2 ) | ( n20843 & n20845 ) | ( ~x2 & n20845 ) ;
  assign n20848 = ( n20846 & ~n20845 ) | ( n20846 & n20847 ) | ( ~n20845 & n20847 ) ;
  assign n20828 = n10015 | n13785 ;
  assign n20829 = n10486 | n13998 ;
  assign n20830 = n20828 &  n20829 ;
  assign n20831 = n10499 &  n14261 ;
  assign n20832 = ( n20830 & ~n10499 ) | ( n20830 & n20831 ) | ( ~n10499 & n20831 ) ;
  assign n20833 = n10017 | n14267 ;
  assign n20834 = n20832 &  n20833 ;
  assign n20835 = x2 &  n20834 ;
  assign n20836 = x2 | n20834 ;
  assign n20837 = ~n20835 & n20836 ;
  assign n20811 = ( n10567 & ~n14001 ) | ( n10567 & 1'b0 ) | ( ~n14001 & 1'b0 ) ;
  assign n20817 = n10567 &  n13790 ;
  assign n20820 = n13785 &  n10499 ;
  assign n20818 = ( n10574 & ~n13787 ) | ( n10574 & 1'b0 ) | ( ~n13787 & 1'b0 ) ;
  assign n20819 = ( x2 & ~n20818 ) | ( x2 & 1'b0 ) | ( ~n20818 & 1'b0 ) ;
  assign n20821 = ( n20820 & ~n10499 ) | ( n20820 & n20819 ) | ( ~n10499 & n20819 ) ;
  assign n20822 = ~n20817 & n20821 ;
  assign n20812 = n10015 | n13787 ;
  assign n20813 = n10486 | n13785 ;
  assign n20814 = n20812 &  n20813 ;
  assign n20815 = n10499 &  n13998 ;
  assign n20816 = ( n20814 & ~n10499 ) | ( n20814 & n20815 ) | ( ~n10499 & n20815 ) ;
  assign n20823 = x2 &  n20816 ;
  assign n20824 = ( n20822 & ~x2 ) | ( n20822 & n20823 ) | ( ~x2 & n20823 ) ;
  assign n20825 = ~n20811 & n20824 ;
  assign n20826 = x0 &  n13787 ;
  assign n20827 = ( n20825 & ~x0 ) | ( n20825 & n20826 ) | ( ~x0 & n20826 ) ;
  assign n20838 = ( n20617 & ~n20837 ) | ( n20617 & n20827 ) | ( ~n20837 & n20827 ) ;
  assign n20849 = x5 &  n20617 ;
  assign n20850 = n20622 &  n20849 ;
  assign n20851 = n20622 | n20849 ;
  assign n20852 = ~n20850 & n20851 ;
  assign n20853 = ( n20848 & ~n20838 ) | ( n20848 & n20852 ) | ( ~n20838 & n20852 ) ;
  assign n20854 = n10015 | n14261 ;
  assign n20855 = n10486 | n14528 ;
  assign n20856 = n20854 &  n20855 ;
  assign n20857 = ( n10499 & ~n14745 ) | ( n10499 & 1'b0 ) | ( ~n14745 & 1'b0 ) ;
  assign n20858 = ( n20856 & ~n10499 ) | ( n20856 & n20857 ) | ( ~n10499 & n20857 ) ;
  assign n20859 = ~n10017 & n14749 ;
  assign n20860 = ( n20858 & ~n20859 ) | ( n20858 & 1'b0 ) | ( ~n20859 & 1'b0 ) ;
  assign n20861 = x2 &  n20860 ;
  assign n20862 = x2 | n20860 ;
  assign n20863 = ~n20861 & n20862 ;
  assign n20864 = ( n20810 & n20853 ) | ( n20810 & n20863 ) | ( n20853 & n20863 ) ;
  assign n20865 = n10015 | n14528 ;
  assign n20866 = ~n10486 & n14745 ;
  assign n20867 = ( n20865 & ~n20866 ) | ( n20865 & 1'b0 ) | ( ~n20866 & 1'b0 ) ;
  assign n20868 = n10499 &  n15322 ;
  assign n20869 = ( n20867 & ~n10499 ) | ( n20867 & n20868 ) | ( ~n10499 & n20868 ) ;
  assign n20870 = ( n10017 & ~n20869 ) | ( n10017 & n15361 ) | ( ~n20869 & n15361 ) ;
  assign n20871 = ( n15361 & ~n20870 ) | ( n15361 & 1'b0 ) | ( ~n20870 & 1'b0 ) ;
  assign n20872 = ( x2 & ~n20869 ) | ( x2 & n20871 ) | ( ~n20869 & n20871 ) ;
  assign n20873 = ( n20869 & ~x2 ) | ( n20869 & n20871 ) | ( ~x2 & n20871 ) ;
  assign n20874 = ( n20872 & ~n20871 ) | ( n20872 & n20873 ) | ( ~n20871 & n20873 ) ;
  assign n20876 = ( n19801 & n20632 ) | ( n19801 & n20642 ) | ( n20632 & n20642 ) ;
  assign n20875 = ( n19801 & ~n20632 ) | ( n19801 & n20642 ) | ( ~n20632 & n20642 ) ;
  assign n20877 = ( n20632 & ~n20876 ) | ( n20632 & n20875 ) | ( ~n20876 & n20875 ) ;
  assign n20878 = ( n20864 & n20874 ) | ( n20864 & n20877 ) | ( n20874 & n20877 ) ;
  assign n20804 = ( n20616 & ~n20606 ) | ( n20616 & n20643 ) | ( ~n20606 & n20643 ) ;
  assign n20805 = ( n20644 & ~n20616 ) | ( n20644 & n20804 ) | ( ~n20616 & n20804 ) ;
  assign n20879 = ~n10015 & n14745 ;
  assign n20880 = n10486 | n15322 ;
  assign n20881 = ~n20879 & n20880 ;
  assign n20882 = n10499 &  n15325 ;
  assign n20883 = ( n20881 & ~n10499 ) | ( n20881 & n20882 ) | ( ~n10499 & n20882 ) ;
  assign n20884 = n10017 | n15346 ;
  assign n20885 = n20883 &  n20884 ;
  assign n20886 = x2 &  n20885 ;
  assign n20887 = x2 | n20885 ;
  assign n20888 = ~n20886 & n20887 ;
  assign n20889 = ( n20878 & ~n20805 ) | ( n20878 & n20888 ) | ( ~n20805 & n20888 ) ;
  assign n20890 = n10015 | n15322 ;
  assign n20891 = n10486 | n15325 ;
  assign n20892 = n20890 &  n20891 ;
  assign n20893 = n10499 &  n15320 ;
  assign n20894 = ( n20892 & ~n10499 ) | ( n20892 & n20893 ) | ( ~n10499 & n20893 ) ;
  assign n20895 = ( n15334 & ~n10017 ) | ( n15334 & n20894 ) | ( ~n10017 & n20894 ) ;
  assign n20896 = ~n15334 & n20895 ;
  assign n20897 = ( x2 & ~n20894 ) | ( x2 & n20896 ) | ( ~n20894 & n20896 ) ;
  assign n20898 = ( n20894 & ~x2 ) | ( n20894 & n20896 ) | ( ~x2 & n20896 ) ;
  assign n20899 = ( n20897 & ~n20896 ) | ( n20897 & n20898 ) | ( ~n20896 & n20898 ) ;
  assign n20900 = ( n20597 & ~n20644 ) | ( n20597 & n20602 ) | ( ~n20644 & n20602 ) ;
  assign n20901 = ( n20602 & ~n20597 ) | ( n20602 & n20644 ) | ( ~n20597 & n20644 ) ;
  assign n20902 = ( n20900 & ~n20602 ) | ( n20900 & n20901 ) | ( ~n20602 & n20901 ) ;
  assign n20903 = ( n20889 & n20899 ) | ( n20889 & n20902 ) | ( n20899 & n20902 ) ;
  assign n20904 = n10015 | n15325 ;
  assign n20905 = n10486 | n15320 ;
  assign n20906 = n20904 &  n20905 ;
  assign n20907 = n10499 &  n15700 ;
  assign n20908 = ( n20906 & ~n10499 ) | ( n20906 & n20907 ) | ( ~n10499 & n20907 ) ;
  assign n20909 = ( n15708 & ~n10017 ) | ( n15708 & n20908 ) | ( ~n10017 & n20908 ) ;
  assign n20910 = ~n15708 & n20909 ;
  assign n20912 = ( x2 & n20908 ) | ( x2 & n20910 ) | ( n20908 & n20910 ) ;
  assign n20911 = ( x2 & ~n20910 ) | ( x2 & n20908 ) | ( ~n20910 & n20908 ) ;
  assign n20913 = ( n20910 & ~n20912 ) | ( n20910 & n20911 ) | ( ~n20912 & n20911 ) ;
  assign n20914 = ( n20587 & ~n20577 ) | ( n20587 & n20645 ) | ( ~n20577 & n20645 ) ;
  assign n20915 = ( n20577 & ~n20645 ) | ( n20577 & n20587 ) | ( ~n20645 & n20587 ) ;
  assign n20916 = ( n20914 & ~n20587 ) | ( n20914 & n20915 ) | ( ~n20587 & n20915 ) ;
  assign n20917 = ( n20903 & n20913 ) | ( n20903 & n20916 ) | ( n20913 & n20916 ) ;
  assign n20928 = ( n20574 & ~n20572 ) | ( n20574 & n20646 ) | ( ~n20572 & n20646 ) ;
  assign n20929 = ( n20572 & ~n20646 ) | ( n20572 & n20574 ) | ( ~n20646 & n20574 ) ;
  assign n20930 = ( n20928 & ~n20574 ) | ( n20928 & n20929 ) | ( ~n20574 & n20929 ) ;
  assign n20918 = n10015 | n15320 ;
  assign n20919 = n10486 | n15700 ;
  assign n20920 = n20918 &  n20919 ;
  assign n20921 = n10499 &  n15897 ;
  assign n20922 = ( n20920 & ~n10499 ) | ( n20920 & n20921 ) | ( ~n10499 & n20921 ) ;
  assign n20923 = ( n15900 & ~n10017 ) | ( n15900 & n20922 ) | ( ~n10017 & n20922 ) ;
  assign n20924 = ~n15900 & n20923 ;
  assign n20925 = ( x2 & ~n20922 ) | ( x2 & n20924 ) | ( ~n20922 & n20924 ) ;
  assign n20926 = ( n20922 & ~x2 ) | ( n20922 & n20924 ) | ( ~x2 & n20924 ) ;
  assign n20927 = ( n20925 & ~n20924 ) | ( n20925 & n20926 ) | ( ~n20924 & n20926 ) ;
  assign n20931 = ( n20917 & ~n20930 ) | ( n20917 & n20927 ) | ( ~n20930 & n20927 ) ;
  assign n20932 = ( n20552 & ~n20562 ) | ( n20552 & n20647 ) | ( ~n20562 & n20647 ) ;
  assign n20933 = ( n20562 & ~n20648 ) | ( n20562 & n20932 ) | ( ~n20648 & n20932 ) ;
  assign n20934 = n10015 | n15700 ;
  assign n20935 = n10486 | n15897 ;
  assign n20936 = n20934 &  n20935 ;
  assign n20937 = n10499 &  n16091 ;
  assign n20938 = ( n20936 & ~n10499 ) | ( n20936 & n20937 ) | ( ~n10499 & n20937 ) ;
  assign n20939 = n10017 | n16094 ;
  assign n20940 = n20938 &  n20939 ;
  assign n20941 = x2 &  n20940 ;
  assign n20942 = x2 | n20940 ;
  assign n20943 = ~n20941 & n20942 ;
  assign n20944 = ( n20931 & n20933 ) | ( n20931 & n20943 ) | ( n20933 & n20943 ) ;
  assign n20945 = ( n20539 & ~n20549 ) | ( n20539 & n20648 ) | ( ~n20549 & n20648 ) ;
  assign n20946 = ( n20549 & ~n20649 ) | ( n20549 & n20945 ) | ( ~n20649 & n20945 ) ;
  assign n20950 = n16591 &  n10499 ;
  assign n20947 = n10015 | n15897 ;
  assign n20948 = n10486 | n16091 ;
  assign n20949 = n20947 &  n20948 ;
  assign n20951 = ( n20950 & ~n10499 ) | ( n20950 & n20949 ) | ( ~n10499 & n20949 ) ;
  assign n20952 = n10017 | n16631 ;
  assign n20953 = n20951 &  n20952 ;
  assign n20954 = x2 &  n20953 ;
  assign n20955 = x2 | n20953 ;
  assign n20956 = ~n20954 & n20955 ;
  assign n20957 = ( n20944 & n20946 ) | ( n20944 & n20956 ) | ( n20946 & n20956 ) ;
  assign n20802 = ( n20526 & ~n20649 ) | ( n20526 & n20536 ) | ( ~n20649 & n20536 ) ;
  assign n20803 = ( n20650 & ~n20536 ) | ( n20650 & n20802 ) | ( ~n20536 & n20802 ) ;
  assign n20958 = n10015 | n16091 ;
  assign n20959 = n10486 | n16591 ;
  assign n20960 = n20958 &  n20959 ;
  assign n20961 = n10499 &  n16595 ;
  assign n20962 = ( n20960 & ~n10499 ) | ( n20960 & n20961 ) | ( ~n10499 & n20961 ) ;
  assign n20963 = n10017 | n16616 ;
  assign n20964 = n20962 &  n20963 ;
  assign n20965 = x2 &  n20964 ;
  assign n20966 = x2 | n20964 ;
  assign n20967 = ~n20965 & n20966 ;
  assign n20968 = ( n20957 & ~n20803 ) | ( n20957 & n20967 ) | ( ~n20803 & n20967 ) ;
  assign n20969 = n10015 | n16591 ;
  assign n20970 = n10486 | n16595 ;
  assign n20971 = n20969 &  n20970 ;
  assign n20972 = n10499 &  n16589 ;
  assign n20973 = ( n20971 & ~n10499 ) | ( n20971 & n20972 ) | ( ~n10499 & n20972 ) ;
  assign n20974 = ( n16604 & ~n10017 ) | ( n16604 & n20973 ) | ( ~n10017 & n20973 ) ;
  assign n20975 = ~n16604 & n20974 ;
  assign n20977 = ( x2 & n20973 ) | ( x2 & n20975 ) | ( n20973 & n20975 ) ;
  assign n20976 = ( x2 & ~n20975 ) | ( x2 & n20973 ) | ( ~n20975 & n20973 ) ;
  assign n20978 = ( n20975 & ~n20977 ) | ( n20975 & n20976 ) | ( ~n20977 & n20976 ) ;
  assign n20979 = ( n20523 & ~n20521 ) | ( n20523 & n20650 ) | ( ~n20521 & n20650 ) ;
  assign n20980 = ( n20521 & ~n20650 ) | ( n20521 & n20523 ) | ( ~n20650 & n20523 ) ;
  assign n20981 = ( n20979 & ~n20523 ) | ( n20979 & n20980 ) | ( ~n20523 & n20980 ) ;
  assign n20982 = ( n20968 & n20978 ) | ( n20968 & n20981 ) | ( n20978 & n20981 ) ;
  assign n20983 = n10015 | n16595 ;
  assign n20984 = n10486 | n16589 ;
  assign n20985 = n20983 &  n20984 ;
  assign n20986 = ( n10499 & ~n17107 ) | ( n10499 & 1'b0 ) | ( ~n17107 & 1'b0 ) ;
  assign n20987 = ( n20985 & ~n10499 ) | ( n20985 & n20986 ) | ( ~n10499 & n20986 ) ;
  assign n20988 = ( n10017 & ~n20987 ) | ( n10017 & n17115 ) | ( ~n20987 & n17115 ) ;
  assign n20989 = ( n17115 & ~n20988 ) | ( n17115 & 1'b0 ) | ( ~n20988 & 1'b0 ) ;
  assign n20990 = ( x2 & ~n20987 ) | ( x2 & n20989 ) | ( ~n20987 & n20989 ) ;
  assign n20991 = ( n20987 & ~x2 ) | ( n20987 & n20989 ) | ( ~x2 & n20989 ) ;
  assign n20992 = ( n20990 & ~n20989 ) | ( n20990 & n20991 ) | ( ~n20989 & n20991 ) ;
  assign n20993 = ( n20511 & ~n20509 ) | ( n20511 & n20651 ) | ( ~n20509 & n20651 ) ;
  assign n20994 = ( n20509 & ~n20651 ) | ( n20509 & n20511 ) | ( ~n20651 & n20511 ) ;
  assign n20995 = ( n20993 & ~n20511 ) | ( n20993 & n20994 ) | ( ~n20511 & n20994 ) ;
  assign n20996 = ( n20982 & n20992 ) | ( n20982 & n20995 ) | ( n20992 & n20995 ) ;
  assign n21007 = ( n20499 & ~n20497 ) | ( n20499 & n20652 ) | ( ~n20497 & n20652 ) ;
  assign n21008 = ( n20497 & ~n20652 ) | ( n20497 & n20499 ) | ( ~n20652 & n20499 ) ;
  assign n21009 = ( n21007 & ~n20499 ) | ( n21007 & n21008 ) | ( ~n20499 & n21008 ) ;
  assign n21000 = n17263 &  n10499 ;
  assign n20997 = n10015 | n16589 ;
  assign n20998 = ~n10486 & n17107 ;
  assign n20999 = ( n20997 & ~n20998 ) | ( n20997 & 1'b0 ) | ( ~n20998 & 1'b0 ) ;
  assign n21001 = ( n21000 & ~n10499 ) | ( n21000 & n20999 ) | ( ~n10499 & n20999 ) ;
  assign n21002 = ( n10017 & ~n21001 ) | ( n10017 & n17271 ) | ( ~n21001 & n17271 ) ;
  assign n21003 = ( n17271 & ~n21002 ) | ( n17271 & 1'b0 ) | ( ~n21002 & 1'b0 ) ;
  assign n21005 = ( x2 & n21001 ) | ( x2 & n21003 ) | ( n21001 & n21003 ) ;
  assign n21004 = ( x2 & ~n21003 ) | ( x2 & n21001 ) | ( ~n21003 & n21001 ) ;
  assign n21006 = ( n21003 & ~n21005 ) | ( n21003 & n21004 ) | ( ~n21005 & n21004 ) ;
  assign n21010 = ( n20996 & ~n21009 ) | ( n20996 & n21006 ) | ( ~n21009 & n21006 ) ;
  assign n21011 = ( n20477 & ~n20487 ) | ( n20477 & n20653 ) | ( ~n20487 & n20653 ) ;
  assign n21012 = ( n20487 & ~n20654 ) | ( n20487 & n21011 ) | ( ~n20654 & n21011 ) ;
  assign n21016 = n17405 &  n10499 ;
  assign n21013 = ~n10015 & n17107 ;
  assign n21014 = n10486 | n17263 ;
  assign n21015 = ~n21013 & n21014 ;
  assign n21017 = ( n21016 & ~n10499 ) | ( n21016 & n21015 ) | ( ~n10499 & n21015 ) ;
  assign n21018 = n10017 | n17413 ;
  assign n21019 = n21017 &  n21018 ;
  assign n21020 = x2 &  n21019 ;
  assign n21021 = x2 | n21019 ;
  assign n21022 = ~n21020 & n21021 ;
  assign n21023 = ( n21010 & n21012 ) | ( n21010 & n21022 ) | ( n21012 & n21022 ) ;
  assign n21024 = ( n20464 & ~n20474 ) | ( n20464 & n20654 ) | ( ~n20474 & n20654 ) ;
  assign n21025 = ( n20474 & ~n20655 ) | ( n20474 & n21024 ) | ( ~n20655 & n21024 ) ;
  assign n21026 = n10015 | n17263 ;
  assign n21027 = n10486 | n17405 ;
  assign n21028 = n21026 &  n21027 ;
  assign n21029 = n10499 &  n17787 ;
  assign n21030 = ( n21028 & ~n10499 ) | ( n21028 & n21029 ) | ( ~n10499 & n21029 ) ;
  assign n21031 = n10017 | n17826 ;
  assign n21032 = n21030 &  n21031 ;
  assign n21033 = x2 &  n21032 ;
  assign n21034 = x2 | n21032 ;
  assign n21035 = ~n21033 & n21034 ;
  assign n21036 = ( n21023 & n21025 ) | ( n21023 & n21035 ) | ( n21025 & n21035 ) ;
  assign n20800 = ( n20451 & ~n20655 ) | ( n20451 & n20461 ) | ( ~n20655 & n20461 ) ;
  assign n20801 = ( n20656 & ~n20461 ) | ( n20656 & n20800 ) | ( ~n20461 & n20800 ) ;
  assign n21037 = n10015 | n17405 ;
  assign n21038 = n10486 | n17787 ;
  assign n21039 = n21037 &  n21038 ;
  assign n21040 = n10499 &  n17791 ;
  assign n21041 = ( n21039 & ~n10499 ) | ( n21039 & n21040 ) | ( ~n10499 & n21040 ) ;
  assign n21042 = n10017 | n17811 ;
  assign n21043 = n21041 &  n21042 ;
  assign n21044 = x2 &  n21043 ;
  assign n21045 = x2 | n21043 ;
  assign n21046 = ~n21044 & n21045 ;
  assign n21047 = ( n21036 & ~n20801 ) | ( n21036 & n21046 ) | ( ~n20801 & n21046 ) ;
  assign n21051 = n17783 &  n10499 ;
  assign n21048 = n10015 | n17787 ;
  assign n21049 = n10486 | n17791 ;
  assign n21050 = n21048 &  n21049 ;
  assign n21052 = ( n21051 & ~n10499 ) | ( n21051 & n21050 ) | ( ~n10499 & n21050 ) ;
  assign n21053 = ( n17799 & ~n10017 ) | ( n17799 & n21052 ) | ( ~n10017 & n21052 ) ;
  assign n21054 = ~n17799 & n21053 ;
  assign n21056 = ( x2 & n21052 ) | ( x2 & n21054 ) | ( n21052 & n21054 ) ;
  assign n21055 = ( x2 & ~n21054 ) | ( x2 & n21052 ) | ( ~n21054 & n21052 ) ;
  assign n21057 = ( n21054 & ~n21056 ) | ( n21054 & n21055 ) | ( ~n21056 & n21055 ) ;
  assign n21058 = ( n20448 & ~n20446 ) | ( n20448 & n20656 ) | ( ~n20446 & n20656 ) ;
  assign n21059 = ( n20446 & ~n20656 ) | ( n20446 & n20448 ) | ( ~n20656 & n20448 ) ;
  assign n21060 = ( n21058 & ~n20448 ) | ( n21058 & n21059 ) | ( ~n20448 & n21059 ) ;
  assign n21061 = ( n21047 & n21057 ) | ( n21047 & n21060 ) | ( n21057 & n21060 ) ;
  assign n21062 = n10015 | n17791 ;
  assign n21063 = n10486 | n17783 ;
  assign n21064 = n21062 &  n21063 ;
  assign n21065 = n10499 &  n18456 ;
  assign n21066 = ( n21064 & ~n10499 ) | ( n21064 & n21065 ) | ( ~n10499 & n21065 ) ;
  assign n21067 = ( n18464 & ~n10017 ) | ( n18464 & n21066 ) | ( ~n10017 & n21066 ) ;
  assign n21068 = ~n18464 & n21067 ;
  assign n21069 = ( x2 & ~n21066 ) | ( x2 & n21068 ) | ( ~n21066 & n21068 ) ;
  assign n21070 = ( n21066 & ~x2 ) | ( n21066 & n21068 ) | ( ~x2 & n21068 ) ;
  assign n21071 = ( n21069 & ~n21068 ) | ( n21069 & n21070 ) | ( ~n21068 & n21070 ) ;
  assign n21072 = ( n20436 & ~n20434 ) | ( n20436 & n20657 ) | ( ~n20434 & n20657 ) ;
  assign n21073 = ( n20434 & ~n20657 ) | ( n20434 & n20436 ) | ( ~n20657 & n20436 ) ;
  assign n21074 = ( n21072 & ~n20436 ) | ( n21072 & n21073 ) | ( ~n20436 & n21073 ) ;
  assign n21075 = ( n21061 & n21071 ) | ( n21061 & n21074 ) | ( n21071 & n21074 ) ;
  assign n21086 = ( n20424 & ~n20422 ) | ( n20424 & n20658 ) | ( ~n20422 & n20658 ) ;
  assign n21087 = ( n20422 & ~n20658 ) | ( n20422 & n20424 ) | ( ~n20658 & n20424 ) ;
  assign n21088 = ( n21086 & ~n20424 ) | ( n21086 & n21087 ) | ( ~n20424 & n21087 ) ;
  assign n21076 = n10015 | n17783 ;
  assign n21077 = n10486 | n18456 ;
  assign n21078 = n21076 &  n21077 ;
  assign n21079 = n10499 &  n18589 ;
  assign n21080 = ( n21078 & ~n10499 ) | ( n21078 & n21079 ) | ( ~n10499 & n21079 ) ;
  assign n21081 = ( n18597 & ~n10017 ) | ( n18597 & n21080 ) | ( ~n10017 & n21080 ) ;
  assign n21082 = ~n18597 & n21081 ;
  assign n21084 = ( x2 & n21080 ) | ( x2 & n21082 ) | ( n21080 & n21082 ) ;
  assign n21083 = ( x2 & ~n21082 ) | ( x2 & n21080 ) | ( ~n21082 & n21080 ) ;
  assign n21085 = ( n21082 & ~n21084 ) | ( n21082 & n21083 ) | ( ~n21084 & n21083 ) ;
  assign n21089 = ( n21075 & ~n21088 ) | ( n21075 & n21085 ) | ( ~n21088 & n21085 ) ;
  assign n21090 = ( n20402 & ~n20412 ) | ( n20402 & n20659 ) | ( ~n20412 & n20659 ) ;
  assign n21091 = ( n20412 & ~n20660 ) | ( n20412 & n21090 ) | ( ~n20660 & n21090 ) ;
  assign n21092 = n10015 | n18456 ;
  assign n21093 = n10486 | n18589 ;
  assign n21094 = n21092 &  n21093 ;
  assign n21095 = n10499 &  n18712 ;
  assign n21096 = ( n21094 & ~n10499 ) | ( n21094 & n21095 ) | ( ~n10499 & n21095 ) ;
  assign n21097 = n10017 | n18720 ;
  assign n21098 = n21096 &  n21097 ;
  assign n21099 = x2 &  n21098 ;
  assign n21100 = x2 | n21098 ;
  assign n21101 = ~n21099 & n21100 ;
  assign n21102 = ( n21089 & n21091 ) | ( n21089 & n21101 ) | ( n21091 & n21101 ) ;
  assign n21103 = ( n20389 & ~n20399 ) | ( n20389 & n20660 ) | ( ~n20399 & n20660 ) ;
  assign n21104 = ( n20399 & ~n20661 ) | ( n20399 & n21103 ) | ( ~n20661 & n21103 ) ;
  assign n21105 = n10015 | n18589 ;
  assign n21106 = n10486 | n18712 ;
  assign n21107 = n21105 &  n21106 ;
  assign n21108 = n10499 &  n19043 ;
  assign n21109 = ( n21107 & ~n10499 ) | ( n21107 & n21108 ) | ( ~n10499 & n21108 ) ;
  assign n21110 = n10017 | n19083 ;
  assign n21111 = n21109 &  n21110 ;
  assign n21112 = x2 &  n21111 ;
  assign n21113 = x2 | n21111 ;
  assign n21114 = ~n21112 & n21113 ;
  assign n21115 = ( n21102 & n21104 ) | ( n21102 & n21114 ) | ( n21104 & n21114 ) ;
  assign n20798 = ( n20376 & ~n20661 ) | ( n20376 & n20386 ) | ( ~n20661 & n20386 ) ;
  assign n20799 = ( n20662 & ~n20386 ) | ( n20662 & n20798 ) | ( ~n20386 & n20798 ) ;
  assign n21116 = n10015 | n18712 ;
  assign n21117 = n10486 | n19043 ;
  assign n21118 = n21116 &  n21117 ;
  assign n21119 = ( n10499 & ~n19047 ) | ( n10499 & 1'b0 ) | ( ~n19047 & 1'b0 ) ;
  assign n21120 = ( n21118 & ~n10499 ) | ( n21118 & n21119 ) | ( ~n10499 & n21119 ) ;
  assign n21121 = ~n10017 & n19068 ;
  assign n21122 = ( n21120 & ~n21121 ) | ( n21120 & 1'b0 ) | ( ~n21121 & 1'b0 ) ;
  assign n21123 = x2 &  n21122 ;
  assign n21124 = x2 | n21122 ;
  assign n21125 = ~n21123 & n21124 ;
  assign n21126 = ( n21115 & ~n20799 ) | ( n21115 & n21125 ) | ( ~n20799 & n21125 ) ;
  assign n21127 = n10015 | n19043 ;
  assign n21128 = ~n10486 & n19047 ;
  assign n21129 = ( n21127 & ~n21128 ) | ( n21127 & 1'b0 ) | ( ~n21128 & 1'b0 ) ;
  assign n21130 = ( n10499 & ~n19040 ) | ( n10499 & 1'b0 ) | ( ~n19040 & 1'b0 ) ;
  assign n21131 = ( n21129 & ~n10499 ) | ( n21129 & n21130 ) | ( ~n10499 & n21130 ) ;
  assign n21132 = ( n19056 & ~n10017 ) | ( n19056 & n21131 ) | ( ~n10017 & n21131 ) ;
  assign n21133 = ~n19056 & n21132 ;
  assign n21135 = ( x2 & n21131 ) | ( x2 & n21133 ) | ( n21131 & n21133 ) ;
  assign n21134 = ( x2 & ~n21133 ) | ( x2 & n21131 ) | ( ~n21133 & n21131 ) ;
  assign n21136 = ( n21133 & ~n21135 ) | ( n21133 & n21134 ) | ( ~n21135 & n21134 ) ;
  assign n21137 = ( n20373 & ~n20371 ) | ( n20373 & n20662 ) | ( ~n20371 & n20662 ) ;
  assign n21138 = ( n20371 & ~n20662 ) | ( n20371 & n20373 ) | ( ~n20662 & n20373 ) ;
  assign n21139 = ( n21137 & ~n20373 ) | ( n21137 & n21138 ) | ( ~n20373 & n21138 ) ;
  assign n21140 = ( n21126 & n21136 ) | ( n21126 & n21139 ) | ( n21136 & n21139 ) ;
  assign n21144 = n10499 &  n19494 ;
  assign n21141 = ~n10015 & n19047 ;
  assign n21142 = ~n10486 & n19040 ;
  assign n21143 = n21141 | n21142 ;
  assign n21145 = ( n10499 & ~n21144 ) | ( n10499 & n21143 ) | ( ~n21144 & n21143 ) ;
  assign n21146 = ( n10017 & ~n19502 ) | ( n10017 & n21145 ) | ( ~n19502 & n21145 ) ;
  assign n21147 = n19502 | n21146 ;
  assign n21149 = ( x2 & n21145 ) | ( x2 & n21147 ) | ( n21145 & n21147 ) ;
  assign n21148 = ( x2 & ~n21147 ) | ( x2 & n21145 ) | ( ~n21147 & n21145 ) ;
  assign n21150 = ( n21147 & ~n21149 ) | ( n21147 & n21148 ) | ( ~n21149 & n21148 ) ;
  assign n21151 = ( n20361 & ~n20359 ) | ( n20361 & n20663 ) | ( ~n20359 & n20663 ) ;
  assign n21152 = ( n20359 & ~n20663 ) | ( n20359 & n20361 ) | ( ~n20663 & n20361 ) ;
  assign n21153 = ( n21151 & ~n20361 ) | ( n21151 & n21152 ) | ( ~n20361 & n21152 ) ;
  assign n21154 = ( n21140 & n21150 ) | ( n21140 & n21153 ) | ( n21150 & n21153 ) ;
  assign n21165 = ( n20349 & ~n20347 ) | ( n20349 & n20664 ) | ( ~n20347 & n20664 ) ;
  assign n21166 = ( n20347 & ~n20664 ) | ( n20347 & n20349 ) | ( ~n20664 & n20349 ) ;
  assign n21167 = ( n21165 & ~n20349 ) | ( n21165 & n21166 ) | ( ~n20349 & n21166 ) ;
  assign n21155 = ~n10015 & n19040 ;
  assign n21156 = n10486 | n19494 ;
  assign n21157 = ~n21155 & n21156 ;
  assign n21158 = n10499 &  n19951 ;
  assign n21159 = ( n21157 & ~n10499 ) | ( n21157 & n21158 ) | ( ~n10499 & n21158 ) ;
  assign n21160 = ( n10017 & ~n21159 ) | ( n10017 & n19959 ) | ( ~n21159 & n19959 ) ;
  assign n21161 = ( n19959 & ~n21160 ) | ( n19959 & 1'b0 ) | ( ~n21160 & 1'b0 ) ;
  assign n21163 = ( x2 & n21159 ) | ( x2 & n21161 ) | ( n21159 & n21161 ) ;
  assign n21162 = ( x2 & ~n21161 ) | ( x2 & n21159 ) | ( ~n21161 & n21159 ) ;
  assign n21164 = ( n21161 & ~n21163 ) | ( n21161 & n21162 ) | ( ~n21163 & n21162 ) ;
  assign n21168 = ( n21154 & ~n21167 ) | ( n21154 & n21164 ) | ( ~n21167 & n21164 ) ;
  assign n21169 = ( n20327 & ~n20337 ) | ( n20327 & n20665 ) | ( ~n20337 & n20665 ) ;
  assign n21170 = ( n20337 & ~n20666 ) | ( n20337 & n21169 ) | ( ~n20666 & n21169 ) ;
  assign n21171 = n10015 | n19494 ;
  assign n21172 = n10486 | n19951 ;
  assign n21173 = n21171 &  n21172 ;
  assign n21174 = n10499 &  n20027 ;
  assign n21175 = ( n21173 & ~n10499 ) | ( n21173 & n21174 ) | ( ~n10499 & n21174 ) ;
  assign n21176 = n10017 | n20035 ;
  assign n21177 = n21175 &  n21176 ;
  assign n21178 = x2 &  n21177 ;
  assign n21179 = x2 | n21177 ;
  assign n21180 = ~n21178 & n21179 ;
  assign n21181 = ( n21168 & n21170 ) | ( n21168 & n21180 ) | ( n21170 & n21180 ) ;
  assign n21182 = n10015 | n19951 ;
  assign n21183 = n10486 | n20027 ;
  assign n21184 = n21182 &  n21183 ;
  assign n21185 = n10499 &  n20241 ;
  assign n21186 = ( n21184 & ~n10499 ) | ( n21184 & n21185 ) | ( ~n10499 & n21185 ) ;
  assign n21187 = n10017 | n20280 ;
  assign n21188 = n21186 &  n21187 ;
  assign n21189 = x2 &  n21188 ;
  assign n21190 = x2 | n21188 ;
  assign n21191 = ~n21189 & n21190 ;
  assign n21192 = ( n20797 & n21181 ) | ( n20797 & n21191 ) | ( n21181 & n21191 ) ;
  assign n21196 = ~n20245 & n10499 ;
  assign n21193 = n10015 | n20027 ;
  assign n21194 = n10486 | n20241 ;
  assign n21195 = n21193 &  n21194 ;
  assign n21197 = ( n21196 & ~n10499 ) | ( n21196 & n21195 ) | ( ~n10499 & n21195 ) ;
  assign n21198 = ( n10017 & ~n21197 ) | ( n10017 & n20265 ) | ( ~n21197 & n20265 ) ;
  assign n21199 = ( n20265 & ~n21198 ) | ( n20265 & 1'b0 ) | ( ~n21198 & 1'b0 ) ;
  assign n21201 = ( x2 & n21197 ) | ( x2 & n21199 ) | ( n21197 & n21199 ) ;
  assign n21200 = ( x2 & ~n21199 ) | ( x2 & n21197 ) | ( ~n21199 & n21197 ) ;
  assign n21202 = ( n21199 & ~n21201 ) | ( n21199 & n21200 ) | ( ~n21201 & n21200 ) ;
  assign n21203 = ( n20311 & ~n20309 ) | ( n20311 & n20667 ) | ( ~n20309 & n20667 ) ;
  assign n21204 = ( n20309 & ~n20667 ) | ( n20309 & n20311 ) | ( ~n20667 & n20311 ) ;
  assign n21205 = ( n21203 & ~n20311 ) | ( n21203 & n21204 ) | ( ~n20311 & n21204 ) ;
  assign n21206 = ( n21192 & n21202 ) | ( n21192 & n21205 ) | ( n21202 & n21205 ) ;
  assign n21217 = ( n20297 & ~n20668 ) | ( n20297 & n20299 ) | ( ~n20668 & n20299 ) ;
  assign n21218 = ( n20299 & ~n20297 ) | ( n20299 & n20668 ) | ( ~n20297 & n20668 ) ;
  assign n21219 = ( n21217 & ~n20299 ) | ( n21217 & n21218 ) | ( ~n20299 & n21218 ) ;
  assign n21210 = ~n20237 & n10499 ;
  assign n21207 = n10015 | n20241 ;
  assign n21208 = ~n10486 & n20245 ;
  assign n21209 = ( n21207 & ~n21208 ) | ( n21207 & 1'b0 ) | ( ~n21208 & 1'b0 ) ;
  assign n21211 = ( n21210 & ~n10499 ) | ( n21210 & n21209 ) | ( ~n10499 & n21209 ) ;
  assign n21212 = ( n10017 & ~n20253 ) | ( n10017 & n21211 ) | ( ~n20253 & n21211 ) ;
  assign n21213 = ~n10017 & n21212 ;
  assign n21215 = ( x2 & n21211 ) | ( x2 & n21213 ) | ( n21211 & n21213 ) ;
  assign n21214 = ( x2 & ~n21213 ) | ( x2 & n21211 ) | ( ~n21213 & n21211 ) ;
  assign n21216 = ( n21213 & ~n21215 ) | ( n21213 & n21214 ) | ( ~n21215 & n21214 ) ;
  assign n21220 = ( n21206 & ~n21219 ) | ( n21206 & n21216 ) | ( ~n21219 & n21216 ) ;
  assign n21224 = n10499 &  n20782 ;
  assign n21221 = ~n10015 & n20245 ;
  assign n21222 = ~n10486 & n20237 ;
  assign n21223 = n21221 | n21222 ;
  assign n21225 = ( n10499 & ~n21224 ) | ( n10499 & n21223 ) | ( ~n21224 & n21223 ) ;
  assign n21226 = ( n20237 & n20782 ) | ( n20237 & n20786 ) | ( n20782 & n20786 ) ;
  assign n21227 = ( n20782 & ~n21226 ) | ( n20782 & n20787 ) | ( ~n21226 & n20787 ) ;
  assign n21228 = ( n21225 & ~n10017 ) | ( n21225 & n21227 ) | ( ~n10017 & n21227 ) ;
  assign n21229 = n10017 | n21228 ;
  assign n21230 = ( x2 & ~n21225 ) | ( x2 & n21229 ) | ( ~n21225 & n21229 ) ;
  assign n21231 = ( n21225 & ~x2 ) | ( n21225 & n21229 ) | ( ~x2 & n21229 ) ;
  assign n21232 = ( n21230 & ~n21229 ) | ( n21230 & n21231 ) | ( ~n21229 & n21231 ) ;
  assign n21233 = ( n20287 & ~n20285 ) | ( n20287 & n20669 ) | ( ~n20285 & n20669 ) ;
  assign n21234 = ( n20285 & ~n20669 ) | ( n20285 & n20287 ) | ( ~n20669 & n20287 ) ;
  assign n21235 = ( n21233 & ~n20287 ) | ( n21233 & n21234 ) | ( ~n20287 & n21234 ) ;
  assign n21236 = ( n21220 & n21232 ) | ( n21220 & n21235 ) | ( n21232 & n21235 ) ;
  assign n21237 = ( n20677 & n20795 ) | ( n20677 & n21236 ) | ( n20795 & n21236 ) ;
  assign n21238 = ( n20687 & n20734 ) | ( n20687 & n20739 ) | ( n20734 & n20739 ) ;
  assign n21239 = ( n20742 & ~n20774 ) | ( n20742 & n20770 ) | ( ~n20774 & n20770 ) ;
  assign n21240 = ( x26 & ~n20700 ) | ( x26 & 1'b0 ) | ( ~n20700 & 1'b0 ) ;
  assign n21241 = ( n20695 & ~x26 ) | ( n20695 & n20700 ) | ( ~x26 & n20700 ) ;
  assign n21242 = ( n20696 & n21240 ) | ( n20696 & n21241 ) | ( n21240 & n21241 ) ;
  assign n21243 = ~n3644 & n14562 ;
  assign n21247 = n14553 | n3653 ;
  assign n21244 = ( n3652 & ~n14071 ) | ( n3652 & 1'b0 ) | ( ~n14071 & 1'b0 ) ;
  assign n21245 = ( n3657 & ~n14355 ) | ( n3657 & 1'b0 ) | ( ~n14355 & 1'b0 ) ;
  assign n21246 = n21244 | n21245 ;
  assign n21248 = ( n21247 & ~n3653 ) | ( n21247 & n21246 ) | ( ~n3653 & n21246 ) ;
  assign n21249 = n21243 | n21248 ;
  assign n21250 = n595 &  n837 ;
  assign n21251 = ( n602 & ~n20689 ) | ( n602 & n21250 ) | ( ~n20689 & n21250 ) ;
  assign n21252 = ~n602 & n21251 ;
  assign n21253 = ( n21242 & n21249 ) | ( n21242 & n21252 ) | ( n21249 & n21252 ) ;
  assign n21254 = ( n21249 & ~n21242 ) | ( n21249 & n21252 ) | ( ~n21242 & n21252 ) ;
  assign n21255 = ( n21242 & ~n21253 ) | ( n21242 & n21254 ) | ( ~n21253 & n21254 ) ;
  assign n21259 = n14800 | n4430 ;
  assign n21256 = n523 | n14803 ;
  assign n21257 = ~n3939 & n14807 ;
  assign n21258 = ( n21256 & ~n21257 ) | ( n21256 & 1'b0 ) | ( ~n21257 & 1'b0 ) ;
  assign n21260 = ( n4430 & ~n21259 ) | ( n4430 & n21258 ) | ( ~n21259 & n21258 ) ;
  assign n21261 = ( n14816 & ~n601 ) | ( n14816 & n21260 ) | ( ~n601 & n21260 ) ;
  assign n21262 = ~n14816 & n21261 ;
  assign n21263 = ( x29 & ~n21260 ) | ( x29 & n21262 ) | ( ~n21260 & n21262 ) ;
  assign n21264 = ( n21260 & ~x29 ) | ( n21260 & n21262 ) | ( ~x29 & n21262 ) ;
  assign n21265 = ( n21263 & ~n21262 ) | ( n21263 & n21264 ) | ( ~n21262 & n21264 ) ;
  assign n21266 = ( n20733 & ~n21255 ) | ( n20733 & n21265 ) | ( ~n21255 & n21265 ) ;
  assign n21267 = ( n20733 & ~n21265 ) | ( n20733 & n21255 ) | ( ~n21265 & n21255 ) ;
  assign n21268 = ( n21266 & ~n20733 ) | ( n21266 & n21267 ) | ( ~n20733 & n21267 ) ;
  assign n21270 = ( n21238 & n21239 ) | ( n21238 & n21268 ) | ( n21239 & n21268 ) ;
  assign n21269 = ( n21239 & ~n21238 ) | ( n21239 & n21268 ) | ( ~n21238 & n21268 ) ;
  assign n21271 = ( n21238 & ~n21270 ) | ( n21238 & n21269 ) | ( ~n21270 & n21269 ) ;
  assign n21277 = ( n20777 & n20789 ) | ( n20777 & n21271 ) | ( n20789 & n21271 ) ;
  assign n21278 = ( n20777 & ~n20789 ) | ( n20777 & n21271 ) | ( ~n20789 & n21271 ) ;
  assign n21279 = ( n20789 & ~n21277 ) | ( n20789 & n21278 ) | ( ~n21277 & n21278 ) ;
  assign n21272 = n10015 | n20782 ;
  assign n21273 = ~n10486 & n20777 ;
  assign n21274 = ( n21272 & ~n21273 ) | ( n21272 & 1'b0 ) | ( ~n21273 & 1'b0 ) ;
  assign n21275 = n10499 &  n21271 ;
  assign n21276 = ( n21274 & ~n10499 ) | ( n21274 & n21275 ) | ( ~n10499 & n21275 ) ;
  assign n21280 = ( n10017 & ~n21279 ) | ( n10017 & n21276 ) | ( ~n21279 & n21276 ) ;
  assign n21281 = ~n10017 & n21280 ;
  assign n21283 = ( x2 & n21276 ) | ( x2 & n21281 ) | ( n21276 & n21281 ) ;
  assign n21282 = ( x2 & ~n21281 ) | ( x2 & n21276 ) | ( ~n21281 & n21276 ) ;
  assign n21284 = ( n21281 & ~n21283 ) | ( n21281 & n21282 ) | ( ~n21283 & n21282 ) ;
  assign n21285 = ( n20674 & ~n21237 ) | ( n20674 & n21284 ) | ( ~n21237 & n21284 ) ;
  assign n21286 = ( n20674 & ~n21284 ) | ( n20674 & n21237 ) | ( ~n21284 & n21237 ) ;
  assign n21287 = ( n21285 & ~n20674 ) | ( n21285 & n21286 ) | ( ~n20674 & n21286 ) ;
  assign n21288 = ( n20677 & ~n20795 ) | ( n20677 & n21236 ) | ( ~n20795 & n21236 ) ;
  assign n21289 = ( n20795 & ~n21237 ) | ( n20795 & n21288 ) | ( ~n21237 & n21288 ) ;
  assign n21290 = n21287 | n21289 ;
  assign n21291 = ( n21287 & ~n21289 ) | ( n21287 & 1'b0 ) | ( ~n21289 & 1'b0 ) ;
  assign n21292 = ( n21290 & ~n21287 ) | ( n21290 & n21291 ) | ( ~n21287 & n21291 ) ;
  assign n21293 = n1345 | n2507 ;
  assign n21294 = ( n6735 & ~n2807 ) | ( n6735 & n21293 ) | ( ~n2807 & n21293 ) ;
  assign n21295 = n2807 | n21294 ;
  assign n21296 = ( n21295 & ~n6859 ) | ( n21295 & n16424 ) | ( ~n6859 & n16424 ) ;
  assign n21297 = n6859 | n21296 ;
  assign n21298 = ( n1184 & n21297 ) | ( n1184 & n1453 ) | ( n21297 & n1453 ) ;
  assign n21299 = ( n1453 & ~n21298 ) | ( n1453 & 1'b0 ) | ( ~n21298 & 1'b0 ) ;
  assign n21300 = ( n21299 & ~n865 ) | ( n21299 & n2484 ) | ( ~n865 & n2484 ) ;
  assign n21301 = ( n21300 & ~n2484 ) | ( n21300 & 1'b0 ) | ( ~n2484 & 1'b0 ) ;
  assign n21302 = ( n70 & n3212 ) | ( n70 & n21301 ) | ( n3212 & n21301 ) ;
  assign n21303 = ~n70 & n21302 ;
  assign n21304 = ( n127 & ~n352 ) | ( n127 & n21303 ) | ( ~n352 & n21303 ) ;
  assign n21305 = ~n127 & n21304 ;
  assign n21306 = ( n460 & ~n150 ) | ( n460 & n21305 ) | ( ~n150 & n21305 ) ;
  assign n21307 = ~n460 & n21306 ;
  assign n21308 = ( n80 & ~n21307 ) | ( n80 & n197 ) | ( ~n21307 & n197 ) ;
  assign n21309 = ( n197 & ~n21308 ) | ( n197 & 1'b0 ) | ( ~n21308 & 1'b0 ) ;
  assign n21310 = ~n358 & n21309 ;
  assign n21311 = ( n331 & ~n14755 ) | ( n331 & n14539 ) | ( ~n14755 & n14539 ) ;
  assign n21317 = n15361 | n3644 ;
  assign n21312 = n3653 | n15322 ;
  assign n21313 = n3657 &  n14745 ;
  assign n21314 = ( n3652 & ~n14528 ) | ( n3652 & 1'b0 ) | ( ~n14528 & 1'b0 ) ;
  assign n21315 = n21313 | n21314 ;
  assign n21316 = ( n21312 & ~n21315 ) | ( n21312 & 1'b0 ) | ( ~n21315 & 1'b0 ) ;
  assign n21318 = ( n3644 & ~n21317 ) | ( n3644 & n21316 ) | ( ~n21317 & n21316 ) ;
  assign n21319 = ( n21310 & ~n21311 ) | ( n21310 & n21318 ) | ( ~n21311 & n21318 ) ;
  assign n21320 = ( n21310 & ~n21318 ) | ( n21310 & n21311 ) | ( ~n21318 & n21311 ) ;
  assign n21321 = ( n21319 & ~n21310 ) | ( n21319 & n21320 ) | ( ~n21310 & n21320 ) ;
  assign n21322 = ( n15339 & ~n14758 ) | ( n15339 & n15426 ) | ( ~n14758 & n15426 ) ;
  assign n21326 = ~n4430 & n15700 ;
  assign n21323 = n523 | n15325 ;
  assign n21324 = n3939 | n15320 ;
  assign n21325 = n21323 &  n21324 ;
  assign n21327 = ( n4430 & n21326 ) | ( n4430 & n21325 ) | ( n21326 & n21325 ) ;
  assign n21328 = ( n15708 & ~n601 ) | ( n15708 & n21327 ) | ( ~n601 & n21327 ) ;
  assign n21329 = ~n15708 & n21328 ;
  assign n21331 = ( x29 & n21327 ) | ( x29 & n21329 ) | ( n21327 & n21329 ) ;
  assign n21330 = ( x29 & ~n21329 ) | ( x29 & n21327 ) | ( ~n21329 & n21327 ) ;
  assign n21332 = ( n21329 & ~n21331 ) | ( n21329 & n21330 ) | ( ~n21331 & n21330 ) ;
  assign n21333 = ( n21321 & ~n21322 ) | ( n21321 & n21332 ) | ( ~n21322 & n21332 ) ;
  assign n21334 = ( n21321 & ~n21332 ) | ( n21321 & n21322 ) | ( ~n21332 & n21322 ) ;
  assign n21335 = ( n21333 & ~n21321 ) | ( n21333 & n21334 ) | ( ~n21321 & n21334 ) ;
  assign n21340 = ~n4962 & n16591 ;
  assign n21337 = n4482 | n15897 ;
  assign n21338 = n4495 | n16091 ;
  assign n21339 = n21337 &  n21338 ;
  assign n21341 = ( n4962 & n21340 ) | ( n4962 & n21339 ) | ( n21340 & n21339 ) ;
  assign n21342 = ( n16631 & ~n4478 ) | ( n16631 & n21341 ) | ( ~n4478 & n21341 ) ;
  assign n21343 = ~n16631 & n21342 ;
  assign n21344 = ( x26 & ~n21341 ) | ( x26 & n21343 ) | ( ~n21341 & n21343 ) ;
  assign n21345 = ( n21341 & ~x26 ) | ( n21341 & n21343 ) | ( ~x26 & n21343 ) ;
  assign n21346 = ( n21344 & ~n21343 ) | ( n21344 & n21345 ) | ( ~n21343 & n21345 ) ;
  assign n21336 = ( n15911 & ~n15429 ) | ( n15911 & n16104 ) | ( ~n15429 & n16104 ) ;
  assign n21347 = ( n21335 & ~n21346 ) | ( n21335 & n21336 ) | ( ~n21346 & n21336 ) ;
  assign n21348 = ( n21335 & ~n21336 ) | ( n21335 & n21346 ) | ( ~n21336 & n21346 ) ;
  assign n21349 = ( n21347 & ~n21335 ) | ( n21347 & n21348 ) | ( ~n21335 & n21348 ) ;
  assign n21353 = n17107 | n5135 ;
  assign n21350 = n5010 | n16595 ;
  assign n21351 = n5067 | n16589 ;
  assign n21352 = n21350 &  n21351 ;
  assign n21354 = ( n5135 & ~n21353 ) | ( n5135 & n21352 ) | ( ~n21353 & n21352 ) ;
  assign n21355 = ~n5012 & n17115 ;
  assign n21356 = ( n21354 & ~n21355 ) | ( n21354 & 1'b0 ) | ( ~n21355 & 1'b0 ) ;
  assign n21357 = x23 &  n21356 ;
  assign n21358 = x23 | n21356 ;
  assign n21359 = ~n21357 & n21358 ;
  assign n21360 = ( n16609 & ~n16107 ) | ( n16609 & n16782 ) | ( ~n16107 & n16782 ) ;
  assign n21361 = ( n21349 & ~n21359 ) | ( n21349 & n21360 ) | ( ~n21359 & n21360 ) ;
  assign n21362 = ( n21349 & ~n21360 ) | ( n21349 & n21359 ) | ( ~n21360 & n21359 ) ;
  assign n21363 = ( n21361 & ~n21349 ) | ( n21361 & n21362 ) | ( ~n21349 & n21362 ) ;
  assign n21365 = ( n5339 & ~n17263 ) | ( n5339 & 1'b0 ) | ( ~n17263 & 1'b0 ) ;
  assign n21366 = n5761 | n17405 ;
  assign n21367 = ~n21365 & n21366 ;
  assign n21368 = ~n5837 & n17787 ;
  assign n21369 = ( n5837 & n21367 ) | ( n5837 & n21368 ) | ( n21367 & n21368 ) ;
  assign n21370 = ( n17826 & ~n5341 ) | ( n17826 & n21369 ) | ( ~n5341 & n21369 ) ;
  assign n21371 = ~n17826 & n21370 ;
  assign n21372 = ( x20 & ~n21369 ) | ( x20 & n21371 ) | ( ~n21369 & n21371 ) ;
  assign n21373 = ( n21369 & ~x20 ) | ( n21369 & n21371 ) | ( ~x20 & n21371 ) ;
  assign n21374 = ( n21372 & ~n21371 ) | ( n21372 & n21373 ) | ( ~n21371 & n21373 ) ;
  assign n21364 = ( n17277 & ~n16785 ) | ( n17277 & n17418 ) | ( ~n16785 & n17418 ) ;
  assign n21375 = ( n21363 & ~n21374 ) | ( n21363 & n21364 ) | ( ~n21374 & n21364 ) ;
  assign n21376 = ( n21363 & ~n21364 ) | ( n21363 & n21374 ) | ( ~n21364 & n21374 ) ;
  assign n21377 = ( n21375 & ~n21363 ) | ( n21375 & n21376 ) | ( ~n21363 & n21376 ) ;
  assign n21381 = ~n6395 & n18456 ;
  assign n21378 = n5970 | n17791 ;
  assign n21379 = n6170 | n17783 ;
  assign n21380 = n21378 &  n21379 ;
  assign n21382 = ( n6395 & n21381 ) | ( n6395 & n21380 ) | ( n21381 & n21380 ) ;
  assign n21383 = n5972 | n18464 ;
  assign n21384 = n21382 &  n21383 ;
  assign n21385 = x17 &  n21384 ;
  assign n21386 = x17 | n21384 ;
  assign n21387 = ~n21385 & n21386 ;
  assign n21388 = ( n17804 & ~n17421 ) | ( n17804 & n18057 ) | ( ~n17421 & n18057 ) ;
  assign n21389 = ( n21377 & ~n21387 ) | ( n21377 & n21388 ) | ( ~n21387 & n21388 ) ;
  assign n21390 = ( n21377 & ~n21388 ) | ( n21377 & n21387 ) | ( ~n21388 & n21387 ) ;
  assign n21391 = ( n21389 & ~n21377 ) | ( n21389 & n21390 ) | ( ~n21377 & n21390 ) ;
  assign n21396 = ~n7097 & n19043 ;
  assign n21393 = n6530 | n18589 ;
  assign n21394 = n6983 | n18712 ;
  assign n21395 = n21393 &  n21394 ;
  assign n21397 = ( n7097 & n21396 ) | ( n7097 & n21395 ) | ( n21396 & n21395 ) ;
  assign n21398 = ( n19083 & ~n6532 ) | ( n19083 & n21397 ) | ( ~n6532 & n21397 ) ;
  assign n21399 = ~n19083 & n21398 ;
  assign n21400 = ( x14 & ~n21397 ) | ( x14 & n21399 ) | ( ~n21397 & n21399 ) ;
  assign n21401 = ( n21397 & ~x14 ) | ( n21397 & n21399 ) | ( ~x14 & n21399 ) ;
  assign n21402 = ( n21400 & ~n21399 ) | ( n21400 & n21401 ) | ( ~n21399 & n21401 ) ;
  assign n21392 = ( n18603 & ~n18060 ) | ( n18603 & n18725 ) | ( ~n18060 & n18725 ) ;
  assign n21403 = ( n21391 & ~n21402 ) | ( n21391 & n21392 ) | ( ~n21402 & n21392 ) ;
  assign n21404 = ( n21391 & ~n21392 ) | ( n21391 & n21402 ) | ( ~n21392 & n21402 ) ;
  assign n21405 = ( n21403 & ~n21391 ) | ( n21403 & n21404 ) | ( ~n21391 & n21404 ) ;
  assign n21406 = n7253 &  n19047 ;
  assign n21407 = ~n7518 & n19040 ;
  assign n21408 = n21406 | n21407 ;
  assign n21409 = ~n7783 & n19494 ;
  assign n21410 = ( n7783 & ~n21408 ) | ( n7783 & n21409 ) | ( ~n21408 & n21409 ) ;
  assign n21411 = n7255 | n19502 ;
  assign n21412 = n21410 &  n21411 ;
  assign n21413 = x11 &  n21412 ;
  assign n21414 = x11 | n21412 ;
  assign n21415 = ~n21413 & n21414 ;
  assign n21416 = ( n19061 & ~n18728 ) | ( n19061 & n19394 ) | ( ~n18728 & n19394 ) ;
  assign n21417 = ( n21405 & ~n21415 ) | ( n21405 & n21416 ) | ( ~n21415 & n21416 ) ;
  assign n21418 = ( n21405 & ~n21416 ) | ( n21405 & n21415 ) | ( ~n21416 & n21415 ) ;
  assign n21419 = ( n21417 & ~n21405 ) | ( n21417 & n21418 ) | ( ~n21405 & n21418 ) ;
  assign n21424 = ~n8764 & n20241 ;
  assign n21421 = ( n8105 & ~n19951 ) | ( n8105 & 1'b0 ) | ( ~n19951 & 1'b0 ) ;
  assign n21422 = n8429 | n20027 ;
  assign n21423 = ~n21421 & n21422 ;
  assign n21425 = ( n8764 & n21424 ) | ( n8764 & n21423 ) | ( n21424 & n21423 ) ;
  assign n21426 = ( n20280 & ~n8107 ) | ( n20280 & n21425 ) | ( ~n8107 & n21425 ) ;
  assign n21427 = ~n20280 & n21426 ;
  assign n21428 = ( x8 & ~n21425 ) | ( x8 & n21427 ) | ( ~n21425 & n21427 ) ;
  assign n21429 = ( n21425 & ~x8 ) | ( n21425 & n21427 ) | ( ~x8 & n21427 ) ;
  assign n21430 = ( n21428 & ~n21427 ) | ( n21428 & n21429 ) | ( ~n21427 & n21429 ) ;
  assign n21420 = ( n19965 & ~n19397 ) | ( n19965 & n20040 ) | ( ~n19397 & n20040 ) ;
  assign n21431 = ( n21419 & ~n21430 ) | ( n21419 & n21420 ) | ( ~n21430 & n21420 ) ;
  assign n21432 = ( n21419 & ~n21420 ) | ( n21419 & n21430 ) | ( ~n21420 & n21430 ) ;
  assign n21433 = ( n21431 & ~n21419 ) | ( n21431 & n21432 ) | ( ~n21419 & n21432 ) ;
  assign n21434 = ~n9160 & n20245 ;
  assign n21435 = ~n9558 & n20237 ;
  assign n21436 = n21434 | n21435 ;
  assign n21437 = ~n9997 & n20782 ;
  assign n21438 = ( n9997 & ~n21436 ) | ( n9997 & n21437 ) | ( ~n21436 & n21437 ) ;
  assign n21439 = n9155 | n21227 ;
  assign n21440 = n21438 &  n21439 ;
  assign n21441 = x5 &  n21440 ;
  assign n21442 = x5 | n21440 ;
  assign n21443 = ~n21441 & n21442 ;
  assign n21444 = ( n20258 & ~n20043 ) | ( n20258 & n20671 ) | ( ~n20043 & n20671 ) ;
  assign n21445 = ( n21433 & ~n21443 ) | ( n21433 & n21444 ) | ( ~n21443 & n21444 ) ;
  assign n21446 = ( n21433 & ~n21444 ) | ( n21433 & n21443 ) | ( ~n21444 & n21443 ) ;
  assign n21447 = ( n21445 & ~n21433 ) | ( n21445 & n21446 ) | ( ~n21433 & n21446 ) ;
  assign n21476 = ~n10015 & n20777 ;
  assign n21477 = n10486 | n21271 ;
  assign n21478 = ~n21476 & n21477 ;
  assign n21449 = ( n20733 & n21255 ) | ( n20733 & n21265 ) | ( n21255 & n21265 ) ;
  assign n21450 = n3939 &  n4430 ;
  assign n21451 = ( n14800 & ~n21450 ) | ( n14800 & 1'b0 ) | ( ~n21450 & 1'b0 ) ;
  assign n21452 = ~n523 & n14807 ;
  assign n21453 = n21451 | n21452 ;
  assign n21454 = ~n601 & n15692 ;
  assign n21455 = n21453 | n21454 ;
  assign n21456 = ( x29 & ~n21455 ) | ( x29 & 1'b0 ) | ( ~n21455 & 1'b0 ) ;
  assign n21457 = ~x29 & n21455 ;
  assign n21458 = n21456 | n21457 ;
  assign n21463 = ~n3644 & n15310 ;
  assign n21464 = ( n3652 & ~n14355 ) | ( n3652 & 1'b0 ) | ( ~n14355 & 1'b0 ) ;
  assign n21465 = n3657 &  n14553 ;
  assign n21466 = n21464 | n21465 ;
  assign n21467 = ~n3653 & n14803 ;
  assign n21468 = ( n3653 & ~n21466 ) | ( n3653 & n21467 ) | ( ~n21466 & n21467 ) ;
  assign n21469 = ~n21463 & n21468 ;
  assign n21459 = n598 &  n662 ;
  assign n21460 = ( n21252 & ~n21459 ) | ( n21252 & n21254 ) | ( ~n21459 & n21254 ) ;
  assign n21461 = ( n21252 & ~n21254 ) | ( n21252 & n21459 ) | ( ~n21254 & n21459 ) ;
  assign n21462 = ( n21460 & ~n21252 ) | ( n21460 & n21461 ) | ( ~n21252 & n21461 ) ;
  assign n21470 = ( n21458 & ~n21469 ) | ( n21458 & n21462 ) | ( ~n21469 & n21462 ) ;
  assign n21471 = ( n21458 & ~n21462 ) | ( n21458 & n21469 ) | ( ~n21462 & n21469 ) ;
  assign n21472 = ( n21470 & ~n21458 ) | ( n21470 & n21471 ) | ( ~n21458 & n21471 ) ;
  assign n21474 = ( n21270 & n21449 ) | ( n21270 & n21472 ) | ( n21449 & n21472 ) ;
  assign n21473 = ( n21270 & ~n21449 ) | ( n21270 & n21472 ) | ( ~n21449 & n21472 ) ;
  assign n21475 = ( n21449 & ~n21474 ) | ( n21449 & n21473 ) | ( ~n21474 & n21473 ) ;
  assign n21479 = ( n10499 & ~n21475 ) | ( n10499 & 1'b0 ) | ( ~n21475 & 1'b0 ) ;
  assign n21480 = ( n21478 & ~n10499 ) | ( n21478 & n21479 ) | ( ~n10499 & n21479 ) ;
  assign n21481 = ( n20777 & ~n21271 ) | ( n20777 & n20789 ) | ( ~n21271 & n20789 ) ;
  assign n21483 = ( n21271 & n21475 ) | ( n21271 & n21481 ) | ( n21475 & n21481 ) ;
  assign n21482 = ( n21271 & ~n21481 ) | ( n21271 & n21475 ) | ( ~n21481 & n21475 ) ;
  assign n21484 = ( n21481 & ~n21483 ) | ( n21481 & n21482 ) | ( ~n21483 & n21482 ) ;
  assign n21485 = ( n10017 & ~n21484 ) | ( n10017 & n21480 ) | ( ~n21484 & n21480 ) ;
  assign n21486 = ~n10017 & n21485 ;
  assign n21487 = ( x2 & ~n21480 ) | ( x2 & n21486 ) | ( ~n21480 & n21486 ) ;
  assign n21488 = ( n21480 & ~x2 ) | ( n21480 & n21486 ) | ( ~x2 & n21486 ) ;
  assign n21489 = ( n21487 & ~n21486 ) | ( n21487 & n21488 ) | ( ~n21486 & n21488 ) ;
  assign n21448 = ( n21237 & ~n20674 ) | ( n21237 & n21284 ) | ( ~n20674 & n21284 ) ;
  assign n21490 = ( n21447 & ~n21489 ) | ( n21447 & n21448 ) | ( ~n21489 & n21448 ) ;
  assign n21491 = ( n21447 & ~n21448 ) | ( n21447 & n21489 ) | ( ~n21448 & n21489 ) ;
  assign n21492 = ( n21490 & ~n21447 ) | ( n21490 & n21491 ) | ( ~n21447 & n21491 ) ;
  assign n21493 = ( n21291 & ~n21492 ) | ( n21291 & 1'b0 ) | ( ~n21492 & 1'b0 ) ;
  assign n21494 = ~n21291 & n21492 ;
  assign n21495 = n21493 | n21494 ;
  assign n21496 = n15927 | n17187 ;
  assign n21497 = ( n6821 & ~n3214 ) | ( n6821 & n21496 ) | ( ~n3214 & n21496 ) ;
  assign n21498 = n3214 | n21497 ;
  assign n21499 = ( n1702 & ~n21498 ) | ( n1702 & n4359 ) | ( ~n21498 & n4359 ) ;
  assign n21500 = ~n1702 & n21499 ;
  assign n21501 = ( n2506 & n4370 ) | ( n2506 & n21500 ) | ( n4370 & n21500 ) ;
  assign n21502 = ~n2506 & n21501 ;
  assign n21503 = ( n886 & ~n2718 ) | ( n886 & n21502 ) | ( ~n2718 & n21502 ) ;
  assign n21504 = ~n886 & n21503 ;
  assign n21505 = ( n906 & ~n779 ) | ( n906 & n21504 ) | ( ~n779 & n21504 ) ;
  assign n21506 = ~n906 & n21505 ;
  assign n21507 = ( n457 & ~n346 ) | ( n457 & n21506 ) | ( ~n346 & n21506 ) ;
  assign n21508 = ~n457 & n21507 ;
  assign n21509 = ( n255 & ~n404 ) | ( n255 & n21508 ) | ( ~n404 & n21508 ) ;
  assign n21510 = ~n255 & n21509 ;
  assign n21511 = ( n205 & ~n149 ) | ( n205 & n21510 ) | ( ~n149 & n21510 ) ;
  assign n21512 = ~n205 & n21511 ;
  assign n21513 = ( n21310 & n21311 ) | ( n21310 & n21318 ) | ( n21311 & n21318 ) ;
  assign n21519 = ~n3644 & n15346 ;
  assign n21514 = n3653 | n15325 ;
  assign n21515 = ( n3657 & ~n15322 ) | ( n3657 & 1'b0 ) | ( ~n15322 & 1'b0 ) ;
  assign n21516 = n3652 &  n14745 ;
  assign n21517 = n21515 | n21516 ;
  assign n21518 = ( n21514 & ~n21517 ) | ( n21514 & 1'b0 ) | ( ~n21517 & 1'b0 ) ;
  assign n21520 = ( n3644 & n21519 ) | ( n3644 & n21518 ) | ( n21519 & n21518 ) ;
  assign n21521 = ( n21512 & ~n21513 ) | ( n21512 & n21520 ) | ( ~n21513 & n21520 ) ;
  assign n21522 = ( n21512 & ~n21520 ) | ( n21512 & n21513 ) | ( ~n21520 & n21513 ) ;
  assign n21523 = ( n21521 & ~n21512 ) | ( n21521 & n21522 ) | ( ~n21512 & n21522 ) ;
  assign n21524 = ( n21321 & n21322 ) | ( n21321 & n21332 ) | ( n21322 & n21332 ) ;
  assign n21528 = ~n4430 & n15897 ;
  assign n21525 = n523 | n15320 ;
  assign n21526 = n3939 | n15700 ;
  assign n21527 = n21525 &  n21526 ;
  assign n21529 = ( n4430 & n21528 ) | ( n4430 & n21527 ) | ( n21528 & n21527 ) ;
  assign n21530 = ( n15900 & ~n601 ) | ( n15900 & n21529 ) | ( ~n601 & n21529 ) ;
  assign n21531 = ~n15900 & n21530 ;
  assign n21532 = ( x29 & ~n21529 ) | ( x29 & n21531 ) | ( ~n21529 & n21531 ) ;
  assign n21533 = ( n21529 & ~x29 ) | ( n21529 & n21531 ) | ( ~x29 & n21531 ) ;
  assign n21534 = ( n21532 & ~n21531 ) | ( n21532 & n21533 ) | ( ~n21531 & n21533 ) ;
  assign n21535 = ( n21523 & ~n21524 ) | ( n21523 & n21534 ) | ( ~n21524 & n21534 ) ;
  assign n21536 = ( n21523 & ~n21534 ) | ( n21523 & n21524 ) | ( ~n21534 & n21524 ) ;
  assign n21537 = ( n21535 & ~n21523 ) | ( n21535 & n21536 ) | ( ~n21523 & n21536 ) ;
  assign n21542 = ~n4962 & n16595 ;
  assign n21539 = n4482 | n16091 ;
  assign n21540 = n4495 | n16591 ;
  assign n21541 = n21539 &  n21540 ;
  assign n21543 = ( n4962 & n21542 ) | ( n4962 & n21541 ) | ( n21542 & n21541 ) ;
  assign n21544 = ( n16616 & ~n4478 ) | ( n16616 & n21543 ) | ( ~n4478 & n21543 ) ;
  assign n21545 = ~n16616 & n21544 ;
  assign n21547 = ( x26 & n21543 ) | ( x26 & n21545 ) | ( n21543 & n21545 ) ;
  assign n21546 = ( x26 & ~n21545 ) | ( x26 & n21543 ) | ( ~n21545 & n21543 ) ;
  assign n21548 = ( n21545 & ~n21547 ) | ( n21545 & n21546 ) | ( ~n21547 & n21546 ) ;
  assign n21538 = ( n21335 & n21336 ) | ( n21335 & n21346 ) | ( n21336 & n21346 ) ;
  assign n21549 = ( n21537 & ~n21548 ) | ( n21537 & n21538 ) | ( ~n21548 & n21538 ) ;
  assign n21550 = ( n21537 & ~n21538 ) | ( n21537 & n21548 ) | ( ~n21538 & n21548 ) ;
  assign n21551 = ( n21549 & ~n21537 ) | ( n21549 & n21550 ) | ( ~n21537 & n21550 ) ;
  assign n21555 = ~n5135 & n17263 ;
  assign n21552 = n5010 | n16589 ;
  assign n21553 = ~n5067 & n17107 ;
  assign n21554 = ( n21552 & ~n21553 ) | ( n21552 & 1'b0 ) | ( ~n21553 & 1'b0 ) ;
  assign n21556 = ( n5135 & n21555 ) | ( n5135 & n21554 ) | ( n21555 & n21554 ) ;
  assign n21557 = ~n5012 & n17271 ;
  assign n21558 = ( n21556 & ~n21557 ) | ( n21556 & 1'b0 ) | ( ~n21557 & 1'b0 ) ;
  assign n21559 = x23 &  n21558 ;
  assign n21560 = x23 | n21558 ;
  assign n21561 = ~n21559 & n21560 ;
  assign n21562 = ( n21349 & n21359 ) | ( n21349 & n21360 ) | ( n21359 & n21360 ) ;
  assign n21563 = ( n21551 & ~n21561 ) | ( n21551 & n21562 ) | ( ~n21561 & n21562 ) ;
  assign n21564 = ( n21551 & ~n21562 ) | ( n21551 & n21561 ) | ( ~n21562 & n21561 ) ;
  assign n21565 = ( n21563 & ~n21551 ) | ( n21563 & n21564 ) | ( ~n21551 & n21564 ) ;
  assign n21570 = ~n5837 & n17791 ;
  assign n21567 = ( n5339 & ~n17405 ) | ( n5339 & 1'b0 ) | ( ~n17405 & 1'b0 ) ;
  assign n21568 = n5761 | n17787 ;
  assign n21569 = ~n21567 & n21568 ;
  assign n21571 = ( n5837 & n21570 ) | ( n5837 & n21569 ) | ( n21570 & n21569 ) ;
  assign n21572 = ( n17811 & ~n5341 ) | ( n17811 & n21571 ) | ( ~n5341 & n21571 ) ;
  assign n21573 = ~n17811 & n21572 ;
  assign n21575 = ( x20 & n21571 ) | ( x20 & n21573 ) | ( n21571 & n21573 ) ;
  assign n21574 = ( x20 & ~n21573 ) | ( x20 & n21571 ) | ( ~n21573 & n21571 ) ;
  assign n21576 = ( n21573 & ~n21575 ) | ( n21573 & n21574 ) | ( ~n21575 & n21574 ) ;
  assign n21566 = ( n21363 & n21364 ) | ( n21363 & n21374 ) | ( n21364 & n21374 ) ;
  assign n21577 = ( n21565 & ~n21576 ) | ( n21565 & n21566 ) | ( ~n21576 & n21566 ) ;
  assign n21578 = ( n21565 & ~n21566 ) | ( n21565 & n21576 ) | ( ~n21566 & n21576 ) ;
  assign n21579 = ( n21577 & ~n21565 ) | ( n21577 & n21578 ) | ( ~n21565 & n21578 ) ;
  assign n21583 = ~n6395 & n18589 ;
  assign n21580 = n5970 | n17783 ;
  assign n21581 = n6170 | n18456 ;
  assign n21582 = n21580 &  n21581 ;
  assign n21584 = ( n6395 & n21583 ) | ( n6395 & n21582 ) | ( n21583 & n21582 ) ;
  assign n21585 = n5972 | n18597 ;
  assign n21586 = n21584 &  n21585 ;
  assign n21587 = x17 &  n21586 ;
  assign n21588 = x17 | n21586 ;
  assign n21589 = ~n21587 & n21588 ;
  assign n21590 = ( n21377 & n21387 ) | ( n21377 & n21388 ) | ( n21387 & n21388 ) ;
  assign n21591 = ( n21579 & ~n21589 ) | ( n21579 & n21590 ) | ( ~n21589 & n21590 ) ;
  assign n21592 = ( n21579 & ~n21590 ) | ( n21579 & n21589 ) | ( ~n21590 & n21589 ) ;
  assign n21593 = ( n21591 & ~n21579 ) | ( n21591 & n21592 ) | ( ~n21579 & n21592 ) ;
  assign n21598 = n19047 | n7097 ;
  assign n21595 = n6530 | n18712 ;
  assign n21596 = n6983 | n19043 ;
  assign n21597 = n21595 &  n21596 ;
  assign n21599 = ( n7097 & ~n21598 ) | ( n7097 & n21597 ) | ( ~n21598 & n21597 ) ;
  assign n21600 = ( n6532 & ~n21599 ) | ( n6532 & n19068 ) | ( ~n21599 & n19068 ) ;
  assign n21601 = ( n19068 & ~n21600 ) | ( n19068 & 1'b0 ) | ( ~n21600 & 1'b0 ) ;
  assign n21603 = ( x14 & n21599 ) | ( x14 & n21601 ) | ( n21599 & n21601 ) ;
  assign n21602 = ( x14 & ~n21601 ) | ( x14 & n21599 ) | ( ~n21601 & n21599 ) ;
  assign n21604 = ( n21601 & ~n21603 ) | ( n21601 & n21602 ) | ( ~n21603 & n21602 ) ;
  assign n21594 = ( n21391 & n21392 ) | ( n21391 & n21402 ) | ( n21392 & n21402 ) ;
  assign n21605 = ( n21593 & ~n21604 ) | ( n21593 & n21594 ) | ( ~n21604 & n21594 ) ;
  assign n21606 = ( n21593 & ~n21594 ) | ( n21593 & n21604 ) | ( ~n21594 & n21604 ) ;
  assign n21607 = ( n21605 & ~n21593 ) | ( n21605 & n21606 ) | ( ~n21593 & n21606 ) ;
  assign n21611 = ~n7783 & n19951 ;
  assign n21608 = n7253 &  n19040 ;
  assign n21609 = n7518 | n19494 ;
  assign n21610 = ~n21608 & n21609 ;
  assign n21612 = ( n7783 & n21611 ) | ( n7783 & n21610 ) | ( n21611 & n21610 ) ;
  assign n21613 = ~n7255 & n19959 ;
  assign n21614 = ( n21612 & ~n21613 ) | ( n21612 & 1'b0 ) | ( ~n21613 & 1'b0 ) ;
  assign n21615 = x11 &  n21614 ;
  assign n21616 = x11 | n21614 ;
  assign n21617 = ~n21615 & n21616 ;
  assign n21618 = ( n21405 & n21415 ) | ( n21405 & n21416 ) | ( n21415 & n21416 ) ;
  assign n21619 = ( n21607 & ~n21617 ) | ( n21607 & n21618 ) | ( ~n21617 & n21618 ) ;
  assign n21620 = ( n21607 & ~n21618 ) | ( n21607 & n21617 ) | ( ~n21618 & n21617 ) ;
  assign n21621 = ( n21619 & ~n21607 ) | ( n21619 & n21620 ) | ( ~n21607 & n21620 ) ;
  assign n21626 = n20245 | n8764 ;
  assign n21623 = ( n8105 & ~n20027 ) | ( n8105 & 1'b0 ) | ( ~n20027 & 1'b0 ) ;
  assign n21624 = n8429 | n20241 ;
  assign n21625 = ~n21623 & n21624 ;
  assign n21627 = ( n8764 & ~n21626 ) | ( n8764 & n21625 ) | ( ~n21626 & n21625 ) ;
  assign n21628 = ( n8107 & ~n21627 ) | ( n8107 & n20265 ) | ( ~n21627 & n20265 ) ;
  assign n21629 = ( n20265 & ~n21628 ) | ( n20265 & 1'b0 ) | ( ~n21628 & 1'b0 ) ;
  assign n21631 = ( x8 & n21627 ) | ( x8 & n21629 ) | ( n21627 & n21629 ) ;
  assign n21630 = ( x8 & ~n21629 ) | ( x8 & n21627 ) | ( ~n21629 & n21627 ) ;
  assign n21632 = ( n21629 & ~n21631 ) | ( n21629 & n21630 ) | ( ~n21631 & n21630 ) ;
  assign n21622 = ( n21419 & n21420 ) | ( n21419 & n21430 ) | ( n21420 & n21430 ) ;
  assign n21633 = ( n21621 & ~n21632 ) | ( n21621 & n21622 ) | ( ~n21632 & n21622 ) ;
  assign n21634 = ( n21621 & ~n21622 ) | ( n21621 & n21632 ) | ( ~n21622 & n21632 ) ;
  assign n21635 = ( n21633 & ~n21621 ) | ( n21633 & n21634 ) | ( ~n21621 & n21634 ) ;
  assign n21636 = n9997 &  n20777 ;
  assign n21637 = ~n9160 & n20237 ;
  assign n21638 = n9558 | n20782 ;
  assign n21639 = ~n21637 & n21638 ;
  assign n21640 = ( n21636 & ~n20777 ) | ( n21636 & n21639 ) | ( ~n20777 & n21639 ) ;
  assign n21641 = n9155 | n20790 ;
  assign n21642 = n21640 &  n21641 ;
  assign n21643 = x5 &  n21642 ;
  assign n21644 = x5 | n21642 ;
  assign n21645 = ~n21643 & n21644 ;
  assign n21646 = ( n21433 & n21443 ) | ( n21433 & n21444 ) | ( n21443 & n21444 ) ;
  assign n21647 = ( n21635 & ~n21645 ) | ( n21635 & n21646 ) | ( ~n21645 & n21646 ) ;
  assign n21648 = ( n21635 & ~n21646 ) | ( n21635 & n21645 ) | ( ~n21646 & n21645 ) ;
  assign n21649 = ( n21647 & ~n21635 ) | ( n21647 & n21648 ) | ( ~n21635 & n21648 ) ;
  assign n21676 = n10015 | n21271 ;
  assign n21677 = ~n10486 & n21475 ;
  assign n21678 = ( n21676 & ~n21677 ) | ( n21676 & 1'b0 ) | ( ~n21677 & 1'b0 ) ;
  assign n21651 = ( n21462 & ~n21458 ) | ( n21462 & n21469 ) | ( ~n21458 & n21469 ) ;
  assign n21652 = ( n21270 & ~n21472 ) | ( n21270 & n21449 ) | ( ~n21472 & n21449 ) ;
  assign n21653 = n14795 &  n21459 ;
  assign n21654 = n14795 | n21459 ;
  assign n21655 = ~n21653 & n21654 ;
  assign n21656 = ( n515 & ~n518 ) | ( n515 & n521 ) | ( ~n518 & n521 ) ;
  assign n21657 = n518 | n21656 ;
  assign n21658 = n14800 &  n21657 ;
  assign n21659 = ( x29 & n21655 ) | ( x29 & n21658 ) | ( n21655 & n21658 ) ;
  assign n21660 = ( n21655 & ~x29 ) | ( n21655 & n21658 ) | ( ~x29 & n21658 ) ;
  assign n21661 = ( x29 & ~n21659 ) | ( x29 & n21660 ) | ( ~n21659 & n21660 ) ;
  assign n21662 = ( n21254 & ~n21252 ) | ( n21254 & n21459 ) | ( ~n21252 & n21459 ) ;
  assign n21663 = ~n3644 & n15294 ;
  assign n21664 = n3652 &  n14553 ;
  assign n21665 = ( n3657 & ~n14803 ) | ( n3657 & 1'b0 ) | ( ~n14803 & 1'b0 ) ;
  assign n21666 = n21664 | n21665 ;
  assign n21667 = n3653 | n14807 ;
  assign n21668 = ( n21666 & ~n3653 ) | ( n21666 & n21667 ) | ( ~n3653 & n21667 ) ;
  assign n21669 = n21663 | n21668 ;
  assign n21670 = ( n21661 & ~n21662 ) | ( n21661 & n21669 ) | ( ~n21662 & n21669 ) ;
  assign n21671 = ( n21662 & ~n21661 ) | ( n21662 & n21669 ) | ( ~n21661 & n21669 ) ;
  assign n21672 = ( n21670 & ~n21669 ) | ( n21670 & n21671 ) | ( ~n21669 & n21671 ) ;
  assign n21673 = ( n21652 & ~n21651 ) | ( n21652 & n21672 ) | ( ~n21651 & n21672 ) ;
  assign n21674 = ( n21651 & n21652 ) | ( n21651 & n21672 ) | ( n21652 & n21672 ) ;
  assign n21675 = ( n21651 & n21673 ) | ( n21651 & ~n21674 ) | ( n21673 & ~n21674 ) ;
  assign n21679 = n10499 &  n21675 ;
  assign n21680 = ( n21678 & ~n10499 ) | ( n21678 & n21679 ) | ( ~n10499 & n21679 ) ;
  assign n21681 = ( n21475 & ~n21271 ) | ( n21475 & n21481 ) | ( ~n21271 & n21481 ) ;
  assign n21682 = ( n21475 & n21675 ) | ( n21475 & n21681 ) | ( n21675 & n21681 ) ;
  assign n21683 = ( n21475 & ~n21675 ) | ( n21475 & n21681 ) | ( ~n21675 & n21681 ) ;
  assign n21684 = ( n21675 & ~n21682 ) | ( n21675 & n21683 ) | ( ~n21682 & n21683 ) ;
  assign n21685 = ( n10017 & ~n21684 ) | ( n10017 & n21680 ) | ( ~n21684 & n21680 ) ;
  assign n21686 = ~n10017 & n21685 ;
  assign n21687 = ( x2 & ~n21680 ) | ( x2 & n21686 ) | ( ~n21680 & n21686 ) ;
  assign n21688 = ( n21680 & ~x2 ) | ( n21680 & n21686 ) | ( ~x2 & n21686 ) ;
  assign n21689 = ( n21687 & ~n21686 ) | ( n21687 & n21688 ) | ( ~n21686 & n21688 ) ;
  assign n21650 = ( n21447 & n21448 ) | ( n21447 & n21489 ) | ( n21448 & n21489 ) ;
  assign n21690 = ( n21649 & ~n21689 ) | ( n21649 & n21650 ) | ( ~n21689 & n21650 ) ;
  assign n21691 = ( n21649 & ~n21650 ) | ( n21649 & n21689 ) | ( ~n21650 & n21689 ) ;
  assign n21692 = ( n21690 & ~n21649 ) | ( n21690 & n21691 ) | ( ~n21649 & n21691 ) ;
  assign n21693 = ( n21493 & ~n21692 ) | ( n21493 & 1'b0 ) | ( ~n21692 & 1'b0 ) ;
  assign n21694 = ~n21493 & n21692 ;
  assign n21695 = n21693 | n21694 ;
  assign n21696 = n1152 | n1426 ;
  assign n21697 = n766 | n21696 ;
  assign n21698 = ( n2571 & ~n2631 ) | ( n2571 & 1'b0 ) | ( ~n2631 & 1'b0 ) ;
  assign n21699 = ( n3214 & ~n21697 ) | ( n3214 & n21698 ) | ( ~n21697 & n21698 ) ;
  assign n21700 = ~n3214 & n21699 ;
  assign n21701 = ( n5196 & n15594 ) | ( n5196 & n21700 ) | ( n15594 & n21700 ) ;
  assign n21702 = ~n5196 & n21701 ;
  assign n21703 = ( n4166 & ~n6836 ) | ( n4166 & n21702 ) | ( ~n6836 & n21702 ) ;
  assign n21704 = n6836 &  n21703 ;
  assign n21705 = ( n1626 & ~n3059 ) | ( n1626 & n21704 ) | ( ~n3059 & n21704 ) ;
  assign n21706 = ~n1626 & n21705 ;
  assign n21707 = ( n1061 & ~n1245 ) | ( n1061 & n21706 ) | ( ~n1245 & n21706 ) ;
  assign n21708 = ~n1061 & n21707 ;
  assign n21709 = ( n334 & ~n21708 ) | ( n334 & n343 ) | ( ~n21708 & n343 ) ;
  assign n21710 = ( n343 & ~n21709 ) | ( n343 & 1'b0 ) | ( ~n21709 & 1'b0 ) ;
  assign n21711 = ( n21512 & n21513 ) | ( n21512 & n21520 ) | ( n21513 & n21520 ) ;
  assign n21717 = ~n3644 & n15334 ;
  assign n21712 = n3653 | n15320 ;
  assign n21713 = ( n3657 & ~n15325 ) | ( n3657 & 1'b0 ) | ( ~n15325 & 1'b0 ) ;
  assign n21714 = ( n3652 & ~n15322 ) | ( n3652 & 1'b0 ) | ( ~n15322 & 1'b0 ) ;
  assign n21715 = n21713 | n21714 ;
  assign n21716 = ( n21712 & ~n21715 ) | ( n21712 & 1'b0 ) | ( ~n21715 & 1'b0 ) ;
  assign n21718 = ( n3644 & n21717 ) | ( n3644 & n21716 ) | ( n21717 & n21716 ) ;
  assign n21719 = ( n21710 & ~n21711 ) | ( n21710 & n21718 ) | ( ~n21711 & n21718 ) ;
  assign n21720 = ( n21710 & ~n21718 ) | ( n21710 & n21711 ) | ( ~n21718 & n21711 ) ;
  assign n21721 = ( n21719 & ~n21710 ) | ( n21719 & n21720 ) | ( ~n21710 & n21720 ) ;
  assign n21722 = ( n21523 & n21524 ) | ( n21523 & n21534 ) | ( n21524 & n21534 ) ;
  assign n21726 = ~n4430 & n16091 ;
  assign n21723 = n523 | n15700 ;
  assign n21724 = n3939 | n15897 ;
  assign n21725 = n21723 &  n21724 ;
  assign n21727 = ( n4430 & n21726 ) | ( n4430 & n21725 ) | ( n21726 & n21725 ) ;
  assign n21728 = ( n16094 & ~n601 ) | ( n16094 & n21727 ) | ( ~n601 & n21727 ) ;
  assign n21729 = ~n16094 & n21728 ;
  assign n21730 = ( x29 & ~n21727 ) | ( x29 & n21729 ) | ( ~n21727 & n21729 ) ;
  assign n21731 = ( n21727 & ~x29 ) | ( n21727 & n21729 ) | ( ~x29 & n21729 ) ;
  assign n21732 = ( n21730 & ~n21729 ) | ( n21730 & n21731 ) | ( ~n21729 & n21731 ) ;
  assign n21733 = ( n21721 & ~n21722 ) | ( n21721 & n21732 ) | ( ~n21722 & n21732 ) ;
  assign n21734 = ( n21721 & ~n21732 ) | ( n21721 & n21722 ) | ( ~n21732 & n21722 ) ;
  assign n21735 = ( n21733 & ~n21721 ) | ( n21733 & n21734 ) | ( ~n21721 & n21734 ) ;
  assign n21740 = ~n4962 & n16589 ;
  assign n21737 = n4482 | n16591 ;
  assign n21738 = n4495 | n16595 ;
  assign n21739 = n21737 &  n21738 ;
  assign n21741 = ( n4962 & n21740 ) | ( n4962 & n21739 ) | ( n21740 & n21739 ) ;
  assign n21742 = ( n16604 & ~n4478 ) | ( n16604 & n21741 ) | ( ~n4478 & n21741 ) ;
  assign n21743 = ~n16604 & n21742 ;
  assign n21745 = ( x26 & n21741 ) | ( x26 & n21743 ) | ( n21741 & n21743 ) ;
  assign n21744 = ( x26 & ~n21743 ) | ( x26 & n21741 ) | ( ~n21743 & n21741 ) ;
  assign n21746 = ( n21743 & ~n21745 ) | ( n21743 & n21744 ) | ( ~n21745 & n21744 ) ;
  assign n21736 = ( n21537 & n21538 ) | ( n21537 & n21548 ) | ( n21538 & n21548 ) ;
  assign n21747 = ( n21735 & ~n21746 ) | ( n21735 & n21736 ) | ( ~n21746 & n21736 ) ;
  assign n21748 = ( n21735 & ~n21736 ) | ( n21735 & n21746 ) | ( ~n21736 & n21746 ) ;
  assign n21749 = ( n21747 & ~n21735 ) | ( n21747 & n21748 ) | ( ~n21735 & n21748 ) ;
  assign n21753 = ~n5135 & n17405 ;
  assign n21750 = ~n5010 & n17107 ;
  assign n21751 = n5067 | n17263 ;
  assign n21752 = ~n21750 & n21751 ;
  assign n21754 = ( n5135 & n21753 ) | ( n5135 & n21752 ) | ( n21753 & n21752 ) ;
  assign n21755 = n5012 | n17413 ;
  assign n21756 = n21754 &  n21755 ;
  assign n21757 = x23 &  n21756 ;
  assign n21758 = x23 | n21756 ;
  assign n21759 = ~n21757 & n21758 ;
  assign n21760 = ( n21551 & n21561 ) | ( n21551 & n21562 ) | ( n21561 & n21562 ) ;
  assign n21761 = ( n21749 & ~n21759 ) | ( n21749 & n21760 ) | ( ~n21759 & n21760 ) ;
  assign n21762 = ( n21749 & ~n21760 ) | ( n21749 & n21759 ) | ( ~n21760 & n21759 ) ;
  assign n21763 = ( n21761 & ~n21749 ) | ( n21761 & n21762 ) | ( ~n21749 & n21762 ) ;
  assign n21768 = ~n5837 & n17783 ;
  assign n21765 = ( n5339 & ~n17787 ) | ( n5339 & 1'b0 ) | ( ~n17787 & 1'b0 ) ;
  assign n21766 = n5761 | n17791 ;
  assign n21767 = ~n21765 & n21766 ;
  assign n21769 = ( n5837 & n21768 ) | ( n5837 & n21767 ) | ( n21768 & n21767 ) ;
  assign n21770 = ( n17799 & ~n5341 ) | ( n17799 & n21769 ) | ( ~n5341 & n21769 ) ;
  assign n21771 = ~n17799 & n21770 ;
  assign n21773 = ( x20 & n21769 ) | ( x20 & n21771 ) | ( n21769 & n21771 ) ;
  assign n21772 = ( x20 & ~n21771 ) | ( x20 & n21769 ) | ( ~n21771 & n21769 ) ;
  assign n21774 = ( n21771 & ~n21773 ) | ( n21771 & n21772 ) | ( ~n21773 & n21772 ) ;
  assign n21764 = ( n21565 & n21566 ) | ( n21565 & n21576 ) | ( n21566 & n21576 ) ;
  assign n21775 = ( n21763 & ~n21774 ) | ( n21763 & n21764 ) | ( ~n21774 & n21764 ) ;
  assign n21776 = ( n21763 & ~n21764 ) | ( n21763 & n21774 ) | ( ~n21764 & n21774 ) ;
  assign n21777 = ( n21775 & ~n21763 ) | ( n21775 & n21776 ) | ( ~n21763 & n21776 ) ;
  assign n21781 = ~n6395 & n18712 ;
  assign n21778 = n5970 | n18456 ;
  assign n21779 = n6170 | n18589 ;
  assign n21780 = n21778 &  n21779 ;
  assign n21782 = ( n6395 & n21781 ) | ( n6395 & n21780 ) | ( n21781 & n21780 ) ;
  assign n21783 = n5972 | n18720 ;
  assign n21784 = n21782 &  n21783 ;
  assign n21785 = x17 &  n21784 ;
  assign n21786 = x17 | n21784 ;
  assign n21787 = ~n21785 & n21786 ;
  assign n21788 = ( n21579 & n21589 ) | ( n21579 & n21590 ) | ( n21589 & n21590 ) ;
  assign n21789 = ( n21777 & ~n21787 ) | ( n21777 & n21788 ) | ( ~n21787 & n21788 ) ;
  assign n21790 = ( n21777 & ~n21788 ) | ( n21777 & n21787 ) | ( ~n21788 & n21787 ) ;
  assign n21791 = ( n21789 & ~n21777 ) | ( n21789 & n21790 ) | ( ~n21777 & n21790 ) ;
  assign n21796 = n19040 | n7097 ;
  assign n21793 = n6530 | n19043 ;
  assign n21794 = ~n6983 & n19047 ;
  assign n21795 = ( n21793 & ~n21794 ) | ( n21793 & 1'b0 ) | ( ~n21794 & 1'b0 ) ;
  assign n21797 = ( n7097 & ~n21796 ) | ( n7097 & n21795 ) | ( ~n21796 & n21795 ) ;
  assign n21798 = ( n19056 & ~n6532 ) | ( n19056 & n21797 ) | ( ~n6532 & n21797 ) ;
  assign n21799 = ~n19056 & n21798 ;
  assign n21801 = ( x14 & n21797 ) | ( x14 & n21799 ) | ( n21797 & n21799 ) ;
  assign n21800 = ( x14 & ~n21799 ) | ( x14 & n21797 ) | ( ~n21799 & n21797 ) ;
  assign n21802 = ( n21799 & ~n21801 ) | ( n21799 & n21800 ) | ( ~n21801 & n21800 ) ;
  assign n21792 = ( n21593 & n21594 ) | ( n21593 & n21604 ) | ( n21594 & n21604 ) ;
  assign n21803 = ( n21791 & ~n21802 ) | ( n21791 & n21792 ) | ( ~n21802 & n21792 ) ;
  assign n21804 = ( n21791 & ~n21792 ) | ( n21791 & n21802 ) | ( ~n21792 & n21802 ) ;
  assign n21805 = ( n21803 & ~n21791 ) | ( n21803 & n21804 ) | ( ~n21791 & n21804 ) ;
  assign n21809 = ~n7783 & n20027 ;
  assign n21806 = ( n7253 & ~n19494 ) | ( n7253 & 1'b0 ) | ( ~n19494 & 1'b0 ) ;
  assign n21807 = n7518 | n19951 ;
  assign n21808 = ~n21806 & n21807 ;
  assign n21810 = ( n7783 & n21809 ) | ( n7783 & n21808 ) | ( n21809 & n21808 ) ;
  assign n21811 = n7255 | n20035 ;
  assign n21812 = n21810 &  n21811 ;
  assign n21813 = x11 &  n21812 ;
  assign n21814 = x11 | n21812 ;
  assign n21815 = ~n21813 & n21814 ;
  assign n21816 = ( n21607 & n21617 ) | ( n21607 & n21618 ) | ( n21617 & n21618 ) ;
  assign n21817 = ( n21805 & ~n21815 ) | ( n21805 & n21816 ) | ( ~n21815 & n21816 ) ;
  assign n21818 = ( n21805 & ~n21816 ) | ( n21805 & n21815 ) | ( ~n21816 & n21815 ) ;
  assign n21819 = ( n21817 & ~n21805 ) | ( n21817 & n21818 ) | ( ~n21805 & n21818 ) ;
  assign n21821 = n8764 &  n20237 ;
  assign n21822 = ( n8105 & ~n20241 ) | ( n8105 & 1'b0 ) | ( ~n20241 & 1'b0 ) ;
  assign n21823 = ~n8429 & n20245 ;
  assign n21824 = n21822 | n21823 ;
  assign n21825 = ( n20237 & ~n21821 ) | ( n20237 & n21824 ) | ( ~n21821 & n21824 ) ;
  assign n21826 = ( n8107 & ~n20253 ) | ( n8107 & n21825 ) | ( ~n20253 & n21825 ) ;
  assign n21827 = n20253 | n21826 ;
  assign n21828 = ( x8 & ~n21825 ) | ( x8 & n21827 ) | ( ~n21825 & n21827 ) ;
  assign n21829 = ( n21825 & ~x8 ) | ( n21825 & n21827 ) | ( ~x8 & n21827 ) ;
  assign n21830 = ( n21828 & ~n21827 ) | ( n21828 & n21829 ) | ( ~n21827 & n21829 ) ;
  assign n21820 = ( n21621 & n21622 ) | ( n21621 & n21632 ) | ( n21622 & n21632 ) ;
  assign n21831 = ( n21819 & ~n21830 ) | ( n21819 & n21820 ) | ( ~n21830 & n21820 ) ;
  assign n21832 = ( n21819 & ~n21820 ) | ( n21819 & n21830 ) | ( ~n21820 & n21830 ) ;
  assign n21833 = ( n21831 & ~n21819 ) | ( n21831 & n21832 ) | ( ~n21819 & n21832 ) ;
  assign n21837 = ~n9997 & n21271 ;
  assign n21834 = n9160 | n20782 ;
  assign n21835 = ~n9558 & n20777 ;
  assign n21836 = ( n21834 & ~n21835 ) | ( n21834 & 1'b0 ) | ( ~n21835 & 1'b0 ) ;
  assign n21838 = ( n9997 & n21837 ) | ( n9997 & n21836 ) | ( n21837 & n21836 ) ;
  assign n21839 = n9155 | n21279 ;
  assign n21840 = n21838 &  n21839 ;
  assign n21841 = x5 &  n21840 ;
  assign n21842 = x5 | n21840 ;
  assign n21843 = ~n21841 & n21842 ;
  assign n21844 = ( n21635 & n21645 ) | ( n21635 & n21646 ) | ( n21645 & n21646 ) ;
  assign n21845 = ( n21833 & ~n21843 ) | ( n21833 & n21844 ) | ( ~n21843 & n21844 ) ;
  assign n21846 = ( n21833 & ~n21844 ) | ( n21833 & n21843 ) | ( ~n21844 & n21843 ) ;
  assign n21847 = ( n21845 & ~n21833 ) | ( n21845 & n21846 ) | ( ~n21833 & n21846 ) ;
  assign n21849 = n3644 | n14816 ;
  assign n21850 = ( n3652 & ~n14803 ) | ( n3652 & 1'b0 ) | ( ~n14803 & 1'b0 ) ;
  assign n21851 = n3657 &  n14807 ;
  assign n21852 = n21850 | n21851 ;
  assign n21853 = n3653 | n14800 ;
  assign n21854 = ( n21852 & ~n3653 ) | ( n21852 & n21853 ) | ( ~n3653 & n21853 ) ;
  assign n21855 = ( n21849 & ~n21854 ) | ( n21849 & 1'b0 ) | ( ~n21854 & 1'b0 ) ;
  assign n21856 = ( x29 & ~n21658 ) | ( x29 & 1'b0 ) | ( ~n21658 & 1'b0 ) ;
  assign n21857 = ( n21653 & ~x29 ) | ( n21653 & n21658 ) | ( ~x29 & n21658 ) ;
  assign n21858 = ( n21654 & n21856 ) | ( n21654 & n21857 ) | ( n21856 & n21857 ) ;
  assign n21859 = ( n21855 & ~n548 ) | ( n21855 & n21858 ) | ( ~n548 & n21858 ) ;
  assign n21860 = ( n548 & ~n21855 ) | ( n548 & n21858 ) | ( ~n21855 & n21858 ) ;
  assign n21861 = ( n21859 & ~n21858 ) | ( n21859 & n21860 ) | ( ~n21858 & n21860 ) ;
  assign n21863 = ( n21671 & n21674 ) | ( n21671 & n21861 ) | ( n21674 & n21861 ) ;
  assign n21862 = ( n21674 & ~n21671 ) | ( n21674 & n21861 ) | ( ~n21671 & n21861 ) ;
  assign n21864 = ( n21671 & ~n21863 ) | ( n21671 & n21862 ) | ( ~n21863 & n21862 ) ;
  assign n21868 = n21864 &  n10499 ;
  assign n21865 = ~n10015 & n21475 ;
  assign n21866 = n10486 | n21675 ;
  assign n21867 = ~n21865 & n21866 ;
  assign n21869 = ( n21868 & ~n10499 ) | ( n21868 & n21867 ) | ( ~n10499 & n21867 ) ;
  assign n21870 = ( n21683 & ~n21675 ) | ( n21683 & n21864 ) | ( ~n21675 & n21864 ) ;
  assign n21871 = ( n21675 & ~n21683 ) | ( n21675 & n21864 ) | ( ~n21683 & n21864 ) ;
  assign n21872 = ( n21870 & ~n21864 ) | ( n21870 & n21871 ) | ( ~n21864 & n21871 ) ;
  assign n21873 = ( n10017 & n21869 ) | ( n10017 & n21872 ) | ( n21869 & n21872 ) ;
  assign n21874 = ~n10017 & n21873 ;
  assign n21876 = ( x2 & n21869 ) | ( x2 & n21874 ) | ( n21869 & n21874 ) ;
  assign n21875 = ( x2 & ~n21874 ) | ( x2 & n21869 ) | ( ~n21874 & n21869 ) ;
  assign n21877 = ( n21874 & ~n21876 ) | ( n21874 & n21875 ) | ( ~n21876 & n21875 ) ;
  assign n21848 = ( n21649 & n21650 ) | ( n21649 & n21689 ) | ( n21650 & n21689 ) ;
  assign n21878 = ( n21847 & ~n21877 ) | ( n21847 & n21848 ) | ( ~n21877 & n21848 ) ;
  assign n21879 = ( n21847 & ~n21848 ) | ( n21847 & n21877 ) | ( ~n21848 & n21877 ) ;
  assign n21880 = ( n21878 & ~n21847 ) | ( n21878 & n21879 ) | ( ~n21847 & n21879 ) ;
  assign n21881 = ( n21693 & ~n21880 ) | ( n21693 & 1'b0 ) | ( ~n21880 & 1'b0 ) ;
  assign n21882 = ~n21693 & n21880 ;
  assign n21883 = n21881 | n21882 ;
  assign n21884 = ( n1437 & ~n2960 ) | ( n1437 & 1'b0 ) | ( ~n2960 & 1'b0 ) ;
  assign n21885 = ( n21884 & ~n1184 ) | ( n21884 & n2484 ) | ( ~n1184 & n2484 ) ;
  assign n21886 = ( n21885 & ~n2484 ) | ( n21885 & 1'b0 ) | ( ~n2484 & 1'b0 ) ;
  assign n21887 = ( n61 & ~n222 ) | ( n61 & n21886 ) | ( ~n222 & n21886 ) ;
  assign n21888 = ~n61 & n21887 ;
  assign n21889 = ( n165 & ~n744 ) | ( n165 & n21888 ) | ( ~n744 & n21888 ) ;
  assign n21890 = ~n165 & n21889 ;
  assign n21891 = ( n561 & ~n404 ) | ( n561 & n21890 ) | ( ~n404 & n21890 ) ;
  assign n21892 = ~n561 & n21891 ;
  assign n21893 = ( n21892 & ~n229 ) | ( n21892 & n266 ) | ( ~n229 & n266 ) ;
  assign n21894 = ( n21893 & ~n266 ) | ( n21893 & 1'b0 ) | ( ~n266 & 1'b0 ) ;
  assign n21895 = n2092 | n2959 ;
  assign n21896 = ( n1209 & ~n2181 ) | ( n1209 & n21895 ) | ( ~n2181 & n21895 ) ;
  assign n21897 = n2181 | n21896 ;
  assign n21898 = ( n998 & ~n629 ) | ( n998 & n21897 ) | ( ~n629 & n21897 ) ;
  assign n21899 = n629 | n21898 ;
  assign n21900 = ( n2610 & ~n21899 ) | ( n2610 & n4322 ) | ( ~n21899 & n4322 ) ;
  assign n21901 = ~n2610 & n21900 ;
  assign n21902 = ( n4911 & ~n2798 ) | ( n4911 & n21901 ) | ( ~n2798 & n21901 ) ;
  assign n21903 = n2798 &  n21902 ;
  assign n21904 = ( n1484 & n21894 ) | ( n1484 & n21903 ) | ( n21894 & n21903 ) ;
  assign n21905 = ~n1484 & n21904 ;
  assign n21906 = ( n477 & ~n912 ) | ( n477 & n21905 ) | ( ~n912 & n21905 ) ;
  assign n21907 = ~n477 & n21906 ;
  assign n21908 = ( n150 & ~n257 ) | ( n150 & n21907 ) | ( ~n257 & n21907 ) ;
  assign n21909 = ~n150 & n21908 ;
  assign n21910 = ( n457 & ~n205 ) | ( n457 & n21909 ) | ( ~n205 & n21909 ) ;
  assign n21911 = ~n457 & n21910 ;
  assign n21912 = ~n432 & n21911 ;
  assign n21913 = ( n21710 & n21711 ) | ( n21710 & n21718 ) | ( n21711 & n21718 ) ;
  assign n21919 = ~n3644 & n15708 ;
  assign n21914 = n3653 | n15700 ;
  assign n21915 = ( n3657 & ~n15320 ) | ( n3657 & 1'b0 ) | ( ~n15320 & 1'b0 ) ;
  assign n21916 = ( n3652 & ~n15325 ) | ( n3652 & 1'b0 ) | ( ~n15325 & 1'b0 ) ;
  assign n21917 = n21915 | n21916 ;
  assign n21918 = ( n21914 & ~n21917 ) | ( n21914 & 1'b0 ) | ( ~n21917 & 1'b0 ) ;
  assign n21920 = ( n3644 & n21919 ) | ( n3644 & n21918 ) | ( n21919 & n21918 ) ;
  assign n21921 = ( n21912 & ~n21913 ) | ( n21912 & n21920 ) | ( ~n21913 & n21920 ) ;
  assign n21922 = ( n21912 & ~n21920 ) | ( n21912 & n21913 ) | ( ~n21920 & n21913 ) ;
  assign n21923 = ( n21921 & ~n21912 ) | ( n21921 & n21922 ) | ( ~n21912 & n21922 ) ;
  assign n21924 = ( n21721 & n21722 ) | ( n21721 & n21732 ) | ( n21722 & n21732 ) ;
  assign n21928 = ~n4430 & n16591 ;
  assign n21925 = n523 | n15897 ;
  assign n21926 = n3939 | n16091 ;
  assign n21927 = n21925 &  n21926 ;
  assign n21929 = ( n4430 & n21928 ) | ( n4430 & n21927 ) | ( n21928 & n21927 ) ;
  assign n21930 = ( n16631 & ~n601 ) | ( n16631 & n21929 ) | ( ~n601 & n21929 ) ;
  assign n21931 = ~n16631 & n21930 ;
  assign n21932 = ( x29 & ~n21929 ) | ( x29 & n21931 ) | ( ~n21929 & n21931 ) ;
  assign n21933 = ( n21929 & ~x29 ) | ( n21929 & n21931 ) | ( ~x29 & n21931 ) ;
  assign n21934 = ( n21932 & ~n21931 ) | ( n21932 & n21933 ) | ( ~n21931 & n21933 ) ;
  assign n21935 = ( n21923 & ~n21924 ) | ( n21923 & n21934 ) | ( ~n21924 & n21934 ) ;
  assign n21936 = ( n21923 & ~n21934 ) | ( n21923 & n21924 ) | ( ~n21934 & n21924 ) ;
  assign n21937 = ( n21935 & ~n21923 ) | ( n21935 & n21936 ) | ( ~n21923 & n21936 ) ;
  assign n21942 = n17107 | n4962 ;
  assign n21939 = n4482 | n16595 ;
  assign n21940 = n4495 | n16589 ;
  assign n21941 = n21939 &  n21940 ;
  assign n21943 = ( n4962 & ~n21942 ) | ( n4962 & n21941 ) | ( ~n21942 & n21941 ) ;
  assign n21944 = ( n4478 & ~n21943 ) | ( n4478 & n17115 ) | ( ~n21943 & n17115 ) ;
  assign n21945 = ( n17115 & ~n21944 ) | ( n17115 & 1'b0 ) | ( ~n21944 & 1'b0 ) ;
  assign n21946 = ( x26 & ~n21943 ) | ( x26 & n21945 ) | ( ~n21943 & n21945 ) ;
  assign n21947 = ( n21943 & ~x26 ) | ( n21943 & n21945 ) | ( ~x26 & n21945 ) ;
  assign n21948 = ( n21946 & ~n21945 ) | ( n21946 & n21947 ) | ( ~n21945 & n21947 ) ;
  assign n21938 = ( n21735 & n21736 ) | ( n21735 & n21746 ) | ( n21736 & n21746 ) ;
  assign n21949 = ( n21937 & ~n21948 ) | ( n21937 & n21938 ) | ( ~n21948 & n21938 ) ;
  assign n21950 = ( n21937 & ~n21938 ) | ( n21937 & n21948 ) | ( ~n21938 & n21948 ) ;
  assign n21951 = ( n21949 & ~n21937 ) | ( n21949 & n21950 ) | ( ~n21937 & n21950 ) ;
  assign n21955 = ~n5135 & n17787 ;
  assign n21952 = n5010 | n17263 ;
  assign n21953 = n5067 | n17405 ;
  assign n21954 = n21952 &  n21953 ;
  assign n21956 = ( n5135 & n21955 ) | ( n5135 & n21954 ) | ( n21955 & n21954 ) ;
  assign n21957 = n5012 | n17826 ;
  assign n21958 = n21956 &  n21957 ;
  assign n21959 = x23 &  n21958 ;
  assign n21960 = x23 | n21958 ;
  assign n21961 = ~n21959 & n21960 ;
  assign n21962 = ( n21749 & n21759 ) | ( n21749 & n21760 ) | ( n21759 & n21760 ) ;
  assign n21963 = ( n21951 & ~n21961 ) | ( n21951 & n21962 ) | ( ~n21961 & n21962 ) ;
  assign n21964 = ( n21951 & ~n21962 ) | ( n21951 & n21961 ) | ( ~n21962 & n21961 ) ;
  assign n21965 = ( n21963 & ~n21951 ) | ( n21963 & n21964 ) | ( ~n21951 & n21964 ) ;
  assign n21970 = ~n5837 & n18456 ;
  assign n21967 = ( n5339 & ~n17791 ) | ( n5339 & 1'b0 ) | ( ~n17791 & 1'b0 ) ;
  assign n21968 = n5761 | n17783 ;
  assign n21969 = ~n21967 & n21968 ;
  assign n21971 = ( n5837 & n21970 ) | ( n5837 & n21969 ) | ( n21970 & n21969 ) ;
  assign n21972 = ( n18464 & ~n5341 ) | ( n18464 & n21971 ) | ( ~n5341 & n21971 ) ;
  assign n21973 = ~n18464 & n21972 ;
  assign n21974 = ( x20 & ~n21971 ) | ( x20 & n21973 ) | ( ~n21971 & n21973 ) ;
  assign n21975 = ( n21971 & ~x20 ) | ( n21971 & n21973 ) | ( ~x20 & n21973 ) ;
  assign n21976 = ( n21974 & ~n21973 ) | ( n21974 & n21975 ) | ( ~n21973 & n21975 ) ;
  assign n21966 = ( n21763 & n21764 ) | ( n21763 & n21774 ) | ( n21764 & n21774 ) ;
  assign n21977 = ( n21965 & ~n21976 ) | ( n21965 & n21966 ) | ( ~n21976 & n21966 ) ;
  assign n21978 = ( n21965 & ~n21966 ) | ( n21965 & n21976 ) | ( ~n21966 & n21976 ) ;
  assign n21979 = ( n21977 & ~n21965 ) | ( n21977 & n21978 ) | ( ~n21965 & n21978 ) ;
  assign n21983 = ~n6395 & n19043 ;
  assign n21980 = n5970 | n18589 ;
  assign n21981 = n6170 | n18712 ;
  assign n21982 = n21980 &  n21981 ;
  assign n21984 = ( n6395 & n21983 ) | ( n6395 & n21982 ) | ( n21983 & n21982 ) ;
  assign n21985 = n5972 | n19083 ;
  assign n21986 = n21984 &  n21985 ;
  assign n21987 = x17 &  n21986 ;
  assign n21988 = x17 | n21986 ;
  assign n21989 = ~n21987 & n21988 ;
  assign n21990 = ( n21777 & n21787 ) | ( n21777 & n21788 ) | ( n21787 & n21788 ) ;
  assign n21991 = ( n21979 & ~n21989 ) | ( n21979 & n21990 ) | ( ~n21989 & n21990 ) ;
  assign n21992 = ( n21979 & ~n21990 ) | ( n21979 & n21989 ) | ( ~n21990 & n21989 ) ;
  assign n21993 = ( n21991 & ~n21979 ) | ( n21991 & n21992 ) | ( ~n21979 & n21992 ) ;
  assign n21995 = ~n6530 & n19047 ;
  assign n21996 = ~n6983 & n19040 ;
  assign n21997 = n21995 | n21996 ;
  assign n21998 = ~n7097 & n19494 ;
  assign n21999 = ( n7097 & ~n21997 ) | ( n7097 & n21998 ) | ( ~n21997 & n21998 ) ;
  assign n22000 = ( n19502 & ~n6532 ) | ( n19502 & n21999 ) | ( ~n6532 & n21999 ) ;
  assign n22001 = ~n19502 & n22000 ;
  assign n22002 = ( x14 & ~n21999 ) | ( x14 & n22001 ) | ( ~n21999 & n22001 ) ;
  assign n22003 = ( n21999 & ~x14 ) | ( n21999 & n22001 ) | ( ~x14 & n22001 ) ;
  assign n22004 = ( n22002 & ~n22001 ) | ( n22002 & n22003 ) | ( ~n22001 & n22003 ) ;
  assign n21994 = ( n21791 & n21792 ) | ( n21791 & n21802 ) | ( n21792 & n21802 ) ;
  assign n22005 = ( n21993 & ~n22004 ) | ( n21993 & n21994 ) | ( ~n22004 & n21994 ) ;
  assign n22006 = ( n21993 & ~n21994 ) | ( n21993 & n22004 ) | ( ~n21994 & n22004 ) ;
  assign n22007 = ( n22005 & ~n21993 ) | ( n22005 & n22006 ) | ( ~n21993 & n22006 ) ;
  assign n22011 = ~n7783 & n20241 ;
  assign n22008 = ( n7253 & ~n19951 ) | ( n7253 & 1'b0 ) | ( ~n19951 & 1'b0 ) ;
  assign n22009 = n7518 | n20027 ;
  assign n22010 = ~n22008 & n22009 ;
  assign n22012 = ( n7783 & n22011 ) | ( n7783 & n22010 ) | ( n22011 & n22010 ) ;
  assign n22013 = n7255 | n20280 ;
  assign n22014 = n22012 &  n22013 ;
  assign n22015 = x11 &  n22014 ;
  assign n22016 = x11 | n22014 ;
  assign n22017 = ~n22015 & n22016 ;
  assign n22018 = ( n21805 & n21815 ) | ( n21805 & n21816 ) | ( n21815 & n21816 ) ;
  assign n22019 = ( n22007 & ~n22017 ) | ( n22007 & n22018 ) | ( ~n22017 & n22018 ) ;
  assign n22020 = ( n22007 & ~n22018 ) | ( n22007 & n22017 ) | ( ~n22018 & n22017 ) ;
  assign n22021 = ( n22019 & ~n22007 ) | ( n22019 & n22020 ) | ( ~n22007 & n22020 ) ;
  assign n22023 = n8105 &  n20245 ;
  assign n22024 = ~n8429 & n20237 ;
  assign n22025 = n22023 | n22024 ;
  assign n22026 = ~n8764 & n20782 ;
  assign n22027 = ( n8764 & ~n22025 ) | ( n8764 & n22026 ) | ( ~n22025 & n22026 ) ;
  assign n22028 = ( n21227 & ~n8107 ) | ( n21227 & n22027 ) | ( ~n8107 & n22027 ) ;
  assign n22029 = ~n21227 & n22028 ;
  assign n22031 = ( x8 & n22027 ) | ( x8 & n22029 ) | ( n22027 & n22029 ) ;
  assign n22030 = ( x8 & ~n22029 ) | ( x8 & n22027 ) | ( ~n22029 & n22027 ) ;
  assign n22032 = ( n22029 & ~n22031 ) | ( n22029 & n22030 ) | ( ~n22031 & n22030 ) ;
  assign n22022 = ( n21819 & n21820 ) | ( n21819 & n21830 ) | ( n21820 & n21830 ) ;
  assign n22033 = ( n22021 & ~n22032 ) | ( n22021 & n22022 ) | ( ~n22032 & n22022 ) ;
  assign n22034 = ( n22021 & ~n22022 ) | ( n22021 & n22032 ) | ( ~n22022 & n22032 ) ;
  assign n22035 = ( n22033 & ~n22021 ) | ( n22033 & n22034 ) | ( ~n22021 & n22034 ) ;
  assign n22039 = n21475 | n9997 ;
  assign n22036 = ~n9160 & n20777 ;
  assign n22037 = n9558 | n21271 ;
  assign n22038 = ~n22036 & n22037 ;
  assign n22040 = ( n9997 & ~n22039 ) | ( n9997 & n22038 ) | ( ~n22039 & n22038 ) ;
  assign n22041 = n9155 | n21484 ;
  assign n22042 = n22040 &  n22041 ;
  assign n22043 = x5 &  n22042 ;
  assign n22044 = x5 | n22042 ;
  assign n22045 = ~n22043 & n22044 ;
  assign n22046 = ( n21833 & n21843 ) | ( n21833 & n21844 ) | ( n21843 & n21844 ) ;
  assign n22047 = ( n22035 & ~n22045 ) | ( n22035 & n22046 ) | ( ~n22045 & n22046 ) ;
  assign n22048 = ( n22035 & ~n22046 ) | ( n22035 & n22045 ) | ( ~n22046 & n22045 ) ;
  assign n22049 = ( n22047 & ~n22035 ) | ( n22047 & n22048 ) | ( ~n22035 & n22048 ) ;
  assign n22064 = n10015 | n21675 ;
  assign n22065 = n10486 | n21864 ;
  assign n22066 = n22064 &  n22065 ;
  assign n22060 = ( n21671 & ~n21674 ) | ( n21671 & n21861 ) | ( ~n21674 & n21861 ) ;
  assign n22051 = ~n3644 & n15692 ;
  assign n22052 = ( n3653 & ~n3657 ) | ( n3653 & 1'b0 ) | ( ~n3657 & 1'b0 ) ;
  assign n22053 = ( n14800 & ~n22052 ) | ( n14800 & 1'b0 ) | ( ~n22052 & 1'b0 ) ;
  assign n22054 = n3652 &  n14807 ;
  assign n22055 = n22053 | n22054 ;
  assign n22056 = n22051 | n22055 ;
  assign n22057 = ( n548 & ~n22056 ) | ( n548 & 1'b0 ) | ( ~n22056 & 1'b0 ) ;
  assign n22058 = ~n548 & n22056 ;
  assign n22059 = n22057 | n22058 ;
  assign n22061 = ( n21859 & ~n22060 ) | ( n21859 & n22059 ) | ( ~n22060 & n22059 ) ;
  assign n22062 = ( n21859 & ~n22059 ) | ( n21859 & n22060 ) | ( ~n22059 & n22060 ) ;
  assign n22063 = ( ~n21859 & n22061 ) | ( ~n21859 & n22062 ) | ( n22061 & n22062 ) ;
  assign n22067 = n10499 &  n22063 ;
  assign n22068 = ( n22066 & ~n10499 ) | ( n22066 & n22067 ) | ( ~n10499 & n22067 ) ;
  assign n22069 = ( n21864 & ~n22063 ) | ( n21864 & n21871 ) | ( ~n22063 & n21871 ) ;
  assign n22070 = ( n21871 & ~n21864 ) | ( n21871 & n22063 ) | ( ~n21864 & n22063 ) ;
  assign n22071 = ( n22069 & ~n21871 ) | ( n22069 & n22070 ) | ( ~n21871 & n22070 ) ;
  assign n22072 = ( n10017 & ~n22071 ) | ( n10017 & n22068 ) | ( ~n22071 & n22068 ) ;
  assign n22073 = ~n10017 & n22072 ;
  assign n22074 = ( x2 & ~n22068 ) | ( x2 & n22073 ) | ( ~n22068 & n22073 ) ;
  assign n22075 = ( n22068 & ~x2 ) | ( n22068 & n22073 ) | ( ~x2 & n22073 ) ;
  assign n22076 = ( n22074 & ~n22073 ) | ( n22074 & n22075 ) | ( ~n22073 & n22075 ) ;
  assign n22050 = ( n21847 & n21848 ) | ( n21847 & n21877 ) | ( n21848 & n21877 ) ;
  assign n22077 = ( n22049 & ~n22076 ) | ( n22049 & n22050 ) | ( ~n22076 & n22050 ) ;
  assign n22078 = ( n22049 & ~n22050 ) | ( n22049 & n22076 ) | ( ~n22050 & n22076 ) ;
  assign n22079 = ( n22077 & ~n22049 ) | ( n22077 & n22078 ) | ( ~n22049 & n22078 ) ;
  assign n22080 = ( n21881 & ~n22079 ) | ( n21881 & 1'b0 ) | ( ~n22079 & 1'b0 ) ;
  assign n22081 = ~n21881 & n22079 ;
  assign n22082 = n22080 | n22081 ;
  assign n22083 = ( n21923 & n21924 ) | ( n21923 & n21934 ) | ( n21924 & n21934 ) ;
  assign n22116 = ~n4430 & n16595 ;
  assign n22113 = n523 | n16091 ;
  assign n22114 = n3939 | n16591 ;
  assign n22115 = n22113 &  n22114 ;
  assign n22117 = ( n4430 & n22116 ) | ( n4430 & n22115 ) | ( n22116 & n22115 ) ;
  assign n22118 = ( n16616 & ~n601 ) | ( n16616 & n22117 ) | ( ~n601 & n22117 ) ;
  assign n22119 = ~n16616 & n22118 ;
  assign n22121 = ( x29 & n22117 ) | ( x29 & n22119 ) | ( n22117 & n22119 ) ;
  assign n22120 = ( x29 & ~n22119 ) | ( x29 & n22117 ) | ( ~n22119 & n22117 ) ;
  assign n22122 = ( n22119 & ~n22121 ) | ( n22119 & n22120 ) | ( ~n22121 & n22120 ) ;
  assign n22084 = ~n1169 & n1249 ;
  assign n22085 = ( n385 & ~n4181 ) | ( n385 & n22084 ) | ( ~n4181 & n22084 ) ;
  assign n22086 = ~n385 & n22085 ;
  assign n22087 = ( n4083 & n14151 ) | ( n4083 & n22086 ) | ( n14151 & n22086 ) ;
  assign n22088 = ~n4083 & n22087 ;
  assign n22089 = ( n163 & n5664 ) | ( n163 & n22088 ) | ( n5664 & n22088 ) ;
  assign n22090 = ~n163 & n22089 ;
  assign n22091 = ( n61 & ~n814 ) | ( n61 & n22090 ) | ( ~n814 & n22090 ) ;
  assign n22092 = ~n61 & n22091 ;
  assign n22093 = ( n475 & ~n72 ) | ( n475 & n22092 ) | ( ~n72 & n22092 ) ;
  assign n22094 = ~n475 & n22093 ;
  assign n22095 = ( n571 & ~n237 ) | ( n571 & n22094 ) | ( ~n237 & n22094 ) ;
  assign n22096 = ~n571 & n22095 ;
  assign n22097 = ( n276 & ~n43 ) | ( n276 & n22096 ) | ( ~n43 & n22096 ) ;
  assign n22098 = ~n276 & n22097 ;
  assign n22099 = ( n617 & ~n86 ) | ( n617 & n22098 ) | ( ~n86 & n22098 ) ;
  assign n22100 = ~n617 & n22099 ;
  assign n22101 = ~n225 & n22100 ;
  assign n22102 = ( n21912 & n21913 ) | ( n21912 & n21920 ) | ( n21913 & n21920 ) ;
  assign n22108 = ~n3644 & n15900 ;
  assign n22103 = n3653 | n15897 ;
  assign n22104 = ( n3657 & ~n15700 ) | ( n3657 & 1'b0 ) | ( ~n15700 & 1'b0 ) ;
  assign n22105 = ( n3652 & ~n15320 ) | ( n3652 & 1'b0 ) | ( ~n15320 & 1'b0 ) ;
  assign n22106 = n22104 | n22105 ;
  assign n22107 = ( n22103 & ~n22106 ) | ( n22103 & 1'b0 ) | ( ~n22106 & 1'b0 ) ;
  assign n22109 = ( n3644 & n22108 ) | ( n3644 & n22107 ) | ( n22108 & n22107 ) ;
  assign n22110 = ( n22101 & ~n22102 ) | ( n22101 & n22109 ) | ( ~n22102 & n22109 ) ;
  assign n22111 = ( n22101 & ~n22109 ) | ( n22101 & n22102 ) | ( ~n22109 & n22102 ) ;
  assign n22112 = ( n22110 & ~n22101 ) | ( n22110 & n22111 ) | ( ~n22101 & n22111 ) ;
  assign n22123 = ( n22083 & ~n22122 ) | ( n22083 & n22112 ) | ( ~n22122 & n22112 ) ;
  assign n22124 = ( n22112 & ~n22083 ) | ( n22112 & n22122 ) | ( ~n22083 & n22122 ) ;
  assign n22125 = ( n22123 & ~n22112 ) | ( n22123 & n22124 ) | ( ~n22112 & n22124 ) ;
  assign n22126 = ( n21937 & n21938 ) | ( n21937 & n21948 ) | ( n21938 & n21948 ) ;
  assign n22130 = ~n4962 & n17263 ;
  assign n22127 = n4482 | n16589 ;
  assign n22128 = ~n4495 & n17107 ;
  assign n22129 = ( n22127 & ~n22128 ) | ( n22127 & 1'b0 ) | ( ~n22128 & 1'b0 ) ;
  assign n22131 = ( n4962 & n22130 ) | ( n4962 & n22129 ) | ( n22130 & n22129 ) ;
  assign n22132 = ( n4478 & ~n22131 ) | ( n4478 & n17271 ) | ( ~n22131 & n17271 ) ;
  assign n22133 = ( n17271 & ~n22132 ) | ( n17271 & 1'b0 ) | ( ~n22132 & 1'b0 ) ;
  assign n22135 = ( x26 & n22131 ) | ( x26 & n22133 ) | ( n22131 & n22133 ) ;
  assign n22134 = ( x26 & ~n22133 ) | ( x26 & n22131 ) | ( ~n22133 & n22131 ) ;
  assign n22136 = ( n22133 & ~n22135 ) | ( n22133 & n22134 ) | ( ~n22135 & n22134 ) ;
  assign n22137 = ( n22125 & ~n22126 ) | ( n22125 & n22136 ) | ( ~n22126 & n22136 ) ;
  assign n22138 = ( n22126 & ~n22125 ) | ( n22126 & n22136 ) | ( ~n22125 & n22136 ) ;
  assign n22139 = ( n22137 & ~n22136 ) | ( n22137 & n22138 ) | ( ~n22136 & n22138 ) ;
  assign n22143 = ~n5135 & n17791 ;
  assign n22140 = n5010 | n17405 ;
  assign n22141 = n5067 | n17787 ;
  assign n22142 = n22140 &  n22141 ;
  assign n22144 = ( n5135 & n22143 ) | ( n5135 & n22142 ) | ( n22143 & n22142 ) ;
  assign n22145 = n5012 | n17811 ;
  assign n22146 = n22144 &  n22145 ;
  assign n22147 = x23 &  n22146 ;
  assign n22148 = x23 | n22146 ;
  assign n22149 = ~n22147 & n22148 ;
  assign n22150 = ( n21951 & n21961 ) | ( n21951 & n21962 ) | ( n21961 & n21962 ) ;
  assign n22151 = ( n22139 & ~n22149 ) | ( n22139 & n22150 ) | ( ~n22149 & n22150 ) ;
  assign n22152 = ( n22139 & ~n22150 ) | ( n22139 & n22149 ) | ( ~n22150 & n22149 ) ;
  assign n22153 = ( n22151 & ~n22139 ) | ( n22151 & n22152 ) | ( ~n22139 & n22152 ) ;
  assign n22158 = ~n5837 & n18589 ;
  assign n22155 = ( n5339 & ~n17783 ) | ( n5339 & 1'b0 ) | ( ~n17783 & 1'b0 ) ;
  assign n22156 = n5761 | n18456 ;
  assign n22157 = ~n22155 & n22156 ;
  assign n22159 = ( n5837 & n22158 ) | ( n5837 & n22157 ) | ( n22158 & n22157 ) ;
  assign n22160 = ( n18597 & ~n5341 ) | ( n18597 & n22159 ) | ( ~n5341 & n22159 ) ;
  assign n22161 = ~n18597 & n22160 ;
  assign n22163 = ( x20 & n22159 ) | ( x20 & n22161 ) | ( n22159 & n22161 ) ;
  assign n22162 = ( x20 & ~n22161 ) | ( x20 & n22159 ) | ( ~n22161 & n22159 ) ;
  assign n22164 = ( n22161 & ~n22163 ) | ( n22161 & n22162 ) | ( ~n22163 & n22162 ) ;
  assign n22154 = ( n21965 & n21966 ) | ( n21965 & n21976 ) | ( n21966 & n21976 ) ;
  assign n22165 = ( n22153 & ~n22164 ) | ( n22153 & n22154 ) | ( ~n22164 & n22154 ) ;
  assign n22166 = ( n22153 & ~n22154 ) | ( n22153 & n22164 ) | ( ~n22154 & n22164 ) ;
  assign n22167 = ( n22165 & ~n22153 ) | ( n22165 & n22166 ) | ( ~n22153 & n22166 ) ;
  assign n22171 = n19047 | n6395 ;
  assign n22168 = n5970 | n18712 ;
  assign n22169 = n6170 | n19043 ;
  assign n22170 = n22168 &  n22169 ;
  assign n22172 = ( n6395 & ~n22171 ) | ( n6395 & n22170 ) | ( ~n22171 & n22170 ) ;
  assign n22173 = ~n5972 & n19068 ;
  assign n22174 = ( n22172 & ~n22173 ) | ( n22172 & 1'b0 ) | ( ~n22173 & 1'b0 ) ;
  assign n22175 = x17 &  n22174 ;
  assign n22176 = x17 | n22174 ;
  assign n22177 = ~n22175 & n22176 ;
  assign n22178 = ( n21979 & n21989 ) | ( n21979 & n21990 ) | ( n21989 & n21990 ) ;
  assign n22179 = ( n22167 & ~n22177 ) | ( n22167 & n22178 ) | ( ~n22177 & n22178 ) ;
  assign n22180 = ( n22167 & ~n22178 ) | ( n22167 & n22177 ) | ( ~n22178 & n22177 ) ;
  assign n22181 = ( n22179 & ~n22167 ) | ( n22179 & n22180 ) | ( ~n22167 & n22180 ) ;
  assign n22186 = ~n7097 & n19951 ;
  assign n22183 = ~n6530 & n19040 ;
  assign n22184 = n6983 | n19494 ;
  assign n22185 = ~n22183 & n22184 ;
  assign n22187 = ( n7097 & n22186 ) | ( n7097 & n22185 ) | ( n22186 & n22185 ) ;
  assign n22188 = ( n6532 & ~n22187 ) | ( n6532 & n19959 ) | ( ~n22187 & n19959 ) ;
  assign n22189 = ( n19959 & ~n22188 ) | ( n19959 & 1'b0 ) | ( ~n22188 & 1'b0 ) ;
  assign n22191 = ( x14 & n22187 ) | ( x14 & n22189 ) | ( n22187 & n22189 ) ;
  assign n22190 = ( x14 & ~n22189 ) | ( x14 & n22187 ) | ( ~n22189 & n22187 ) ;
  assign n22192 = ( n22189 & ~n22191 ) | ( n22189 & n22190 ) | ( ~n22191 & n22190 ) ;
  assign n22182 = ( n21993 & n21994 ) | ( n21993 & n22004 ) | ( n21994 & n22004 ) ;
  assign n22193 = ( n22181 & ~n22192 ) | ( n22181 & n22182 ) | ( ~n22192 & n22182 ) ;
  assign n22194 = ( n22181 & ~n22182 ) | ( n22181 & n22192 ) | ( ~n22182 & n22192 ) ;
  assign n22195 = ( n22193 & ~n22181 ) | ( n22193 & n22194 ) | ( ~n22181 & n22194 ) ;
  assign n22199 = n20245 | n7783 ;
  assign n22196 = ( n7253 & ~n20027 ) | ( n7253 & 1'b0 ) | ( ~n20027 & 1'b0 ) ;
  assign n22197 = n7518 | n20241 ;
  assign n22198 = ~n22196 & n22197 ;
  assign n22200 = ( n7783 & ~n22199 ) | ( n7783 & n22198 ) | ( ~n22199 & n22198 ) ;
  assign n22201 = ~n7255 & n20265 ;
  assign n22202 = ( n22200 & ~n22201 ) | ( n22200 & 1'b0 ) | ( ~n22201 & 1'b0 ) ;
  assign n22203 = x11 &  n22202 ;
  assign n22204 = x11 | n22202 ;
  assign n22205 = ~n22203 & n22204 ;
  assign n22206 = ( n22007 & n22017 ) | ( n22007 & n22018 ) | ( n22017 & n22018 ) ;
  assign n22207 = ( n22195 & ~n22205 ) | ( n22195 & n22206 ) | ( ~n22205 & n22206 ) ;
  assign n22208 = ( n22195 & ~n22206 ) | ( n22195 & n22205 ) | ( ~n22206 & n22205 ) ;
  assign n22209 = ( n22207 & ~n22195 ) | ( n22207 & n22208 ) | ( ~n22195 & n22208 ) ;
  assign n22214 = n8764 | n20777 ;
  assign n22211 = n8105 &  n20237 ;
  assign n22212 = n8429 | n20782 ;
  assign n22213 = ~n22211 & n22212 ;
  assign n22215 = ( n8764 & ~n22214 ) | ( n8764 & n22213 ) | ( ~n22214 & n22213 ) ;
  assign n22216 = ( n20790 & ~n8107 ) | ( n20790 & n22215 ) | ( ~n8107 & n22215 ) ;
  assign n22217 = ~n20790 & n22216 ;
  assign n22219 = ( x8 & n22215 ) | ( x8 & n22217 ) | ( n22215 & n22217 ) ;
  assign n22218 = ( x8 & ~n22217 ) | ( x8 & n22215 ) | ( ~n22217 & n22215 ) ;
  assign n22220 = ( n22217 & ~n22219 ) | ( n22217 & n22218 ) | ( ~n22219 & n22218 ) ;
  assign n22210 = ( n22021 & n22022 ) | ( n22021 & n22032 ) | ( n22022 & n22032 ) ;
  assign n22221 = ( n22209 & ~n22220 ) | ( n22209 & n22210 ) | ( ~n22220 & n22210 ) ;
  assign n22222 = ( n22209 & ~n22210 ) | ( n22209 & n22220 ) | ( ~n22210 & n22220 ) ;
  assign n22223 = ( n22221 & ~n22209 ) | ( n22221 & n22222 ) | ( ~n22209 & n22222 ) ;
  assign n22227 = ~n9997 & n21675 ;
  assign n22224 = n9160 | n21271 ;
  assign n22225 = ~n9558 & n21475 ;
  assign n22226 = ( n22224 & ~n22225 ) | ( n22224 & 1'b0 ) | ( ~n22225 & 1'b0 ) ;
  assign n22228 = ( n9997 & n22227 ) | ( n9997 & n22226 ) | ( n22227 & n22226 ) ;
  assign n22229 = n9155 | n21684 ;
  assign n22230 = n22228 &  n22229 ;
  assign n22231 = x5 &  n22230 ;
  assign n22232 = x5 | n22230 ;
  assign n22233 = ~n22231 & n22232 ;
  assign n22234 = ( n22035 & n22045 ) | ( n22035 & n22046 ) | ( n22045 & n22046 ) ;
  assign n22235 = ( n22223 & ~n22233 ) | ( n22223 & n22234 ) | ( ~n22233 & n22234 ) ;
  assign n22236 = ( n22223 & ~n22234 ) | ( n22223 & n22233 ) | ( ~n22234 & n22233 ) ;
  assign n22237 = ( n22235 & ~n22223 ) | ( n22235 & n22236 ) | ( ~n22223 & n22236 ) ;
  assign n22245 = n10015 | n21864 ;
  assign n22246 = n10486 | n22063 ;
  assign n22247 = n22245 &  n22246 ;
  assign n22241 = ( n22059 & ~n21859 ) | ( n22059 & n22060 ) | ( ~n21859 & n22060 ) ;
  assign n22239 = x31 | n41 ;
  assign n22240 = n14800 &  n22239 ;
  assign n22242 = ( n22057 & ~n22241 ) | ( n22057 & n22240 ) | ( ~n22241 & n22240 ) ;
  assign n22243 = ( n22057 & ~n22240 ) | ( n22057 & n22241 ) | ( ~n22240 & n22241 ) ;
  assign n22244 = ( n22242 & ~n22057 ) | ( n22242 & n22243 ) | ( ~n22057 & n22243 ) ;
  assign n22248 = ( n10499 & ~n22244 ) | ( n10499 & 1'b0 ) | ( ~n22244 & 1'b0 ) ;
  assign n22249 = ( n22247 & ~n10499 ) | ( n22247 & n22248 ) | ( ~n10499 & n22248 ) ;
  assign n22250 = ( n21864 & n21871 ) | ( n21864 & n22063 ) | ( n21871 & n22063 ) ;
  assign n22252 = ( n22063 & n22244 ) | ( n22063 & n22250 ) | ( n22244 & n22250 ) ;
  assign n22251 = ( n22063 & ~n22244 ) | ( n22063 & n22250 ) | ( ~n22244 & n22250 ) ;
  assign n22253 = ( n22244 & ~n22252 ) | ( n22244 & n22251 ) | ( ~n22252 & n22251 ) ;
  assign n22254 = ( n10017 & n22249 ) | ( n10017 & n22253 ) | ( n22249 & n22253 ) ;
  assign n22255 = ~n10017 & n22254 ;
  assign n22257 = ( x2 & n22249 ) | ( x2 & n22255 ) | ( n22249 & n22255 ) ;
  assign n22256 = ( x2 & ~n22255 ) | ( x2 & n22249 ) | ( ~n22255 & n22249 ) ;
  assign n22258 = ( n22255 & ~n22257 ) | ( n22255 & n22256 ) | ( ~n22257 & n22256 ) ;
  assign n22238 = ( n22049 & n22050 ) | ( n22049 & n22076 ) | ( n22050 & n22076 ) ;
  assign n22259 = ( n22237 & ~n22258 ) | ( n22237 & n22238 ) | ( ~n22258 & n22238 ) ;
  assign n22260 = ( n22237 & ~n22238 ) | ( n22237 & n22258 ) | ( ~n22238 & n22258 ) ;
  assign n22261 = ( n22259 & ~n22237 ) | ( n22259 & n22260 ) | ( ~n22237 & n22260 ) ;
  assign n22262 = ( n22080 & ~n22261 ) | ( n22080 & 1'b0 ) | ( ~n22261 & 1'b0 ) ;
  assign n22263 = ~n22080 & n22261 ;
  assign n22264 = n22262 | n22263 ;
  assign n22265 = ( n22223 & n22233 ) | ( n22223 & n22234 ) | ( n22233 & n22234 ) ;
  assign n22266 = ( n22083 & n22112 ) | ( n22083 & n22122 ) | ( n22112 & n22122 ) ;
  assign n22274 = n1513 | n21697 ;
  assign n22275 = ( n998 & ~n462 ) | ( n998 & n22274 ) | ( ~n462 & n22274 ) ;
  assign n22276 = n462 | n22275 ;
  assign n22267 = ~n2462 & n2594 ;
  assign n22268 = ( n493 & ~n453 ) | ( n493 & n22267 ) | ( ~n453 & n22267 ) ;
  assign n22269 = ~n493 & n22268 ;
  assign n22270 = ( n343 & ~n22269 ) | ( n343 & n529 ) | ( ~n22269 & n529 ) ;
  assign n22271 = ( n343 & ~n22270 ) | ( n343 & 1'b0 ) | ( ~n22270 & 1'b0 ) ;
  assign n22272 = ( n617 & ~n252 ) | ( n617 & n22271 ) | ( ~n252 & n22271 ) ;
  assign n22273 = ~n617 & n22272 ;
  assign n22277 = ( n17191 & ~n22276 ) | ( n17191 & n22273 ) | ( ~n22276 & n22273 ) ;
  assign n22278 = ~n17191 & n22277 ;
  assign n22279 = ( n5424 & ~n15923 ) | ( n5424 & n22278 ) | ( ~n15923 & n22278 ) ;
  assign n22280 = ~n5424 & n22279 ;
  assign n22281 = ( n1625 & ~n912 ) | ( n1625 & n22280 ) | ( ~n912 & n22280 ) ;
  assign n22282 = ~n1625 & n22281 ;
  assign n22283 = ( n1490 & n3212 ) | ( n1490 & n22282 ) | ( n3212 & n22282 ) ;
  assign n22284 = ~n1490 & n22283 ;
  assign n22285 = ( n62 & ~n490 ) | ( n62 & n22284 ) | ( ~n490 & n22284 ) ;
  assign n22286 = ~n62 & n22285 ;
  assign n22287 = ( n162 & n197 ) | ( n162 & n22286 ) | ( n197 & n22286 ) ;
  assign n22288 = ~n162 & n22287 ;
  assign n22289 = ( n340 & ~n137 ) | ( n340 & n22288 ) | ( ~n137 & n22288 ) ;
  assign n22290 = ~n340 & n22289 ;
  assign n22291 = ( n229 & ~n22290 ) | ( n229 & n354 ) | ( ~n22290 & n354 ) ;
  assign n22292 = ( n354 & ~n22291 ) | ( n354 & 1'b0 ) | ( ~n22291 & 1'b0 ) ;
  assign n22293 = ~n39 & n22292 ;
  assign n22299 = ~n3644 & n16094 ;
  assign n22294 = n3653 | n16091 ;
  assign n22295 = ( n3657 & ~n15897 ) | ( n3657 & 1'b0 ) | ( ~n15897 & 1'b0 ) ;
  assign n22296 = ( n3652 & ~n15700 ) | ( n3652 & 1'b0 ) | ( ~n15700 & 1'b0 ) ;
  assign n22297 = n22295 | n22296 ;
  assign n22298 = ( n22294 & ~n22297 ) | ( n22294 & 1'b0 ) | ( ~n22297 & 1'b0 ) ;
  assign n22300 = ( n3644 & n22299 ) | ( n3644 & n22298 ) | ( n22299 & n22298 ) ;
  assign n22301 = n22293 | n22300 ;
  assign n22302 = ( n22293 & ~n22300 ) | ( n22293 & 1'b0 ) | ( ~n22300 & 1'b0 ) ;
  assign n22303 = ( n22301 & ~n22293 ) | ( n22301 & n22302 ) | ( ~n22293 & n22302 ) ;
  assign n22308 = ~n4430 & n16589 ;
  assign n22305 = n523 | n16591 ;
  assign n22306 = n3939 | n16595 ;
  assign n22307 = n22305 &  n22306 ;
  assign n22309 = ( n4430 & n22308 ) | ( n4430 & n22307 ) | ( n22308 & n22307 ) ;
  assign n22310 = ( n16604 & ~n601 ) | ( n16604 & n22309 ) | ( ~n601 & n22309 ) ;
  assign n22311 = ~n16604 & n22310 ;
  assign n22313 = ( x29 & n22309 ) | ( x29 & n22311 ) | ( n22309 & n22311 ) ;
  assign n22312 = ( x29 & ~n22311 ) | ( x29 & n22309 ) | ( ~n22311 & n22309 ) ;
  assign n22314 = ( n22311 & ~n22313 ) | ( n22311 & n22312 ) | ( ~n22313 & n22312 ) ;
  assign n22304 = ( n22101 & n22102 ) | ( n22101 & n22109 ) | ( n22102 & n22109 ) ;
  assign n22315 = ( n22303 & ~n22314 ) | ( n22303 & n22304 ) | ( ~n22314 & n22304 ) ;
  assign n22316 = ( n22303 & ~n22304 ) | ( n22303 & n22314 ) | ( ~n22304 & n22314 ) ;
  assign n22317 = ( n22315 & ~n22303 ) | ( n22315 & n22316 ) | ( ~n22303 & n22316 ) ;
  assign n22318 = ~n22266 & n22317 ;
  assign n22319 = ( n22266 & ~n22317 ) | ( n22266 & 1'b0 ) | ( ~n22317 & 1'b0 ) ;
  assign n22320 = n22318 | n22319 ;
  assign n22325 = ~n4962 & n17405 ;
  assign n22322 = ~n4482 & n17107 ;
  assign n22323 = n4495 | n17263 ;
  assign n22324 = ~n22322 & n22323 ;
  assign n22326 = ( n4962 & n22325 ) | ( n4962 & n22324 ) | ( n22325 & n22324 ) ;
  assign n22327 = ( n17413 & ~n4478 ) | ( n17413 & n22326 ) | ( ~n4478 & n22326 ) ;
  assign n22328 = ~n17413 & n22327 ;
  assign n22330 = ( x26 & n22326 ) | ( x26 & n22328 ) | ( n22326 & n22328 ) ;
  assign n22329 = ( x26 & ~n22328 ) | ( x26 & n22326 ) | ( ~n22328 & n22326 ) ;
  assign n22331 = ( n22328 & ~n22330 ) | ( n22328 & n22329 ) | ( ~n22330 & n22329 ) ;
  assign n22321 = ( n22125 & n22126 ) | ( n22125 & n22136 ) | ( n22126 & n22136 ) ;
  assign n22332 = ( n22320 & ~n22331 ) | ( n22320 & n22321 ) | ( ~n22331 & n22321 ) ;
  assign n22333 = ( n22320 & ~n22321 ) | ( n22320 & n22331 ) | ( ~n22321 & n22331 ) ;
  assign n22334 = ( n22332 & ~n22320 ) | ( n22332 & n22333 ) | ( ~n22320 & n22333 ) ;
  assign n22345 = ( n22139 & n22149 ) | ( n22139 & n22150 ) | ( n22149 & n22150 ) ;
  assign n22335 = ( n5135 & ~n17783 ) | ( n5135 & 1'b0 ) | ( ~n17783 & 1'b0 ) ;
  assign n22336 = n5010 | n17787 ;
  assign n22337 = n5067 | n17791 ;
  assign n22338 = n22336 &  n22337 ;
  assign n22339 = ( n17783 & n22335 ) | ( n17783 & n22338 ) | ( n22335 & n22338 ) ;
  assign n22340 = n5012 | n17799 ;
  assign n22341 = n22339 &  n22340 ;
  assign n22342 = x23 &  n22341 ;
  assign n22343 = x23 | n22341 ;
  assign n22344 = ~n22342 & n22343 ;
  assign n22346 = ( n22334 & ~n22345 ) | ( n22334 & n22344 ) | ( ~n22345 & n22344 ) ;
  assign n22347 = ( n22334 & ~n22344 ) | ( n22334 & n22345 ) | ( ~n22344 & n22345 ) ;
  assign n22348 = ( n22346 & ~n22334 ) | ( n22346 & n22347 ) | ( ~n22334 & n22347 ) ;
  assign n22353 = ~n5837 & n18712 ;
  assign n22350 = ( n5339 & ~n18456 ) | ( n5339 & 1'b0 ) | ( ~n18456 & 1'b0 ) ;
  assign n22351 = n5761 | n18589 ;
  assign n22352 = ~n22350 & n22351 ;
  assign n22354 = ( n5837 & n22353 ) | ( n5837 & n22352 ) | ( n22353 & n22352 ) ;
  assign n22355 = ( n18720 & ~n5341 ) | ( n18720 & n22354 ) | ( ~n5341 & n22354 ) ;
  assign n22356 = ~n18720 & n22355 ;
  assign n22358 = ( x20 & n22354 ) | ( x20 & n22356 ) | ( n22354 & n22356 ) ;
  assign n22357 = ( x20 & ~n22356 ) | ( x20 & n22354 ) | ( ~n22356 & n22354 ) ;
  assign n22359 = ( n22356 & ~n22358 ) | ( n22356 & n22357 ) | ( ~n22358 & n22357 ) ;
  assign n22349 = ( n22153 & n22154 ) | ( n22153 & n22164 ) | ( n22154 & n22164 ) ;
  assign n22360 = ( n22348 & ~n22359 ) | ( n22348 & n22349 ) | ( ~n22359 & n22349 ) ;
  assign n22361 = ( n22348 & ~n22349 ) | ( n22348 & n22359 ) | ( ~n22349 & n22359 ) ;
  assign n22362 = ( n22360 & ~n22348 ) | ( n22360 & n22361 ) | ( ~n22348 & n22361 ) ;
  assign n22373 = ( n22167 & n22177 ) | ( n22167 & n22178 ) | ( n22177 & n22178 ) ;
  assign n22366 = n19040 | n6395 ;
  assign n22363 = n5970 | n19043 ;
  assign n22364 = ~n6170 & n19047 ;
  assign n22365 = ( n22363 & ~n22364 ) | ( n22363 & 1'b0 ) | ( ~n22364 & 1'b0 ) ;
  assign n22367 = ( n6395 & ~n22366 ) | ( n6395 & n22365 ) | ( ~n22366 & n22365 ) ;
  assign n22368 = n5972 | n19056 ;
  assign n22369 = n22367 &  n22368 ;
  assign n22370 = x17 &  n22369 ;
  assign n22371 = x17 | n22369 ;
  assign n22372 = ~n22370 & n22371 ;
  assign n22374 = ( n22362 & ~n22373 ) | ( n22362 & n22372 ) | ( ~n22373 & n22372 ) ;
  assign n22375 = ( n22362 & ~n22372 ) | ( n22362 & n22373 ) | ( ~n22372 & n22373 ) ;
  assign n22376 = ( n22374 & ~n22362 ) | ( n22374 & n22375 ) | ( ~n22362 & n22375 ) ;
  assign n22381 = ~n7097 & n20027 ;
  assign n22378 = n6530 | n19494 ;
  assign n22379 = n6983 | n19951 ;
  assign n22380 = n22378 &  n22379 ;
  assign n22382 = ( n7097 & n22381 ) | ( n7097 & n22380 ) | ( n22381 & n22380 ) ;
  assign n22383 = ( n20035 & ~n6532 ) | ( n20035 & n22382 ) | ( ~n6532 & n22382 ) ;
  assign n22384 = ~n20035 & n22383 ;
  assign n22386 = ( x14 & n22382 ) | ( x14 & n22384 ) | ( n22382 & n22384 ) ;
  assign n22385 = ( x14 & ~n22384 ) | ( x14 & n22382 ) | ( ~n22384 & n22382 ) ;
  assign n22387 = ( n22384 & ~n22386 ) | ( n22384 & n22385 ) | ( ~n22386 & n22385 ) ;
  assign n22377 = ( n22181 & n22182 ) | ( n22181 & n22192 ) | ( n22182 & n22192 ) ;
  assign n22388 = ( n22376 & ~n22387 ) | ( n22376 & n22377 ) | ( ~n22387 & n22377 ) ;
  assign n22389 = ( n22376 & ~n22377 ) | ( n22376 & n22387 ) | ( ~n22377 & n22387 ) ;
  assign n22390 = ( n22388 & ~n22376 ) | ( n22388 & n22389 ) | ( ~n22376 & n22389 ) ;
  assign n22401 = ( n22195 & n22205 ) | ( n22195 & n22206 ) | ( n22205 & n22206 ) ;
  assign n22391 = n7783 &  n20237 ;
  assign n22392 = ( n7253 & ~n20241 ) | ( n7253 & 1'b0 ) | ( ~n20241 & 1'b0 ) ;
  assign n22393 = ~n7518 & n20245 ;
  assign n22394 = n22392 | n22393 ;
  assign n22395 = ( n20237 & ~n22391 ) | ( n20237 & n22394 ) | ( ~n22391 & n22394 ) ;
  assign n22396 = n7255 | n20253 ;
  assign n22397 = ~n22395 & n22396 ;
  assign n22398 = x11 &  n22397 ;
  assign n22399 = x11 | n22397 ;
  assign n22400 = ~n22398 & n22399 ;
  assign n22402 = ( n22390 & ~n22401 ) | ( n22390 & n22400 ) | ( ~n22401 & n22400 ) ;
  assign n22403 = ( n22390 & ~n22400 ) | ( n22390 & n22401 ) | ( ~n22400 & n22401 ) ;
  assign n22404 = ( n22402 & ~n22390 ) | ( n22402 & n22403 ) | ( ~n22390 & n22403 ) ;
  assign n22406 = ( n8105 & ~n20782 ) | ( n8105 & 1'b0 ) | ( ~n20782 & 1'b0 ) ;
  assign n22407 = ~n8429 & n20777 ;
  assign n22408 = n22406 | n22407 ;
  assign n22409 = ~n8764 & n21271 ;
  assign n22410 = ( n8764 & ~n22408 ) | ( n8764 & n22409 ) | ( ~n22408 & n22409 ) ;
  assign n22411 = ( n21279 & ~n8107 ) | ( n21279 & n22410 ) | ( ~n8107 & n22410 ) ;
  assign n22412 = ~n21279 & n22411 ;
  assign n22414 = ( x8 & n22410 ) | ( x8 & n22412 ) | ( n22410 & n22412 ) ;
  assign n22413 = ( x8 & ~n22412 ) | ( x8 & n22410 ) | ( ~n22412 & n22410 ) ;
  assign n22415 = ( n22412 & ~n22414 ) | ( n22412 & n22413 ) | ( ~n22414 & n22413 ) ;
  assign n22405 = ( n22209 & n22210 ) | ( n22209 & n22220 ) | ( n22210 & n22220 ) ;
  assign n22416 = ( n22404 & ~n22415 ) | ( n22404 & n22405 ) | ( ~n22415 & n22405 ) ;
  assign n22417 = ( n22404 & ~n22405 ) | ( n22404 & n22415 ) | ( ~n22405 & n22415 ) ;
  assign n22418 = ( n22416 & ~n22404 ) | ( n22416 & n22417 ) | ( ~n22404 & n22417 ) ;
  assign n22432 = ~n10017 & n22251 ;
  assign n22429 = ~n15688 & n22244 ;
  assign n22430 = n10015 | n22063 ;
  assign n22431 = ~n22429 & n22430 ;
  assign n22433 = ( n10017 & n22432 ) | ( n10017 & n22431 ) | ( n22432 & n22431 ) ;
  assign n22434 = x2 | n22433 ;
  assign n22435 = ( x2 & ~n22433 ) | ( x2 & 1'b0 ) | ( ~n22433 & 1'b0 ) ;
  assign n22436 = ( n22434 & ~x2 ) | ( n22434 & n22435 ) | ( ~x2 & n22435 ) ;
  assign n22419 = ( n9997 & ~n21864 ) | ( n9997 & 1'b0 ) | ( ~n21864 & 1'b0 ) ;
  assign n22420 = ~n9160 & n21475 ;
  assign n22421 = n9558 | n21675 ;
  assign n22422 = ~n22420 & n22421 ;
  assign n22423 = ( n21864 & n22419 ) | ( n21864 & n22422 ) | ( n22419 & n22422 ) ;
  assign n22424 = ~n9155 & n21872 ;
  assign n22425 = ( n22423 & ~n22424 ) | ( n22423 & 1'b0 ) | ( ~n22424 & 1'b0 ) ;
  assign n22426 = x5 &  n22425 ;
  assign n22427 = x5 | n22425 ;
  assign n22428 = ~n22426 & n22427 ;
  assign n22437 = ( n22418 & ~n22436 ) | ( n22418 & n22428 ) | ( ~n22436 & n22428 ) ;
  assign n22438 = ( n22418 & ~n22428 ) | ( n22418 & n22436 ) | ( ~n22428 & n22436 ) ;
  assign n22439 = ( n22437 & ~n22418 ) | ( n22437 & n22438 ) | ( ~n22418 & n22438 ) ;
  assign n22440 = ( n22237 & n22238 ) | ( n22237 & n22258 ) | ( n22238 & n22258 ) ;
  assign n22441 = ( n22265 & ~n22439 ) | ( n22265 & n22440 ) | ( ~n22439 & n22440 ) ;
  assign n22442 = ( n22265 & ~n22440 ) | ( n22265 & n22439 ) | ( ~n22440 & n22439 ) ;
  assign n22443 = ( n22441 & ~n22265 ) | ( n22441 & n22442 ) | ( ~n22265 & n22442 ) ;
  assign n22444 = ( n22262 & ~n22443 ) | ( n22262 & 1'b0 ) | ( ~n22443 & 1'b0 ) ;
  assign n22445 = ~n22262 & n22443 ;
  assign n22446 = n22444 | n22445 ;
  assign n22450 = ~n9997 & n22063 ;
  assign n22447 = n9160 | n21675 ;
  assign n22448 = n9558 | n21864 ;
  assign n22449 = n22447 &  n22448 ;
  assign n22451 = ( n9997 & n22450 ) | ( n9997 & n22449 ) | ( n22450 & n22449 ) ;
  assign n22452 = n9155 | n22071 ;
  assign n22453 = n22451 &  n22452 ;
  assign n22454 = x5 &  n22453 ;
  assign n22455 = x5 | n22453 ;
  assign n22456 = ~n22454 & n22455 ;
  assign n22602 = n8764 | n21475 ;
  assign n22599 = n8105 &  n20777 ;
  assign n22600 = n8429 | n21271 ;
  assign n22601 = ~n22599 & n22600 ;
  assign n22603 = ( n8764 & ~n22602 ) | ( n8764 & n22601 ) | ( ~n22602 & n22601 ) ;
  assign n22604 = n8107 | n21484 ;
  assign n22605 = n22603 &  n22604 ;
  assign n22606 = x8 &  n22605 ;
  assign n22607 = x8 | n22605 ;
  assign n22608 = ~n22606 & n22607 ;
  assign n22585 = n7253 &  n20245 ;
  assign n22586 = ~n7518 & n20237 ;
  assign n22587 = n22585 | n22586 ;
  assign n22588 = ~n7783 & n20782 ;
  assign n22589 = ( n7783 & ~n22587 ) | ( n7783 & n22588 ) | ( ~n22587 & n22588 ) ;
  assign n22590 = n7255 | n21227 ;
  assign n22591 = n22589 &  n22590 ;
  assign n22592 = x11 &  n22591 ;
  assign n22593 = x11 | n22591 ;
  assign n22594 = ~n22592 & n22593 ;
  assign n22574 = ~n7097 & n20241 ;
  assign n22571 = n6530 | n19951 ;
  assign n22572 = n6983 | n20027 ;
  assign n22573 = n22571 &  n22572 ;
  assign n22575 = ( n7097 & n22574 ) | ( n7097 & n22573 ) | ( n22574 & n22573 ) ;
  assign n22576 = n6532 | n20280 ;
  assign n22577 = n22575 &  n22576 ;
  assign n22578 = x14 &  n22577 ;
  assign n22579 = x14 | n22577 ;
  assign n22580 = ~n22578 & n22579 ;
  assign n22557 = ~n5970 & n19047 ;
  assign n22558 = ~n6170 & n19040 ;
  assign n22559 = n22557 | n22558 ;
  assign n22560 = ~n6395 & n19494 ;
  assign n22561 = ( n6395 & ~n22559 ) | ( n6395 & n22560 ) | ( ~n22559 & n22560 ) ;
  assign n22562 = n5972 | n19502 ;
  assign n22563 = n22561 &  n22562 ;
  assign n22564 = x17 &  n22563 ;
  assign n22565 = x17 | n22563 ;
  assign n22566 = ~n22564 & n22565 ;
  assign n22546 = ~n5837 & n19043 ;
  assign n22543 = ( n5339 & ~n18589 ) | ( n5339 & 1'b0 ) | ( ~n18589 & 1'b0 ) ;
  assign n22544 = n5761 | n18712 ;
  assign n22545 = ~n22543 & n22544 ;
  assign n22547 = ( n5837 & n22546 ) | ( n5837 & n22545 ) | ( n22546 & n22545 ) ;
  assign n22548 = n5341 | n19083 ;
  assign n22549 = n22547 &  n22548 ;
  assign n22550 = x20 &  n22549 ;
  assign n22551 = x20 | n22549 ;
  assign n22552 = ~n22550 & n22551 ;
  assign n22532 = ~n5135 & n18456 ;
  assign n22529 = n5010 | n17791 ;
  assign n22530 = n5067 | n17783 ;
  assign n22531 = n22529 &  n22530 ;
  assign n22533 = ( n5135 & n22532 ) | ( n5135 & n22531 ) | ( n22532 & n22531 ) ;
  assign n22534 = n5012 | n18464 ;
  assign n22535 = n22533 &  n22534 ;
  assign n22536 = x23 &  n22535 ;
  assign n22537 = x23 | n22535 ;
  assign n22538 = ~n22536 & n22537 ;
  assign n22518 = ~n4962 & n17787 ;
  assign n22515 = n4482 | n17263 ;
  assign n22516 = n4495 | n17405 ;
  assign n22517 = n22515 &  n22516 ;
  assign n22519 = ( n4962 & n22518 ) | ( n4962 & n22517 ) | ( n22518 & n22517 ) ;
  assign n22520 = n4478 | n17826 ;
  assign n22521 = n22519 &  n22520 ;
  assign n22522 = x26 &  n22521 ;
  assign n22523 = x26 | n22521 ;
  assign n22524 = ~n22522 & n22523 ;
  assign n22457 = ( n22303 & ~n22304 ) | ( n22303 & 1'b0 ) | ( ~n22304 & 1'b0 ) ;
  assign n22458 = ( n22304 & ~n22303 ) | ( n22304 & n22314 ) | ( ~n22303 & n22314 ) ;
  assign n22459 = ( n22457 & ~n22318 ) | ( n22457 & n22458 ) | ( ~n22318 & n22458 ) ;
  assign n22481 = n3644 | n16631 ;
  assign n22482 = ( n3652 & ~n15897 ) | ( n3652 & 1'b0 ) | ( ~n15897 & 1'b0 ) ;
  assign n22483 = ( n3657 & ~n16091 ) | ( n3657 & 1'b0 ) | ( ~n16091 & 1'b0 ) ;
  assign n22484 = n22482 | n22483 ;
  assign n22485 = ~n3653 & n16591 ;
  assign n22486 = ( n3653 & ~n22484 ) | ( n3653 & n22485 ) | ( ~n22484 & n22485 ) ;
  assign n22487 = n22481 &  n22486 ;
  assign n22488 = n2945 | n3222 ;
  assign n22489 = ( n22488 & ~n6838 ) | ( n22488 & n18867 ) | ( ~n6838 & n18867 ) ;
  assign n22490 = n6838 | n22489 ;
  assign n22491 = ( n1343 & ~n18935 ) | ( n1343 & n22490 ) | ( ~n18935 & n22490 ) ;
  assign n22492 = ( n1343 & ~n22491 ) | ( n1343 & 1'b0 ) | ( ~n22491 & 1'b0 ) ;
  assign n22493 = ( n843 & n989 ) | ( n843 & n22492 ) | ( n989 & n22492 ) ;
  assign n22494 = ~n843 & n22493 ;
  assign n22495 = ( n1185 & ~n2757 ) | ( n1185 & n22494 ) | ( ~n2757 & n22494 ) ;
  assign n22496 = ~n1185 & n22495 ;
  assign n22497 = ( n785 & ~n22496 ) | ( n785 & n3280 ) | ( ~n22496 & n3280 ) ;
  assign n22498 = ( n3280 & ~n22497 ) | ( n3280 & 1'b0 ) | ( ~n22497 & 1'b0 ) ;
  assign n22499 = ( n194 & ~n218 ) | ( n194 & n22498 ) | ( ~n218 & n22498 ) ;
  assign n22500 = ~n194 & n22499 ;
  assign n22501 = ( n237 & ~n274 ) | ( n237 & n22500 ) | ( ~n274 & n22500 ) ;
  assign n22502 = ~n237 & n22501 ;
  assign n22503 = ( n148 & ~n405 ) | ( n148 & n22502 ) | ( ~n405 & n22502 ) ;
  assign n22504 = ~n148 & n22503 ;
  assign n22505 = ~n104 & n22504 ;
  assign n22506 = n22487 | n22505 ;
  assign n22507 = ~n22487 & n22505 ;
  assign n22508 = ( n22506 & ~n22505 ) | ( n22506 & n22507 ) | ( ~n22505 & n22507 ) ;
  assign n22470 = ~n22057 & n22240 ;
  assign n22471 = ( n22057 & ~n22240 ) | ( n22057 & 1'b0 ) | ( ~n22240 & 1'b0 ) ;
  assign n22472 = n22470 | n22471 ;
  assign n22474 = ( n15737 & n22241 ) | ( n15737 & n22472 ) | ( n22241 & n22472 ) ;
  assign n22473 = n22241 &  n22472 ;
  assign n22475 = ( x2 & ~n22474 ) | ( x2 & n22473 ) | ( ~n22474 & n22473 ) ;
  assign n22476 = ( n22241 & ~x2 ) | ( n22241 & n22472 ) | ( ~x2 & n22472 ) ;
  assign n22477 = ( n22241 & ~n15737 ) | ( n22241 & n22472 ) | ( ~n15737 & n22472 ) ;
  assign n22478 = ( n22476 & ~n22477 ) | ( n22476 & 1'b0 ) | ( ~n22477 & 1'b0 ) ;
  assign n22479 = n22475 | n22478 ;
  assign n22480 = ( n22293 & n22300 ) | ( n22293 & n22304 ) | ( n22300 & n22304 ) ;
  assign n22510 = ( n22479 & n22480 ) | ( n22479 & n22508 ) | ( n22480 & n22508 ) ;
  assign n22509 = ( n22479 & ~n22508 ) | ( n22479 & n22480 ) | ( ~n22508 & n22480 ) ;
  assign n22511 = ( n22508 & ~n22510 ) | ( n22508 & n22509 ) | ( ~n22510 & n22509 ) ;
  assign n22465 = n17115 | n601 ;
  assign n22463 = n17107 | n4430 ;
  assign n22460 = n523 | n16595 ;
  assign n22461 = n3939 | n16589 ;
  assign n22462 = n22460 &  n22461 ;
  assign n22464 = ( n4430 & ~n22463 ) | ( n4430 & n22462 ) | ( ~n22463 & n22462 ) ;
  assign n22466 = ( n601 & ~n22465 ) | ( n601 & n22464 ) | ( ~n22465 & n22464 ) ;
  assign n22467 = x29 &  n22466 ;
  assign n22468 = x29 | n22466 ;
  assign n22469 = ~n22467 & n22468 ;
  assign n22512 = ( n22459 & ~n22511 ) | ( n22459 & n22469 ) | ( ~n22511 & n22469 ) ;
  assign n22513 = ( n22459 & ~n22469 ) | ( n22459 & n22511 ) | ( ~n22469 & n22511 ) ;
  assign n22514 = ( n22512 & ~n22459 ) | ( n22512 & n22513 ) | ( ~n22459 & n22513 ) ;
  assign n22525 = ( n22320 & n22321 ) | ( n22320 & n22331 ) | ( n22321 & n22331 ) ;
  assign n22526 = ( n22524 & ~n22514 ) | ( n22524 & n22525 ) | ( ~n22514 & n22525 ) ;
  assign n22527 = ( n22514 & ~n22524 ) | ( n22514 & n22525 ) | ( ~n22524 & n22525 ) ;
  assign n22528 = ( n22526 & ~n22525 ) | ( n22526 & n22527 ) | ( ~n22525 & n22527 ) ;
  assign n22539 = ( n22334 & n22344 ) | ( n22334 & n22345 ) | ( n22344 & n22345 ) ;
  assign n22540 = ( n22538 & ~n22528 ) | ( n22538 & n22539 ) | ( ~n22528 & n22539 ) ;
  assign n22541 = ( n22528 & ~n22538 ) | ( n22528 & n22539 ) | ( ~n22538 & n22539 ) ;
  assign n22542 = ( n22540 & ~n22539 ) | ( n22540 & n22541 ) | ( ~n22539 & n22541 ) ;
  assign n22553 = ( n22348 & n22349 ) | ( n22348 & n22359 ) | ( n22349 & n22359 ) ;
  assign n22554 = ( n22552 & ~n22542 ) | ( n22552 & n22553 ) | ( ~n22542 & n22553 ) ;
  assign n22555 = ( n22542 & ~n22552 ) | ( n22542 & n22553 ) | ( ~n22552 & n22553 ) ;
  assign n22556 = ( n22554 & ~n22553 ) | ( n22554 & n22555 ) | ( ~n22553 & n22555 ) ;
  assign n22567 = ( n22362 & n22372 ) | ( n22362 & n22373 ) | ( n22372 & n22373 ) ;
  assign n22568 = ( n22566 & ~n22556 ) | ( n22566 & n22567 ) | ( ~n22556 & n22567 ) ;
  assign n22569 = ( n22556 & ~n22566 ) | ( n22556 & n22567 ) | ( ~n22566 & n22567 ) ;
  assign n22570 = ( n22568 & ~n22567 ) | ( n22568 & n22569 ) | ( ~n22567 & n22569 ) ;
  assign n22581 = ( n22376 & n22377 ) | ( n22376 & n22387 ) | ( n22377 & n22387 ) ;
  assign n22582 = ( n22580 & ~n22570 ) | ( n22580 & n22581 ) | ( ~n22570 & n22581 ) ;
  assign n22583 = ( n22570 & ~n22580 ) | ( n22570 & n22581 ) | ( ~n22580 & n22581 ) ;
  assign n22584 = ( n22582 & ~n22581 ) | ( n22582 & n22583 ) | ( ~n22581 & n22583 ) ;
  assign n22595 = ( n22390 & n22400 ) | ( n22390 & n22401 ) | ( n22400 & n22401 ) ;
  assign n22596 = ( n22594 & ~n22584 ) | ( n22594 & n22595 ) | ( ~n22584 & n22595 ) ;
  assign n22597 = ( n22584 & ~n22594 ) | ( n22584 & n22595 ) | ( ~n22594 & n22595 ) ;
  assign n22598 = ( n22596 & ~n22595 ) | ( n22596 & n22597 ) | ( ~n22595 & n22597 ) ;
  assign n22609 = ( n22404 & n22405 ) | ( n22404 & n22415 ) | ( n22405 & n22415 ) ;
  assign n22610 = ( n22608 & ~n22598 ) | ( n22608 & n22609 ) | ( ~n22598 & n22609 ) ;
  assign n22611 = ( n22598 & ~n22608 ) | ( n22598 & n22609 ) | ( ~n22608 & n22609 ) ;
  assign n22612 = ( n22610 & ~n22609 ) | ( n22610 & n22611 ) | ( ~n22609 & n22611 ) ;
  assign n22613 = ( n22418 & n22428 ) | ( n22418 & n22436 ) | ( n22428 & n22436 ) ;
  assign n22614 = ( n22456 & n22612 ) | ( n22456 & n22613 ) | ( n22612 & n22613 ) ;
  assign n22615 = ( n22612 & ~n22456 ) | ( n22612 & n22613 ) | ( ~n22456 & n22613 ) ;
  assign n22616 = ( n22456 & ~n22614 ) | ( n22456 & n22615 ) | ( ~n22614 & n22615 ) ;
  assign n22617 = ( n22265 & n22439 ) | ( n22265 & n22440 ) | ( n22439 & n22440 ) ;
  assign n22619 = ( n22444 & n22616 ) | ( n22444 & n22617 ) | ( n22616 & n22617 ) ;
  assign n22618 = ( n22444 & ~n22616 ) | ( n22444 & n22617 ) | ( ~n22616 & n22617 ) ;
  assign n22620 = ( n22616 & ~n22619 ) | ( n22616 & n22618 ) | ( ~n22619 & n22618 ) ;
  assign n22621 = ( n22616 & ~n22262 ) | ( n22616 & n22617 ) | ( ~n22262 & n22617 ) ;
  assign n22622 = ( n22616 & ~n22443 ) | ( n22616 & n22617 ) | ( ~n22443 & n22617 ) ;
  assign n22623 = ~n22621 & n22622 ;
  assign n22646 = ( n22487 & ~n22479 ) | ( n22487 & n22505 ) | ( ~n22479 & n22505 ) ;
  assign n22657 = ( n22479 & ~n22487 ) | ( n22479 & n22505 ) | ( ~n22487 & n22505 ) ;
  assign n22658 = ( n22646 & ~n22505 ) | ( n22646 & n22657 ) | ( ~n22505 & n22657 ) ;
  assign n22659 = ( n22469 & ~n22658 ) | ( n22469 & n22480 ) | ( ~n22658 & n22480 ) ;
  assign n22624 = ( n645 & ~n11283 ) | ( n645 & 1'b0 ) | ( ~n11283 & 1'b0 ) ;
  assign n22625 = ( n374 & ~n722 ) | ( n374 & n22624 ) | ( ~n722 & n22624 ) ;
  assign n22626 = ~n374 & n22625 ;
  assign n22627 = ~n229 & n22626 ;
  assign n22628 = n736 | n14010 ;
  assign n22629 = ( n3214 & ~n2346 ) | ( n3214 & n22628 ) | ( ~n2346 & n22628 ) ;
  assign n22630 = n2346 | n22629 ;
  assign n22631 = ( n11353 & ~n22627 ) | ( n11353 & n22630 ) | ( ~n22627 & n22630 ) ;
  assign n22632 = ( n11353 & ~n22631 ) | ( n11353 & 1'b0 ) | ( ~n22631 & 1'b0 ) ;
  assign n22633 = ( n2247 & ~n2687 ) | ( n2247 & n22632 ) | ( ~n2687 & n22632 ) ;
  assign n22634 = ( n22633 & ~n2247 ) | ( n22633 & 1'b0 ) | ( ~n2247 & 1'b0 ) ;
  assign n22635 = ( n1876 & ~n675 ) | ( n1876 & n22634 ) | ( ~n675 & n22634 ) ;
  assign n22636 = ~n1876 & n22635 ;
  assign n22637 = ( n1567 & ~n865 ) | ( n1567 & n22636 ) | ( ~n865 & n22636 ) ;
  assign n22638 = ~n1567 & n22637 ;
  assign n22639 = ( n22638 & ~n414 ) | ( n22638 & n2936 ) | ( ~n414 & n2936 ) ;
  assign n22640 = ( n22639 & ~n2936 ) | ( n22639 & 1'b0 ) | ( ~n2936 & 1'b0 ) ;
  assign n22641 = ( n273 & ~n357 ) | ( n273 & n22640 ) | ( ~n357 & n22640 ) ;
  assign n22642 = ~n273 & n22641 ;
  assign n22643 = ( n279 & ~n646 ) | ( n279 & n22642 ) | ( ~n646 & n22642 ) ;
  assign n22644 = ~n279 & n22643 ;
  assign n22645 = ~n83 & n22644 ;
  assign n22647 = ( n22479 & ~n22645 ) | ( n22479 & n22646 ) | ( ~n22645 & n22646 ) ;
  assign n22648 = ( n22645 & ~n22479 ) | ( n22645 & n22646 ) | ( ~n22479 & n22646 ) ;
  assign n22649 = ( n22647 & ~n22646 ) | ( n22647 & n22648 ) | ( ~n22646 & n22648 ) ;
  assign n22650 = n3644 | n16616 ;
  assign n22651 = ( n3652 & ~n16091 ) | ( n3652 & 1'b0 ) | ( ~n16091 & 1'b0 ) ;
  assign n22652 = ( n3657 & ~n16591 ) | ( n3657 & 1'b0 ) | ( ~n16591 & 1'b0 ) ;
  assign n22653 = n22651 | n22652 ;
  assign n22654 = ~n3653 & n16595 ;
  assign n22655 = ( n3653 & ~n22653 ) | ( n3653 & n22654 ) | ( ~n22653 & n22654 ) ;
  assign n22656 = n22650 &  n22655 ;
  assign n22660 = ( n22649 & n22656 ) | ( n22649 & n22659 ) | ( n22656 & n22659 ) ;
  assign n22661 = ( n22649 & ~n22659 ) | ( n22649 & n22656 ) | ( ~n22659 & n22656 ) ;
  assign n22662 = ( n22659 & ~n22660 ) | ( n22659 & n22661 ) | ( ~n22660 & n22661 ) ;
  assign n22666 = ~n4962 & n17791 ;
  assign n22663 = n4482 | n17405 ;
  assign n22664 = n4495 | n17787 ;
  assign n22665 = n22663 &  n22664 ;
  assign n22667 = ( n4962 & n22666 ) | ( n4962 & n22665 ) | ( n22666 & n22665 ) ;
  assign n22668 = n4478 | n17811 ;
  assign n22669 = n22667 &  n22668 ;
  assign n22670 = x26 &  n22669 ;
  assign n22671 = x26 | n22669 ;
  assign n22672 = ~n22670 & n22671 ;
  assign n22676 = ~n4430 & n17263 ;
  assign n22673 = n523 | n16589 ;
  assign n22674 = ~n3939 & n17107 ;
  assign n22675 = ( n22673 & ~n22674 ) | ( n22673 & 1'b0 ) | ( ~n22674 & 1'b0 ) ;
  assign n22677 = ( n4430 & n22676 ) | ( n4430 & n22675 ) | ( n22676 & n22675 ) ;
  assign n22678 = ~n601 & n17271 ;
  assign n22679 = ( n22677 & ~n22678 ) | ( n22677 & 1'b0 ) | ( ~n22678 & 1'b0 ) ;
  assign n22680 = x29 &  n22679 ;
  assign n22681 = x29 | n22679 ;
  assign n22682 = ~n22680 & n22681 ;
  assign n22683 = ( n22662 & n22672 ) | ( n22662 & n22682 ) | ( n22672 & n22682 ) ;
  assign n22684 = ( n22672 & ~n22662 ) | ( n22672 & n22682 ) | ( ~n22662 & n22682 ) ;
  assign n22685 = ( n22662 & ~n22683 ) | ( n22662 & n22684 ) | ( ~n22683 & n22684 ) ;
  assign n22686 = n22469 &  n22511 ;
  assign n22687 = n22469 | n22511 ;
  assign n22688 = ~n22686 & n22687 ;
  assign n22689 = ( n22459 & ~n22688 ) | ( n22459 & n22524 ) | ( ~n22688 & n22524 ) ;
  assign n22693 = ~n5135 & n18589 ;
  assign n22690 = n5010 | n17783 ;
  assign n22691 = n5067 | n18456 ;
  assign n22692 = n22690 &  n22691 ;
  assign n22694 = ( n5135 & n22693 ) | ( n5135 & n22692 ) | ( n22693 & n22692 ) ;
  assign n22695 = n5012 | n18597 ;
  assign n22696 = n22694 &  n22695 ;
  assign n22697 = x23 &  n22696 ;
  assign n22698 = x23 | n22696 ;
  assign n22699 = ~n22697 & n22698 ;
  assign n22701 = ( n22685 & n22689 ) | ( n22685 & n22699 ) | ( n22689 & n22699 ) ;
  assign n22700 = ( n22689 & ~n22685 ) | ( n22689 & n22699 ) | ( ~n22685 & n22699 ) ;
  assign n22702 = ( n22685 & ~n22701 ) | ( n22685 & n22700 ) | ( ~n22701 & n22700 ) ;
  assign n22703 = n22514 &  n22524 ;
  assign n22704 = n22514 | n22524 ;
  assign n22705 = ~n22703 & n22704 ;
  assign n22706 = ( n22525 & ~n22705 ) | ( n22525 & n22538 ) | ( ~n22705 & n22538 ) ;
  assign n22710 = n19047 | n5837 ;
  assign n22707 = ( n5339 & ~n18712 ) | ( n5339 & 1'b0 ) | ( ~n18712 & 1'b0 ) ;
  assign n22708 = n5761 | n19043 ;
  assign n22709 = ~n22707 & n22708 ;
  assign n22711 = ( n5837 & ~n22710 ) | ( n5837 & n22709 ) | ( ~n22710 & n22709 ) ;
  assign n22712 = ~n5341 & n19068 ;
  assign n22713 = ( n22711 & ~n22712 ) | ( n22711 & 1'b0 ) | ( ~n22712 & 1'b0 ) ;
  assign n22714 = x20 &  n22713 ;
  assign n22715 = x20 | n22713 ;
  assign n22716 = ~n22714 & n22715 ;
  assign n22718 = ( n22702 & n22706 ) | ( n22702 & n22716 ) | ( n22706 & n22716 ) ;
  assign n22717 = ( n22706 & ~n22702 ) | ( n22706 & n22716 ) | ( ~n22702 & n22716 ) ;
  assign n22719 = ( n22702 & ~n22718 ) | ( n22702 & n22717 ) | ( ~n22718 & n22717 ) ;
  assign n22723 = ~n6395 & n19951 ;
  assign n22720 = ~n5970 & n19040 ;
  assign n22721 = n6170 | n19494 ;
  assign n22722 = ~n22720 & n22721 ;
  assign n22724 = ( n6395 & n22723 ) | ( n6395 & n22722 ) | ( n22723 & n22722 ) ;
  assign n22725 = ~n5972 & n19959 ;
  assign n22726 = ( n22724 & ~n22725 ) | ( n22724 & 1'b0 ) | ( ~n22725 & 1'b0 ) ;
  assign n22727 = x17 &  n22726 ;
  assign n22728 = x17 | n22726 ;
  assign n22729 = ~n22727 & n22728 ;
  assign n22730 = ~n22528 & n22538 ;
  assign n22731 = ( n22528 & ~n22538 ) | ( n22528 & 1'b0 ) | ( ~n22538 & 1'b0 ) ;
  assign n22732 = n22730 | n22731 ;
  assign n22733 = ( n22539 & ~n22732 ) | ( n22539 & n22552 ) | ( ~n22732 & n22552 ) ;
  assign n22735 = ( n22719 & n22729 ) | ( n22719 & n22733 ) | ( n22729 & n22733 ) ;
  assign n22734 = ( n22729 & ~n22719 ) | ( n22729 & n22733 ) | ( ~n22719 & n22733 ) ;
  assign n22736 = ( n22719 & ~n22735 ) | ( n22719 & n22734 ) | ( ~n22735 & n22734 ) ;
  assign n22740 = n20245 | n7097 ;
  assign n22737 = n6530 | n20027 ;
  assign n22738 = n6983 | n20241 ;
  assign n22739 = n22737 &  n22738 ;
  assign n22741 = ( n7097 & ~n22740 ) | ( n7097 & n22739 ) | ( ~n22740 & n22739 ) ;
  assign n22742 = ~n6532 & n20265 ;
  assign n22743 = ( n22741 & ~n22742 ) | ( n22741 & 1'b0 ) | ( ~n22742 & 1'b0 ) ;
  assign n22744 = x14 &  n22743 ;
  assign n22745 = x14 | n22743 ;
  assign n22746 = ~n22744 & n22745 ;
  assign n22748 = ( x20 & n22542 ) | ( x20 & n22549 ) | ( n22542 & n22549 ) ;
  assign n22747 = ( n22542 & ~x20 ) | ( n22542 & n22549 ) | ( ~x20 & n22549 ) ;
  assign n22749 = ( x20 & ~n22748 ) | ( x20 & n22747 ) | ( ~n22748 & n22747 ) ;
  assign n22750 = ( n22553 & ~n22749 ) | ( n22553 & n22566 ) | ( ~n22749 & n22566 ) ;
  assign n22752 = ( n22736 & n22746 ) | ( n22736 & n22750 ) | ( n22746 & n22750 ) ;
  assign n22751 = ( n22746 & ~n22736 ) | ( n22746 & n22750 ) | ( ~n22736 & n22750 ) ;
  assign n22753 = ( n22736 & ~n22752 ) | ( n22736 & n22751 ) | ( ~n22752 & n22751 ) ;
  assign n22757 = n7783 | n20777 ;
  assign n22754 = n7253 &  n20237 ;
  assign n22755 = n7518 | n20782 ;
  assign n22756 = ~n22754 & n22755 ;
  assign n22758 = ( n7783 & ~n22757 ) | ( n7783 & n22756 ) | ( ~n22757 & n22756 ) ;
  assign n22759 = n7255 | n20790 ;
  assign n22760 = n22758 &  n22759 ;
  assign n22761 = x11 &  n22760 ;
  assign n22762 = x11 | n22760 ;
  assign n22763 = ~n22761 & n22762 ;
  assign n22765 = ( x17 & n22556 ) | ( x17 & n22563 ) | ( n22556 & n22563 ) ;
  assign n22764 = ( n22556 & ~x17 ) | ( n22556 & n22563 ) | ( ~x17 & n22563 ) ;
  assign n22766 = ( x17 & ~n22765 ) | ( x17 & n22764 ) | ( ~n22765 & n22764 ) ;
  assign n22767 = ( n22567 & ~n22766 ) | ( n22567 & n22580 ) | ( ~n22766 & n22580 ) ;
  assign n22769 = ( n22753 & n22763 ) | ( n22753 & n22767 ) | ( n22763 & n22767 ) ;
  assign n22768 = ( n22763 & ~n22753 ) | ( n22763 & n22767 ) | ( ~n22753 & n22767 ) ;
  assign n22770 = ( n22753 & ~n22769 ) | ( n22753 & n22768 ) | ( ~n22769 & n22768 ) ;
  assign n22771 = ( n8105 & ~n21271 ) | ( n8105 & 1'b0 ) | ( ~n21271 & 1'b0 ) ;
  assign n22772 = ~n8429 & n21475 ;
  assign n22773 = n22771 | n22772 ;
  assign n22774 = ~n8764 & n21675 ;
  assign n22775 = ( n8764 & ~n22773 ) | ( n8764 & n22774 ) | ( ~n22773 & n22774 ) ;
  assign n22776 = n8107 | n21684 ;
  assign n22777 = n22775 &  n22776 ;
  assign n22778 = x8 &  n22777 ;
  assign n22779 = x8 | n22777 ;
  assign n22780 = ~n22778 & n22779 ;
  assign n22782 = ( x14 & n22570 ) | ( x14 & n22577 ) | ( n22570 & n22577 ) ;
  assign n22781 = ( n22570 & ~x14 ) | ( n22570 & n22577 ) | ( ~x14 & n22577 ) ;
  assign n22783 = ( x14 & ~n22782 ) | ( x14 & n22781 ) | ( ~n22782 & n22781 ) ;
  assign n22784 = ( n22581 & ~n22783 ) | ( n22581 & n22594 ) | ( ~n22783 & n22594 ) ;
  assign n22786 = ( n22770 & n22780 ) | ( n22770 & n22784 ) | ( n22780 & n22784 ) ;
  assign n22785 = ( n22780 & ~n22770 ) | ( n22780 & n22784 ) | ( ~n22770 & n22784 ) ;
  assign n22787 = ( n22770 & ~n22786 ) | ( n22770 & n22785 ) | ( ~n22786 & n22785 ) ;
  assign n22791 = n22244 | n9997 ;
  assign n22788 = n9160 | n21864 ;
  assign n22789 = n9558 | n22063 ;
  assign n22790 = n22788 &  n22789 ;
  assign n22792 = ( n9997 & ~n22791 ) | ( n9997 & n22790 ) | ( ~n22791 & n22790 ) ;
  assign n22793 = ~n9155 & n22253 ;
  assign n22794 = ( n22792 & ~n22793 ) | ( n22792 & 1'b0 ) | ( ~n22793 & 1'b0 ) ;
  assign n22795 = x5 &  n22794 ;
  assign n22796 = x5 | n22794 ;
  assign n22797 = ~n22795 & n22796 ;
  assign n22799 = ( x11 & n22584 ) | ( x11 & n22591 ) | ( n22584 & n22591 ) ;
  assign n22798 = ( n22584 & ~x11 ) | ( n22584 & n22591 ) | ( ~x11 & n22591 ) ;
  assign n22800 = ( x11 & ~n22799 ) | ( x11 & n22798 ) | ( ~n22799 & n22798 ) ;
  assign n22801 = ( n22595 & ~n22800 ) | ( n22595 & n22608 ) | ( ~n22800 & n22608 ) ;
  assign n22803 = ( n22787 & n22797 ) | ( n22787 & n22801 ) | ( n22797 & n22801 ) ;
  assign n22802 = ( n22797 & ~n22787 ) | ( n22797 & n22801 ) | ( ~n22787 & n22801 ) ;
  assign n22804 = ( n22787 & ~n22803 ) | ( n22787 & n22802 ) | ( ~n22803 & n22802 ) ;
  assign n22806 = ( x8 & n22598 ) | ( x8 & n22605 ) | ( n22598 & n22605 ) ;
  assign n22805 = ( n22598 & ~x8 ) | ( n22598 & n22605 ) | ( ~x8 & n22605 ) ;
  assign n22807 = ( x8 & ~n22806 ) | ( x8 & n22805 ) | ( ~n22806 & n22805 ) ;
  assign n22808 = ~n22609 & n22807 ;
  assign n22809 = n22456 | n22612 ;
  assign n22810 = ~n22808 & n22809 ;
  assign n22811 = ~n22456 & n22612 ;
  assign n22812 = ( n22456 & ~n22612 ) | ( n22456 & 1'b0 ) | ( ~n22612 & 1'b0 ) ;
  assign n22813 = n22811 | n22812 ;
  assign n22814 = ( n22613 & ~n22813 ) | ( n22613 & n22617 ) | ( ~n22813 & n22617 ) ;
  assign n22816 = ( n22804 & n22810 ) | ( n22804 & n22814 ) | ( n22810 & n22814 ) ;
  assign n22815 = ( n22810 & ~n22804 ) | ( n22810 & n22814 ) | ( ~n22804 & n22814 ) ;
  assign n22817 = ( n22804 & ~n22816 ) | ( n22804 & n22815 ) | ( ~n22816 & n22815 ) ;
  assign n22818 = n22623 &  n22817 ;
  assign n22819 = n22623 | n22817 ;
  assign n22820 = ~n22818 & n22819 ;
  assign n22958 = ~n9155 & n22251 ;
  assign n22955 = ~n16564 & n22244 ;
  assign n22956 = n9160 | n22063 ;
  assign n22957 = ~n22955 & n22956 ;
  assign n22959 = ( n9155 & n22958 ) | ( n9155 & n22957 ) | ( n22958 & n22957 ) ;
  assign n22960 = ( x5 & ~n22785 ) | ( x5 & n22959 ) | ( ~n22785 & n22959 ) ;
  assign n22961 = ( x5 & ~n22959 ) | ( x5 & n22785 ) | ( ~n22959 & n22785 ) ;
  assign n22962 = ( n22960 & ~x5 ) | ( n22960 & n22961 ) | ( ~x5 & n22961 ) ;
  assign n22821 = ( n7253 & ~n20782 ) | ( n7253 & 1'b0 ) | ( ~n20782 & 1'b0 ) ;
  assign n22822 = ~n7518 & n20777 ;
  assign n22823 = n22821 | n22822 ;
  assign n22824 = ~n7783 & n21271 ;
  assign n22825 = ( n7783 & ~n22823 ) | ( n7783 & n22824 ) | ( ~n22823 & n22824 ) ;
  assign n22826 = n7255 | n21279 ;
  assign n22827 = n22825 &  n22826 ;
  assign n22828 = x11 &  n22827 ;
  assign n22829 = x11 | n22827 ;
  assign n22830 = ~n22828 & n22829 ;
  assign n22926 = n7097 &  n20237 ;
  assign n22927 = n6530 | n20241 ;
  assign n22928 = ~n6983 & n20245 ;
  assign n22929 = ( n22927 & ~n22928 ) | ( n22927 & 1'b0 ) | ( ~n22928 & 1'b0 ) ;
  assign n22930 = ( n22926 & ~n20237 ) | ( n22926 & n22929 ) | ( ~n20237 & n22929 ) ;
  assign n22931 = n6532 | n20253 ;
  assign n22932 = n22930 &  n22931 ;
  assign n22933 = x14 &  n22932 ;
  assign n22934 = x14 | n22932 ;
  assign n22935 = ~n22933 & n22934 ;
  assign n22831 = ( n4962 & ~n17783 ) | ( n4962 & 1'b0 ) | ( ~n17783 & 1'b0 ) ;
  assign n22832 = n4482 | n17787 ;
  assign n22833 = n4495 | n17791 ;
  assign n22834 = n22832 &  n22833 ;
  assign n22835 = ( n17783 & n22831 ) | ( n17783 & n22834 ) | ( n22831 & n22834 ) ;
  assign n22836 = n4478 | n17799 ;
  assign n22837 = n22835 &  n22836 ;
  assign n22838 = x26 &  n22837 ;
  assign n22839 = x26 | n22837 ;
  assign n22840 = ~n22838 & n22839 ;
  assign n22841 = n3228 | n15940 ;
  assign n22842 = ( n3569 & ~n2062 ) | ( n3569 & n22841 ) | ( ~n2062 & n22841 ) ;
  assign n22843 = n2062 | n22842 ;
  assign n22844 = ( n5582 & ~n4118 ) | ( n5582 & n22843 ) | ( ~n4118 & n22843 ) ;
  assign n22845 = n4118 | n22844 ;
  assign n22846 = ( n1579 & ~n22845 ) | ( n1579 & n1794 ) | ( ~n22845 & n1794 ) ;
  assign n22847 = ( n22846 & ~n1579 ) | ( n22846 & 1'b0 ) | ( ~n1579 & 1'b0 ) ;
  assign n22848 = ( n1061 & ~n3245 ) | ( n1061 & n22847 ) | ( ~n3245 & n22847 ) ;
  assign n22849 = ~n1061 & n22848 ;
  assign n22850 = ( n947 & ~n3009 ) | ( n947 & n22849 ) | ( ~n3009 & n22849 ) ;
  assign n22851 = ~n947 & n22850 ;
  assign n22852 = ( n362 & ~n425 ) | ( n362 & n22851 ) | ( ~n425 & n22851 ) ;
  assign n22853 = ~n362 & n22852 ;
  assign n22854 = ( n22853 & ~n676 ) | ( n22853 & n796 ) | ( ~n676 & n796 ) ;
  assign n22855 = ( n22854 & ~n796 ) | ( n22854 & 1'b0 ) | ( ~n796 & 1'b0 ) ;
  assign n22856 = ~n285 & n22855 ;
  assign n22857 = ( n22479 & ~n22856 ) | ( n22479 & 1'b0 ) | ( ~n22856 & 1'b0 ) ;
  assign n22858 = ~n22479 & n22856 ;
  assign n22859 = n22857 | n22858 ;
  assign n22860 = n3644 | n16604 ;
  assign n22861 = ( n3652 & ~n16591 ) | ( n3652 & 1'b0 ) | ( ~n16591 & 1'b0 ) ;
  assign n22862 = ( n3657 & ~n16595 ) | ( n3657 & 1'b0 ) | ( ~n16595 & 1'b0 ) ;
  assign n22863 = n22861 | n22862 ;
  assign n22864 = ~n3653 & n16589 ;
  assign n22865 = ( n3653 & ~n22863 ) | ( n3653 & n22864 ) | ( ~n22863 & n22864 ) ;
  assign n22866 = n22860 &  n22865 ;
  assign n22867 = ( n22648 & ~n22859 ) | ( n22648 & n22866 ) | ( ~n22859 & n22866 ) ;
  assign n22868 = ( n22859 & ~n22648 ) | ( n22859 & n22866 ) | ( ~n22648 & n22866 ) ;
  assign n22869 = ( n22867 & ~n22866 ) | ( n22867 & n22868 ) | ( ~n22866 & n22868 ) ;
  assign n22873 = ~n4430 & n17405 ;
  assign n22870 = ~n523 & n17107 ;
  assign n22871 = n3939 | n17263 ;
  assign n22872 = ~n22870 & n22871 ;
  assign n22874 = ( n4430 & n22873 ) | ( n4430 & n22872 ) | ( n22873 & n22872 ) ;
  assign n22875 = n601 | n17413 ;
  assign n22876 = n22874 &  n22875 ;
  assign n22877 = x29 &  n22876 ;
  assign n22878 = x29 | n22876 ;
  assign n22879 = ~n22877 & n22878 ;
  assign n22880 = ( n22656 & ~n22649 ) | ( n22656 & n22659 ) | ( ~n22649 & n22659 ) ;
  assign n22881 = ( n22869 & n22879 ) | ( n22869 & n22880 ) | ( n22879 & n22880 ) ;
  assign n22882 = ( n22879 & ~n22869 ) | ( n22879 & n22880 ) | ( ~n22869 & n22880 ) ;
  assign n22883 = ( n22869 & ~n22881 ) | ( n22869 & n22882 ) | ( ~n22881 & n22882 ) ;
  assign n22884 = ( n22684 & n22840 ) | ( n22684 & n22883 ) | ( n22840 & n22883 ) ;
  assign n22885 = ( n22840 & ~n22684 ) | ( n22840 & n22883 ) | ( ~n22684 & n22883 ) ;
  assign n22886 = ( n22684 & ~n22884 ) | ( n22684 & n22885 ) | ( ~n22884 & n22885 ) ;
  assign n22890 = ~n5135 & n18712 ;
  assign n22887 = n5010 | n18456 ;
  assign n22888 = n5067 | n18589 ;
  assign n22889 = n22887 &  n22888 ;
  assign n22891 = ( n5135 & n22890 ) | ( n5135 & n22889 ) | ( n22890 & n22889 ) ;
  assign n22892 = n5012 | n18720 ;
  assign n22893 = n22891 &  n22892 ;
  assign n22894 = x23 &  n22893 ;
  assign n22895 = x23 | n22893 ;
  assign n22896 = ~n22894 & n22895 ;
  assign n22897 = ( n22700 & ~n22886 ) | ( n22700 & n22896 ) | ( ~n22886 & n22896 ) ;
  assign n22898 = ( n22700 & ~n22896 ) | ( n22700 & n22886 ) | ( ~n22896 & n22886 ) ;
  assign n22899 = ( n22897 & ~n22700 ) | ( n22897 & n22898 ) | ( ~n22700 & n22898 ) ;
  assign n22903 = n19040 | n5837 ;
  assign n22900 = ( n5339 & ~n19043 ) | ( n5339 & 1'b0 ) | ( ~n19043 & 1'b0 ) ;
  assign n22901 = ~n5761 & n19047 ;
  assign n22902 = n22900 | n22901 ;
  assign n22904 = ( n22903 & ~n5837 ) | ( n22903 & n22902 ) | ( ~n5837 & n22902 ) ;
  assign n22905 = n5341 | n19056 ;
  assign n22906 = ~n22904 & n22905 ;
  assign n22907 = x20 &  n22906 ;
  assign n22908 = x20 | n22906 ;
  assign n22909 = ~n22907 & n22908 ;
  assign n22910 = ( n22717 & ~n22899 ) | ( n22717 & n22909 ) | ( ~n22899 & n22909 ) ;
  assign n22911 = ( n22717 & ~n22909 ) | ( n22717 & n22899 ) | ( ~n22909 & n22899 ) ;
  assign n22912 = ( n22910 & ~n22717 ) | ( n22910 & n22911 ) | ( ~n22717 & n22911 ) ;
  assign n22916 = ~n6395 & n20027 ;
  assign n22913 = n5970 | n19494 ;
  assign n22914 = n6170 | n19951 ;
  assign n22915 = n22913 &  n22914 ;
  assign n22917 = ( n6395 & n22916 ) | ( n6395 & n22915 ) | ( n22916 & n22915 ) ;
  assign n22918 = n5972 | n20035 ;
  assign n22919 = n22917 &  n22918 ;
  assign n22920 = x17 &  n22919 ;
  assign n22921 = x17 | n22919 ;
  assign n22922 = ~n22920 & n22921 ;
  assign n22923 = ( n22734 & ~n22912 ) | ( n22734 & n22922 ) | ( ~n22912 & n22922 ) ;
  assign n22924 = ( n22734 & ~n22922 ) | ( n22734 & n22912 ) | ( ~n22922 & n22912 ) ;
  assign n22925 = ( n22923 & ~n22734 ) | ( n22923 & n22924 ) | ( ~n22734 & n22924 ) ;
  assign n22937 = n22925 &  n22935 ;
  assign n22936 = ( n22925 & ~n22935 ) | ( n22925 & 1'b0 ) | ( ~n22935 & 1'b0 ) ;
  assign n22938 = ( n22935 & ~n22937 ) | ( n22935 & n22936 ) | ( ~n22937 & n22936 ) ;
  assign n22939 = ( n22830 & ~n22751 ) | ( n22830 & n22938 ) | ( ~n22751 & n22938 ) ;
  assign n22940 = ( n22751 & ~n22830 ) | ( n22751 & n22938 ) | ( ~n22830 & n22938 ) ;
  assign n22941 = ( n22939 & ~n22938 ) | ( n22939 & n22940 ) | ( ~n22938 & n22940 ) ;
  assign n22945 = ~n8764 & n21864 ;
  assign n22942 = n8105 &  n21475 ;
  assign n22943 = n8429 | n21675 ;
  assign n22944 = ~n22942 & n22943 ;
  assign n22946 = ( n8764 & n22945 ) | ( n8764 & n22944 ) | ( n22945 & n22944 ) ;
  assign n22947 = ~n8107 & n21872 ;
  assign n22948 = ( n22946 & ~n22947 ) | ( n22946 & 1'b0 ) | ( ~n22947 & 1'b0 ) ;
  assign n22949 = x8 &  n22948 ;
  assign n22950 = x8 | n22948 ;
  assign n22951 = ~n22949 & n22950 ;
  assign n22953 = ( n22768 & n22941 ) | ( n22768 & n22951 ) | ( n22941 & n22951 ) ;
  assign n22952 = ( n22768 & ~n22941 ) | ( n22768 & n22951 ) | ( ~n22941 & n22951 ) ;
  assign n22954 = ( n22941 & ~n22953 ) | ( n22941 & n22952 ) | ( ~n22953 & n22952 ) ;
  assign n22964 = n22954 &  n22962 ;
  assign n22963 = ( n22954 & ~n22962 ) | ( n22954 & 1'b0 ) | ( ~n22962 & 1'b0 ) ;
  assign n22965 = ( n22962 & ~n22964 ) | ( n22962 & n22963 ) | ( ~n22964 & n22963 ) ;
  assign n22966 = ( n22815 & ~n22802 ) | ( n22815 & n22965 ) | ( ~n22802 & n22965 ) ;
  assign n22967 = ( n22802 & ~n22815 ) | ( n22802 & n22965 ) | ( ~n22815 & n22965 ) ;
  assign n22968 = ( n22966 & ~n22965 ) | ( n22966 & n22967 ) | ( ~n22965 & n22967 ) ;
  assign n22969 = n22818 &  n22968 ;
  assign n22970 = n22818 | n22968 ;
  assign n22971 = ~n22969 & n22970 ;
  assign n22972 = ~n22954 & n22962 ;
  assign n22973 = n22963 | n22972 ;
  assign n22974 = ( n22802 & ~n22973 ) | ( n22802 & n22815 ) | ( ~n22973 & n22815 ) ;
  assign n22975 = ( x5 & ~n22959 ) | ( x5 & 1'b0 ) | ( ~n22959 & 1'b0 ) ;
  assign n22976 = ~x5 & n22959 ;
  assign n22977 = n22975 | n22976 ;
  assign n22978 = ( n22785 & ~n22954 ) | ( n22785 & n22977 ) | ( ~n22954 & n22977 ) ;
  assign n23124 = ( x14 & n22925 ) | ( x14 & n22932 ) | ( n22925 & n22932 ) ;
  assign n23123 = ( n22925 & ~x14 ) | ( n22925 & n22932 ) | ( ~x14 & n22932 ) ;
  assign n23125 = ( x14 & ~n23124 ) | ( x14 & n23123 ) | ( ~n23124 & n23123 ) ;
  assign n23126 = ( n22751 & ~n23125 ) | ( n22751 & n22830 ) | ( ~n23125 & n22830 ) ;
  assign n23090 = ( x20 & n22899 ) | ( x20 & n22906 ) | ( n22899 & n22906 ) ;
  assign n23089 = ( n22899 & ~x20 ) | ( n22899 & n22906 ) | ( ~x20 & n22906 ) ;
  assign n23091 = ( x20 & ~n23090 ) | ( x20 & n23089 ) | ( ~n23090 & n23089 ) ;
  assign n23092 = ( n22717 & ~n23091 ) | ( n22717 & n22922 ) | ( ~n23091 & n22922 ) ;
  assign n23073 = ( x23 & n22886 ) | ( x23 & n22893 ) | ( n22886 & n22893 ) ;
  assign n23072 = ( n22886 & ~x23 ) | ( n22886 & n22893 ) | ( ~x23 & n22893 ) ;
  assign n23074 = ( x23 & ~n23073 ) | ( x23 & n23072 ) | ( ~n23073 & n23072 ) ;
  assign n23075 = ( n22700 & ~n23074 ) | ( n22700 & n22909 ) | ( ~n23074 & n22909 ) ;
  assign n23055 = ( x26 & ~n22837 ) | ( x26 & n22883 ) | ( ~n22837 & n22883 ) ;
  assign n23056 = ( x26 & ~n22883 ) | ( x26 & n22837 ) | ( ~n22883 & n22837 ) ;
  assign n23057 = ( n23055 & ~x26 ) | ( n23055 & n23056 ) | ( ~x26 & n23056 ) ;
  assign n23058 = ( n22684 & ~n23057 ) | ( n22684 & n22896 ) | ( ~n23057 & n22896 ) ;
  assign n22979 = n22869 | n22880 ;
  assign n22980 = ( n22869 & ~n22880 ) | ( n22869 & 1'b0 ) | ( ~n22880 & 1'b0 ) ;
  assign n22981 = ( n22979 & ~n22869 ) | ( n22979 & n22980 ) | ( ~n22869 & n22980 ) ;
  assign n22982 = ( n22840 & ~n22981 ) | ( n22840 & n22879 ) | ( ~n22981 & n22879 ) ;
  assign n22993 = ( n22479 & ~n22856 ) | ( n22479 & n22648 ) | ( ~n22856 & n22648 ) ;
  assign n22994 = ( n22648 & ~n22479 ) | ( n22648 & n22856 ) | ( ~n22479 & n22856 ) ;
  assign n22995 = ( n22993 & ~n22648 ) | ( n22993 & n22994 ) | ( ~n22648 & n22994 ) ;
  assign n22996 = ( n22866 & ~n22995 ) | ( n22866 & n22880 ) | ( ~n22995 & n22880 ) ;
  assign n23000 = ~n4430 & n17787 ;
  assign n22997 = n523 | n17263 ;
  assign n22998 = n3939 | n17405 ;
  assign n22999 = n22997 &  n22998 ;
  assign n23001 = ( n4430 & n23000 ) | ( n4430 & n22999 ) | ( n23000 & n22999 ) ;
  assign n23002 = n601 | n17826 ;
  assign n23003 = n23001 &  n23002 ;
  assign n23004 = x29 &  n23003 ;
  assign n23005 = x29 | n23003 ;
  assign n23006 = ~n23004 & n23005 ;
  assign n23011 = ( n2733 & ~n4842 ) | ( n2733 & 1'b0 ) | ( ~n4842 & 1'b0 ) ;
  assign n23012 = ( n2036 & ~n4859 ) | ( n2036 & n23011 ) | ( ~n4859 & n23011 ) ;
  assign n23013 = ~n2036 & n23012 ;
  assign n23014 = ( n629 & ~n1949 ) | ( n629 & n23013 ) | ( ~n1949 & n23013 ) ;
  assign n23015 = ~n629 & n23014 ;
  assign n23016 = ( n18541 & ~n4242 ) | ( n18541 & n23015 ) | ( ~n4242 & n23015 ) ;
  assign n23017 = n4242 &  n23016 ;
  assign n23018 = ( n102 & ~n884 ) | ( n102 & n23017 ) | ( ~n884 & n23017 ) ;
  assign n23019 = ~n102 & n23018 ;
  assign n23020 = ( n555 & ~n474 ) | ( n555 & n23019 ) | ( ~n474 & n23019 ) ;
  assign n23021 = ~n555 & n23020 ;
  assign n23022 = ( n23021 & ~n789 ) | ( n23021 & n800 ) | ( ~n789 & n800 ) ;
  assign n23023 = ( n23022 & ~n800 ) | ( n23022 & 1'b0 ) | ( ~n800 & 1'b0 ) ;
  assign n23024 = ( n140 & ~n166 ) | ( n140 & n23023 ) | ( ~n166 & n23023 ) ;
  assign n23025 = ~n140 & n23024 ;
  assign n23007 = n16263 &  n22244 ;
  assign n23008 = ~x5 & n23007 ;
  assign n23009 = ( x5 & ~n23007 ) | ( x5 & 1'b0 ) | ( ~n23007 & 1'b0 ) ;
  assign n23010 = n23008 | n23009 ;
  assign n23026 = ( n22479 & ~n23025 ) | ( n22479 & n23010 ) | ( ~n23025 & n23010 ) ;
  assign n23027 = ( n22479 & ~n23010 ) | ( n22479 & n23025 ) | ( ~n23010 & n23025 ) ;
  assign n23028 = ( n23026 & ~n22479 ) | ( n23026 & n23027 ) | ( ~n22479 & n23027 ) ;
  assign n23029 = ~n3644 & n17115 ;
  assign n23033 = n17107 | n3653 ;
  assign n23030 = ( n3652 & ~n16595 ) | ( n3652 & 1'b0 ) | ( ~n16595 & 1'b0 ) ;
  assign n23031 = ( n3657 & ~n16589 ) | ( n3657 & 1'b0 ) | ( ~n16589 & 1'b0 ) ;
  assign n23032 = n23030 | n23031 ;
  assign n23034 = ( n23033 & ~n3653 ) | ( n23033 & n23032 ) | ( ~n3653 & n23032 ) ;
  assign n23035 = n23029 | n23034 ;
  assign n23037 = ( n22994 & n23028 ) | ( n22994 & n23035 ) | ( n23028 & n23035 ) ;
  assign n23036 = ( n22994 & ~n23028 ) | ( n22994 & n23035 ) | ( ~n23028 & n23035 ) ;
  assign n23038 = ( n23028 & ~n23037 ) | ( n23028 & n23036 ) | ( ~n23037 & n23036 ) ;
  assign n23039 = ( n22996 & n23006 ) | ( n22996 & n23038 ) | ( n23006 & n23038 ) ;
  assign n23040 = ( n23006 & ~n22996 ) | ( n23006 & n23038 ) | ( ~n22996 & n23038 ) ;
  assign n23041 = ( n22996 & ~n23039 ) | ( n22996 & n23040 ) | ( ~n23039 & n23040 ) ;
  assign n22986 = ~n4962 & n18456 ;
  assign n22983 = n4482 | n17791 ;
  assign n22984 = n4495 | n17783 ;
  assign n22985 = n22983 &  n22984 ;
  assign n22987 = ( n4962 & n22986 ) | ( n4962 & n22985 ) | ( n22986 & n22985 ) ;
  assign n22988 = n4478 | n18464 ;
  assign n22989 = n22987 &  n22988 ;
  assign n22990 = x26 &  n22989 ;
  assign n22991 = x26 | n22989 ;
  assign n22992 = ~n22990 & n22991 ;
  assign n23042 = ( n22982 & ~n23041 ) | ( n22982 & n22992 ) | ( ~n23041 & n22992 ) ;
  assign n23043 = ( n22982 & ~n22992 ) | ( n22982 & n23041 ) | ( ~n22992 & n23041 ) ;
  assign n23044 = ( n23042 & ~n22982 ) | ( n23042 & n23043 ) | ( ~n22982 & n23043 ) ;
  assign n23048 = ~n5135 & n19043 ;
  assign n23045 = n5010 | n18589 ;
  assign n23046 = n5067 | n18712 ;
  assign n23047 = n23045 &  n23046 ;
  assign n23049 = ( n5135 & n23048 ) | ( n5135 & n23047 ) | ( n23048 & n23047 ) ;
  assign n23050 = n5012 | n19083 ;
  assign n23051 = n23049 &  n23050 ;
  assign n23052 = x23 &  n23051 ;
  assign n23053 = x23 | n23051 ;
  assign n23054 = ~n23052 & n23053 ;
  assign n23059 = ( n23044 & n23054 ) | ( n23044 & n23058 ) | ( n23054 & n23058 ) ;
  assign n23060 = ( n23044 & ~n23058 ) | ( n23044 & n23054 ) | ( ~n23058 & n23054 ) ;
  assign n23061 = ( n23058 & ~n23059 ) | ( n23058 & n23060 ) | ( ~n23059 & n23060 ) ;
  assign n23062 = n5339 &  n19047 ;
  assign n23063 = ~n5761 & n19040 ;
  assign n23064 = n23062 | n23063 ;
  assign n23065 = ~n5837 & n19494 ;
  assign n23066 = ( n5837 & ~n23064 ) | ( n5837 & n23065 ) | ( ~n23064 & n23065 ) ;
  assign n23067 = n5341 | n19502 ;
  assign n23068 = n23066 &  n23067 ;
  assign n23069 = x20 &  n23068 ;
  assign n23070 = x20 | n23068 ;
  assign n23071 = ~n23069 & n23070 ;
  assign n23076 = ( n23061 & n23071 ) | ( n23061 & n23075 ) | ( n23071 & n23075 ) ;
  assign n23077 = ( n23061 & ~n23075 ) | ( n23061 & n23071 ) | ( ~n23075 & n23071 ) ;
  assign n23078 = ( n23075 & ~n23076 ) | ( n23075 & n23077 ) | ( ~n23076 & n23077 ) ;
  assign n23082 = ~n6395 & n20241 ;
  assign n23079 = n5970 | n19951 ;
  assign n23080 = n6170 | n20027 ;
  assign n23081 = n23079 &  n23080 ;
  assign n23083 = ( n6395 & n23082 ) | ( n6395 & n23081 ) | ( n23082 & n23081 ) ;
  assign n23084 = n5972 | n20280 ;
  assign n23085 = n23083 &  n23084 ;
  assign n23086 = x17 &  n23085 ;
  assign n23087 = x17 | n23085 ;
  assign n23088 = ~n23086 & n23087 ;
  assign n23093 = ( n23078 & n23088 ) | ( n23078 & n23092 ) | ( n23088 & n23092 ) ;
  assign n23094 = ( n23078 & ~n23092 ) | ( n23078 & n23088 ) | ( ~n23092 & n23088 ) ;
  assign n23095 = ( n23092 & ~n23093 ) | ( n23092 & n23094 ) | ( ~n23093 & n23094 ) ;
  assign n23096 = ~n6530 & n20245 ;
  assign n23097 = ~n6983 & n20237 ;
  assign n23098 = n23096 | n23097 ;
  assign n23099 = ~n7097 & n20782 ;
  assign n23100 = ( n7097 & ~n23098 ) | ( n7097 & n23099 ) | ( ~n23098 & n23099 ) ;
  assign n23101 = n6532 | n21227 ;
  assign n23102 = n23100 &  n23101 ;
  assign n23103 = x14 &  n23102 ;
  assign n23104 = x14 | n23102 ;
  assign n23105 = ~n23103 & n23104 ;
  assign n23107 = ( x17 & n22912 ) | ( x17 & n22919 ) | ( n22912 & n22919 ) ;
  assign n23106 = ( n22912 & ~x17 ) | ( n22912 & n22919 ) | ( ~x17 & n22919 ) ;
  assign n23108 = ( x17 & ~n23107 ) | ( x17 & n23106 ) | ( ~n23107 & n23106 ) ;
  assign n23109 = ( n22734 & ~n23108 ) | ( n22734 & n22935 ) | ( ~n23108 & n22935 ) ;
  assign n23110 = ( n23095 & n23105 ) | ( n23095 & n23109 ) | ( n23105 & n23109 ) ;
  assign n23111 = ( n23105 & ~n23095 ) | ( n23105 & n23109 ) | ( ~n23095 & n23109 ) ;
  assign n23112 = ( n23095 & ~n23110 ) | ( n23095 & n23111 ) | ( ~n23110 & n23111 ) ;
  assign n23116 = n7783 | n21475 ;
  assign n23113 = n7253 &  n20777 ;
  assign n23114 = n7518 | n21271 ;
  assign n23115 = ~n23113 & n23114 ;
  assign n23117 = ( n7783 & ~n23116 ) | ( n7783 & n23115 ) | ( ~n23116 & n23115 ) ;
  assign n23118 = n7255 | n21484 ;
  assign n23119 = n23117 &  n23118 ;
  assign n23120 = x11 &  n23119 ;
  assign n23121 = x11 | n23119 ;
  assign n23122 = ~n23120 & n23121 ;
  assign n23127 = ( n23112 & n23122 ) | ( n23112 & n23126 ) | ( n23122 & n23126 ) ;
  assign n23128 = ( n23112 & ~n23126 ) | ( n23112 & n23122 ) | ( ~n23126 & n23122 ) ;
  assign n23129 = ( n23126 & ~n23127 ) | ( n23126 & n23128 ) | ( ~n23127 & n23128 ) ;
  assign n23133 = ~n8764 & n22063 ;
  assign n23130 = ( n8105 & ~n21675 ) | ( n8105 & 1'b0 ) | ( ~n21675 & 1'b0 ) ;
  assign n23131 = n8429 | n21864 ;
  assign n23132 = ~n23130 & n23131 ;
  assign n23134 = ( n8764 & n23133 ) | ( n8764 & n23132 ) | ( n23133 & n23132 ) ;
  assign n23135 = n8107 | n22071 ;
  assign n23136 = n23134 &  n23135 ;
  assign n23137 = x8 &  n23136 ;
  assign n23138 = x8 | n23136 ;
  assign n23139 = ~n23137 & n23138 ;
  assign n23140 = ( n22952 & n23129 ) | ( n22952 & n23139 ) | ( n23129 & n23139 ) ;
  assign n23141 = ( n22952 & ~n23129 ) | ( n22952 & n23139 ) | ( ~n23129 & n23139 ) ;
  assign n23142 = ( n23129 & ~n23140 ) | ( n23129 & n23141 ) | ( ~n23140 & n23141 ) ;
  assign n23143 = ( n22974 & n22978 ) | ( n22974 & n23142 ) | ( n22978 & n23142 ) ;
  assign n23144 = ( n22978 & ~n22974 ) | ( n22978 & n23142 ) | ( ~n22974 & n23142 ) ;
  assign n23145 = ( n22974 & ~n23143 ) | ( n22974 & n23144 ) | ( ~n23143 & n23144 ) ;
  assign n23146 = n22969 | n23145 ;
  assign n23147 = n22969 &  n23145 ;
  assign n23148 = ( n23146 & ~n23147 ) | ( n23146 & 1'b0 ) | ( ~n23147 & 1'b0 ) ;
  assign n23149 = ( n22974 & ~n23142 ) | ( n22974 & n22978 ) | ( ~n23142 & n22978 ) ;
  assign n23150 = ( n23122 & ~n23112 ) | ( n23122 & n23126 ) | ( ~n23112 & n23126 ) ;
  assign n23151 = ( n7253 & ~n21271 ) | ( n7253 & 1'b0 ) | ( ~n21271 & 1'b0 ) ;
  assign n23152 = ~n7518 & n21475 ;
  assign n23153 = n23151 | n23152 ;
  assign n23154 = ~n7783 & n21675 ;
  assign n23155 = ( n7783 & ~n23153 ) | ( n7783 & n23154 ) | ( ~n23153 & n23154 ) ;
  assign n23156 = n7255 | n21684 ;
  assign n23157 = n23155 &  n23156 ;
  assign n23158 = x11 &  n23157 ;
  assign n23159 = x11 | n23157 ;
  assign n23160 = ~n23158 & n23159 ;
  assign n23171 = ( n23088 & ~n23078 ) | ( n23088 & n23092 ) | ( ~n23078 & n23092 ) ;
  assign n23182 = ( n23071 & ~n23061 ) | ( n23071 & n23075 ) | ( ~n23061 & n23075 ) ;
  assign n23193 = ( n23054 & ~n23044 ) | ( n23054 & n23058 ) | ( ~n23044 & n23058 ) ;
  assign n23207 = ~n4962 & n18589 ;
  assign n23204 = n4482 | n17783 ;
  assign n23205 = n4495 | n18456 ;
  assign n23206 = n23204 &  n23205 ;
  assign n23208 = ( n4962 & n23207 ) | ( n4962 & n23206 ) | ( n23207 & n23206 ) ;
  assign n23209 = n4478 | n18597 ;
  assign n23210 = n23208 &  n23209 ;
  assign n23211 = x26 &  n23210 ;
  assign n23212 = x26 | n23210 ;
  assign n23213 = ~n23211 & n23212 ;
  assign n23214 = ( n22996 & ~n23038 ) | ( n22996 & n23006 ) | ( ~n23038 & n23006 ) ;
  assign n23215 = ~n2248 & n6258 ;
  assign n23216 = ( n2149 & ~n2279 ) | ( n2149 & n23215 ) | ( ~n2279 & n23215 ) ;
  assign n23217 = ~n2149 & n23216 ;
  assign n23218 = ( n1703 & ~n6811 ) | ( n1703 & n23217 ) | ( ~n6811 & n23217 ) ;
  assign n23219 = ~n1703 & n23218 ;
  assign n23220 = ( n1876 & ~n1277 ) | ( n1876 & n23219 ) | ( ~n1277 & n23219 ) ;
  assign n23221 = ~n1876 & n23220 ;
  assign n23222 = ( n126 & ~n948 ) | ( n126 & n23221 ) | ( ~n948 & n23221 ) ;
  assign n23223 = ~n126 & n23222 ;
  assign n23224 = ( n273 & ~n231 ) | ( n273 & n23223 ) | ( ~n231 & n23223 ) ;
  assign n23225 = ~n273 & n23224 ;
  assign n23226 = ~n165 & n23225 ;
  assign n23227 = n1429 | n2626 ;
  assign n23228 = ( n6861 & ~n254 ) | ( n6861 & n23227 ) | ( ~n254 & n23227 ) ;
  assign n23229 = n254 | n23228 ;
  assign n23230 = ( n2307 & ~n23226 ) | ( n2307 & n23229 ) | ( ~n23226 & n23229 ) ;
  assign n23231 = ( n2307 & ~n23230 ) | ( n2307 & 1'b0 ) | ( ~n23230 & 1'b0 ) ;
  assign n23232 = ( n1677 & ~n23231 ) | ( n1677 & n3568 ) | ( ~n23231 & n3568 ) ;
  assign n23233 = ( n1677 & ~n23232 ) | ( n1677 & 1'b0 ) | ( ~n23232 & 1'b0 ) ;
  assign n23234 = ( n1427 & ~n1461 ) | ( n1427 & n23233 ) | ( ~n1461 & n23233 ) ;
  assign n23235 = ( n23234 & ~n1427 ) | ( n23234 & n1616 ) | ( ~n1427 & n1616 ) ;
  assign n23236 = ( n23235 & ~n1616 ) | ( n23235 & 1'b0 ) | ( ~n1616 & 1'b0 ) ;
  assign n23237 = ( n425 & ~n352 ) | ( n425 & n23236 ) | ( ~n352 & n23236 ) ;
  assign n23238 = ~n425 & n23237 ;
  assign n23239 = ( n765 & ~n127 ) | ( n765 & n23238 ) | ( ~n127 & n23238 ) ;
  assign n23240 = ~n765 & n23239 ;
  assign n23241 = ( n561 & ~n905 ) | ( n561 & n23240 ) | ( ~n905 & n23240 ) ;
  assign n23242 = ~n561 & n23241 ;
  assign n23243 = ( n43 & ~n666 ) | ( n43 & n23242 ) | ( ~n666 & n23242 ) ;
  assign n23244 = ~n43 & n23243 ;
  assign n23245 = ~n3644 & n17271 ;
  assign n23246 = ( n3652 & ~n16589 ) | ( n3652 & 1'b0 ) | ( ~n16589 & 1'b0 ) ;
  assign n23247 = n3657 &  n17107 ;
  assign n23248 = n23246 | n23247 ;
  assign n23249 = ~n3653 & n17263 ;
  assign n23250 = ( n3653 & ~n23248 ) | ( n3653 & n23249 ) | ( ~n23248 & n23249 ) ;
  assign n23251 = ~n23245 & n23250 ;
  assign n23252 = ( n22479 & n23010 ) | ( n22479 & n23025 ) | ( n23010 & n23025 ) ;
  assign n23253 = ( n23244 & ~n23251 ) | ( n23244 & n23252 ) | ( ~n23251 & n23252 ) ;
  assign n23254 = ( n23244 & ~n23252 ) | ( n23244 & n23251 ) | ( ~n23252 & n23251 ) ;
  assign n23255 = ( n23253 & ~n23244 ) | ( n23253 & n23254 ) | ( ~n23244 & n23254 ) ;
  assign n23261 = ~n601 & n17811 ;
  assign n23259 = ~n4430 & n17791 ;
  assign n23256 = n523 | n17405 ;
  assign n23257 = n3939 | n17787 ;
  assign n23258 = n23256 &  n23257 ;
  assign n23260 = ( n4430 & n23259 ) | ( n4430 & n23258 ) | ( n23259 & n23258 ) ;
  assign n23262 = ( n601 & n23261 ) | ( n601 & n23260 ) | ( n23261 & n23260 ) ;
  assign n23263 = x29 &  n23262 ;
  assign n23264 = x29 | n23262 ;
  assign n23265 = ~n23263 & n23264 ;
  assign n23266 = ( n22994 & ~n23035 ) | ( n22994 & n23028 ) | ( ~n23035 & n23028 ) ;
  assign n23268 = ( n23255 & n23265 ) | ( n23255 & n23266 ) | ( n23265 & n23266 ) ;
  assign n23267 = ( n23265 & ~n23255 ) | ( n23265 & n23266 ) | ( ~n23255 & n23266 ) ;
  assign n23269 = ( n23255 & ~n23268 ) | ( n23255 & n23267 ) | ( ~n23268 & n23267 ) ;
  assign n23270 = n23214 | n23269 ;
  assign n23271 = ~n23214 & n23269 ;
  assign n23272 = ( n23270 & ~n23269 ) | ( n23270 & n23271 ) | ( ~n23269 & n23271 ) ;
  assign n23273 = ( n23213 & ~n23042 ) | ( n23213 & n23272 ) | ( ~n23042 & n23272 ) ;
  assign n23274 = ( n23042 & ~n23213 ) | ( n23042 & n23272 ) | ( ~n23213 & n23272 ) ;
  assign n23275 = ( n23273 & ~n23272 ) | ( n23273 & n23274 ) | ( ~n23272 & n23274 ) ;
  assign n23197 = n19047 | n5135 ;
  assign n23194 = n5010 | n18712 ;
  assign n23195 = n5067 | n19043 ;
  assign n23196 = n23194 &  n23195 ;
  assign n23198 = ( n5135 & ~n23197 ) | ( n5135 & n23196 ) | ( ~n23197 & n23196 ) ;
  assign n23199 = ~n5012 & n19068 ;
  assign n23200 = ( n23198 & ~n23199 ) | ( n23198 & 1'b0 ) | ( ~n23199 & 1'b0 ) ;
  assign n23201 = x23 &  n23200 ;
  assign n23202 = x23 | n23200 ;
  assign n23203 = ~n23201 & n23202 ;
  assign n23276 = ( n23193 & ~n23275 ) | ( n23193 & n23203 ) | ( ~n23275 & n23203 ) ;
  assign n23277 = ( n23193 & ~n23203 ) | ( n23193 & n23275 ) | ( ~n23203 & n23275 ) ;
  assign n23278 = ( n23276 & ~n23193 ) | ( n23276 & n23277 ) | ( ~n23193 & n23277 ) ;
  assign n23186 = ~n5837 & n19951 ;
  assign n23183 = n5339 &  n19040 ;
  assign n23184 = n5761 | n19494 ;
  assign n23185 = ~n23183 & n23184 ;
  assign n23187 = ( n5837 & n23186 ) | ( n5837 & n23185 ) | ( n23186 & n23185 ) ;
  assign n23188 = ~n5341 & n19959 ;
  assign n23189 = ( n23187 & ~n23188 ) | ( n23187 & 1'b0 ) | ( ~n23188 & 1'b0 ) ;
  assign n23190 = x20 &  n23189 ;
  assign n23191 = x20 | n23189 ;
  assign n23192 = ~n23190 & n23191 ;
  assign n23279 = ( n23182 & ~n23278 ) | ( n23182 & n23192 ) | ( ~n23278 & n23192 ) ;
  assign n23280 = ( n23182 & ~n23192 ) | ( n23182 & n23278 ) | ( ~n23192 & n23278 ) ;
  assign n23281 = ( n23279 & ~n23182 ) | ( n23279 & n23280 ) | ( ~n23182 & n23280 ) ;
  assign n23175 = n20245 | n6395 ;
  assign n23172 = n5970 | n20027 ;
  assign n23173 = n6170 | n20241 ;
  assign n23174 = n23172 &  n23173 ;
  assign n23176 = ( n6395 & ~n23175 ) | ( n6395 & n23174 ) | ( ~n23175 & n23174 ) ;
  assign n23177 = ~n5972 & n20265 ;
  assign n23178 = ( n23176 & ~n23177 ) | ( n23176 & 1'b0 ) | ( ~n23177 & 1'b0 ) ;
  assign n23179 = x17 &  n23178 ;
  assign n23180 = x17 | n23178 ;
  assign n23181 = ~n23179 & n23180 ;
  assign n23282 = ( n23171 & ~n23281 ) | ( n23171 & n23181 ) | ( ~n23281 & n23181 ) ;
  assign n23283 = ( n23171 & ~n23181 ) | ( n23171 & n23281 ) | ( ~n23181 & n23281 ) ;
  assign n23284 = ( n23282 & ~n23171 ) | ( n23282 & n23283 ) | ( ~n23171 & n23283 ) ;
  assign n23161 = n7097 &  n20777 ;
  assign n23162 = ~n6530 & n20237 ;
  assign n23163 = n6983 | n20782 ;
  assign n23164 = ~n23162 & n23163 ;
  assign n23165 = ( n23161 & ~n20777 ) | ( n23161 & n23164 ) | ( ~n20777 & n23164 ) ;
  assign n23166 = n6532 | n20790 ;
  assign n23167 = n23165 &  n23166 ;
  assign n23168 = x14 &  n23167 ;
  assign n23169 = x14 | n23167 ;
  assign n23170 = ~n23168 & n23169 ;
  assign n23285 = ( n23111 & ~n23284 ) | ( n23111 & n23170 ) | ( ~n23284 & n23170 ) ;
  assign n23286 = ( n23111 & ~n23170 ) | ( n23111 & n23284 ) | ( ~n23170 & n23284 ) ;
  assign n23287 = ( n23285 & ~n23111 ) | ( n23285 & n23286 ) | ( ~n23111 & n23286 ) ;
  assign n23288 = ( n23150 & n23160 ) | ( n23150 & n23287 ) | ( n23160 & n23287 ) ;
  assign n23289 = ( n23160 & ~n23150 ) | ( n23160 & n23287 ) | ( ~n23150 & n23287 ) ;
  assign n23290 = ( n23150 & ~n23288 ) | ( n23150 & n23289 ) | ( ~n23288 & n23289 ) ;
  assign n23294 = n8764 | n22244 ;
  assign n23291 = ( n8105 & ~n21864 ) | ( n8105 & 1'b0 ) | ( ~n21864 & 1'b0 ) ;
  assign n23292 = n8429 | n22063 ;
  assign n23293 = ~n23291 & n23292 ;
  assign n23295 = ( n8764 & ~n23294 ) | ( n8764 & n23293 ) | ( ~n23294 & n23293 ) ;
  assign n23296 = ~n8107 & n22253 ;
  assign n23297 = ( n23295 & ~n23296 ) | ( n23295 & 1'b0 ) | ( ~n23296 & 1'b0 ) ;
  assign n23298 = x8 &  n23297 ;
  assign n23299 = x8 | n23297 ;
  assign n23300 = ~n23298 & n23299 ;
  assign n23301 = ~n23290 & n23300 ;
  assign n23302 = ( n23290 & ~n23300 ) | ( n23290 & 1'b0 ) | ( ~n23300 & 1'b0 ) ;
  assign n23303 = n23301 | n23302 ;
  assign n23304 = ( n23141 & ~n23149 ) | ( n23141 & n23303 ) | ( ~n23149 & n23303 ) ;
  assign n23305 = ( n23141 & ~n23303 ) | ( n23141 & n23149 ) | ( ~n23303 & n23149 ) ;
  assign n23306 = ( n23304 & ~n23141 ) | ( n23304 & n23305 ) | ( ~n23141 & n23305 ) ;
  assign n23307 = n23147 | n23306 ;
  assign n23308 = ( n23147 & ~n23306 ) | ( n23147 & 1'b0 ) | ( ~n23306 & 1'b0 ) ;
  assign n23309 = ( n23307 & ~n23147 ) | ( n23307 & n23308 ) | ( ~n23147 & n23308 ) ;
  assign n23310 = n23147 &  n23306 ;
  assign n23311 = ( n23213 & ~n23269 ) | ( n23213 & n23214 ) | ( ~n23269 & n23214 ) ;
  assign n23312 = ( n4430 & ~n17783 ) | ( n4430 & 1'b0 ) | ( ~n17783 & 1'b0 ) ;
  assign n23313 = n523 | n17787 ;
  assign n23314 = n3939 | n17791 ;
  assign n23315 = n23313 &  n23314 ;
  assign n23316 = ( n17783 & n23312 ) | ( n17783 & n23315 ) | ( n23312 & n23315 ) ;
  assign n23317 = n601 | n17799 ;
  assign n23318 = n23316 &  n23317 ;
  assign n23319 = x29 &  n23318 ;
  assign n23320 = x29 | n23318 ;
  assign n23321 = ~n23319 & n23320 ;
  assign n23322 = ( n23251 & ~n23244 ) | ( n23251 & n23252 ) | ( ~n23244 & n23252 ) ;
  assign n23335 = n676 | n778 ;
  assign n23336 = ( n101 & ~n714 ) | ( n101 & n23335 ) | ( ~n714 & n23335 ) ;
  assign n23337 = n714 | n23336 ;
  assign n23338 = ( n549 & ~n561 ) | ( n549 & n23337 ) | ( ~n561 & n23337 ) ;
  assign n23339 = n561 | n23338 ;
  assign n23340 = ( n353 & ~n603 ) | ( n353 & n23339 ) | ( ~n603 & n23339 ) ;
  assign n23341 = n603 | n23340 ;
  assign n23342 = n670 | n23341 ;
  assign n23343 = ( n17653 & ~n18857 ) | ( n17653 & 1'b0 ) | ( ~n18857 & 1'b0 ) ;
  assign n23323 = n3244 | n3828 ;
  assign n23324 = ( n3213 & ~n134 ) | ( n3213 & n23323 ) | ( ~n134 & n23323 ) ;
  assign n23325 = ( n134 & ~n1920 ) | ( n134 & n23324 ) | ( ~n1920 & n23324 ) ;
  assign n23326 = n1920 | n23325 ;
  assign n23327 = ( n163 & ~n23326 ) | ( n163 & n3221 ) | ( ~n23326 & n3221 ) ;
  assign n23328 = ~n163 & n23327 ;
  assign n23329 = ( n243 & ~n461 ) | ( n243 & n23328 ) | ( ~n461 & n23328 ) ;
  assign n23330 = ~n243 & n23329 ;
  assign n23331 = ( n644 & n735 ) | ( n644 & n23330 ) | ( n735 & n23330 ) ;
  assign n23332 = ~n735 & n23331 ;
  assign n23333 = ( n205 & ~n23332 ) | ( n205 & n343 ) | ( ~n23332 & n343 ) ;
  assign n23334 = ( n343 & ~n23333 ) | ( n343 & 1'b0 ) | ( ~n23333 & 1'b0 ) ;
  assign n23344 = ( n23342 & ~n23343 ) | ( n23342 & n23334 ) | ( ~n23343 & n23334 ) ;
  assign n23345 = ( n6662 & ~n23344 ) | ( n6662 & n23334 ) | ( ~n23344 & n23334 ) ;
  assign n23346 = ~n6662 & n23345 ;
  assign n23347 = ( n4147 & ~n23346 ) | ( n4147 & n4250 ) | ( ~n23346 & n4250 ) ;
  assign n23348 = ( n4250 & ~n23347 ) | ( n4250 & 1'b0 ) | ( ~n23347 & 1'b0 ) ;
  assign n23349 = ( n23348 & ~n138 ) | ( n23348 & n376 ) | ( ~n138 & n376 ) ;
  assign n23350 = ( n23349 & ~n376 ) | ( n23349 & 1'b0 ) | ( ~n376 & 1'b0 ) ;
  assign n23351 = ( n74 & ~n232 ) | ( n74 & n23350 ) | ( ~n232 & n23350 ) ;
  assign n23352 = ~n74 & n23351 ;
  assign n23353 = ( n89 & ~n405 ) | ( n89 & n23352 ) | ( ~n405 & n23352 ) ;
  assign n23354 = ~n89 & n23353 ;
  assign n23355 = ( n252 & ~n213 ) | ( n252 & n23354 ) | ( ~n213 & n23354 ) ;
  assign n23356 = ~n252 & n23355 ;
  assign n23357 = ( n23322 & ~n23244 ) | ( n23322 & n23356 ) | ( ~n23244 & n23356 ) ;
  assign n23358 = ( n23244 & ~n23356 ) | ( n23244 & n23322 ) | ( ~n23356 & n23322 ) ;
  assign n23359 = ( n23357 & ~n23322 ) | ( n23357 & n23358 ) | ( ~n23322 & n23358 ) ;
  assign n23360 = n3644 | n17413 ;
  assign n23361 = n3652 &  n17107 ;
  assign n23362 = ( n3657 & ~n17263 ) | ( n3657 & 1'b0 ) | ( ~n17263 & 1'b0 ) ;
  assign n23363 = n23361 | n23362 ;
  assign n23364 = ~n3653 & n17405 ;
  assign n23365 = ( n3653 & ~n23363 ) | ( n3653 & n23364 ) | ( ~n23363 & n23364 ) ;
  assign n23366 = n23360 &  n23365 ;
  assign n23367 = ( n23267 & n23359 ) | ( n23267 & n23366 ) | ( n23359 & n23366 ) ;
  assign n23368 = ( n23359 & ~n23267 ) | ( n23359 & n23366 ) | ( ~n23267 & n23366 ) ;
  assign n23369 = ( n23267 & ~n23367 ) | ( n23267 & n23368 ) | ( ~n23367 & n23368 ) ;
  assign n23373 = ~n4962 & n18712 ;
  assign n23370 = n4482 | n18456 ;
  assign n23371 = n4495 | n18589 ;
  assign n23372 = n23370 &  n23371 ;
  assign n23374 = ( n4962 & n23373 ) | ( n4962 & n23372 ) | ( n23373 & n23372 ) ;
  assign n23375 = n4478 | n18720 ;
  assign n23376 = n23374 &  n23375 ;
  assign n23377 = x26 &  n23376 ;
  assign n23378 = x26 | n23376 ;
  assign n23379 = ~n23377 & n23378 ;
  assign n23380 = ( n23321 & ~n23369 ) | ( n23321 & n23379 ) | ( ~n23369 & n23379 ) ;
  assign n23381 = ( n23321 & ~n23379 ) | ( n23321 & n23369 ) | ( ~n23379 & n23369 ) ;
  assign n23382 = ( n23380 & ~n23321 ) | ( n23380 & n23381 ) | ( ~n23321 & n23381 ) ;
  assign n23386 = n19040 | n5135 ;
  assign n23383 = n5010 | n19043 ;
  assign n23384 = ~n5067 & n19047 ;
  assign n23385 = ( n23383 & ~n23384 ) | ( n23383 & 1'b0 ) | ( ~n23384 & 1'b0 ) ;
  assign n23387 = ( n5135 & ~n23386 ) | ( n5135 & n23385 ) | ( ~n23386 & n23385 ) ;
  assign n23388 = n5012 | n19056 ;
  assign n23389 = n23387 &  n23388 ;
  assign n23390 = x23 &  n23389 ;
  assign n23391 = x23 | n23389 ;
  assign n23392 = ~n23390 & n23391 ;
  assign n23393 = ( n23311 & n23382 ) | ( n23311 & n23392 ) | ( n23382 & n23392 ) ;
  assign n23394 = ( n23382 & ~n23311 ) | ( n23382 & n23392 ) | ( ~n23311 & n23392 ) ;
  assign n23395 = ( n23311 & ~n23393 ) | ( n23311 & n23394 ) | ( ~n23393 & n23394 ) ;
  assign n23399 = ~n5837 & n20027 ;
  assign n23396 = ( n5339 & ~n19494 ) | ( n5339 & 1'b0 ) | ( ~n19494 & 1'b0 ) ;
  assign n23397 = n5761 | n19951 ;
  assign n23398 = ~n23396 & n23397 ;
  assign n23400 = ( n5837 & n23399 ) | ( n5837 & n23398 ) | ( n23399 & n23398 ) ;
  assign n23401 = n5341 | n20035 ;
  assign n23402 = n23400 &  n23401 ;
  assign n23403 = x20 &  n23402 ;
  assign n23404 = x20 | n23402 ;
  assign n23405 = ~n23403 & n23404 ;
  assign n23406 = ( n23213 & ~n23214 ) | ( n23213 & n23269 ) | ( ~n23214 & n23269 ) ;
  assign n23407 = ( n23214 & ~n23213 ) | ( n23214 & n23269 ) | ( ~n23213 & n23269 ) ;
  assign n23408 = ( n23406 & ~n23269 ) | ( n23406 & n23407 ) | ( ~n23269 & n23407 ) ;
  assign n23409 = ( n23042 & ~n23408 ) | ( n23042 & n23203 ) | ( ~n23408 & n23203 ) ;
  assign n23411 = ( n23395 & n23405 ) | ( n23395 & n23409 ) | ( n23405 & n23409 ) ;
  assign n23410 = ( n23405 & ~n23395 ) | ( n23405 & n23409 ) | ( ~n23395 & n23409 ) ;
  assign n23412 = ( n23395 & ~n23411 ) | ( n23395 & n23410 ) | ( ~n23411 & n23410 ) ;
  assign n23413 = n6395 &  n20237 ;
  assign n23414 = n5970 | n20241 ;
  assign n23415 = ~n6170 & n20245 ;
  assign n23416 = ( n23414 & ~n23415 ) | ( n23414 & 1'b0 ) | ( ~n23415 & 1'b0 ) ;
  assign n23417 = ( n23413 & ~n20237 ) | ( n23413 & n23416 ) | ( ~n20237 & n23416 ) ;
  assign n23418 = n5972 | n20253 ;
  assign n23419 = n23417 &  n23418 ;
  assign n23420 = x17 &  n23419 ;
  assign n23421 = x17 | n23419 ;
  assign n23422 = ~n23420 & n23421 ;
  assign n23424 = ( x23 & n23200 ) | ( x23 & n23275 ) | ( n23200 & n23275 ) ;
  assign n23423 = ( n23200 & ~x23 ) | ( n23200 & n23275 ) | ( ~x23 & n23275 ) ;
  assign n23425 = ( x23 & ~n23424 ) | ( x23 & n23423 ) | ( ~n23424 & n23423 ) ;
  assign n23426 = ( n23192 & ~n23425 ) | ( n23192 & n23193 ) | ( ~n23425 & n23193 ) ;
  assign n23428 = ( n23412 & n23422 ) | ( n23412 & n23426 ) | ( n23422 & n23426 ) ;
  assign n23427 = ( n23422 & ~n23412 ) | ( n23422 & n23426 ) | ( ~n23412 & n23426 ) ;
  assign n23429 = ( n23412 & ~n23428 ) | ( n23412 & n23427 ) | ( ~n23428 & n23427 ) ;
  assign n23433 = ~n7097 & n21271 ;
  assign n23430 = n6530 | n20782 ;
  assign n23431 = ~n6983 & n20777 ;
  assign n23432 = ( n23430 & ~n23431 ) | ( n23430 & 1'b0 ) | ( ~n23431 & 1'b0 ) ;
  assign n23434 = ( n7097 & n23433 ) | ( n7097 & n23432 ) | ( n23433 & n23432 ) ;
  assign n23435 = n6532 | n21279 ;
  assign n23436 = n23434 &  n23435 ;
  assign n23437 = x14 &  n23436 ;
  assign n23438 = x14 | n23436 ;
  assign n23439 = ~n23437 & n23438 ;
  assign n23441 = ( x20 & n23189 ) | ( x20 & n23278 ) | ( n23189 & n23278 ) ;
  assign n23440 = ( n23189 & ~x20 ) | ( n23189 & n23278 ) | ( ~x20 & n23278 ) ;
  assign n23442 = ( x20 & ~n23441 ) | ( x20 & n23440 ) | ( ~n23441 & n23440 ) ;
  assign n23443 = ( n23181 & ~n23442 ) | ( n23181 & n23182 ) | ( ~n23442 & n23182 ) ;
  assign n23445 = ( n23429 & n23439 ) | ( n23429 & n23443 ) | ( n23439 & n23443 ) ;
  assign n23444 = ( n23439 & ~n23429 ) | ( n23439 & n23443 ) | ( ~n23429 & n23443 ) ;
  assign n23446 = ( n23429 & ~n23445 ) | ( n23429 & n23444 ) | ( ~n23445 & n23444 ) ;
  assign n23450 = ~n7783 & n21864 ;
  assign n23447 = n7253 &  n21475 ;
  assign n23448 = n7518 | n21675 ;
  assign n23449 = ~n23447 & n23448 ;
  assign n23451 = ( n7783 & n23450 ) | ( n7783 & n23449 ) | ( n23450 & n23449 ) ;
  assign n23452 = ~n7255 & n21872 ;
  assign n23453 = ( n23451 & ~n23452 ) | ( n23451 & 1'b0 ) | ( ~n23452 & 1'b0 ) ;
  assign n23454 = x11 &  n23453 ;
  assign n23455 = x11 | n23453 ;
  assign n23456 = ~n23454 & n23455 ;
  assign n23458 = ( x17 & n23178 ) | ( x17 & n23281 ) | ( n23178 & n23281 ) ;
  assign n23457 = ( n23178 & ~x17 ) | ( n23178 & n23281 ) | ( ~x17 & n23281 ) ;
  assign n23459 = ( x17 & ~n23458 ) | ( x17 & n23457 ) | ( ~n23458 & n23457 ) ;
  assign n23460 = ( n23170 & ~n23459 ) | ( n23170 & n23171 ) | ( ~n23459 & n23171 ) ;
  assign n23462 = ( n23446 & n23456 ) | ( n23446 & n23460 ) | ( n23456 & n23460 ) ;
  assign n23461 = ( n23456 & ~n23446 ) | ( n23456 & n23460 ) | ( ~n23446 & n23460 ) ;
  assign n23463 = ( n23446 & ~n23462 ) | ( n23446 & n23461 ) | ( ~n23462 & n23461 ) ;
  assign n23468 = ~n17092 & n22244 ;
  assign n23469 = ( n8105 & ~n22063 ) | ( n8105 & 1'b0 ) | ( ~n22063 & 1'b0 ) ;
  assign n23470 = n23468 | n23469 ;
  assign n23471 = ~n8107 & n22251 ;
  assign n23472 = ( n8107 & ~n23470 ) | ( n8107 & n23471 ) | ( ~n23470 & n23471 ) ;
  assign n23474 = x8 &  n23472 ;
  assign n23473 = ~x8 & n23472 ;
  assign n23475 = ( x8 & ~n23474 ) | ( x8 & n23473 ) | ( ~n23474 & n23473 ) ;
  assign n23465 = ( x14 & n23167 ) | ( x14 & n23284 ) | ( n23167 & n23284 ) ;
  assign n23464 = ( n23167 & ~x14 ) | ( n23167 & n23284 ) | ( ~x14 & n23284 ) ;
  assign n23466 = ( x14 & ~n23465 ) | ( x14 & n23464 ) | ( ~n23465 & n23464 ) ;
  assign n23467 = ( n23111 & ~n23466 ) | ( n23111 & n23160 ) | ( ~n23466 & n23160 ) ;
  assign n23476 = ( n23463 & ~n23475 ) | ( n23463 & n23467 ) | ( ~n23475 & n23467 ) ;
  assign n23477 = ( n23467 & ~n23463 ) | ( n23467 & n23475 ) | ( ~n23463 & n23475 ) ;
  assign n23478 = ( n23476 & ~n23467 ) | ( n23476 & n23477 ) | ( ~n23467 & n23477 ) ;
  assign n23479 = ( x11 & ~n23157 ) | ( x11 & n23287 ) | ( ~n23157 & n23287 ) ;
  assign n23480 = ( x11 & ~n23287 ) | ( x11 & n23157 ) | ( ~n23287 & n23157 ) ;
  assign n23481 = ( n23479 & ~x11 ) | ( n23479 & n23480 ) | ( ~x11 & n23480 ) ;
  assign n23482 = ( n23150 & ~n23481 ) | ( n23150 & n23300 ) | ( ~n23481 & n23300 ) ;
  assign n23483 = ( n23478 & ~n23305 ) | ( n23478 & n23482 ) | ( ~n23305 & n23482 ) ;
  assign n23484 = ( n23305 & ~n23478 ) | ( n23305 & n23482 ) | ( ~n23478 & n23482 ) ;
  assign n23485 = ( n23483 & ~n23482 ) | ( n23483 & n23484 ) | ( ~n23482 & n23484 ) ;
  assign n23486 = n23310 &  n23485 ;
  assign n23487 = n23310 | n23485 ;
  assign n23488 = ~n23486 & n23487 ;
  assign n23492 = ~n5837 & n20241 ;
  assign n23489 = ( n5339 & ~n19951 ) | ( n5339 & 1'b0 ) | ( ~n19951 & 1'b0 ) ;
  assign n23490 = n5761 | n20027 ;
  assign n23491 = ~n23489 & n23490 ;
  assign n23493 = ( n5837 & n23492 ) | ( n5837 & n23491 ) | ( n23492 & n23491 ) ;
  assign n23494 = n5341 | n20280 ;
  assign n23495 = n23493 &  n23494 ;
  assign n23496 = x20 &  n23495 ;
  assign n23497 = x20 | n23495 ;
  assign n23498 = ~n23496 & n23497 ;
  assign n23499 = ~n5010 & n19047 ;
  assign n23500 = ~n5067 & n19040 ;
  assign n23501 = n23499 | n23500 ;
  assign n23502 = ~n5135 & n19494 ;
  assign n23503 = ( n5135 & ~n23501 ) | ( n5135 & n23502 ) | ( ~n23501 & n23502 ) ;
  assign n23504 = n5012 | n19502 ;
  assign n23505 = n23503 &  n23504 ;
  assign n23506 = x23 &  n23505 ;
  assign n23507 = x23 | n23505 ;
  assign n23508 = ~n23506 & n23507 ;
  assign n23512 = ~n4962 & n19043 ;
  assign n23509 = n4482 | n18589 ;
  assign n23510 = n4495 | n18712 ;
  assign n23511 = n23509 &  n23510 ;
  assign n23513 = ( n4962 & n23512 ) | ( n4962 & n23511 ) | ( n23512 & n23511 ) ;
  assign n23514 = n4478 | n19083 ;
  assign n23515 = n23513 &  n23514 ;
  assign n23516 = x26 &  n23515 ;
  assign n23517 = x26 | n23515 ;
  assign n23518 = ~n23516 & n23517 ;
  assign n23522 = ~n4430 & n18456 ;
  assign n23519 = n523 | n17791 ;
  assign n23520 = n3939 | n17783 ;
  assign n23521 = n23519 &  n23520 ;
  assign n23523 = ( n4430 & n23522 ) | ( n4430 & n23521 ) | ( n23522 & n23521 ) ;
  assign n23524 = n601 | n18464 ;
  assign n23525 = n23523 &  n23524 ;
  assign n23526 = x29 &  n23525 ;
  assign n23527 = x29 | n23525 ;
  assign n23528 = ~n23526 & n23527 ;
  assign n23551 = n3644 | n17826 ;
  assign n23552 = ( n3652 & ~n17263 ) | ( n3652 & 1'b0 ) | ( ~n17263 & 1'b0 ) ;
  assign n23553 = ( n3657 & ~n17405 ) | ( n3657 & 1'b0 ) | ( ~n17405 & 1'b0 ) ;
  assign n23554 = n23552 | n23553 ;
  assign n23555 = ~n3653 & n17787 ;
  assign n23556 = ( n3653 & ~n23554 ) | ( n3653 & n23555 ) | ( ~n23554 & n23555 ) ;
  assign n23557 = n23551 &  n23556 ;
  assign n23534 = n1286 | n1949 ;
  assign n23535 = ( n2345 & ~n1063 ) | ( n2345 & n23534 ) | ( ~n1063 & n23534 ) ;
  assign n23536 = n1063 | n23535 ;
  assign n23537 = ( n265 & n23536 ) | ( n265 & n2796 ) | ( n23536 & n2796 ) ;
  assign n23538 = ( n2796 & ~n23537 ) | ( n2796 & 1'b0 ) | ( ~n23537 & 1'b0 ) ;
  assign n23539 = ( n3565 & n2484 ) | ( n3565 & n23538 ) | ( n2484 & n23538 ) ;
  assign n23540 = ~n2484 & n23539 ;
  assign n23541 = ( n1493 & ~n1414 ) | ( n1493 & n23540 ) | ( ~n1414 & n23540 ) ;
  assign n23542 = ~n1493 & n23541 ;
  assign n23543 = ( n575 & ~n3281 ) | ( n575 & n23542 ) | ( ~n3281 & n23542 ) ;
  assign n23544 = ~n575 & n23543 ;
  assign n23545 = ( n1152 & ~n679 ) | ( n1152 & n23544 ) | ( ~n679 & n23544 ) ;
  assign n23546 = ~n1152 & n23545 ;
  assign n23547 = ~n406 & n23546 ;
  assign n23530 = n17184 &  n22472 ;
  assign n23529 = n17184 &  n22241 ;
  assign n23532 = ( x8 & n23529 ) | ( x8 & n23530 ) | ( n23529 & n23530 ) ;
  assign n23531 = ( x8 & ~n23530 ) | ( x8 & n23529 ) | ( ~n23530 & n23529 ) ;
  assign n23533 = ( n23530 & ~n23532 ) | ( n23530 & n23531 ) | ( ~n23532 & n23531 ) ;
  assign n23548 = ( n23244 & ~n23547 ) | ( n23244 & n23533 ) | ( ~n23547 & n23533 ) ;
  assign n23549 = ( n23533 & ~n23244 ) | ( n23533 & n23547 ) | ( ~n23244 & n23547 ) ;
  assign n23550 = ( n23548 & ~n23533 ) | ( n23548 & n23549 ) | ( ~n23533 & n23549 ) ;
  assign n23559 = ( n23357 & n23550 ) | ( n23357 & n23557 ) | ( n23550 & n23557 ) ;
  assign n23558 = ( n23357 & ~n23557 ) | ( n23357 & n23550 ) | ( ~n23557 & n23550 ) ;
  assign n23560 = ( n23557 & ~n23559 ) | ( n23557 & n23558 ) | ( ~n23559 & n23558 ) ;
  assign n23561 = ( n23267 & ~n23359 ) | ( n23267 & n23366 ) | ( ~n23359 & n23366 ) ;
  assign n23562 = ( n23528 & ~n23560 ) | ( n23528 & n23561 ) | ( ~n23560 & n23561 ) ;
  assign n23563 = ( n23528 & ~n23561 ) | ( n23528 & n23560 ) | ( ~n23561 & n23560 ) ;
  assign n23564 = ( n23562 & ~n23528 ) | ( n23562 & n23563 ) | ( ~n23528 & n23563 ) ;
  assign n23565 = ( n23380 & n23518 ) | ( n23380 & n23564 ) | ( n23518 & n23564 ) ;
  assign n23566 = ( n23380 & ~n23518 ) | ( n23380 & n23564 ) | ( ~n23518 & n23564 ) ;
  assign n23567 = ( n23518 & ~n23565 ) | ( n23518 & n23566 ) | ( ~n23565 & n23566 ) ;
  assign n23568 = ( n23311 & ~n23382 ) | ( n23311 & n23392 ) | ( ~n23382 & n23392 ) ;
  assign n23569 = ( n23508 & n23567 ) | ( n23508 & n23568 ) | ( n23567 & n23568 ) ;
  assign n23570 = ( n23567 & ~n23508 ) | ( n23567 & n23568 ) | ( ~n23508 & n23568 ) ;
  assign n23571 = ( n23508 & ~n23569 ) | ( n23508 & n23570 ) | ( ~n23569 & n23570 ) ;
  assign n23572 = ( n23410 & n23498 ) | ( n23410 & n23571 ) | ( n23498 & n23571 ) ;
  assign n23573 = ( n23410 & ~n23498 ) | ( n23410 & n23571 ) | ( ~n23498 & n23571 ) ;
  assign n23574 = ( n23498 & ~n23572 ) | ( n23498 & n23573 ) | ( ~n23572 & n23573 ) ;
  assign n23575 = ~n5970 & n20245 ;
  assign n23576 = ~n6170 & n20237 ;
  assign n23577 = n23575 | n23576 ;
  assign n23578 = ~n6395 & n20782 ;
  assign n23579 = ( n6395 & ~n23577 ) | ( n6395 & n23578 ) | ( ~n23577 & n23578 ) ;
  assign n23580 = n5972 | n21227 ;
  assign n23581 = n23579 &  n23580 ;
  assign n23582 = x17 &  n23581 ;
  assign n23583 = x17 | n23581 ;
  assign n23584 = ~n23582 & n23583 ;
  assign n23586 = ( n23427 & n23574 ) | ( n23427 & n23584 ) | ( n23574 & n23584 ) ;
  assign n23585 = ( n23427 & ~n23574 ) | ( n23427 & n23584 ) | ( ~n23574 & n23584 ) ;
  assign n23587 = ( n23574 & ~n23586 ) | ( n23574 & n23585 ) | ( ~n23586 & n23585 ) ;
  assign n23591 = n21475 | n7097 ;
  assign n23588 = ~n6530 & n20777 ;
  assign n23589 = n6983 | n21271 ;
  assign n23590 = ~n23588 & n23589 ;
  assign n23592 = ( n7097 & ~n23591 ) | ( n7097 & n23590 ) | ( ~n23591 & n23590 ) ;
  assign n23593 = n6532 | n21484 ;
  assign n23594 = n23592 &  n23593 ;
  assign n23595 = x14 &  n23594 ;
  assign n23596 = x14 | n23594 ;
  assign n23597 = ~n23595 & n23596 ;
  assign n23598 = ( n23444 & ~n23587 ) | ( n23444 & n23597 ) | ( ~n23587 & n23597 ) ;
  assign n23599 = ( n23444 & ~n23597 ) | ( n23444 & n23587 ) | ( ~n23597 & n23587 ) ;
  assign n23600 = ( n23598 & ~n23444 ) | ( n23598 & n23599 ) | ( ~n23444 & n23599 ) ;
  assign n23604 = ~n7783 & n22063 ;
  assign n23601 = ( n7253 & ~n21675 ) | ( n7253 & 1'b0 ) | ( ~n21675 & 1'b0 ) ;
  assign n23602 = n7518 | n21864 ;
  assign n23603 = ~n23601 & n23602 ;
  assign n23605 = ( n7783 & n23604 ) | ( n7783 & n23603 ) | ( n23604 & n23603 ) ;
  assign n23606 = n7255 | n22071 ;
  assign n23607 = n23605 &  n23606 ;
  assign n23608 = ( x11 & ~n23607 ) | ( x11 & n23461 ) | ( ~n23607 & n23461 ) ;
  assign n23609 = ( x11 & ~n23461 ) | ( x11 & n23607 ) | ( ~n23461 & n23607 ) ;
  assign n23610 = ( n23608 & ~x11 ) | ( n23608 & n23609 ) | ( ~x11 & n23609 ) ;
  assign n23611 = ( n23600 & ~n23610 ) | ( n23600 & 1'b0 ) | ( ~n23610 & 1'b0 ) ;
  assign n23612 = ~n23600 & n23610 ;
  assign n23613 = n23611 | n23612 ;
  assign n23614 = ( n23477 & ~n23613 ) | ( n23477 & n23484 ) | ( ~n23613 & n23484 ) ;
  assign n23615 = ( n23484 & ~n23477 ) | ( n23484 & n23613 ) | ( ~n23477 & n23613 ) ;
  assign n23616 = ( n23614 & ~n23484 ) | ( n23614 & n23615 ) | ( ~n23484 & n23615 ) ;
  assign n23617 = ~n23486 & n23616 ;
  assign n23618 = ( n23486 & ~n23616 ) | ( n23486 & 1'b0 ) | ( ~n23616 & 1'b0 ) ;
  assign n23619 = n23617 | n23618 ;
  assign n23630 = ( n23444 & n23587 ) | ( n23444 & n23597 ) | ( n23587 & n23597 ) ;
  assign n23623 = ~n7097 & n21675 ;
  assign n23620 = n6530 | n21271 ;
  assign n23621 = ~n6983 & n21475 ;
  assign n23622 = ( n23620 & ~n23621 ) | ( n23620 & 1'b0 ) | ( ~n23621 & 1'b0 ) ;
  assign n23624 = ( n7097 & n23623 ) | ( n7097 & n23622 ) | ( n23623 & n23622 ) ;
  assign n23625 = n6532 | n21684 ;
  assign n23626 = n23624 &  n23625 ;
  assign n23627 = x14 &  n23626 ;
  assign n23628 = x14 | n23626 ;
  assign n23629 = ~n23627 & n23628 ;
  assign n23631 = ( n23244 & n23533 ) | ( n23244 & n23547 ) | ( n23533 & n23547 ) ;
  assign n23632 = n3644 | n17811 ;
  assign n23633 = ( n3652 & ~n17405 ) | ( n3652 & 1'b0 ) | ( ~n17405 & 1'b0 ) ;
  assign n23634 = ( n3657 & ~n17787 ) | ( n3657 & 1'b0 ) | ( ~n17787 & 1'b0 ) ;
  assign n23635 = n23633 | n23634 ;
  assign n23636 = ~n3653 & n17791 ;
  assign n23637 = ( n3653 & ~n23635 ) | ( n3653 & n23636 ) | ( ~n23635 & n23636 ) ;
  assign n23638 = n23632 &  n23637 ;
  assign n23639 = n1064 | n2405 ;
  assign n23640 = ( n389 & n23639 ) | ( n389 & n17595 ) | ( n23639 & n17595 ) ;
  assign n23641 = ( n17595 & ~n23640 ) | ( n17595 & 1'b0 ) | ( ~n23640 & 1'b0 ) ;
  assign n23642 = ( n5216 & ~n3777 ) | ( n5216 & n23641 ) | ( ~n3777 & n23641 ) ;
  assign n23643 = ~n5216 & n23642 ;
  assign n23644 = ( n23643 & ~n171 ) | ( n23643 & n1206 ) | ( ~n171 & n1206 ) ;
  assign n23645 = ( n2620 & ~n23644 ) | ( n2620 & n1206 ) | ( ~n23644 & n1206 ) ;
  assign n23646 = ( n2620 & ~n23645 ) | ( n2620 & 1'b0 ) | ( ~n23645 & 1'b0 ) ;
  assign n23647 = ( n23646 & ~n72 ) | ( n23646 & n796 ) | ( ~n72 & n796 ) ;
  assign n23648 = ( n23647 & ~n796 ) | ( n23647 & 1'b0 ) | ( ~n796 & 1'b0 ) ;
  assign n23649 = ( n255 & ~n905 ) | ( n255 & n23648 ) | ( ~n905 & n23648 ) ;
  assign n23650 = ~n255 & n23649 ;
  assign n23651 = ( n452 & ~n135 ) | ( n452 & n23650 ) | ( ~n135 & n23650 ) ;
  assign n23652 = ~n452 & n23651 ;
  assign n23653 = ~n670 & n23652 ;
  assign n23654 = ( n23631 & ~n23638 ) | ( n23631 & n23653 ) | ( ~n23638 & n23653 ) ;
  assign n23655 = ( n23631 & ~n23653 ) | ( n23631 & n23638 ) | ( ~n23653 & n23638 ) ;
  assign n23656 = ( n23654 & ~n23631 ) | ( n23654 & n23655 ) | ( ~n23631 & n23655 ) ;
  assign n23660 = ~n4430 & n18589 ;
  assign n23657 = n523 | n17783 ;
  assign n23658 = n3939 | n18456 ;
  assign n23659 = n23657 &  n23658 ;
  assign n23661 = ( n4430 & n23660 ) | ( n4430 & n23659 ) | ( n23660 & n23659 ) ;
  assign n23662 = ( n18597 & ~n601 ) | ( n18597 & n23661 ) | ( ~n601 & n23661 ) ;
  assign n23663 = ~n18597 & n23662 ;
  assign n23665 = ( x29 & n23661 ) | ( x29 & n23663 ) | ( n23661 & n23663 ) ;
  assign n23664 = ( x29 & ~n23663 ) | ( x29 & n23661 ) | ( ~n23663 & n23661 ) ;
  assign n23666 = ( n23663 & ~n23665 ) | ( n23663 & n23664 ) | ( ~n23665 & n23664 ) ;
  assign n23667 = ( n23559 & n23656 ) | ( n23559 & n23666 ) | ( n23656 & n23666 ) ;
  assign n23668 = ( n23656 & ~n23559 ) | ( n23656 & n23666 ) | ( ~n23559 & n23666 ) ;
  assign n23669 = ( n23559 & ~n23667 ) | ( n23559 & n23668 ) | ( ~n23667 & n23668 ) ;
  assign n23670 = ( n23528 & n23560 ) | ( n23528 & n23561 ) | ( n23560 & n23561 ) ;
  assign n23674 = n19047 | n4962 ;
  assign n23671 = n4482 | n18712 ;
  assign n23672 = n4495 | n19043 ;
  assign n23673 = n23671 &  n23672 ;
  assign n23675 = ( n4962 & ~n23674 ) | ( n4962 & n23673 ) | ( ~n23674 & n23673 ) ;
  assign n23676 = ~n4478 & n19068 ;
  assign n23677 = ( n23675 & ~n23676 ) | ( n23675 & 1'b0 ) | ( ~n23676 & 1'b0 ) ;
  assign n23678 = x26 &  n23677 ;
  assign n23679 = x26 | n23677 ;
  assign n23680 = ~n23678 & n23679 ;
  assign n23681 = ( n23669 & ~n23670 ) | ( n23669 & n23680 ) | ( ~n23670 & n23680 ) ;
  assign n23682 = ( n23669 & ~n23680 ) | ( n23669 & n23670 ) | ( ~n23680 & n23670 ) ;
  assign n23683 = ( n23681 & ~n23669 ) | ( n23681 & n23682 ) | ( ~n23669 & n23682 ) ;
  assign n23687 = ~n5135 & n19951 ;
  assign n23684 = ~n5010 & n19040 ;
  assign n23685 = n5067 | n19494 ;
  assign n23686 = ~n23684 & n23685 ;
  assign n23688 = ( n5135 & n23687 ) | ( n5135 & n23686 ) | ( n23687 & n23686 ) ;
  assign n23689 = ~n5012 & n19959 ;
  assign n23690 = ( n23688 & ~n23689 ) | ( n23688 & 1'b0 ) | ( ~n23689 & 1'b0 ) ;
  assign n23691 = x23 &  n23690 ;
  assign n23692 = x23 | n23690 ;
  assign n23693 = ~n23691 & n23692 ;
  assign n23694 = ( n23565 & n23683 ) | ( n23565 & n23693 ) | ( n23683 & n23693 ) ;
  assign n23695 = ( n23683 & ~n23565 ) | ( n23683 & n23693 ) | ( ~n23565 & n23693 ) ;
  assign n23696 = ( n23565 & ~n23694 ) | ( n23565 & n23695 ) | ( ~n23694 & n23695 ) ;
  assign n23700 = n20245 | n5837 ;
  assign n23697 = ( n5339 & ~n20027 ) | ( n5339 & 1'b0 ) | ( ~n20027 & 1'b0 ) ;
  assign n23698 = n5761 | n20241 ;
  assign n23699 = ~n23697 & n23698 ;
  assign n23701 = ( n5837 & ~n23700 ) | ( n5837 & n23699 ) | ( ~n23700 & n23699 ) ;
  assign n23702 = ~n5341 & n20265 ;
  assign n23703 = ( n23701 & ~n23702 ) | ( n23701 & 1'b0 ) | ( ~n23702 & 1'b0 ) ;
  assign n23704 = x20 &  n23703 ;
  assign n23705 = x20 | n23703 ;
  assign n23706 = ~n23704 & n23705 ;
  assign n23707 = ( n23569 & n23696 ) | ( n23569 & n23706 ) | ( n23696 & n23706 ) ;
  assign n23708 = ( n23696 & ~n23569 ) | ( n23696 & n23706 ) | ( ~n23569 & n23706 ) ;
  assign n23709 = ( n23569 & ~n23707 ) | ( n23569 & n23708 ) | ( ~n23707 & n23708 ) ;
  assign n23713 = n20777 | n6395 ;
  assign n23710 = ~n5970 & n20237 ;
  assign n23711 = n6170 | n20782 ;
  assign n23712 = ~n23710 & n23711 ;
  assign n23714 = ( n6395 & ~n23713 ) | ( n6395 & n23712 ) | ( ~n23713 & n23712 ) ;
  assign n23715 = n5972 | n20790 ;
  assign n23716 = n23714 &  n23715 ;
  assign n23717 = x17 &  n23716 ;
  assign n23718 = x17 | n23716 ;
  assign n23719 = ~n23717 & n23718 ;
  assign n23720 = ( n23572 & n23709 ) | ( n23572 & n23719 ) | ( n23709 & n23719 ) ;
  assign n23721 = ( n23709 & ~n23572 ) | ( n23709 & n23719 ) | ( ~n23572 & n23719 ) ;
  assign n23722 = ( n23572 & ~n23720 ) | ( n23572 & n23721 ) | ( ~n23720 & n23721 ) ;
  assign n23724 = n23586 &  n23722 ;
  assign n23723 = ~n23586 & n23722 ;
  assign n23725 = ( n23586 & ~n23724 ) | ( n23586 & n23723 ) | ( ~n23724 & n23723 ) ;
  assign n23726 = ( n23630 & ~n23629 ) | ( n23630 & n23725 ) | ( ~n23629 & n23725 ) ;
  assign n23727 = ( n23629 & ~n23630 ) | ( n23629 & n23725 ) | ( ~n23630 & n23725 ) ;
  assign n23728 = ( n23726 & ~n23725 ) | ( n23726 & n23727 ) | ( ~n23725 & n23727 ) ;
  assign n23732 = n7783 | n22244 ;
  assign n23729 = ( n7253 & ~n21864 ) | ( n7253 & 1'b0 ) | ( ~n21864 & 1'b0 ) ;
  assign n23730 = n7518 | n22063 ;
  assign n23731 = ~n23729 & n23730 ;
  assign n23733 = ( n7783 & ~n23732 ) | ( n7783 & n23731 ) | ( ~n23732 & n23731 ) ;
  assign n23734 = ~n7255 & n22253 ;
  assign n23735 = ( n23733 & ~n23734 ) | ( n23733 & 1'b0 ) | ( ~n23734 & 1'b0 ) ;
  assign n23736 = x11 &  n23735 ;
  assign n23737 = x11 | n23735 ;
  assign n23738 = ~n23736 & n23737 ;
  assign n23739 = ~n23728 & n23738 ;
  assign n23740 = ( n23728 & ~n23738 ) | ( n23728 & 1'b0 ) | ( ~n23738 & 1'b0 ) ;
  assign n23741 = n23739 | n23740 ;
  assign n23742 = ( n23477 & n23484 ) | ( n23477 & n23613 ) | ( n23484 & n23613 ) ;
  assign n23743 = x11 &  n23607 ;
  assign n23744 = x11 | n23607 ;
  assign n23745 = ~n23743 & n23744 ;
  assign n23746 = ( n23461 & n23600 ) | ( n23461 & n23745 ) | ( n23600 & n23745 ) ;
  assign n23747 = ( n23741 & ~n23742 ) | ( n23741 & n23746 ) | ( ~n23742 & n23746 ) ;
  assign n23748 = ( n23742 & ~n23741 ) | ( n23742 & n23746 ) | ( ~n23741 & n23746 ) ;
  assign n23749 = ( n23747 & ~n23746 ) | ( n23747 & n23748 ) | ( ~n23746 & n23748 ) ;
  assign n23750 = n23618 | n23749 ;
  assign n23751 = ( n23618 & ~n23749 ) | ( n23618 & 1'b0 ) | ( ~n23749 & 1'b0 ) ;
  assign n23752 = ( n23750 & ~n23618 ) | ( n23750 & n23751 ) | ( ~n23618 & n23751 ) ;
  assign n23753 = ( n23572 & ~n23709 ) | ( n23572 & n23719 ) | ( ~n23709 & n23719 ) ;
  assign n23754 = ( n23569 & ~n23696 ) | ( n23569 & n23706 ) | ( ~n23696 & n23706 ) ;
  assign n23755 = ( n23565 & ~n23683 ) | ( n23565 & n23693 ) | ( ~n23683 & n23693 ) ;
  assign n23756 = ( n23670 & ~n23669 ) | ( n23670 & n23680 ) | ( ~n23669 & n23680 ) ;
  assign n23757 = n3644 | n17799 ;
  assign n23758 = ( n3652 & ~n17787 ) | ( n3652 & 1'b0 ) | ( ~n17787 & 1'b0 ) ;
  assign n23759 = ( n3657 & ~n17791 ) | ( n3657 & 1'b0 ) | ( ~n17791 & 1'b0 ) ;
  assign n23760 = n23758 | n23759 ;
  assign n23761 = ~n3653 & n17783 ;
  assign n23762 = ( n3653 & ~n23760 ) | ( n3653 & n23761 ) | ( ~n23760 & n23761 ) ;
  assign n23763 = n23757 &  n23762 ;
  assign n23764 = ( n3529 & ~n3570 ) | ( n3529 & 1'b0 ) | ( ~n3570 & 1'b0 ) ;
  assign n23765 = ( n1963 & ~n1192 ) | ( n1963 & n23764 ) | ( ~n1192 & n23764 ) ;
  assign n23766 = ~n1963 & n23765 ;
  assign n23767 = ( n1877 & ~n18614 ) | ( n1877 & n23766 ) | ( ~n18614 & n23766 ) ;
  assign n23768 = ~n1877 & n23767 ;
  assign n23769 = ( n5664 & ~n23768 ) | ( n5664 & n14900 ) | ( ~n23768 & n14900 ) ;
  assign n23770 = ( n5664 & ~n23769 ) | ( n5664 & 1'b0 ) | ( ~n23769 & 1'b0 ) ;
  assign n23771 = ( n1093 & ~n1360 ) | ( n1093 & n23770 ) | ( ~n1360 & n23770 ) ;
  assign n23772 = ( n23771 & ~n1093 ) | ( n23771 & 1'b0 ) | ( ~n1093 & 1'b0 ) ;
  assign n23773 = ( n1244 & n23226 ) | ( n1244 & n23772 ) | ( n23226 & n23772 ) ;
  assign n23774 = ~n1244 & n23773 ;
  assign n23775 = ( n1762 & ~n2187 ) | ( n1762 & n23774 ) | ( ~n2187 & n23774 ) ;
  assign n23776 = ~n1762 & n23775 ;
  assign n23777 = ( n734 & ~n792 ) | ( n734 & n23776 ) | ( ~n792 & n23776 ) ;
  assign n23778 = ~n734 & n23777 ;
  assign n23779 = ( n456 & ~n49 ) | ( n456 & n23778 ) | ( ~n49 & n23778 ) ;
  assign n23780 = ~n456 & n23779 ;
  assign n23781 = ~n104 & n23780 ;
  assign n23782 = ( n23653 & ~n23781 ) | ( n23653 & n23655 ) | ( ~n23781 & n23655 ) ;
  assign n23783 = ( n23653 & ~n23655 ) | ( n23653 & n23781 ) | ( ~n23655 & n23781 ) ;
  assign n23784 = ( n23782 & ~n23653 ) | ( n23782 & n23783 ) | ( ~n23653 & n23783 ) ;
  assign n23788 = ~n4430 & n18712 ;
  assign n23785 = n523 | n18456 ;
  assign n23786 = n3939 | n18589 ;
  assign n23787 = n23785 &  n23786 ;
  assign n23789 = ( n4430 & n23788 ) | ( n4430 & n23787 ) | ( n23788 & n23787 ) ;
  assign n23790 = ( n18720 & ~n601 ) | ( n18720 & n23789 ) | ( ~n601 & n23789 ) ;
  assign n23791 = ~n18720 & n23790 ;
  assign n23793 = ( x29 & n23789 ) | ( x29 & n23791 ) | ( n23789 & n23791 ) ;
  assign n23792 = ( x29 & ~n23791 ) | ( x29 & n23789 ) | ( ~n23791 & n23789 ) ;
  assign n23794 = ( n23791 & ~n23793 ) | ( n23791 & n23792 ) | ( ~n23793 & n23792 ) ;
  assign n23795 = ( n23763 & n23784 ) | ( n23763 & n23794 ) | ( n23784 & n23794 ) ;
  assign n23796 = ( n23784 & ~n23763 ) | ( n23784 & n23794 ) | ( ~n23763 & n23794 ) ;
  assign n23797 = ( n23763 & ~n23795 ) | ( n23763 & n23796 ) | ( ~n23795 & n23796 ) ;
  assign n23798 = ( n23559 & ~n23656 ) | ( n23559 & n23666 ) | ( ~n23656 & n23666 ) ;
  assign n23802 = n19040 | n4962 ;
  assign n23799 = n4482 | n19043 ;
  assign n23800 = ~n4495 & n19047 ;
  assign n23801 = ( n23799 & ~n23800 ) | ( n23799 & 1'b0 ) | ( ~n23800 & 1'b0 ) ;
  assign n23803 = ( n4962 & ~n23802 ) | ( n4962 & n23801 ) | ( ~n23802 & n23801 ) ;
  assign n23804 = n4478 | n19056 ;
  assign n23805 = n23803 &  n23804 ;
  assign n23806 = x26 &  n23805 ;
  assign n23807 = x26 | n23805 ;
  assign n23808 = ~n23806 & n23807 ;
  assign n23809 = ( n23797 & ~n23798 ) | ( n23797 & n23808 ) | ( ~n23798 & n23808 ) ;
  assign n23810 = ( n23797 & ~n23808 ) | ( n23797 & n23798 ) | ( ~n23808 & n23798 ) ;
  assign n23811 = ( n23809 & ~n23797 ) | ( n23809 & n23810 ) | ( ~n23797 & n23810 ) ;
  assign n23815 = ~n5135 & n20027 ;
  assign n23812 = n5010 | n19494 ;
  assign n23813 = n5067 | n19951 ;
  assign n23814 = n23812 &  n23813 ;
  assign n23816 = ( n5135 & n23815 ) | ( n5135 & n23814 ) | ( n23815 & n23814 ) ;
  assign n23817 = n5012 | n20035 ;
  assign n23818 = n23816 &  n23817 ;
  assign n23819 = x23 &  n23818 ;
  assign n23820 = x23 | n23818 ;
  assign n23821 = ~n23819 & n23820 ;
  assign n23822 = ( n23756 & n23811 ) | ( n23756 & n23821 ) | ( n23811 & n23821 ) ;
  assign n23823 = ( n23811 & ~n23756 ) | ( n23811 & n23821 ) | ( ~n23756 & n23821 ) ;
  assign n23824 = ( n23756 & ~n23822 ) | ( n23756 & n23823 ) | ( ~n23822 & n23823 ) ;
  assign n23825 = n5837 &  n20237 ;
  assign n23826 = ( n5339 & ~n20241 ) | ( n5339 & 1'b0 ) | ( ~n20241 & 1'b0 ) ;
  assign n23827 = ~n5761 & n20245 ;
  assign n23828 = n23826 | n23827 ;
  assign n23829 = ( n20237 & ~n23825 ) | ( n20237 & n23828 ) | ( ~n23825 & n23828 ) ;
  assign n23830 = n5341 | n20253 ;
  assign n23831 = ~n23829 & n23830 ;
  assign n23832 = x20 &  n23831 ;
  assign n23833 = x20 | n23831 ;
  assign n23834 = ~n23832 & n23833 ;
  assign n23835 = ( n23755 & n23824 ) | ( n23755 & n23834 ) | ( n23824 & n23834 ) ;
  assign n23836 = ( n23824 & ~n23755 ) | ( n23824 & n23834 ) | ( ~n23755 & n23834 ) ;
  assign n23837 = ( n23755 & ~n23835 ) | ( n23755 & n23836 ) | ( ~n23835 & n23836 ) ;
  assign n23841 = ~n6395 & n21271 ;
  assign n23838 = n5970 | n20782 ;
  assign n23839 = ~n6170 & n20777 ;
  assign n23840 = ( n23838 & ~n23839 ) | ( n23838 & 1'b0 ) | ( ~n23839 & 1'b0 ) ;
  assign n23842 = ( n6395 & n23841 ) | ( n6395 & n23840 ) | ( n23841 & n23840 ) ;
  assign n23843 = n5972 | n21279 ;
  assign n23844 = n23842 &  n23843 ;
  assign n23845 = x17 &  n23844 ;
  assign n23846 = x17 | n23844 ;
  assign n23847 = ~n23845 & n23846 ;
  assign n23848 = ( n23754 & n23837 ) | ( n23754 & n23847 ) | ( n23837 & n23847 ) ;
  assign n23849 = ( n23837 & ~n23754 ) | ( n23837 & n23847 ) | ( ~n23754 & n23847 ) ;
  assign n23850 = ( n23754 & ~n23848 ) | ( n23754 & n23849 ) | ( ~n23848 & n23849 ) ;
  assign n23851 = ( n7097 & ~n21864 ) | ( n7097 & 1'b0 ) | ( ~n21864 & 1'b0 ) ;
  assign n23852 = ~n6530 & n21475 ;
  assign n23853 = n6983 | n21675 ;
  assign n23854 = ~n23852 & n23853 ;
  assign n23855 = ( n21864 & n23851 ) | ( n21864 & n23854 ) | ( n23851 & n23854 ) ;
  assign n23856 = ~n6532 & n21872 ;
  assign n23857 = ( n23855 & ~n23856 ) | ( n23855 & 1'b0 ) | ( ~n23856 & 1'b0 ) ;
  assign n23858 = x14 &  n23857 ;
  assign n23859 = x14 | n23857 ;
  assign n23860 = ~n23858 & n23859 ;
  assign n23861 = ( n23753 & n23850 ) | ( n23753 & n23860 ) | ( n23850 & n23860 ) ;
  assign n23862 = ( n23850 & ~n23753 ) | ( n23850 & n23860 ) | ( ~n23753 & n23860 ) ;
  assign n23863 = ( n23753 & ~n23861 ) | ( n23753 & n23862 ) | ( ~n23861 & n23862 ) ;
  assign n23865 = ~n17759 & n22244 ;
  assign n23866 = ( n7253 & ~n22063 ) | ( n7253 & 1'b0 ) | ( ~n22063 & 1'b0 ) ;
  assign n23867 = n23865 | n23866 ;
  assign n23868 = ~n7255 & n22251 ;
  assign n23869 = ( n7255 & ~n23867 ) | ( n7255 & n23868 ) | ( ~n23867 & n23868 ) ;
  assign n23871 = x11 &  n23869 ;
  assign n23870 = ~x11 & n23869 ;
  assign n23872 = ( x11 & ~n23871 ) | ( x11 & n23870 ) | ( ~n23871 & n23870 ) ;
  assign n23864 = ( n23586 & ~n23722 ) | ( n23586 & n23629 ) | ( ~n23722 & n23629 ) ;
  assign n23873 = ( n23863 & ~n23872 ) | ( n23863 & n23864 ) | ( ~n23872 & n23864 ) ;
  assign n23874 = ( n23864 & ~n23863 ) | ( n23864 & n23872 ) | ( ~n23863 & n23872 ) ;
  assign n23875 = ( n23873 & ~n23864 ) | ( n23873 & n23874 ) | ( ~n23864 & n23874 ) ;
  assign n23876 = ( n23586 & n23629 ) | ( n23586 & n23722 ) | ( n23629 & n23722 ) ;
  assign n23877 = ( n23629 & ~n23586 ) | ( n23629 & n23722 ) | ( ~n23586 & n23722 ) ;
  assign n23878 = ( n23586 & ~n23876 ) | ( n23586 & n23877 ) | ( ~n23876 & n23877 ) ;
  assign n23879 = ( n23630 & ~n23878 ) | ( n23630 & n23738 ) | ( ~n23878 & n23738 ) ;
  assign n23880 = ( n23875 & ~n23748 ) | ( n23875 & n23879 ) | ( ~n23748 & n23879 ) ;
  assign n23881 = ( n23748 & ~n23875 ) | ( n23748 & n23879 ) | ( ~n23875 & n23879 ) ;
  assign n23882 = ( n23880 & ~n23879 ) | ( n23880 & n23881 ) | ( ~n23879 & n23881 ) ;
  assign n23883 = n23618 &  n23749 ;
  assign n23884 = n23882 &  n23883 ;
  assign n23885 = n23882 | n23883 ;
  assign n23886 = ~n23884 & n23885 ;
  assign n23887 = ( n23753 & ~n23850 ) | ( n23753 & n23860 ) | ( ~n23850 & n23860 ) ;
  assign n23891 = n21475 | n6395 ;
  assign n23888 = ~n5970 & n20777 ;
  assign n23889 = n6170 | n21271 ;
  assign n23890 = ~n23888 & n23889 ;
  assign n23892 = ( n6395 & ~n23891 ) | ( n6395 & n23890 ) | ( ~n23891 & n23890 ) ;
  assign n23893 = n5972 | n21484 ;
  assign n23894 = n23892 &  n23893 ;
  assign n23895 = x17 &  n23894 ;
  assign n23896 = x17 | n23894 ;
  assign n23897 = ~n23895 & n23896 ;
  assign n23898 = ( n23755 & ~n23824 ) | ( n23755 & n23834 ) | ( ~n23824 & n23834 ) ;
  assign n23902 = ~n5135 & n20241 ;
  assign n23899 = n5010 | n19951 ;
  assign n23900 = n5067 | n20027 ;
  assign n23901 = n23899 &  n23900 ;
  assign n23903 = ( n5135 & n23902 ) | ( n5135 & n23901 ) | ( n23902 & n23901 ) ;
  assign n23904 = n5012 | n20280 ;
  assign n23905 = n23903 &  n23904 ;
  assign n23906 = x23 &  n23905 ;
  assign n23907 = x23 | n23905 ;
  assign n23908 = ~n23906 & n23907 ;
  assign n23909 = ~n4482 & n19047 ;
  assign n23910 = ~n4495 & n19040 ;
  assign n23911 = n23909 | n23910 ;
  assign n23912 = ~n4962 & n19494 ;
  assign n23913 = ( n4962 & ~n23911 ) | ( n4962 & n23912 ) | ( ~n23911 & n23912 ) ;
  assign n23914 = n4478 | n19502 ;
  assign n23915 = n23913 &  n23914 ;
  assign n23916 = x26 &  n23915 ;
  assign n23917 = x26 | n23915 ;
  assign n23918 = ~n23916 & n23917 ;
  assign n23935 = n17590 &  n22244 ;
  assign n23936 = x11 | n23935 ;
  assign n23937 = ( x11 & ~n23935 ) | ( x11 & 1'b0 ) | ( ~n23935 & 1'b0 ) ;
  assign n23938 = ( n23936 & ~x11 ) | ( n23936 & n23937 ) | ( ~x11 & n23937 ) ;
  assign n23919 = ~n1715 & n3013 ;
  assign n23920 = ( n377 & ~n5426 ) | ( n377 & n23919 ) | ( ~n5426 & n23919 ) ;
  assign n23921 = ( n23920 & ~n377 ) | ( n23920 & 1'b0 ) | ( ~n377 & 1'b0 ) ;
  assign n23922 = ( n2331 & ~n23921 ) | ( n2331 & n5397 ) | ( ~n23921 & n5397 ) ;
  assign n23923 = ( n2331 & ~n23922 ) | ( n2331 & 1'b0 ) | ( ~n23922 & 1'b0 ) ;
  assign n23924 = ( n1495 & ~n1340 ) | ( n1495 & n23923 ) | ( ~n1340 & n23923 ) ;
  assign n23925 = ~n1495 & n23924 ;
  assign n23926 = ( n23925 & ~n1278 ) | ( n23925 & n2357 ) | ( ~n1278 & n2357 ) ;
  assign n23927 = ( n23926 & ~n2357 ) | ( n23926 & 1'b0 ) | ( ~n2357 & 1'b0 ) ;
  assign n23928 = ( n2191 & ~n884 ) | ( n2191 & n23927 ) | ( ~n884 & n23927 ) ;
  assign n23929 = ~n2191 & n23928 ;
  assign n23930 = ( n72 & ~n434 ) | ( n72 & n23929 ) | ( ~n434 & n23929 ) ;
  assign n23931 = ~n72 & n23930 ;
  assign n23932 = ( n232 & ~n256 ) | ( n232 & n23931 ) | ( ~n256 & n23931 ) ;
  assign n23933 = ~n232 & n23932 ;
  assign n23934 = ~n83 & n23933 ;
  assign n23939 = ( n23653 & n23934 ) | ( n23653 & n23938 ) | ( n23934 & n23938 ) ;
  assign n23940 = ( n23653 & ~n23938 ) | ( n23653 & n23934 ) | ( ~n23938 & n23934 ) ;
  assign n23941 = ( n23938 & ~n23939 ) | ( n23938 & n23940 ) | ( ~n23939 & n23940 ) ;
  assign n23942 = ( n23655 & ~n23653 ) | ( n23655 & n23781 ) | ( ~n23653 & n23781 ) ;
  assign n23943 = n3644 | n18464 ;
  assign n23944 = ( n3652 & ~n17791 ) | ( n3652 & 1'b0 ) | ( ~n17791 & 1'b0 ) ;
  assign n23945 = ( n3657 & ~n17783 ) | ( n3657 & 1'b0 ) | ( ~n17783 & 1'b0 ) ;
  assign n23946 = n23944 | n23945 ;
  assign n23947 = ~n3653 & n18456 ;
  assign n23948 = ( n3653 & ~n23946 ) | ( n3653 & n23947 ) | ( ~n23946 & n23947 ) ;
  assign n23949 = n23943 &  n23948 ;
  assign n23950 = ( n23941 & ~n23942 ) | ( n23941 & n23949 ) | ( ~n23942 & n23949 ) ;
  assign n23951 = ( n23941 & ~n23949 ) | ( n23941 & n23942 ) | ( ~n23949 & n23942 ) ;
  assign n23952 = ( n23950 & ~n23941 ) | ( n23950 & n23951 ) | ( ~n23941 & n23951 ) ;
  assign n23953 = ( n23763 & ~n23784 ) | ( n23763 & n23794 ) | ( ~n23784 & n23794 ) ;
  assign n23957 = ~n4430 & n19043 ;
  assign n23954 = n523 | n18589 ;
  assign n23955 = n3939 | n18712 ;
  assign n23956 = n23954 &  n23955 ;
  assign n23958 = ( n4430 & n23957 ) | ( n4430 & n23956 ) | ( n23957 & n23956 ) ;
  assign n23959 = n601 | n19083 ;
  assign n23960 = n23958 &  n23959 ;
  assign n23961 = x29 &  n23960 ;
  assign n23962 = x29 | n23960 ;
  assign n23963 = ~n23961 & n23962 ;
  assign n23964 = ( n23952 & ~n23953 ) | ( n23952 & n23963 ) | ( ~n23953 & n23963 ) ;
  assign n23965 = ( n23952 & ~n23963 ) | ( n23952 & n23953 ) | ( ~n23963 & n23953 ) ;
  assign n23966 = ( n23964 & ~n23952 ) | ( n23964 & n23965 ) | ( ~n23952 & n23965 ) ;
  assign n23967 = ( n23798 & ~n23797 ) | ( n23798 & n23808 ) | ( ~n23797 & n23808 ) ;
  assign n23968 = ( n23918 & ~n23966 ) | ( n23918 & n23967 ) | ( ~n23966 & n23967 ) ;
  assign n23969 = ( n23918 & ~n23967 ) | ( n23918 & n23966 ) | ( ~n23967 & n23966 ) ;
  assign n23970 = ( n23968 & ~n23918 ) | ( n23968 & n23969 ) | ( ~n23918 & n23969 ) ;
  assign n23971 = ( n23756 & ~n23811 ) | ( n23756 & n23821 ) | ( ~n23811 & n23821 ) ;
  assign n23972 = ( n23908 & n23970 ) | ( n23908 & n23971 ) | ( n23970 & n23971 ) ;
  assign n23973 = ( n23970 & ~n23908 ) | ( n23970 & n23971 ) | ( ~n23908 & n23971 ) ;
  assign n23974 = ( n23908 & ~n23972 ) | ( n23908 & n23973 ) | ( ~n23972 & n23973 ) ;
  assign n23975 = n5339 &  n20245 ;
  assign n23976 = ~n5761 & n20237 ;
  assign n23977 = n23975 | n23976 ;
  assign n23978 = ~n5837 & n20782 ;
  assign n23979 = ( n5837 & ~n23977 ) | ( n5837 & n23978 ) | ( ~n23977 & n23978 ) ;
  assign n23980 = n5341 | n21227 ;
  assign n23981 = n23979 &  n23980 ;
  assign n23982 = x20 &  n23981 ;
  assign n23983 = x20 | n23981 ;
  assign n23984 = ~n23982 & n23983 ;
  assign n23985 = ( n23898 & n23974 ) | ( n23898 & n23984 ) | ( n23974 & n23984 ) ;
  assign n23986 = ( n23974 & ~n23898 ) | ( n23974 & n23984 ) | ( ~n23898 & n23984 ) ;
  assign n23987 = ( n23898 & ~n23985 ) | ( n23898 & n23986 ) | ( ~n23985 & n23986 ) ;
  assign n23988 = ( n23754 & ~n23837 ) | ( n23754 & n23847 ) | ( ~n23837 & n23847 ) ;
  assign n23989 = ( n23897 & n23987 ) | ( n23897 & n23988 ) | ( n23987 & n23988 ) ;
  assign n23990 = ( n23987 & ~n23897 ) | ( n23987 & n23988 ) | ( ~n23897 & n23988 ) ;
  assign n23991 = ( n23897 & ~n23989 ) | ( n23897 & n23990 ) | ( ~n23989 & n23990 ) ;
  assign n23995 = ~n7097 & n22063 ;
  assign n23992 = n6530 | n21675 ;
  assign n23993 = n6983 | n21864 ;
  assign n23994 = n23992 &  n23993 ;
  assign n23996 = ( n7097 & n23995 ) | ( n7097 & n23994 ) | ( n23995 & n23994 ) ;
  assign n23997 = n6532 | n22071 ;
  assign n23998 = n23996 &  n23997 ;
  assign n23999 = x14 &  n23998 ;
  assign n24000 = x14 | n23998 ;
  assign n24001 = ~n23999 & n24000 ;
  assign n24002 = ( n23887 & n23991 ) | ( n23887 & n24001 ) | ( n23991 & n24001 ) ;
  assign n24003 = ( n23991 & ~n23887 ) | ( n23991 & n24001 ) | ( ~n23887 & n24001 ) ;
  assign n24004 = ( n23887 & ~n24002 ) | ( n23887 & n24003 ) | ( ~n24002 & n24003 ) ;
  assign n24005 = ( n23874 & ~n24004 ) | ( n23874 & n23881 ) | ( ~n24004 & n23881 ) ;
  assign n24006 = ( n23881 & ~n23874 ) | ( n23881 & n24004 ) | ( ~n23874 & n24004 ) ;
  assign n24007 = ( n24005 & ~n23881 ) | ( n24005 & n24006 ) | ( ~n23881 & n24006 ) ;
  assign n24008 = ~n23884 & n24007 ;
  assign n24009 = ( n23884 & ~n24007 ) | ( n23884 & 1'b0 ) | ( ~n24007 & 1'b0 ) ;
  assign n24010 = n24008 | n24009 ;
  assign n24011 = ( n23918 & n23966 ) | ( n23918 & n23967 ) | ( n23966 & n23967 ) ;
  assign n24012 = ( n23941 & n23942 ) | ( n23941 & n23949 ) | ( n23942 & n23949 ) ;
  assign n24013 = n3644 | n18597 ;
  assign n24014 = ( n3652 & ~n17783 ) | ( n3652 & 1'b0 ) | ( ~n17783 & 1'b0 ) ;
  assign n24015 = ( n3657 & ~n18456 ) | ( n3657 & 1'b0 ) | ( ~n18456 & 1'b0 ) ;
  assign n24016 = n24014 | n24015 ;
  assign n24017 = ~n3653 & n18589 ;
  assign n24018 = ( n3653 & ~n24016 ) | ( n3653 & n24017 ) | ( ~n24016 & n24017 ) ;
  assign n24019 = n24013 &  n24018 ;
  assign n24020 = n246 | n2414 ;
  assign n24021 = ( n791 & ~n1810 ) | ( n791 & n24020 ) | ( ~n1810 & n24020 ) ;
  assign n24022 = n1810 | n24021 ;
  assign n24023 = ( n19433 & ~n24022 ) | ( n19433 & n21894 ) | ( ~n24022 & n21894 ) ;
  assign n24024 = ~n19433 & n24023 ;
  assign n24025 = ( n14912 & ~n22273 ) | ( n14912 & n24024 ) | ( ~n22273 & n24024 ) ;
  assign n24026 = ( n22273 & ~n19898 ) | ( n22273 & n24025 ) | ( ~n19898 & n24025 ) ;
  assign n24027 = n19898 &  n24026 ;
  assign n24028 = ( n339 & ~n2309 ) | ( n339 & n24027 ) | ( ~n2309 & n24027 ) ;
  assign n24029 = ~n339 & n24028 ;
  assign n24030 = ( n814 & ~n789 ) | ( n814 & n24029 ) | ( ~n789 & n24029 ) ;
  assign n24031 = ~n814 & n24030 ;
  assign n24032 = ( n271 & ~n793 ) | ( n271 & n24031 ) | ( ~n793 & n24031 ) ;
  assign n24033 = ~n271 & n24032 ;
  assign n24034 = ~n149 & n24033 ;
  assign n24035 = ( n23939 & ~n24019 ) | ( n23939 & n24034 ) | ( ~n24019 & n24034 ) ;
  assign n24036 = ( n23939 & ~n24034 ) | ( n23939 & n24019 ) | ( ~n24034 & n24019 ) ;
  assign n24037 = ( n24035 & ~n23939 ) | ( n24035 & n24036 ) | ( ~n23939 & n24036 ) ;
  assign n24041 = n19047 | n4430 ;
  assign n24038 = n523 | n18712 ;
  assign n24039 = n3939 | n19043 ;
  assign n24040 = n24038 &  n24039 ;
  assign n24042 = ( n4430 & ~n24041 ) | ( n4430 & n24040 ) | ( ~n24041 & n24040 ) ;
  assign n24043 = ( n601 & ~n24042 ) | ( n601 & n19068 ) | ( ~n24042 & n19068 ) ;
  assign n24044 = ( n19068 & ~n24043 ) | ( n19068 & 1'b0 ) | ( ~n24043 & 1'b0 ) ;
  assign n24046 = ( x29 & n24042 ) | ( x29 & n24044 ) | ( n24042 & n24044 ) ;
  assign n24045 = ( x29 & ~n24044 ) | ( x29 & n24042 ) | ( ~n24044 & n24042 ) ;
  assign n24047 = ( n24044 & ~n24046 ) | ( n24044 & n24045 ) | ( ~n24046 & n24045 ) ;
  assign n24048 = ( n24012 & n24037 ) | ( n24012 & n24047 ) | ( n24037 & n24047 ) ;
  assign n24049 = ( n24037 & ~n24012 ) | ( n24037 & n24047 ) | ( ~n24012 & n24047 ) ;
  assign n24050 = ( n24012 & ~n24048 ) | ( n24012 & n24049 ) | ( ~n24048 & n24049 ) ;
  assign n24051 = ( n23952 & n23953 ) | ( n23952 & n23963 ) | ( n23953 & n23963 ) ;
  assign n24055 = ~n4962 & n19951 ;
  assign n24052 = ~n4482 & n19040 ;
  assign n24053 = n4495 | n19494 ;
  assign n24054 = ~n24052 & n24053 ;
  assign n24056 = ( n4962 & n24055 ) | ( n4962 & n24054 ) | ( n24055 & n24054 ) ;
  assign n24057 = ~n4478 & n19959 ;
  assign n24058 = ( n24056 & ~n24057 ) | ( n24056 & 1'b0 ) | ( ~n24057 & 1'b0 ) ;
  assign n24059 = x26 &  n24058 ;
  assign n24060 = x26 | n24058 ;
  assign n24061 = ~n24059 & n24060 ;
  assign n24062 = ( n24050 & ~n24051 ) | ( n24050 & n24061 ) | ( ~n24051 & n24061 ) ;
  assign n24063 = ( n24050 & ~n24061 ) | ( n24050 & n24051 ) | ( ~n24061 & n24051 ) ;
  assign n24064 = ( n24062 & ~n24050 ) | ( n24062 & n24063 ) | ( ~n24050 & n24063 ) ;
  assign n24068 = n20245 | n5135 ;
  assign n24065 = n5010 | n20027 ;
  assign n24066 = n5067 | n20241 ;
  assign n24067 = n24065 &  n24066 ;
  assign n24069 = ( n5135 & ~n24068 ) | ( n5135 & n24067 ) | ( ~n24068 & n24067 ) ;
  assign n24070 = ~n5012 & n20265 ;
  assign n24071 = ( n24069 & ~n24070 ) | ( n24069 & 1'b0 ) | ( ~n24070 & 1'b0 ) ;
  assign n24072 = x23 &  n24071 ;
  assign n24073 = x23 | n24071 ;
  assign n24074 = ~n24072 & n24073 ;
  assign n24075 = ( n24011 & n24064 ) | ( n24011 & n24074 ) | ( n24064 & n24074 ) ;
  assign n24076 = ( n24064 & ~n24011 ) | ( n24064 & n24074 ) | ( ~n24011 & n24074 ) ;
  assign n24077 = ( n24011 & ~n24075 ) | ( n24011 & n24076 ) | ( ~n24075 & n24076 ) ;
  assign n24081 = n5837 | n20777 ;
  assign n24078 = n5339 &  n20237 ;
  assign n24079 = n5761 | n20782 ;
  assign n24080 = ~n24078 & n24079 ;
  assign n24082 = ( n5837 & ~n24081 ) | ( n5837 & n24080 ) | ( ~n24081 & n24080 ) ;
  assign n24083 = n5341 | n20790 ;
  assign n24084 = n24082 &  n24083 ;
  assign n24085 = x20 &  n24084 ;
  assign n24086 = x20 | n24084 ;
  assign n24087 = ~n24085 & n24086 ;
  assign n24088 = ( n23972 & n24077 ) | ( n23972 & n24087 ) | ( n24077 & n24087 ) ;
  assign n24089 = ( n24077 & ~n23972 ) | ( n24077 & n24087 ) | ( ~n23972 & n24087 ) ;
  assign n24090 = ( n23972 & ~n24088 ) | ( n23972 & n24089 ) | ( ~n24088 & n24089 ) ;
  assign n24094 = ~n6395 & n21675 ;
  assign n24091 = n5970 | n21271 ;
  assign n24092 = ~n6170 & n21475 ;
  assign n24093 = ( n24091 & ~n24092 ) | ( n24091 & 1'b0 ) | ( ~n24092 & 1'b0 ) ;
  assign n24095 = ( n6395 & n24094 ) | ( n6395 & n24093 ) | ( n24094 & n24093 ) ;
  assign n24096 = n5972 | n21684 ;
  assign n24097 = n24095 &  n24096 ;
  assign n24098 = x17 &  n24097 ;
  assign n24099 = x17 | n24097 ;
  assign n24100 = ~n24098 & n24099 ;
  assign n24101 = ( n23985 & n24090 ) | ( n23985 & n24100 ) | ( n24090 & n24100 ) ;
  assign n24102 = ( n24090 & ~n23985 ) | ( n24090 & n24100 ) | ( ~n23985 & n24100 ) ;
  assign n24103 = ( n23985 & ~n24101 ) | ( n23985 & n24102 ) | ( ~n24101 & n24102 ) ;
  assign n24107 = n22244 | n7097 ;
  assign n24104 = n6530 | n21864 ;
  assign n24105 = n6983 | n22063 ;
  assign n24106 = n24104 &  n24105 ;
  assign n24108 = ( n7097 & ~n24107 ) | ( n7097 & n24106 ) | ( ~n24107 & n24106 ) ;
  assign n24109 = ~n6532 & n22253 ;
  assign n24110 = ( n24108 & ~n24109 ) | ( n24108 & 1'b0 ) | ( ~n24109 & 1'b0 ) ;
  assign n24111 = x14 &  n24110 ;
  assign n24112 = x14 | n24110 ;
  assign n24113 = ~n24111 & n24112 ;
  assign n24114 = ( n23989 & n24103 ) | ( n23989 & n24113 ) | ( n24103 & n24113 ) ;
  assign n24115 = ( n24103 & ~n23989 ) | ( n24103 & n24113 ) | ( ~n23989 & n24113 ) ;
  assign n24116 = ( n23989 & ~n24114 ) | ( n23989 & n24115 ) | ( ~n24114 & n24115 ) ;
  assign n24117 = n24002 | n24116 ;
  assign n24118 = n24002 &  n24116 ;
  assign n24119 = ( n24117 & ~n24118 ) | ( n24117 & 1'b0 ) | ( ~n24118 & 1'b0 ) ;
  assign n24120 = ( n23874 & n23881 ) | ( n23874 & n24004 ) | ( n23881 & n24004 ) ;
  assign n24121 = ( n24009 & n24119 ) | ( n24009 & n24120 ) | ( n24119 & n24120 ) ;
  assign n24122 = ( n24009 & ~n24119 ) | ( n24009 & n24120 ) | ( ~n24119 & n24120 ) ;
  assign n24123 = ( n24119 & ~n24121 ) | ( n24119 & n24122 ) | ( ~n24121 & n24122 ) ;
  assign n24124 = ( n24119 & ~n23884 ) | ( n24119 & n24120 ) | ( ~n23884 & n24120 ) ;
  assign n24125 = ( n24119 & ~n24007 ) | ( n24119 & n24120 ) | ( ~n24007 & n24120 ) ;
  assign n24126 = ~n24124 & n24125 ;
  assign n24127 = ( n23972 & ~n24077 ) | ( n23972 & n24087 ) | ( ~n24077 & n24087 ) ;
  assign n24128 = ( n24011 & ~n24064 ) | ( n24011 & n24074 ) | ( ~n24064 & n24074 ) ;
  assign n24129 = ( n24051 & ~n24050 ) | ( n24051 & n24061 ) | ( ~n24050 & n24061 ) ;
  assign n24133 = n19040 | n4430 ;
  assign n24130 = n523 | n19043 ;
  assign n24131 = ~n3939 & n19047 ;
  assign n24132 = ( n24130 & ~n24131 ) | ( n24130 & 1'b0 ) | ( ~n24131 & 1'b0 ) ;
  assign n24134 = ( n4430 & ~n24133 ) | ( n4430 & n24132 ) | ( ~n24133 & n24132 ) ;
  assign n24135 = n601 | n19056 ;
  assign n24136 = n24134 &  n24135 ;
  assign n24137 = x29 &  n24136 ;
  assign n24138 = x29 | n24136 ;
  assign n24139 = ~n24137 & n24138 ;
  assign n24140 = n3644 | n18720 ;
  assign n24141 = ( n3652 & ~n18456 ) | ( n3652 & 1'b0 ) | ( ~n18456 & 1'b0 ) ;
  assign n24142 = ( n3657 & ~n18589 ) | ( n3657 & 1'b0 ) | ( ~n18589 & 1'b0 ) ;
  assign n24143 = n24141 | n24142 ;
  assign n24144 = ~n3653 & n18712 ;
  assign n24145 = ( n3653 & ~n24143 ) | ( n3653 & n24144 ) | ( ~n24143 & n24144 ) ;
  assign n24146 = n24140 &  n24145 ;
  assign n24147 = n1732 | n3017 ;
  assign n24148 = n3854 | n24147 ;
  assign n24149 = ( n24148 & ~n3738 ) | ( n24148 & n3784 ) | ( ~n3738 & n3784 ) ;
  assign n24150 = ( n3738 & n24149 ) | ( n3738 & n4304 ) | ( n24149 & n4304 ) ;
  assign n24151 = ( n4304 & ~n24150 ) | ( n4304 & 1'b0 ) | ( ~n24150 & 1'b0 ) ;
  assign n24152 = ( n1104 & n3303 ) | ( n1104 & n24151 ) | ( n3303 & n24151 ) ;
  assign n24153 = ~n3303 & n24152 ;
  assign n24154 = ( n717 & n5576 ) | ( n717 & n24153 ) | ( n5576 & n24153 ) ;
  assign n24155 = ~n717 & n24154 ;
  assign n24156 = ( n125 & ~n793 ) | ( n125 & n24155 ) | ( ~n793 & n24155 ) ;
  assign n24157 = ~n125 & n24156 ;
  assign n24158 = ( n735 & ~n231 ) | ( n735 & n24157 ) | ( ~n231 & n24157 ) ;
  assign n24159 = ~n735 & n24158 ;
  assign n24160 = ( n190 & ~n905 ) | ( n190 & n24159 ) | ( ~n905 & n24159 ) ;
  assign n24161 = ~n190 & n24160 ;
  assign n24162 = ( n664 & ~n77 ) | ( n664 & n24161 ) | ( ~n77 & n24161 ) ;
  assign n24163 = ~n664 & n24162 ;
  assign n24164 = ( n24146 & ~n24034 ) | ( n24146 & n24163 ) | ( ~n24034 & n24163 ) ;
  assign n24165 = ( n24034 & ~n24146 ) | ( n24034 & n24163 ) | ( ~n24146 & n24163 ) ;
  assign n24166 = ( n24164 & ~n24163 ) | ( n24164 & n24165 ) | ( ~n24163 & n24165 ) ;
  assign n24167 = ( n24012 & ~n24037 ) | ( n24012 & n24047 ) | ( ~n24037 & n24047 ) ;
  assign n24168 = ( n24036 & n24166 ) | ( n24036 & n24167 ) | ( n24166 & n24167 ) ;
  assign n24169 = ( n24166 & ~n24036 ) | ( n24166 & n24167 ) | ( ~n24036 & n24167 ) ;
  assign n24170 = ( n24036 & ~n24168 ) | ( n24036 & n24169 ) | ( ~n24168 & n24169 ) ;
  assign n24174 = ~n4962 & n20027 ;
  assign n24171 = n4482 | n19494 ;
  assign n24172 = n4495 | n19951 ;
  assign n24173 = n24171 &  n24172 ;
  assign n24175 = ( n4962 & n24174 ) | ( n4962 & n24173 ) | ( n24174 & n24173 ) ;
  assign n24176 = n4478 | n20035 ;
  assign n24177 = n24175 &  n24176 ;
  assign n24178 = x26 &  n24177 ;
  assign n24179 = x26 | n24177 ;
  assign n24180 = ~n24178 & n24179 ;
  assign n24181 = ( n24139 & ~n24170 ) | ( n24139 & n24180 ) | ( ~n24170 & n24180 ) ;
  assign n24182 = ( n24139 & ~n24180 ) | ( n24139 & n24170 ) | ( ~n24180 & n24170 ) ;
  assign n24183 = ( n24181 & ~n24139 ) | ( n24181 & n24182 ) | ( ~n24139 & n24182 ) ;
  assign n24184 = n5135 &  n20237 ;
  assign n24185 = n5010 | n20241 ;
  assign n24186 = ~n5067 & n20245 ;
  assign n24187 = ( n24185 & ~n24186 ) | ( n24185 & 1'b0 ) | ( ~n24186 & 1'b0 ) ;
  assign n24188 = ( n24184 & ~n20237 ) | ( n24184 & n24187 ) | ( ~n20237 & n24187 ) ;
  assign n24189 = n5012 | n20253 ;
  assign n24190 = n24188 &  n24189 ;
  assign n24191 = x23 &  n24190 ;
  assign n24192 = x23 | n24190 ;
  assign n24193 = ~n24191 & n24192 ;
  assign n24194 = ( n24129 & n24183 ) | ( n24129 & n24193 ) | ( n24183 & n24193 ) ;
  assign n24195 = ( n24183 & ~n24129 ) | ( n24183 & n24193 ) | ( ~n24129 & n24193 ) ;
  assign n24196 = ( n24129 & ~n24194 ) | ( n24129 & n24195 ) | ( ~n24194 & n24195 ) ;
  assign n24197 = ( n5339 & ~n20782 ) | ( n5339 & 1'b0 ) | ( ~n20782 & 1'b0 ) ;
  assign n24198 = ~n5761 & n20777 ;
  assign n24199 = n24197 | n24198 ;
  assign n24200 = ~n5837 & n21271 ;
  assign n24201 = ( n5837 & ~n24199 ) | ( n5837 & n24200 ) | ( ~n24199 & n24200 ) ;
  assign n24202 = n5341 | n21279 ;
  assign n24203 = n24201 &  n24202 ;
  assign n24204 = x20 &  n24203 ;
  assign n24205 = x20 | n24203 ;
  assign n24206 = ~n24204 & n24205 ;
  assign n24207 = ( n24128 & n24196 ) | ( n24128 & n24206 ) | ( n24196 & n24206 ) ;
  assign n24208 = ( n24196 & ~n24128 ) | ( n24196 & n24206 ) | ( ~n24128 & n24206 ) ;
  assign n24209 = ( n24128 & ~n24207 ) | ( n24128 & n24208 ) | ( ~n24207 & n24208 ) ;
  assign n24210 = ( n6395 & ~n21864 ) | ( n6395 & 1'b0 ) | ( ~n21864 & 1'b0 ) ;
  assign n24211 = ~n5970 & n21475 ;
  assign n24212 = n6170 | n21675 ;
  assign n24213 = ~n24211 & n24212 ;
  assign n24214 = ( n21864 & n24210 ) | ( n21864 & n24213 ) | ( n24210 & n24213 ) ;
  assign n24215 = ~n5972 & n21872 ;
  assign n24216 = ( n24214 & ~n24215 ) | ( n24214 & 1'b0 ) | ( ~n24215 & 1'b0 ) ;
  assign n24217 = x17 &  n24216 ;
  assign n24218 = x17 | n24216 ;
  assign n24219 = ~n24217 & n24218 ;
  assign n24220 = ( n24127 & n24209 ) | ( n24127 & n24219 ) | ( n24209 & n24219 ) ;
  assign n24221 = ( n24209 & ~n24127 ) | ( n24209 & n24219 ) | ( ~n24127 & n24219 ) ;
  assign n24222 = ( n24127 & ~n24220 ) | ( n24127 & n24221 ) | ( ~n24220 & n24221 ) ;
  assign n24223 = ( n23985 & ~n24090 ) | ( n23985 & n24100 ) | ( ~n24090 & n24100 ) ;
  assign n24227 = ~n6532 & n22251 ;
  assign n24224 = ~n18327 & n22244 ;
  assign n24225 = n6530 | n22063 ;
  assign n24226 = ~n24224 & n24225 ;
  assign n24228 = ( n6532 & n24227 ) | ( n6532 & n24226 ) | ( n24227 & n24226 ) ;
  assign n24229 = ( x14 & ~n24223 ) | ( x14 & n24228 ) | ( ~n24223 & n24228 ) ;
  assign n24230 = ( x14 & ~n24228 ) | ( x14 & n24223 ) | ( ~n24228 & n24223 ) ;
  assign n24231 = ( n24229 & ~x14 ) | ( n24229 & n24230 ) | ( ~x14 & n24230 ) ;
  assign n24232 = ( n24222 & ~n24231 ) | ( n24222 & 1'b0 ) | ( ~n24231 & 1'b0 ) ;
  assign n24233 = ~n24222 & n24231 ;
  assign n24234 = n24232 | n24233 ;
  assign n24235 = ( n24002 & ~n24116 ) | ( n24002 & n24120 ) | ( ~n24116 & n24120 ) ;
  assign n24236 = ( n23989 & ~n24103 ) | ( n23989 & n24113 ) | ( ~n24103 & n24113 ) ;
  assign n24237 = ( n24234 & ~n24235 ) | ( n24234 & n24236 ) | ( ~n24235 & n24236 ) ;
  assign n24238 = ( n24235 & ~n24234 ) | ( n24235 & n24236 ) | ( ~n24234 & n24236 ) ;
  assign n24239 = ( n24237 & ~n24236 ) | ( n24237 & n24238 ) | ( ~n24236 & n24238 ) ;
  assign n24240 = n24126 &  n24239 ;
  assign n24241 = n24126 | n24239 ;
  assign n24242 = ~n24240 & n24241 ;
  assign n24247 = ( n24127 & ~n24209 ) | ( n24127 & n24219 ) | ( ~n24209 & n24219 ) ;
  assign n24251 = n5837 | n21475 ;
  assign n24248 = n5339 &  n20777 ;
  assign n24249 = n5761 | n21271 ;
  assign n24250 = ~n24248 & n24249 ;
  assign n24252 = ( n5837 & ~n24251 ) | ( n5837 & n24250 ) | ( ~n24251 & n24250 ) ;
  assign n24253 = n5341 | n21484 ;
  assign n24254 = n24252 &  n24253 ;
  assign n24255 = x20 &  n24254 ;
  assign n24256 = x20 | n24254 ;
  assign n24257 = ~n24255 & n24256 ;
  assign n24258 = ( n24129 & ~n24183 ) | ( n24129 & n24193 ) | ( ~n24183 & n24193 ) ;
  assign n24262 = ~n4962 & n20241 ;
  assign n24259 = n4482 | n19951 ;
  assign n24260 = n4495 | n20027 ;
  assign n24261 = n24259 &  n24260 ;
  assign n24263 = ( n4962 & n24262 ) | ( n4962 & n24261 ) | ( n24262 & n24261 ) ;
  assign n24264 = n4478 | n20280 ;
  assign n24265 = n24263 &  n24264 ;
  assign n24266 = x26 &  n24265 ;
  assign n24267 = x26 | n24265 ;
  assign n24268 = ~n24266 & n24267 ;
  assign n24269 = ~n523 & n19047 ;
  assign n24270 = ~n3939 & n19040 ;
  assign n24271 = n24269 | n24270 ;
  assign n24272 = ~n4430 & n19494 ;
  assign n24273 = ( n4430 & ~n24271 ) | ( n4430 & n24272 ) | ( ~n24271 & n24272 ) ;
  assign n24274 = n601 | n19502 ;
  assign n24275 = n24273 &  n24274 ;
  assign n24276 = x29 &  n24275 ;
  assign n24277 = x29 | n24275 ;
  assign n24278 = ~n24276 & n24277 ;
  assign n24298 = n3644 | n19083 ;
  assign n24299 = ( n3652 & ~n18589 ) | ( n3652 & 1'b0 ) | ( ~n18589 & 1'b0 ) ;
  assign n24300 = ( n3657 & ~n18712 ) | ( n3657 & 1'b0 ) | ( ~n18712 & 1'b0 ) ;
  assign n24301 = n24299 | n24300 ;
  assign n24302 = ~n3653 & n19043 ;
  assign n24303 = ( n3653 & ~n24301 ) | ( n3653 & n24302 ) | ( ~n24301 & n24302 ) ;
  assign n24304 = n24298 &  n24303 ;
  assign n24283 = ~n3340 & n4230 ;
  assign n24284 = ( n2764 & ~n11265 ) | ( n2764 & n24283 ) | ( ~n11265 & n24283 ) ;
  assign n24285 = ( n24284 & ~n2764 ) | ( n24284 & 1'b0 ) | ( ~n2764 & 1'b0 ) ;
  assign n24286 = ( n18362 & ~n6818 ) | ( n18362 & n24285 ) | ( ~n6818 & n24285 ) ;
  assign n24287 = n6818 &  n24286 ;
  assign n24288 = ( n2227 & n1948 ) | ( n2227 & n24287 ) | ( n1948 & n24287 ) ;
  assign n24289 = ~n1948 & n24288 ;
  assign n24290 = ( n2091 & ~n1380 ) | ( n2091 & n24289 ) | ( ~n1380 & n24289 ) ;
  assign n24291 = ~n2091 & n24290 ;
  assign n24292 = ( n269 & ~n905 ) | ( n269 & n24291 ) | ( ~n905 & n24291 ) ;
  assign n24293 = ~n269 & n24292 ;
  assign n24294 = ~n281 & n24293 ;
  assign n24279 = n18535 &  n22244 ;
  assign n24280 = ~x14 & n24279 ;
  assign n24281 = ( x14 & ~n24279 ) | ( x14 & 1'b0 ) | ( ~n24279 & 1'b0 ) ;
  assign n24282 = n24280 | n24281 ;
  assign n24295 = ( n24034 & ~n24294 ) | ( n24034 & n24282 ) | ( ~n24294 & n24282 ) ;
  assign n24296 = ( n24282 & ~n24034 ) | ( n24282 & n24294 ) | ( ~n24034 & n24294 ) ;
  assign n24297 = ( n24295 & ~n24282 ) | ( n24295 & n24296 ) | ( ~n24282 & n24296 ) ;
  assign n24306 = ( n24164 & n24297 ) | ( n24164 & n24304 ) | ( n24297 & n24304 ) ;
  assign n24305 = ( n24164 & ~n24304 ) | ( n24164 & n24297 ) | ( ~n24304 & n24297 ) ;
  assign n24307 = ( n24304 & ~n24306 ) | ( n24304 & n24305 ) | ( ~n24306 & n24305 ) ;
  assign n24308 = ( n24036 & ~n24166 ) | ( n24036 & n24167 ) | ( ~n24166 & n24167 ) ;
  assign n24309 = ( n24278 & ~n24307 ) | ( n24278 & n24308 ) | ( ~n24307 & n24308 ) ;
  assign n24310 = ( n24278 & ~n24308 ) | ( n24278 & n24307 ) | ( ~n24308 & n24307 ) ;
  assign n24311 = ( n24309 & ~n24278 ) | ( n24309 & n24310 ) | ( ~n24278 & n24310 ) ;
  assign n24312 = ( n24181 & n24268 ) | ( n24181 & n24311 ) | ( n24268 & n24311 ) ;
  assign n24313 = ( n24181 & ~n24268 ) | ( n24181 & n24311 ) | ( ~n24268 & n24311 ) ;
  assign n24314 = ( n24268 & ~n24312 ) | ( n24268 & n24313 ) | ( ~n24312 & n24313 ) ;
  assign n24315 = ~n5010 & n20245 ;
  assign n24316 = ~n5067 & n20237 ;
  assign n24317 = n24315 | n24316 ;
  assign n24318 = ~n5135 & n20782 ;
  assign n24319 = ( n5135 & ~n24317 ) | ( n5135 & n24318 ) | ( ~n24317 & n24318 ) ;
  assign n24320 = n5012 | n21227 ;
  assign n24321 = n24319 &  n24320 ;
  assign n24322 = x23 &  n24321 ;
  assign n24323 = x23 | n24321 ;
  assign n24324 = ~n24322 & n24323 ;
  assign n24325 = ( n24258 & n24314 ) | ( n24258 & n24324 ) | ( n24314 & n24324 ) ;
  assign n24326 = ( n24314 & ~n24258 ) | ( n24314 & n24324 ) | ( ~n24258 & n24324 ) ;
  assign n24327 = ( n24258 & ~n24325 ) | ( n24258 & n24326 ) | ( ~n24325 & n24326 ) ;
  assign n24328 = ( n24128 & ~n24196 ) | ( n24128 & n24206 ) | ( ~n24196 & n24206 ) ;
  assign n24329 = ( n24257 & n24327 ) | ( n24257 & n24328 ) | ( n24327 & n24328 ) ;
  assign n24330 = ( n24327 & ~n24257 ) | ( n24327 & n24328 ) | ( ~n24257 & n24328 ) ;
  assign n24331 = ( n24257 & ~n24329 ) | ( n24257 & n24330 ) | ( ~n24329 & n24330 ) ;
  assign n24335 = ~n6395 & n22063 ;
  assign n24332 = n5970 | n21675 ;
  assign n24333 = n6170 | n21864 ;
  assign n24334 = n24332 &  n24333 ;
  assign n24336 = ( n6395 & n24335 ) | ( n6395 & n24334 ) | ( n24335 & n24334 ) ;
  assign n24337 = n5972 | n22071 ;
  assign n24338 = n24336 &  n24337 ;
  assign n24339 = x17 &  n24338 ;
  assign n24340 = x17 | n24338 ;
  assign n24341 = ~n24339 & n24340 ;
  assign n24342 = ( n24247 & n24331 ) | ( n24247 & n24341 ) | ( n24331 & n24341 ) ;
  assign n24343 = ( n24331 & ~n24247 ) | ( n24331 & n24341 ) | ( ~n24247 & n24341 ) ;
  assign n24344 = ( n24247 & ~n24342 ) | ( n24247 & n24343 ) | ( ~n24342 & n24343 ) ;
  assign n24243 = x14 | n24228 ;
  assign n24244 = x14 &  n24228 ;
  assign n24245 = ( n24243 & ~n24244 ) | ( n24243 & 1'b0 ) | ( ~n24244 & 1'b0 ) ;
  assign n24246 = ( n24223 & ~n24222 ) | ( n24223 & n24245 ) | ( ~n24222 & n24245 ) ;
  assign n24345 = ( n24238 & ~n24344 ) | ( n24238 & n24246 ) | ( ~n24344 & n24246 ) ;
  assign n24346 = ( n24238 & ~n24246 ) | ( n24238 & n24344 ) | ( ~n24246 & n24344 ) ;
  assign n24347 = ( n24345 & ~n24238 ) | ( n24345 & n24346 ) | ( ~n24238 & n24346 ) ;
  assign n24348 = ~n24240 & n24347 ;
  assign n24349 = ( n24240 & ~n24347 ) | ( n24240 & 1'b0 ) | ( ~n24347 & 1'b0 ) ;
  assign n24350 = n24348 | n24349 ;
  assign n24351 = ( n24034 & n24282 ) | ( n24034 & n24294 ) | ( n24282 & n24294 ) ;
  assign n24352 = ~n3644 & n19068 ;
  assign n24356 = n19047 | n3653 ;
  assign n24353 = ( n3652 & ~n18712 ) | ( n3652 & 1'b0 ) | ( ~n18712 & 1'b0 ) ;
  assign n24354 = ( n3657 & ~n19043 ) | ( n3657 & 1'b0 ) | ( ~n19043 & 1'b0 ) ;
  assign n24355 = n24353 | n24354 ;
  assign n24357 = ( n24356 & ~n3653 ) | ( n24356 & n24355 ) | ( ~n3653 & n24355 ) ;
  assign n24358 = n24352 | n24357 ;
  assign n24359 = ~n1109 & n2298 ;
  assign n24360 = ( n1047 & ~n16414 ) | ( n1047 & n24359 ) | ( ~n16414 & n24359 ) ;
  assign n24361 = ~n1047 & n24360 ;
  assign n24362 = ( n5412 & ~n6082 ) | ( n5412 & n24361 ) | ( ~n6082 & n24361 ) ;
  assign n24363 = ( n24362 & ~n5412 ) | ( n24362 & 1'b0 ) | ( ~n5412 & 1'b0 ) ;
  assign n24364 = ( n1044 & ~n1955 ) | ( n1044 & n24363 ) | ( ~n1955 & n24363 ) ;
  assign n24365 = ( n24364 & ~n1044 ) | ( n24364 & 1'b0 ) | ( ~n1044 & 1'b0 ) ;
  assign n24366 = ( n2128 & ~n570 ) | ( n2128 & n24365 ) | ( ~n570 & n24365 ) ;
  assign n24367 = ~n2128 & n24366 ;
  assign n24368 = ( n604 & n3565 ) | ( n604 & n24367 ) | ( n3565 & n24367 ) ;
  assign n24369 = ~n604 & n24368 ;
  assign n24370 = ( n65 & ~n2687 ) | ( n65 & n24369 ) | ( ~n2687 & n24369 ) ;
  assign n24371 = ~n65 & n24370 ;
  assign n24372 = ( n24371 & ~n276 ) | ( n24371 & n745 ) | ( ~n276 & n745 ) ;
  assign n24373 = ( n24372 & ~n745 ) | ( n24372 & 1'b0 ) | ( ~n745 & 1'b0 ) ;
  assign n24374 = ~n166 & n24373 ;
  assign n24375 = ( n24351 & n24358 ) | ( n24351 & n24374 ) | ( n24358 & n24374 ) ;
  assign n24376 = ( n24358 & ~n24351 ) | ( n24358 & n24374 ) | ( ~n24351 & n24374 ) ;
  assign n24377 = ( n24351 & ~n24375 ) | ( n24351 & n24376 ) | ( ~n24375 & n24376 ) ;
  assign n24381 = ~n4430 & n19951 ;
  assign n24378 = ~n523 & n19040 ;
  assign n24379 = n3939 | n19494 ;
  assign n24380 = ~n24378 & n24379 ;
  assign n24382 = ( n4430 & n24381 ) | ( n4430 & n24380 ) | ( n24381 & n24380 ) ;
  assign n24383 = ( n601 & ~n24382 ) | ( n601 & n19959 ) | ( ~n24382 & n19959 ) ;
  assign n24384 = ( n19959 & ~n24383 ) | ( n19959 & 1'b0 ) | ( ~n24383 & 1'b0 ) ;
  assign n24386 = ( x29 & n24382 ) | ( x29 & n24384 ) | ( n24382 & n24384 ) ;
  assign n24385 = ( x29 & ~n24384 ) | ( x29 & n24382 ) | ( ~n24384 & n24382 ) ;
  assign n24387 = ( n24384 & ~n24386 ) | ( n24384 & n24385 ) | ( ~n24386 & n24385 ) ;
  assign n24388 = ( n24306 & ~n24377 ) | ( n24306 & n24387 ) | ( ~n24377 & n24387 ) ;
  assign n24389 = ( n24306 & ~n24387 ) | ( n24306 & n24377 ) | ( ~n24387 & n24377 ) ;
  assign n24390 = ( n24388 & ~n24306 ) | ( n24388 & n24389 ) | ( ~n24306 & n24389 ) ;
  assign n24395 = n20245 | n4962 ;
  assign n24392 = n4482 | n20027 ;
  assign n24393 = n4495 | n20241 ;
  assign n24394 = n24392 &  n24393 ;
  assign n24396 = ( n4962 & ~n24395 ) | ( n4962 & n24394 ) | ( ~n24395 & n24394 ) ;
  assign n24397 = ~n4478 & n20265 ;
  assign n24398 = ( n24396 & ~n24397 ) | ( n24396 & 1'b0 ) | ( ~n24397 & 1'b0 ) ;
  assign n24399 = x26 &  n24398 ;
  assign n24400 = x26 | n24398 ;
  assign n24401 = ~n24399 & n24400 ;
  assign n24391 = ( n24278 & n24307 ) | ( n24278 & n24308 ) | ( n24307 & n24308 ) ;
  assign n24402 = ( n24390 & ~n24401 ) | ( n24390 & n24391 ) | ( ~n24401 & n24391 ) ;
  assign n24403 = ( n24390 & ~n24391 ) | ( n24390 & n24401 ) | ( ~n24391 & n24401 ) ;
  assign n24404 = ( n24402 & ~n24390 ) | ( n24402 & n24403 ) | ( ~n24390 & n24403 ) ;
  assign n24408 = n20777 | n5135 ;
  assign n24405 = ~n5010 & n20237 ;
  assign n24406 = n5067 | n20782 ;
  assign n24407 = ~n24405 & n24406 ;
  assign n24409 = ( n5135 & ~n24408 ) | ( n5135 & n24407 ) | ( ~n24408 & n24407 ) ;
  assign n24410 = n5012 | n20790 ;
  assign n24411 = n24409 &  n24410 ;
  assign n24412 = x23 &  n24411 ;
  assign n24413 = x23 | n24411 ;
  assign n24414 = ~n24412 & n24413 ;
  assign n24415 = ( n24312 & ~n24404 ) | ( n24312 & n24414 ) | ( ~n24404 & n24414 ) ;
  assign n24416 = ( n24312 & ~n24414 ) | ( n24312 & n24404 ) | ( ~n24414 & n24404 ) ;
  assign n24417 = ( n24415 & ~n24312 ) | ( n24415 & n24416 ) | ( ~n24312 & n24416 ) ;
  assign n24418 = ( n5339 & ~n21271 ) | ( n5339 & 1'b0 ) | ( ~n21271 & 1'b0 ) ;
  assign n24419 = ~n5761 & n21475 ;
  assign n24420 = n24418 | n24419 ;
  assign n24421 = ~n5837 & n21675 ;
  assign n24422 = ( n5837 & ~n24420 ) | ( n5837 & n24421 ) | ( ~n24420 & n24421 ) ;
  assign n24423 = n5341 | n21684 ;
  assign n24424 = n24422 &  n24423 ;
  assign n24425 = x20 &  n24424 ;
  assign n24426 = x20 | n24424 ;
  assign n24427 = ~n24425 & n24426 ;
  assign n24428 = ( n24325 & ~n24417 ) | ( n24325 & n24427 ) | ( ~n24417 & n24427 ) ;
  assign n24429 = ( n24325 & ~n24427 ) | ( n24325 & n24417 ) | ( ~n24427 & n24417 ) ;
  assign n24430 = ( n24428 & ~n24325 ) | ( n24428 & n24429 ) | ( ~n24325 & n24429 ) ;
  assign n24434 = n22244 | n6395 ;
  assign n24431 = n5970 | n21864 ;
  assign n24432 = n6170 | n22063 ;
  assign n24433 = n24431 &  n24432 ;
  assign n24435 = ( n6395 & ~n24434 ) | ( n6395 & n24433 ) | ( ~n24434 & n24433 ) ;
  assign n24436 = ~n5972 & n22253 ;
  assign n24437 = ( n24435 & ~n24436 ) | ( n24435 & 1'b0 ) | ( ~n24436 & 1'b0 ) ;
  assign n24438 = x17 &  n24437 ;
  assign n24439 = x17 | n24437 ;
  assign n24440 = ~n24438 & n24439 ;
  assign n24441 = ( n24329 & ~n24430 ) | ( n24329 & n24440 ) | ( ~n24430 & n24440 ) ;
  assign n24442 = ( n24329 & ~n24440 ) | ( n24329 & n24430 ) | ( ~n24440 & n24430 ) ;
  assign n24443 = ( n24441 & ~n24329 ) | ( n24441 & n24442 ) | ( ~n24329 & n24442 ) ;
  assign n24444 = ~n24342 & n24443 ;
  assign n24445 = ( n24342 & ~n24443 ) | ( n24342 & 1'b0 ) | ( ~n24443 & 1'b0 ) ;
  assign n24446 = n24444 | n24445 ;
  assign n24447 = ( n24238 & n24246 ) | ( n24238 & n24344 ) | ( n24246 & n24344 ) ;
  assign n24449 = ( n24349 & n24446 ) | ( n24349 & n24447 ) | ( n24446 & n24447 ) ;
  assign n24448 = ( n24349 & ~n24446 ) | ( n24349 & n24447 ) | ( ~n24446 & n24447 ) ;
  assign n24450 = ( n24446 & ~n24449 ) | ( n24446 & n24448 ) | ( ~n24449 & n24448 ) ;
  assign n24547 = ( n24329 & n24430 ) | ( n24329 & n24440 ) | ( n24430 & n24440 ) ;
  assign n24534 = ( n24325 & n24417 ) | ( n24325 & n24427 ) | ( n24417 & n24427 ) ;
  assign n24451 = ( n24312 & n24404 ) | ( n24312 & n24414 ) | ( n24404 & n24414 ) ;
  assign n24452 = ( n24390 & n24391 ) | ( n24390 & n24401 ) | ( n24391 & n24401 ) ;
  assign n24453 = n3644 | n19056 ;
  assign n24457 = n19040 | n3653 ;
  assign n24454 = ( n3652 & ~n19043 ) | ( n3652 & 1'b0 ) | ( ~n19043 & 1'b0 ) ;
  assign n24455 = n3657 &  n19047 ;
  assign n24456 = n24454 | n24455 ;
  assign n24458 = ( n24457 & ~n3653 ) | ( n24457 & n24456 ) | ( ~n3653 & n24456 ) ;
  assign n24459 = ( n24453 & ~n24458 ) | ( n24453 & 1'b0 ) | ( ~n24458 & 1'b0 ) ;
  assign n24460 = n72 | n2192 ;
  assign n24461 = n280 | n24460 ;
  assign n24462 = n1550 | n2808 ;
  assign n24463 = ( n24461 & ~n1429 ) | ( n24461 & n24462 ) | ( ~n1429 & n24462 ) ;
  assign n24464 = n1429 | n24463 ;
  assign n24465 = ( n5567 & n3885 ) | ( n5567 & n24464 ) | ( n3885 & n24464 ) ;
  assign n24466 = ( n5567 & ~n24465 ) | ( n5567 & 1'b0 ) | ( ~n24465 & 1'b0 ) ;
  assign n24467 = ( n3287 & ~n2666 ) | ( n3287 & n24466 ) | ( ~n2666 & n24466 ) ;
  assign n24468 = ( n2059 & ~n24467 ) | ( n2059 & n3287 ) | ( ~n24467 & n3287 ) ;
  assign n24469 = ( n2059 & ~n24468 ) | ( n2059 & 1'b0 ) | ( ~n24468 & 1'b0 ) ;
  assign n24470 = ( n2309 & ~n959 ) | ( n2309 & n24469 ) | ( ~n959 & n24469 ) ;
  assign n24471 = ~n2309 & n24470 ;
  assign n24472 = ( n734 & ~n260 ) | ( n734 & n24471 ) | ( ~n260 & n24471 ) ;
  assign n24473 = ~n734 & n24472 ;
  assign n24474 = ( n236 & ~n560 ) | ( n236 & n24473 ) | ( ~n560 & n24473 ) ;
  assign n24475 = ~n236 & n24474 ;
  assign n24476 = ( n24475 & ~n628 ) | ( n24475 & n643 ) | ( ~n628 & n643 ) ;
  assign n24477 = ( n24476 & ~n643 ) | ( n24476 & 1'b0 ) | ( ~n643 & 1'b0 ) ;
  assign n24479 = ( n24374 & n24376 ) | ( n24374 & n24477 ) | ( n24376 & n24477 ) ;
  assign n24478 = ( n24374 & ~n24376 ) | ( n24374 & n24477 ) | ( ~n24376 & n24477 ) ;
  assign n24480 = ( n24376 & ~n24479 ) | ( n24376 & n24478 ) | ( ~n24479 & n24478 ) ;
  assign n24484 = ~n4430 & n20027 ;
  assign n24481 = n523 | n19494 ;
  assign n24482 = n3939 | n19951 ;
  assign n24483 = n24481 &  n24482 ;
  assign n24485 = ( n4430 & n24484 ) | ( n4430 & n24483 ) | ( n24484 & n24483 ) ;
  assign n24486 = ( n20035 & ~n601 ) | ( n20035 & n24485 ) | ( ~n601 & n24485 ) ;
  assign n24487 = ~n20035 & n24486 ;
  assign n24489 = ( x29 & n24485 ) | ( x29 & n24487 ) | ( n24485 & n24487 ) ;
  assign n24488 = ( x29 & ~n24487 ) | ( x29 & n24485 ) | ( ~n24487 & n24485 ) ;
  assign n24490 = ( n24487 & ~n24489 ) | ( n24487 & n24488 ) | ( ~n24489 & n24488 ) ;
  assign n24491 = ( n24459 & ~n24480 ) | ( n24459 & n24490 ) | ( ~n24480 & n24490 ) ;
  assign n24492 = ( n24459 & ~n24490 ) | ( n24459 & n24480 ) | ( ~n24490 & n24480 ) ;
  assign n24493 = ( n24491 & ~n24459 ) | ( n24491 & n24492 ) | ( ~n24459 & n24492 ) ;
  assign n24495 = n4962 &  n20237 ;
  assign n24496 = n4482 | n20241 ;
  assign n24497 = ~n4495 & n20245 ;
  assign n24498 = ( n24496 & ~n24497 ) | ( n24496 & 1'b0 ) | ( ~n24497 & 1'b0 ) ;
  assign n24499 = ( n24495 & ~n20237 ) | ( n24495 & n24498 ) | ( ~n20237 & n24498 ) ;
  assign n24500 = n4478 | n20253 ;
  assign n24501 = n24499 &  n24500 ;
  assign n24502 = x26 &  n24501 ;
  assign n24503 = x26 | n24501 ;
  assign n24504 = ~n24502 & n24503 ;
  assign n24494 = ( n24306 & n24377 ) | ( n24306 & n24387 ) | ( n24377 & n24387 ) ;
  assign n24505 = ( n24493 & ~n24504 ) | ( n24493 & n24494 ) | ( ~n24504 & n24494 ) ;
  assign n24506 = ( n24493 & ~n24494 ) | ( n24493 & n24504 ) | ( ~n24494 & n24504 ) ;
  assign n24507 = ( n24505 & ~n24493 ) | ( n24505 & n24506 ) | ( ~n24493 & n24506 ) ;
  assign n24511 = ~n5135 & n21271 ;
  assign n24508 = n5010 | n20782 ;
  assign n24509 = ~n5067 & n20777 ;
  assign n24510 = ( n24508 & ~n24509 ) | ( n24508 & 1'b0 ) | ( ~n24509 & 1'b0 ) ;
  assign n24512 = ( n5135 & n24511 ) | ( n5135 & n24510 ) | ( n24511 & n24510 ) ;
  assign n24513 = n5012 | n21279 ;
  assign n24514 = n24512 &  n24513 ;
  assign n24515 = x23 &  n24514 ;
  assign n24516 = x23 | n24514 ;
  assign n24517 = ~n24515 & n24516 ;
  assign n24518 = ( n24452 & ~n24507 ) | ( n24452 & n24517 ) | ( ~n24507 & n24517 ) ;
  assign n24519 = ( n24452 & ~n24517 ) | ( n24452 & n24507 ) | ( ~n24517 & n24507 ) ;
  assign n24520 = ( n24518 & ~n24452 ) | ( n24518 & n24519 ) | ( ~n24452 & n24519 ) ;
  assign n24524 = ~n5837 & n21864 ;
  assign n24521 = n5339 &  n21475 ;
  assign n24522 = n5761 | n21675 ;
  assign n24523 = ~n24521 & n24522 ;
  assign n24525 = ( n5837 & n24524 ) | ( n5837 & n24523 ) | ( n24524 & n24523 ) ;
  assign n24526 = ~n5341 & n21872 ;
  assign n24527 = ( n24525 & ~n24526 ) | ( n24525 & 1'b0 ) | ( ~n24526 & 1'b0 ) ;
  assign n24528 = x20 &  n24527 ;
  assign n24529 = x20 | n24527 ;
  assign n24530 = ~n24528 & n24529 ;
  assign n24531 = ( n24451 & ~n24520 ) | ( n24451 & n24530 ) | ( ~n24520 & n24530 ) ;
  assign n24532 = ( n24451 & ~n24530 ) | ( n24451 & n24520 ) | ( ~n24530 & n24520 ) ;
  assign n24533 = ( n24531 & ~n24451 ) | ( n24531 & n24532 ) | ( ~n24451 & n24532 ) ;
  assign n24535 = ( n5972 & ~n22251 ) | ( n5972 & 1'b0 ) | ( ~n22251 & 1'b0 ) ;
  assign n24536 = ~n19016 & n22244 ;
  assign n24537 = n5970 | n22063 ;
  assign n24538 = ~n24536 & n24537 ;
  assign n24539 = ( n22251 & n24535 ) | ( n22251 & n24538 ) | ( n24535 & n24538 ) ;
  assign n24541 = x17 &  n24539 ;
  assign n24540 = ~x17 & n24539 ;
  assign n24542 = ( x17 & ~n24541 ) | ( x17 & n24540 ) | ( ~n24541 & n24540 ) ;
  assign n24543 = ( n24533 & n24534 ) | ( n24533 & n24542 ) | ( n24534 & n24542 ) ;
  assign n24544 = ( n24533 & ~n24534 ) | ( n24533 & n24542 ) | ( ~n24534 & n24542 ) ;
  assign n24545 = ( n24534 & ~n24543 ) | ( n24534 & n24544 ) | ( ~n24543 & n24544 ) ;
  assign n24546 = ( n24342 & n24443 ) | ( n24342 & n24447 ) | ( n24443 & n24447 ) ;
  assign n24549 = ( n24545 & n24546 ) | ( n24545 & n24547 ) | ( n24546 & n24547 ) ;
  assign n24548 = ( n24545 & ~n24547 ) | ( n24545 & n24546 ) | ( ~n24547 & n24546 ) ;
  assign n24550 = ( n24547 & ~n24549 ) | ( n24547 & n24548 ) | ( ~n24549 & n24548 ) ;
  assign n24551 = ( n24240 & ~n24447 ) | ( n24240 & n24446 ) | ( ~n24447 & n24446 ) ;
  assign n24552 = ( n24347 & ~n24447 ) | ( n24347 & n24446 ) | ( ~n24447 & n24446 ) ;
  assign n24553 = ( n24551 & ~n24552 ) | ( n24551 & 1'b0 ) | ( ~n24552 & 1'b0 ) ;
  assign n24554 = ~n24550 & n24553 ;
  assign n24555 = ( n24550 & ~n24553 ) | ( n24550 & 1'b0 ) | ( ~n24553 & 1'b0 ) ;
  assign n24556 = n24554 | n24555 ;
  assign n24630 = ( n24451 & n24520 ) | ( n24451 & n24530 ) | ( n24520 & n24530 ) ;
  assign n24557 = ~n4482 & n20245 ;
  assign n24558 = ~n4495 & n20237 ;
  assign n24559 = n24557 | n24558 ;
  assign n24560 = ~n4962 & n20782 ;
  assign n24561 = ( n4962 & ~n24559 ) | ( n4962 & n24560 ) | ( ~n24559 & n24560 ) ;
  assign n24562 = n4478 | n21227 ;
  assign n24563 = n24561 &  n24562 ;
  assign n24564 = x26 &  n24563 ;
  assign n24565 = x26 | n24563 ;
  assign n24566 = ~n24564 & n24565 ;
  assign n24567 = ( n24493 & n24494 ) | ( n24493 & n24504 ) | ( n24494 & n24504 ) ;
  assign n24588 = ( n24376 & ~n24374 ) | ( n24376 & n24477 ) | ( ~n24374 & n24477 ) ;
  assign n24572 = n2094 | n14031 ;
  assign n24573 = ( n3584 & ~n24572 ) | ( n3584 & n5210 ) | ( ~n24572 & n5210 ) ;
  assign n24574 = ~n3584 & n24573 ;
  assign n24575 = ( n4559 & ~n24574 ) | ( n4559 & n18923 ) | ( ~n24574 & n18923 ) ;
  assign n24576 = ( n4559 & ~n24575 ) | ( n4559 & 1'b0 ) | ( ~n24575 & 1'b0 ) ;
  assign n24577 = ( n1594 & ~n1882 ) | ( n1594 & n24576 ) | ( ~n1882 & n24576 ) ;
  assign n24578 = ( n24577 & ~n1594 ) | ( n24577 & 1'b0 ) | ( ~n1594 & 1'b0 ) ;
  assign n24579 = ( n126 & ~n357 ) | ( n126 & n24578 ) | ( ~n357 & n24578 ) ;
  assign n24580 = ~n126 & n24579 ;
  assign n24581 = ( n24580 & ~n359 ) | ( n24580 & n714 ) | ( ~n359 & n714 ) ;
  assign n24582 = ( n24581 & ~n714 ) | ( n24581 & 1'b0 ) | ( ~n714 & 1'b0 ) ;
  assign n24583 = ( n628 & ~n358 ) | ( n628 & n24582 ) | ( ~n358 & n24582 ) ;
  assign n24584 = ~n628 & n24583 ;
  assign n24568 = n18852 &  n22244 ;
  assign n24569 = ~x17 & n24568 ;
  assign n24570 = ( x17 & ~n24568 ) | ( x17 & 1'b0 ) | ( ~n24568 & 1'b0 ) ;
  assign n24571 = n24569 | n24570 ;
  assign n24585 = ( n24477 & ~n24584 ) | ( n24477 & n24571 ) | ( ~n24584 & n24571 ) ;
  assign n24586 = ( n24571 & ~n24477 ) | ( n24571 & n24584 ) | ( ~n24477 & n24584 ) ;
  assign n24587 = ( n24585 & ~n24571 ) | ( n24585 & n24586 ) | ( ~n24571 & n24586 ) ;
  assign n24589 = n3644 | n19502 ;
  assign n24590 = n3652 &  n19047 ;
  assign n24591 = n3657 &  n19040 ;
  assign n24592 = n24590 | n24591 ;
  assign n24593 = ~n3653 & n19494 ;
  assign n24594 = ( n3653 & ~n24592 ) | ( n3653 & n24593 ) | ( ~n24592 & n24593 ) ;
  assign n24595 = n24589 &  n24594 ;
  assign n24596 = ( n24588 & ~n24587 ) | ( n24588 & n24595 ) | ( ~n24587 & n24595 ) ;
  assign n24597 = ( n24587 & ~n24588 ) | ( n24587 & n24595 ) | ( ~n24588 & n24595 ) ;
  assign n24598 = ( n24596 & ~n24595 ) | ( n24596 & n24597 ) | ( ~n24595 & n24597 ) ;
  assign n24603 = ~n4430 & n20241 ;
  assign n24600 = n523 | n19951 ;
  assign n24601 = n3939 | n20027 ;
  assign n24602 = n24600 &  n24601 ;
  assign n24604 = ( n4430 & n24603 ) | ( n4430 & n24602 ) | ( n24603 & n24602 ) ;
  assign n24605 = n601 | n20280 ;
  assign n24606 = n24604 &  n24605 ;
  assign n24607 = x29 &  n24606 ;
  assign n24608 = x29 | n24606 ;
  assign n24609 = ~n24607 & n24608 ;
  assign n24599 = ( n24459 & n24480 ) | ( n24459 & n24490 ) | ( n24480 & n24490 ) ;
  assign n24610 = ( n24598 & ~n24609 ) | ( n24598 & n24599 ) | ( ~n24609 & n24599 ) ;
  assign n24611 = ( n24598 & ~n24599 ) | ( n24598 & n24609 ) | ( ~n24599 & n24609 ) ;
  assign n24612 = ( n24610 & ~n24598 ) | ( n24610 & n24611 ) | ( ~n24598 & n24611 ) ;
  assign n24614 = ( n24566 & n24567 ) | ( n24566 & n24612 ) | ( n24567 & n24612 ) ;
  assign n24613 = ( n24567 & ~n24566 ) | ( n24567 & n24612 ) | ( ~n24566 & n24612 ) ;
  assign n24615 = ( n24566 & ~n24614 ) | ( n24566 & n24613 ) | ( ~n24614 & n24613 ) ;
  assign n24620 = n21475 | n5135 ;
  assign n24617 = ~n5010 & n20777 ;
  assign n24618 = n5067 | n21271 ;
  assign n24619 = ~n24617 & n24618 ;
  assign n24621 = ( n5135 & ~n24620 ) | ( n5135 & n24619 ) | ( ~n24620 & n24619 ) ;
  assign n24622 = n5012 | n21484 ;
  assign n24623 = n24621 &  n24622 ;
  assign n24624 = x23 &  n24623 ;
  assign n24625 = x23 | n24623 ;
  assign n24626 = ~n24624 & n24625 ;
  assign n24616 = ( n24452 & n24507 ) | ( n24452 & n24517 ) | ( n24507 & n24517 ) ;
  assign n24627 = ( n24615 & ~n24626 ) | ( n24615 & n24616 ) | ( ~n24626 & n24616 ) ;
  assign n24628 = ( n24615 & ~n24616 ) | ( n24615 & n24626 ) | ( ~n24616 & n24626 ) ;
  assign n24629 = ( n24627 & ~n24615 ) | ( n24627 & n24628 ) | ( ~n24615 & n24628 ) ;
  assign n24634 = ~n5837 & n22063 ;
  assign n24631 = ( n5339 & ~n21675 ) | ( n5339 & 1'b0 ) | ( ~n21675 & 1'b0 ) ;
  assign n24632 = n5761 | n21864 ;
  assign n24633 = ~n24631 & n24632 ;
  assign n24635 = ( n5837 & n24634 ) | ( n5837 & n24633 ) | ( n24634 & n24633 ) ;
  assign n24636 = n5341 | n22071 ;
  assign n24637 = n24635 &  n24636 ;
  assign n24638 = x20 &  n24637 ;
  assign n24639 = x20 | n24637 ;
  assign n24640 = ~n24638 & n24639 ;
  assign n24642 = ( n24629 & n24630 ) | ( n24629 & n24640 ) | ( n24630 & n24640 ) ;
  assign n24641 = ( n24629 & ~n24630 ) | ( n24629 & n24640 ) | ( ~n24630 & n24640 ) ;
  assign n24643 = ( n24630 & ~n24642 ) | ( n24630 & n24641 ) | ( ~n24642 & n24641 ) ;
  assign n24644 = ( n24543 & n24549 ) | ( n24543 & n24643 ) | ( n24549 & n24643 ) ;
  assign n24645 = ( n24543 & ~n24549 ) | ( n24543 & n24643 ) | ( ~n24549 & n24643 ) ;
  assign n24646 = ( n24549 & ~n24644 ) | ( n24549 & n24645 ) | ( ~n24644 & n24645 ) ;
  assign n24647 = n24554 | n24646 ;
  assign n24648 = n24554 &  n24646 ;
  assign n24649 = ( n24647 & ~n24648 ) | ( n24647 & 1'b0 ) | ( ~n24648 & 1'b0 ) ;
  assign n24650 = ( n24616 & ~n24615 ) | ( n24616 & n24626 ) | ( ~n24615 & n24626 ) ;
  assign n24651 = ( n24566 & ~n24612 ) | ( n24566 & n24567 ) | ( ~n24612 & n24567 ) ;
  assign n24652 = ( n24477 & n24571 ) | ( n24477 & n24584 ) | ( n24571 & n24584 ) ;
  assign n24653 = ~n3644 & n19959 ;
  assign n24654 = n3652 &  n19040 ;
  assign n24655 = ( n3657 & ~n19494 ) | ( n3657 & 1'b0 ) | ( ~n19494 & 1'b0 ) ;
  assign n24656 = n24654 | n24655 ;
  assign n24657 = ~n3653 & n19951 ;
  assign n24658 = ( n3653 & ~n24656 ) | ( n3653 & n24657 ) | ( ~n24656 & n24657 ) ;
  assign n24659 = ~n24653 & n24658 ;
  assign n24660 = n1687 | n14763 ;
  assign n24661 = ( n3445 & n6627 ) | ( n3445 & n24660 ) | ( n6627 & n24660 ) ;
  assign n24662 = ( n3445 & ~n24661 ) | ( n3445 & 1'b0 ) | ( ~n24661 & 1'b0 ) ;
  assign n24663 = ( n1324 & ~n24662 ) | ( n1324 & n3346 ) | ( ~n24662 & n3346 ) ;
  assign n24664 = ( n3346 & ~n24663 ) | ( n3346 & 1'b0 ) | ( ~n24663 & 1'b0 ) ;
  assign n24665 = ( n23334 & n1580 ) | ( n23334 & n24664 ) | ( n1580 & n24664 ) ;
  assign n24666 = ~n1580 & n24665 ;
  assign n24667 = ( n409 & ~n383 ) | ( n409 & n24666 ) | ( ~n383 & n24666 ) ;
  assign n24668 = ~n409 & n24667 ;
  assign n24669 = ( n429 & ~n150 ) | ( n429 & n24668 ) | ( ~n150 & n24668 ) ;
  assign n24670 = ~n429 & n24669 ;
  assign n24671 = ( n217 & ~n800 ) | ( n217 & n24670 ) | ( ~n800 & n24670 ) ;
  assign n24672 = ~n217 & n24671 ;
  assign n24673 = ( n136 & ~n274 ) | ( n136 & n24672 ) | ( ~n274 & n24672 ) ;
  assign n24674 = ~n136 & n24673 ;
  assign n24675 = ( n24652 & ~n24659 ) | ( n24652 & n24674 ) | ( ~n24659 & n24674 ) ;
  assign n24676 = ( n24652 & ~n24674 ) | ( n24652 & n24659 ) | ( ~n24674 & n24659 ) ;
  assign n24677 = ( n24675 & ~n24652 ) | ( n24675 & n24676 ) | ( ~n24652 & n24676 ) ;
  assign n24681 = n20245 | n4430 ;
  assign n24678 = n523 | n20027 ;
  assign n24679 = n3939 | n20241 ;
  assign n24680 = n24678 &  n24679 ;
  assign n24682 = ( n4430 & ~n24681 ) | ( n4430 & n24680 ) | ( ~n24681 & n24680 ) ;
  assign n24683 = ( n601 & ~n24682 ) | ( n601 & n20265 ) | ( ~n24682 & n20265 ) ;
  assign n24684 = ( n20265 & ~n24683 ) | ( n20265 & 1'b0 ) | ( ~n24683 & 1'b0 ) ;
  assign n24686 = ( x29 & n24682 ) | ( x29 & n24684 ) | ( n24682 & n24684 ) ;
  assign n24685 = ( x29 & ~n24684 ) | ( x29 & n24682 ) | ( ~n24684 & n24682 ) ;
  assign n24687 = ( n24684 & ~n24686 ) | ( n24684 & n24685 ) | ( ~n24686 & n24685 ) ;
  assign n24688 = ( n24597 & n24677 ) | ( n24597 & n24687 ) | ( n24677 & n24687 ) ;
  assign n24689 = ( n24677 & ~n24597 ) | ( n24677 & n24687 ) | ( ~n24597 & n24687 ) ;
  assign n24690 = ( n24597 & ~n24688 ) | ( n24597 & n24689 ) | ( ~n24688 & n24689 ) ;
  assign n24691 = ( n24599 & ~n24598 ) | ( n24599 & n24609 ) | ( ~n24598 & n24609 ) ;
  assign n24692 = n4962 &  n20777 ;
  assign n24693 = ~n4482 & n20237 ;
  assign n24694 = n4495 | n20782 ;
  assign n24695 = ~n24693 & n24694 ;
  assign n24696 = ( n24692 & ~n20777 ) | ( n24692 & n24695 ) | ( ~n20777 & n24695 ) ;
  assign n24697 = n4478 | n20790 ;
  assign n24698 = n24696 &  n24697 ;
  assign n24699 = x26 &  n24698 ;
  assign n24700 = x26 | n24698 ;
  assign n24701 = ~n24699 & n24700 ;
  assign n24702 = ( n24690 & ~n24691 ) | ( n24690 & n24701 ) | ( ~n24691 & n24701 ) ;
  assign n24703 = ( n24690 & ~n24701 ) | ( n24690 & n24691 ) | ( ~n24701 & n24691 ) ;
  assign n24704 = ( n24702 & ~n24690 ) | ( n24702 & n24703 ) | ( ~n24690 & n24703 ) ;
  assign n24708 = ~n5135 & n21675 ;
  assign n24705 = n5010 | n21271 ;
  assign n24706 = ~n5067 & n21475 ;
  assign n24707 = ( n24705 & ~n24706 ) | ( n24705 & 1'b0 ) | ( ~n24706 & 1'b0 ) ;
  assign n24709 = ( n5135 & n24708 ) | ( n5135 & n24707 ) | ( n24708 & n24707 ) ;
  assign n24710 = n5012 | n21684 ;
  assign n24711 = n24709 &  n24710 ;
  assign n24712 = x23 &  n24711 ;
  assign n24713 = x23 | n24711 ;
  assign n24714 = ~n24712 & n24713 ;
  assign n24715 = ( n24651 & n24704 ) | ( n24651 & n24714 ) | ( n24704 & n24714 ) ;
  assign n24716 = ( n24704 & ~n24651 ) | ( n24704 & n24714 ) | ( ~n24651 & n24714 ) ;
  assign n24717 = ( n24651 & ~n24715 ) | ( n24651 & n24716 ) | ( ~n24715 & n24716 ) ;
  assign n24721 = n5837 | n22244 ;
  assign n24718 = ( n5339 & ~n21864 ) | ( n5339 & 1'b0 ) | ( ~n21864 & 1'b0 ) ;
  assign n24719 = n5761 | n22063 ;
  assign n24720 = ~n24718 & n24719 ;
  assign n24722 = ( n5837 & ~n24721 ) | ( n5837 & n24720 ) | ( ~n24721 & n24720 ) ;
  assign n24723 = ~n5341 & n22253 ;
  assign n24724 = ( n24722 & ~n24723 ) | ( n24722 & 1'b0 ) | ( ~n24723 & 1'b0 ) ;
  assign n24725 = x20 &  n24724 ;
  assign n24726 = x20 | n24724 ;
  assign n24727 = ~n24725 & n24726 ;
  assign n24728 = ( n24650 & n24717 ) | ( n24650 & n24727 ) | ( n24717 & n24727 ) ;
  assign n24729 = ( n24717 & ~n24650 ) | ( n24717 & n24727 ) | ( ~n24650 & n24727 ) ;
  assign n24730 = ( n24650 & ~n24728 ) | ( n24650 & n24729 ) | ( ~n24728 & n24729 ) ;
  assign n24731 = ( n24630 & ~n24629 ) | ( n24630 & n24640 ) | ( ~n24629 & n24640 ) ;
  assign n24732 = ( n24543 & ~n24643 ) | ( n24543 & n24549 ) | ( ~n24643 & n24549 ) ;
  assign n24734 = ( n24730 & n24731 ) | ( n24730 & n24732 ) | ( n24731 & n24732 ) ;
  assign n24733 = ( n24731 & ~n24730 ) | ( n24731 & n24732 ) | ( ~n24730 & n24732 ) ;
  assign n24735 = ( n24730 & ~n24734 ) | ( n24730 & n24733 ) | ( ~n24734 & n24733 ) ;
  assign n24736 = n24648 | n24735 ;
  assign n24737 = ( n24648 & ~n24735 ) | ( n24648 & 1'b0 ) | ( ~n24735 & 1'b0 ) ;
  assign n24738 = ( n24736 & ~n24648 ) | ( n24736 & n24737 ) | ( ~n24648 & n24737 ) ;
  assign n24739 = n24648 &  n24735 ;
  assign n24740 = ( n24691 & ~n24690 ) | ( n24691 & n24701 ) | ( ~n24690 & n24701 ) ;
  assign n24741 = n4430 &  n20237 ;
  assign n24742 = n523 | n20241 ;
  assign n24743 = ~n3939 & n20245 ;
  assign n24744 = ( n24742 & ~n24743 ) | ( n24742 & 1'b0 ) | ( ~n24743 & 1'b0 ) ;
  assign n24745 = ( n24741 & ~n20237 ) | ( n24741 & n24744 ) | ( ~n20237 & n24744 ) ;
  assign n24746 = n601 | n20253 ;
  assign n24747 = n24745 &  n24746 ;
  assign n24748 = x29 &  n24747 ;
  assign n24749 = x29 | n24747 ;
  assign n24750 = ~n24748 & n24749 ;
  assign n24751 = n3644 | n20035 ;
  assign n24752 = ( n3652 & ~n19494 ) | ( n3652 & 1'b0 ) | ( ~n19494 & 1'b0 ) ;
  assign n24753 = ( n3657 & ~n19951 ) | ( n3657 & 1'b0 ) | ( ~n19951 & 1'b0 ) ;
  assign n24754 = n24752 | n24753 ;
  assign n24755 = ~n3653 & n20027 ;
  assign n24756 = ( n3653 & ~n24754 ) | ( n3653 & n24755 ) | ( ~n24754 & n24755 ) ;
  assign n24757 = n24751 &  n24756 ;
  assign n24758 = n18932 | n24461 ;
  assign n24759 = ( n4868 & ~n6675 ) | ( n4868 & n24758 ) | ( ~n6675 & n24758 ) ;
  assign n24760 = ( n4868 & ~n24759 ) | ( n4868 & 1'b0 ) | ( ~n24759 & 1'b0 ) ;
  assign n24761 = ( n1360 & n4540 ) | ( n1360 & n24760 ) | ( n4540 & n24760 ) ;
  assign n24762 = ~n1360 & n24761 ;
  assign n24763 = ( n1491 & ~n227 ) | ( n1491 & n24762 ) | ( ~n227 & n24762 ) ;
  assign n24764 = ~n1491 & n24763 ;
  assign n24765 = ( n22627 & n1616 ) | ( n22627 & n24764 ) | ( n1616 & n24764 ) ;
  assign n24766 = ~n1616 & n24765 ;
  assign n24767 = ( n257 & ~n52 ) | ( n257 & n24766 ) | ( ~n52 & n24766 ) ;
  assign n24768 = ~n257 & n24767 ;
  assign n24769 = ( n95 & ~n417 ) | ( n95 & n24768 ) | ( ~n417 & n24768 ) ;
  assign n24770 = ~n95 & n24769 ;
  assign n24771 = ( n24757 & ~n24674 ) | ( n24757 & n24770 ) | ( ~n24674 & n24770 ) ;
  assign n24772 = ( n24674 & ~n24757 ) | ( n24674 & n24770 ) | ( ~n24757 & n24770 ) ;
  assign n24773 = ( n24771 & ~n24770 ) | ( n24771 & n24772 ) | ( ~n24770 & n24772 ) ;
  assign n24774 = ( n24597 & ~n24677 ) | ( n24597 & n24687 ) | ( ~n24677 & n24687 ) ;
  assign n24775 = ( n24676 & n24773 ) | ( n24676 & n24774 ) | ( n24773 & n24774 ) ;
  assign n24776 = ( n24773 & ~n24676 ) | ( n24773 & n24774 ) | ( ~n24676 & n24774 ) ;
  assign n24777 = ( n24676 & ~n24775 ) | ( n24676 & n24776 ) | ( ~n24775 & n24776 ) ;
  assign n24781 = ~n4962 & n21271 ;
  assign n24778 = n4482 | n20782 ;
  assign n24779 = ~n4495 & n20777 ;
  assign n24780 = ( n24778 & ~n24779 ) | ( n24778 & 1'b0 ) | ( ~n24779 & 1'b0 ) ;
  assign n24782 = ( n4962 & n24781 ) | ( n4962 & n24780 ) | ( n24781 & n24780 ) ;
  assign n24783 = n4478 | n21279 ;
  assign n24784 = n24782 &  n24783 ;
  assign n24785 = x26 | n24784 ;
  assign n24786 = ( x26 & ~n24784 ) | ( x26 & 1'b0 ) | ( ~n24784 & 1'b0 ) ;
  assign n24787 = ( n24785 & ~x26 ) | ( n24785 & n24786 ) | ( ~x26 & n24786 ) ;
  assign n24788 = ( n24750 & ~n24777 ) | ( n24750 & n24787 ) | ( ~n24777 & n24787 ) ;
  assign n24789 = ( n24750 & ~n24787 ) | ( n24750 & n24777 ) | ( ~n24787 & n24777 ) ;
  assign n24790 = ( n24788 & ~n24750 ) | ( n24788 & n24789 ) | ( ~n24750 & n24789 ) ;
  assign n24791 = ( n5135 & ~n21864 ) | ( n5135 & 1'b0 ) | ( ~n21864 & 1'b0 ) ;
  assign n24792 = ~n5010 & n21475 ;
  assign n24793 = n5067 | n21675 ;
  assign n24794 = ~n24792 & n24793 ;
  assign n24795 = ( n21864 & n24791 ) | ( n21864 & n24794 ) | ( n24791 & n24794 ) ;
  assign n24796 = ~n5012 & n21872 ;
  assign n24797 = ( n24795 & ~n24796 ) | ( n24795 & 1'b0 ) | ( ~n24796 & 1'b0 ) ;
  assign n24798 = x23 &  n24797 ;
  assign n24799 = x23 | n24797 ;
  assign n24800 = ~n24798 & n24799 ;
  assign n24801 = ( n24740 & n24790 ) | ( n24740 & n24800 ) | ( n24790 & n24800 ) ;
  assign n24802 = ( n24790 & ~n24740 ) | ( n24790 & n24800 ) | ( ~n24740 & n24800 ) ;
  assign n24803 = ( n24740 & ~n24801 ) | ( n24740 & n24802 ) | ( ~n24801 & n24802 ) ;
  assign n24804 = ( n24651 & ~n24704 ) | ( n24651 & n24714 ) | ( ~n24704 & n24714 ) ;
  assign n24805 = ~n19402 & n22244 ;
  assign n24806 = ( n5339 & ~n22063 ) | ( n5339 & 1'b0 ) | ( ~n22063 & 1'b0 ) ;
  assign n24807 = n24805 | n24806 ;
  assign n24808 = ~n5341 & n22251 ;
  assign n24809 = ( n5341 & ~n24807 ) | ( n5341 & n24808 ) | ( ~n24807 & n24808 ) ;
  assign n24811 = ( x20 & n24804 ) | ( x20 & n24809 ) | ( n24804 & n24809 ) ;
  assign n24810 = ( x20 & ~n24804 ) | ( x20 & n24809 ) | ( ~n24804 & n24809 ) ;
  assign n24812 = ( n24804 & ~n24811 ) | ( n24804 & n24810 ) | ( ~n24811 & n24810 ) ;
  assign n24813 = ( n24803 & ~n24812 ) | ( n24803 & 1'b0 ) | ( ~n24812 & 1'b0 ) ;
  assign n24814 = ~n24803 & n24812 ;
  assign n24815 = n24813 | n24814 ;
  assign n24816 = ( n24650 & ~n24717 ) | ( n24650 & n24727 ) | ( ~n24717 & n24727 ) ;
  assign n24817 = ( n24815 & ~n24733 ) | ( n24815 & n24816 ) | ( ~n24733 & n24816 ) ;
  assign n24818 = ( n24733 & ~n24815 ) | ( n24733 & n24816 ) | ( ~n24815 & n24816 ) ;
  assign n24819 = ( n24817 & ~n24816 ) | ( n24817 & n24818 ) | ( ~n24816 & n24818 ) ;
  assign n24820 = n24739 &  n24819 ;
  assign n24821 = n24739 | n24819 ;
  assign n24822 = ~n24820 & n24821 ;
  assign n24827 = ( n24740 & ~n24790 ) | ( n24740 & n24800 ) | ( ~n24790 & n24800 ) ;
  assign n24838 = ( n24676 & ~n24773 ) | ( n24676 & n24774 ) | ( ~n24773 & n24774 ) ;
  assign n24863 = n3644 | n20280 ;
  assign n24864 = ( n3652 & ~n19951 ) | ( n3652 & 1'b0 ) | ( ~n19951 & 1'b0 ) ;
  assign n24865 = ( n3657 & ~n20027 ) | ( n3657 & 1'b0 ) | ( ~n20027 & 1'b0 ) ;
  assign n24866 = n24864 | n24865 ;
  assign n24867 = ~n3653 & n20241 ;
  assign n24868 = ( n3653 & ~n24866 ) | ( n3653 & n24867 ) | ( ~n24866 & n24867 ) ;
  assign n24869 = n24863 &  n24868 ;
  assign n24843 = n1051 | n3474 ;
  assign n24844 = ( n15926 & ~n1357 ) | ( n15926 & n24843 ) | ( ~n1357 & n24843 ) ;
  assign n24845 = n1357 | n24844 ;
  assign n24846 = ( n4832 & ~n14128 ) | ( n4832 & n24845 ) | ( ~n14128 & n24845 ) ;
  assign n24847 = ( n4832 & ~n24846 ) | ( n4832 & 1'b0 ) | ( ~n24846 & 1'b0 ) ;
  assign n24848 = ( n1820 & n2009 ) | ( n1820 & n24847 ) | ( n2009 & n24847 ) ;
  assign n24849 = ~n1820 & n24848 ;
  assign n24850 = ( n528 & ~n3287 ) | ( n528 & n24849 ) | ( ~n3287 & n24849 ) ;
  assign n24851 = ~n528 & n24850 ;
  assign n24852 = ( n1185 & ~n24851 ) | ( n1185 & n1279 ) | ( ~n24851 & n1279 ) ;
  assign n24853 = ( n1279 & ~n24852 ) | ( n1279 & 1'b0 ) | ( ~n24852 & 1'b0 ) ;
  assign n24854 = ( n712 & ~n125 ) | ( n712 & n24853 ) | ( ~n125 & n24853 ) ;
  assign n24855 = ~n712 & n24854 ;
  assign n24856 = ( n333 & ~n531 ) | ( n333 & n24855 ) | ( ~n531 & n24855 ) ;
  assign n24857 = ~n333 & n24856 ;
  assign n24858 = ( n169 & ~n281 ) | ( n169 & n24857 ) | ( ~n281 & n24857 ) ;
  assign n24859 = ~n169 & n24858 ;
  assign n24839 = n19919 &  n22244 ;
  assign n24840 = ~x20 & n24839 ;
  assign n24841 = ( x20 & ~n24839 ) | ( x20 & 1'b0 ) | ( ~n24839 & 1'b0 ) ;
  assign n24842 = n24840 | n24841 ;
  assign n24860 = ( n24674 & ~n24859 ) | ( n24674 & n24842 ) | ( ~n24859 & n24842 ) ;
  assign n24861 = ( n24842 & ~n24674 ) | ( n24842 & n24859 ) | ( ~n24674 & n24859 ) ;
  assign n24862 = ( n24860 & ~n24842 ) | ( n24860 & n24861 ) | ( ~n24842 & n24861 ) ;
  assign n24871 = ( n24771 & n24862 ) | ( n24771 & n24869 ) | ( n24862 & n24869 ) ;
  assign n24870 = ( n24771 & ~n24869 ) | ( n24771 & n24862 ) | ( ~n24869 & n24862 ) ;
  assign n24872 = ( n24869 & ~n24871 ) | ( n24869 & n24870 ) | ( ~n24871 & n24870 ) ;
  assign n24873 = ~n523 & n20245 ;
  assign n24874 = ~n3939 & n20237 ;
  assign n24875 = n24873 | n24874 ;
  assign n24876 = ~n4430 & n20782 ;
  assign n24877 = ( n4430 & ~n24875 ) | ( n4430 & n24876 ) | ( ~n24875 & n24876 ) ;
  assign n24878 = n601 | n21227 ;
  assign n24879 = n24877 &  n24878 ;
  assign n24880 = x29 &  n24879 ;
  assign n24881 = x29 | n24879 ;
  assign n24882 = ~n24880 & n24881 ;
  assign n24883 = ( n24838 & ~n24872 ) | ( n24838 & n24882 ) | ( ~n24872 & n24882 ) ;
  assign n24884 = ( n24838 & ~n24882 ) | ( n24838 & n24872 ) | ( ~n24882 & n24872 ) ;
  assign n24885 = ( n24883 & ~n24838 ) | ( n24883 & n24884 ) | ( ~n24838 & n24884 ) ;
  assign n24831 = n21475 | n4962 ;
  assign n24828 = ~n4482 & n20777 ;
  assign n24829 = n4495 | n21271 ;
  assign n24830 = ~n24828 & n24829 ;
  assign n24832 = ( n4962 & ~n24831 ) | ( n4962 & n24830 ) | ( ~n24831 & n24830 ) ;
  assign n24833 = n4478 | n21484 ;
  assign n24834 = n24832 &  n24833 ;
  assign n24835 = x26 &  n24834 ;
  assign n24836 = x26 | n24834 ;
  assign n24837 = ~n24835 & n24836 ;
  assign n24886 = ( n24788 & ~n24885 ) | ( n24788 & n24837 ) | ( ~n24885 & n24837 ) ;
  assign n24887 = ( n24837 & ~n24788 ) | ( n24837 & n24885 ) | ( ~n24788 & n24885 ) ;
  assign n24888 = ( n24886 & ~n24837 ) | ( n24886 & n24887 ) | ( ~n24837 & n24887 ) ;
  assign n24892 = ~n5135 & n22063 ;
  assign n24889 = n5010 | n21675 ;
  assign n24890 = n5067 | n21864 ;
  assign n24891 = n24889 &  n24890 ;
  assign n24893 = ( n5135 & n24892 ) | ( n5135 & n24891 ) | ( n24892 & n24891 ) ;
  assign n24894 = n5012 | n22071 ;
  assign n24895 = n24893 &  n24894 ;
  assign n24896 = x23 &  n24895 ;
  assign n24897 = x23 | n24895 ;
  assign n24898 = ~n24896 & n24897 ;
  assign n24899 = ( n24827 & n24888 ) | ( n24827 & n24898 ) | ( n24888 & n24898 ) ;
  assign n24900 = ( n24888 & ~n24827 ) | ( n24888 & n24898 ) | ( ~n24827 & n24898 ) ;
  assign n24901 = ( n24827 & ~n24899 ) | ( n24827 & n24900 ) | ( ~n24899 & n24900 ) ;
  assign n24823 = x20 &  n24809 ;
  assign n24824 = x20 | n24809 ;
  assign n24825 = ~n24823 & n24824 ;
  assign n24826 = ( n24804 & ~n24803 ) | ( n24804 & n24825 ) | ( ~n24803 & n24825 ) ;
  assign n24902 = ( n24818 & ~n24901 ) | ( n24818 & n24826 ) | ( ~n24901 & n24826 ) ;
  assign n24903 = ( n24818 & ~n24826 ) | ( n24818 & n24901 ) | ( ~n24826 & n24901 ) ;
  assign n24904 = ( n24902 & ~n24818 ) | ( n24902 & n24903 ) | ( ~n24818 & n24903 ) ;
  assign n24905 = ~n24820 & n24904 ;
  assign n24906 = ( n24820 & ~n24904 ) | ( n24820 & 1'b0 ) | ( ~n24904 & 1'b0 ) ;
  assign n24907 = n24905 | n24906 ;
  assign n24909 = ( n24788 & n24837 ) | ( n24788 & n24885 ) | ( n24837 & n24885 ) ;
  assign n24910 = ( n24674 & n24842 ) | ( n24674 & n24859 ) | ( n24842 & n24859 ) ;
  assign n24911 = ~n3644 & n20265 ;
  assign n24915 = n20245 | n3653 ;
  assign n24912 = ( n3652 & ~n20027 ) | ( n3652 & 1'b0 ) | ( ~n20027 & 1'b0 ) ;
  assign n24913 = ( n3657 & ~n20241 ) | ( n3657 & 1'b0 ) | ( ~n20241 & 1'b0 ) ;
  assign n24914 = n24912 | n24913 ;
  assign n24916 = ( n24915 & ~n3653 ) | ( n24915 & n24914 ) | ( ~n3653 & n24914 ) ;
  assign n24917 = n24911 | n24916 ;
  assign n24918 = n2633 | n5247 ;
  assign n24919 = ( n2544 & ~n2508 ) | ( n2544 & n24918 ) | ( ~n2508 & n24918 ) ;
  assign n24920 = n2508 | n24919 ;
  assign n24921 = ( n24920 & ~n1270 ) | ( n24920 & n16407 ) | ( ~n1270 & n16407 ) ;
  assign n24922 = n1270 | n24921 ;
  assign n24923 = ( n2588 & ~n24922 ) | ( n2588 & n4559 ) | ( ~n24922 & n4559 ) ;
  assign n24924 = ~n2588 & n24923 ;
  assign n24925 = ( n4226 & ~n11336 ) | ( n4226 & n24924 ) | ( ~n11336 & n24924 ) ;
  assign n24926 = ~n4226 & n24925 ;
  assign n24927 = ( n127 & ~n2191 ) | ( n127 & n24926 ) | ( ~n2191 & n24926 ) ;
  assign n24928 = ~n127 & n24927 ;
  assign n24929 = ( n558 & ~n257 ) | ( n558 & n24928 ) | ( ~n257 & n24928 ) ;
  assign n24930 = ~n558 & n24929 ;
  assign n24931 = ( n225 & ~n267 ) | ( n225 & n24930 ) | ( ~n267 & n24930 ) ;
  assign n24932 = ~n225 & n24931 ;
  assign n24933 = ( n24910 & n24917 ) | ( n24910 & n24932 ) | ( n24917 & n24932 ) ;
  assign n24934 = ( n24917 & ~n24910 ) | ( n24917 & n24932 ) | ( ~n24910 & n24932 ) ;
  assign n24935 = ( n24910 & ~n24933 ) | ( n24910 & n24934 ) | ( ~n24933 & n24934 ) ;
  assign n24936 = n4430 &  n20777 ;
  assign n24937 = ~n523 & n20237 ;
  assign n24938 = n3939 | n20782 ;
  assign n24939 = ~n24937 & n24938 ;
  assign n24940 = ( n24936 & ~n20777 ) | ( n24936 & n24939 ) | ( ~n20777 & n24939 ) ;
  assign n24941 = ( n20790 & ~n601 ) | ( n20790 & n24940 ) | ( ~n601 & n24940 ) ;
  assign n24942 = ~n20790 & n24941 ;
  assign n24944 = ( x29 & n24940 ) | ( x29 & n24942 ) | ( n24940 & n24942 ) ;
  assign n24943 = ( x29 & ~n24942 ) | ( x29 & n24940 ) | ( ~n24942 & n24940 ) ;
  assign n24945 = ( n24942 & ~n24944 ) | ( n24942 & n24943 ) | ( ~n24944 & n24943 ) ;
  assign n24946 = ( n24871 & ~n24935 ) | ( n24871 & n24945 ) | ( ~n24935 & n24945 ) ;
  assign n24947 = ( n24871 & ~n24945 ) | ( n24871 & n24935 ) | ( ~n24945 & n24935 ) ;
  assign n24948 = ( n24946 & ~n24871 ) | ( n24946 & n24947 ) | ( ~n24871 & n24947 ) ;
  assign n24953 = ~n4962 & n21675 ;
  assign n24950 = n4482 | n21271 ;
  assign n24951 = ~n4495 & n21475 ;
  assign n24952 = ( n24950 & ~n24951 ) | ( n24950 & 1'b0 ) | ( ~n24951 & 1'b0 ) ;
  assign n24954 = ( n4962 & n24953 ) | ( n4962 & n24952 ) | ( n24953 & n24952 ) ;
  assign n24955 = n4478 | n21684 ;
  assign n24956 = n24954 &  n24955 ;
  assign n24957 = x26 &  n24956 ;
  assign n24958 = x26 | n24956 ;
  assign n24959 = ~n24957 & n24958 ;
  assign n24949 = ( n24838 & n24872 ) | ( n24838 & n24882 ) | ( n24872 & n24882 ) ;
  assign n24960 = ( n24948 & ~n24959 ) | ( n24948 & n24949 ) | ( ~n24959 & n24949 ) ;
  assign n24961 = ( n24948 & ~n24949 ) | ( n24948 & n24959 ) | ( ~n24949 & n24959 ) ;
  assign n24962 = ( n24960 & ~n24948 ) | ( n24960 & n24961 ) | ( ~n24948 & n24961 ) ;
  assign n24966 = n22244 | n5135 ;
  assign n24963 = n5010 | n21864 ;
  assign n24964 = n5067 | n22063 ;
  assign n24965 = n24963 &  n24964 ;
  assign n24967 = ( n5135 & ~n24966 ) | ( n5135 & n24965 ) | ( ~n24966 & n24965 ) ;
  assign n24968 = ~n5012 & n22253 ;
  assign n24969 = ( n24967 & ~n24968 ) | ( n24967 & 1'b0 ) | ( ~n24968 & 1'b0 ) ;
  assign n24970 = x23 &  n24969 ;
  assign n24971 = x23 | n24969 ;
  assign n24972 = ~n24970 & n24971 ;
  assign n24973 = ( n24909 & ~n24962 ) | ( n24909 & n24972 ) | ( ~n24962 & n24972 ) ;
  assign n24974 = ( n24909 & ~n24972 ) | ( n24909 & n24962 ) | ( ~n24972 & n24962 ) ;
  assign n24975 = ( n24973 & ~n24909 ) | ( n24973 & n24974 ) | ( ~n24909 & n24974 ) ;
  assign n24908 = ( n24818 & n24826 ) | ( n24818 & n24901 ) | ( n24826 & n24901 ) ;
  assign n24976 = ( n24899 & n24908 ) | ( n24899 & n24975 ) | ( n24908 & n24975 ) ;
  assign n24977 = ( n24899 & ~n24975 ) | ( n24899 & n24908 ) | ( ~n24975 & n24908 ) ;
  assign n24978 = ( n24975 & ~n24976 ) | ( n24975 & n24977 ) | ( ~n24976 & n24977 ) ;
  assign n24980 = n24906 &  n24978 ;
  assign n24979 = ~n24906 & n24978 ;
  assign n24981 = ( n24906 & ~n24980 ) | ( n24906 & n24979 ) | ( ~n24980 & n24979 ) ;
  assign n25046 = ( n24909 & n24962 ) | ( n24909 & n24972 ) | ( n24962 & n24972 ) ;
  assign n24985 = ~n4430 & n21271 ;
  assign n24982 = n523 | n20782 ;
  assign n24983 = ~n3939 & n20777 ;
  assign n24984 = ( n24982 & ~n24983 ) | ( n24982 & 1'b0 ) | ( ~n24983 & 1'b0 ) ;
  assign n24986 = ( n4430 & n24985 ) | ( n4430 & n24984 ) | ( n24985 & n24984 ) ;
  assign n24987 = n601 | n21279 ;
  assign n24988 = n24986 &  n24987 ;
  assign n24989 = x29 &  n24988 ;
  assign n24990 = x29 | n24988 ;
  assign n24991 = ~n24989 & n24990 ;
  assign n25010 = n3644 | n20253 ;
  assign n25011 = ( n3652 & ~n20241 ) | ( n3652 & 1'b0 ) | ( ~n20241 & 1'b0 ) ;
  assign n25012 = n3657 &  n20245 ;
  assign n25013 = n25011 | n25012 ;
  assign n25014 = n3653 | n20237 ;
  assign n25015 = ( n25013 & ~n3653 ) | ( n25013 & n25014 ) | ( ~n3653 & n25014 ) ;
  assign n25016 = ( n25010 & ~n25015 ) | ( n25010 & 1'b0 ) | ( ~n25015 & 1'b0 ) ;
  assign n24992 = n142 | n14765 ;
  assign n24993 = ( n14642 & ~n2035 ) | ( n14642 & n24992 ) | ( ~n2035 & n24992 ) ;
  assign n24994 = n2035 | n24993 ;
  assign n24995 = ( n3679 & n20159 ) | ( n3679 & n24994 ) | ( n20159 & n24994 ) ;
  assign n24996 = ( n3679 & ~n24995 ) | ( n3679 & 1'b0 ) | ( ~n24995 & 1'b0 ) ;
  assign n24997 = ( n1360 & ~n23342 ) | ( n1360 & n24996 ) | ( ~n23342 & n24996 ) ;
  assign n24998 = ~n1360 & n24997 ;
  assign n24999 = ( n1511 & ~n2191 ) | ( n1511 & n24998 ) | ( ~n2191 & n24998 ) ;
  assign n25000 = ~n1511 & n24999 ;
  assign n25001 = ( n450 & ~n645 ) | ( n450 & n25000 ) | ( ~n645 & n25000 ) ;
  assign n25002 = n645 &  n25001 ;
  assign n25003 = ( n720 & ~n105 ) | ( n720 & n25002 ) | ( ~n105 & n25002 ) ;
  assign n25004 = ~n720 & n25003 ;
  assign n25005 = ( n909 & ~n559 ) | ( n909 & n25004 ) | ( ~n559 & n25004 ) ;
  assign n25006 = ~n909 & n25005 ;
  assign n25007 = ( n24932 & ~n25006 ) | ( n24932 & n24934 ) | ( ~n25006 & n24934 ) ;
  assign n25008 = ( n24934 & ~n24932 ) | ( n24934 & n25006 ) | ( ~n24932 & n25006 ) ;
  assign n25009 = ( n25007 & ~n24934 ) | ( n25007 & n25008 ) | ( ~n24934 & n25008 ) ;
  assign n25017 = ( n24871 & n24935 ) | ( n24871 & n24945 ) | ( n24935 & n24945 ) ;
  assign n25018 = ( n25016 & ~n25009 ) | ( n25016 & n25017 ) | ( ~n25009 & n25017 ) ;
  assign n25019 = ( n25009 & ~n25016 ) | ( n25009 & n25017 ) | ( ~n25016 & n25017 ) ;
  assign n25020 = ( n25018 & ~n25017 ) | ( n25018 & n25019 ) | ( ~n25017 & n25019 ) ;
  assign n25021 = ( n4962 & ~n21864 ) | ( n4962 & 1'b0 ) | ( ~n21864 & 1'b0 ) ;
  assign n25022 = ~n4482 & n21475 ;
  assign n25023 = n4495 | n21675 ;
  assign n25024 = ~n25022 & n25023 ;
  assign n25025 = ( n21864 & n25021 ) | ( n21864 & n25024 ) | ( n25021 & n25024 ) ;
  assign n25026 = ~n4478 & n21872 ;
  assign n25027 = ( n25025 & ~n25026 ) | ( n25025 & 1'b0 ) | ( ~n25026 & 1'b0 ) ;
  assign n25028 = x26 &  n25027 ;
  assign n25029 = x26 | n25027 ;
  assign n25030 = ~n25028 & n25029 ;
  assign n25031 = ( n24991 & n25020 ) | ( n24991 & n25030 ) | ( n25020 & n25030 ) ;
  assign n25032 = ( n25020 & ~n24991 ) | ( n25020 & n25030 ) | ( ~n24991 & n25030 ) ;
  assign n25033 = ( n24991 & ~n25031 ) | ( n24991 & n25032 ) | ( ~n25031 & n25032 ) ;
  assign n25034 = ( n24948 & n24949 ) | ( n24948 & n24959 ) | ( n24949 & n24959 ) ;
  assign n25035 = ( n5012 & ~n22251 ) | ( n5012 & 1'b0 ) | ( ~n22251 & 1'b0 ) ;
  assign n25036 = ~n20215 & n22244 ;
  assign n25037 = n5010 | n22063 ;
  assign n25038 = ~n25036 & n25037 ;
  assign n25039 = ( n22251 & n25035 ) | ( n22251 & n25038 ) | ( n25035 & n25038 ) ;
  assign n25041 = ( x23 & n25034 ) | ( x23 & n25039 ) | ( n25034 & n25039 ) ;
  assign n25040 = ( x23 & ~n25034 ) | ( x23 & n25039 ) | ( ~n25034 & n25039 ) ;
  assign n25042 = ( n25034 & ~n25041 ) | ( n25034 & n25040 ) | ( ~n25041 & n25040 ) ;
  assign n25043 = n25033 | n25042 ;
  assign n25044 = n25033 &  n25042 ;
  assign n25045 = ( n25043 & ~n25044 ) | ( n25043 & 1'b0 ) | ( ~n25044 & 1'b0 ) ;
  assign n25048 = ( n24976 & n25045 ) | ( n24976 & n25046 ) | ( n25045 & n25046 ) ;
  assign n25047 = ( n24976 & ~n25046 ) | ( n24976 & n25045 ) | ( ~n25046 & n25045 ) ;
  assign n25049 = ( n25046 & ~n25048 ) | ( n25046 & n25047 ) | ( ~n25048 & n25047 ) ;
  assign n25050 = ( n24906 & ~n24978 ) | ( n24906 & 1'b0 ) | ( ~n24978 & 1'b0 ) ;
  assign n25051 = ~n25049 & n25050 ;
  assign n25052 = ( n25049 & ~n25050 ) | ( n25049 & 1'b0 ) | ( ~n25050 & 1'b0 ) ;
  assign n25053 = n25051 | n25052 ;
  assign n25061 = ~n4962 & n22063 ;
  assign n25058 = n4482 | n21675 ;
  assign n25059 = n4495 | n21864 ;
  assign n25060 = n25058 &  n25059 ;
  assign n25062 = ( n4962 & n25061 ) | ( n4962 & n25060 ) | ( n25061 & n25060 ) ;
  assign n25063 = n4478 | n22071 ;
  assign n25064 = n25062 &  n25063 ;
  assign n25065 = x26 &  n25064 ;
  assign n25066 = x26 | n25064 ;
  assign n25067 = ~n25065 & n25066 ;
  assign n25068 = ( n25009 & n25016 ) | ( n25009 & n25017 ) | ( n25016 & n25017 ) ;
  assign n25073 = ~n5230 & n13803 ;
  assign n25074 = ( n619 & n760 ) | ( n619 & n25073 ) | ( n760 & n25073 ) ;
  assign n25075 = ~n619 & n25074 ;
  assign n25076 = ( n1428 & ~n691 ) | ( n1428 & n25075 ) | ( ~n691 & n25075 ) ;
  assign n25077 = ~n1428 & n25076 ;
  assign n25078 = ( n947 & ~n777 ) | ( n947 & n25077 ) | ( ~n777 & n25077 ) ;
  assign n25079 = ~n947 & n25078 ;
  assign n25080 = ( n525 & ~n25079 ) | ( n525 & n788 ) | ( ~n25079 & n788 ) ;
  assign n25081 = ( n525 & ~n25080 ) | ( n525 & 1'b0 ) | ( ~n25080 & 1'b0 ) ;
  assign n25082 = ( n453 & ~n425 ) | ( n453 & n25081 ) | ( ~n425 & n25081 ) ;
  assign n25083 = ~n453 & n25082 ;
  assign n25084 = ( n192 & ~n485 ) | ( n192 & n25083 ) | ( ~n485 & n25083 ) ;
  assign n25085 = ~n192 & n25084 ;
  assign n25086 = ~n88 & n25085 ;
  assign n25069 = n20124 &  n22244 ;
  assign n25070 = ~x23 & n25069 ;
  assign n25071 = ( x23 & ~n25069 ) | ( x23 & 1'b0 ) | ( ~n25069 & 1'b0 ) ;
  assign n25072 = n25070 | n25071 ;
  assign n25087 = ( n25006 & ~n25086 ) | ( n25006 & n25072 ) | ( ~n25086 & n25072 ) ;
  assign n25088 = ( n25072 & ~n25006 ) | ( n25072 & n25086 ) | ( ~n25006 & n25086 ) ;
  assign n25089 = ( n25087 & ~n25072 ) | ( n25087 & n25088 ) | ( ~n25072 & n25088 ) ;
  assign n25090 = n3644 | n21227 ;
  assign n25091 = n3652 &  n20245 ;
  assign n25092 = n3657 &  n20237 ;
  assign n25093 = n25091 | n25092 ;
  assign n25094 = ~n3653 & n20782 ;
  assign n25095 = ( n3653 & ~n25093 ) | ( n3653 & n25094 ) | ( ~n25093 & n25094 ) ;
  assign n25096 = n25090 &  n25095 ;
  assign n25097 = ( n25008 & ~n25089 ) | ( n25008 & n25096 ) | ( ~n25089 & n25096 ) ;
  assign n25098 = ( n25089 & ~n25008 ) | ( n25089 & n25096 ) | ( ~n25008 & n25096 ) ;
  assign n25099 = ( n25097 & ~n25096 ) | ( n25097 & n25098 ) | ( ~n25096 & n25098 ) ;
  assign n25103 = n21475 | n4430 ;
  assign n25100 = ~n523 & n20777 ;
  assign n25101 = n3939 | n21271 ;
  assign n25102 = ~n25100 & n25101 ;
  assign n25104 = ( n4430 & ~n25103 ) | ( n4430 & n25102 ) | ( ~n25103 & n25102 ) ;
  assign n25105 = n601 | n21484 ;
  assign n25106 = n25104 &  n25105 ;
  assign n25107 = x29 &  n25106 ;
  assign n25108 = x29 | n25106 ;
  assign n25109 = ~n25107 & n25108 ;
  assign n25110 = ( n25068 & n25099 ) | ( n25068 & n25109 ) | ( n25099 & n25109 ) ;
  assign n25111 = ( n25099 & ~n25068 ) | ( n25099 & n25109 ) | ( ~n25068 & n25109 ) ;
  assign n25112 = ( n25068 & ~n25110 ) | ( n25068 & n25111 ) | ( ~n25110 & n25111 ) ;
  assign n25114 = ( n25031 & n25067 ) | ( n25031 & n25112 ) | ( n25067 & n25112 ) ;
  assign n25113 = ( n25031 & ~n25067 ) | ( n25031 & n25112 ) | ( ~n25067 & n25112 ) ;
  assign n25115 = ( n25067 & ~n25114 ) | ( n25067 & n25113 ) | ( ~n25114 & n25113 ) ;
  assign n25054 = x23 &  n25039 ;
  assign n25055 = x23 | n25039 ;
  assign n25056 = ~n25054 & n25055 ;
  assign n25057 = ( n25033 & n25034 ) | ( n25033 & n25056 ) | ( n25034 & n25056 ) ;
  assign n25116 = ( n25048 & ~n25115 ) | ( n25048 & n25057 ) | ( ~n25115 & n25057 ) ;
  assign n25117 = ( n25048 & ~n25057 ) | ( n25048 & n25115 ) | ( ~n25057 & n25115 ) ;
  assign n25118 = ( n25116 & ~n25048 ) | ( n25116 & n25117 ) | ( ~n25048 & n25117 ) ;
  assign n25119 = n25051 | n25118 ;
  assign n25120 = n25051 &  n25118 ;
  assign n25121 = ( n25119 & ~n25120 ) | ( n25119 & 1'b0 ) | ( ~n25120 & 1'b0 ) ;
  assign n25122 = ( n25031 & ~n25112 ) | ( n25031 & n25067 ) | ( ~n25112 & n25067 ) ;
  assign n25123 = ( n25068 & ~n25099 ) | ( n25068 & n25109 ) | ( ~n25099 & n25109 ) ;
  assign n25167 = n22244 | n4962 ;
  assign n25164 = n4482 | n21864 ;
  assign n25165 = n4495 | n22063 ;
  assign n25166 = n25164 &  n25165 ;
  assign n25168 = ( n4962 & ~n25167 ) | ( n4962 & n25166 ) | ( ~n25167 & n25166 ) ;
  assign n25169 = ~n4478 & n22253 ;
  assign n25170 = ( n25168 & ~n25169 ) | ( n25168 & 1'b0 ) | ( ~n25169 & 1'b0 ) ;
  assign n25171 = x26 &  n25170 ;
  assign n25172 = x26 | n25170 ;
  assign n25173 = ~n25171 & n25172 ;
  assign n25124 = ( n25006 & n25072 ) | ( n25006 & n25086 ) | ( n25072 & n25086 ) ;
  assign n25125 = n3644 | n20790 ;
  assign n25126 = n3652 &  n20237 ;
  assign n25127 = ( n3657 & ~n20782 ) | ( n3657 & 1'b0 ) | ( ~n20782 & 1'b0 ) ;
  assign n25128 = n25126 | n25127 ;
  assign n25129 = n3653 | n20777 ;
  assign n25130 = ( n25128 & ~n3653 ) | ( n25128 & n25129 ) | ( ~n3653 & n25129 ) ;
  assign n25131 = ( n25125 & ~n25130 ) | ( n25125 & 1'b0 ) | ( ~n25130 & 1'b0 ) ;
  assign n25132 = n2632 | n16973 ;
  assign n25133 = ( n25132 & ~n1130 ) | ( n25132 & n6714 ) | ( ~n1130 & n6714 ) ;
  assign n25134 = n1130 | n25133 ;
  assign n25135 = ( n20689 & n14632 ) | ( n20689 & n25134 ) | ( n14632 & n25134 ) ;
  assign n25136 = ( n14632 & ~n25135 ) | ( n14632 & 1'b0 ) | ( ~n25135 & 1'b0 ) ;
  assign n25137 = ( n25136 & ~n754 ) | ( n25136 & n874 ) | ( ~n754 & n874 ) ;
  assign n25138 = ~n874 & n25137 ;
  assign n25139 = ( n2128 & ~n647 ) | ( n2128 & n25138 ) | ( ~n647 & n25138 ) ;
  assign n25140 = ~n2128 & n25139 ;
  assign n25141 = ( n238 & ~n715 ) | ( n238 & n25140 ) | ( ~n715 & n25140 ) ;
  assign n25142 = ~n238 & n25141 ;
  assign n25143 = ( n355 & ~n25142 ) | ( n355 & n712 ) | ( ~n25142 & n712 ) ;
  assign n25144 = ( n355 & ~n25143 ) | ( n355 & 1'b0 ) | ( ~n25143 & 1'b0 ) ;
  assign n25145 = ( n267 & ~n89 ) | ( n267 & n25144 ) | ( ~n89 & n25144 ) ;
  assign n25146 = ~n267 & n25145 ;
  assign n25147 = ~n86 & n25146 ;
  assign n25148 = ( n25124 & ~n25131 ) | ( n25124 & n25147 ) | ( ~n25131 & n25147 ) ;
  assign n25149 = ( n25124 & ~n25147 ) | ( n25124 & n25131 ) | ( ~n25147 & n25131 ) ;
  assign n25150 = ( n25148 & ~n25124 ) | ( n25148 & n25149 ) | ( ~n25124 & n25149 ) ;
  assign n25154 = ~n4430 & n21675 ;
  assign n25151 = n523 | n21271 ;
  assign n25152 = ~n3939 & n21475 ;
  assign n25153 = ( n25151 & ~n25152 ) | ( n25151 & 1'b0 ) | ( ~n25152 & 1'b0 ) ;
  assign n25155 = ( n4430 & n25154 ) | ( n4430 & n25153 ) | ( n25154 & n25153 ) ;
  assign n25156 = ( n21684 & ~n601 ) | ( n21684 & n25155 ) | ( ~n601 & n25155 ) ;
  assign n25157 = ~n21684 & n25156 ;
  assign n25158 = ( x29 & ~n25155 ) | ( x29 & n25157 ) | ( ~n25155 & n25157 ) ;
  assign n25159 = ( n25155 & ~x29 ) | ( n25155 & n25157 ) | ( ~x29 & n25157 ) ;
  assign n25160 = ( n25158 & ~n25157 ) | ( n25158 & n25159 ) | ( ~n25157 & n25159 ) ;
  assign n25161 = ( n25098 & n25150 ) | ( n25098 & n25160 ) | ( n25150 & n25160 ) ;
  assign n25162 = ( n25150 & ~n25098 ) | ( n25150 & n25160 ) | ( ~n25098 & n25160 ) ;
  assign n25163 = ( n25098 & ~n25161 ) | ( n25098 & n25162 ) | ( ~n25161 & n25162 ) ;
  assign n25174 = ( n25123 & ~n25173 ) | ( n25123 & n25163 ) | ( ~n25173 & n25163 ) ;
  assign n25175 = ( n25163 & ~n25123 ) | ( n25163 & n25173 ) | ( ~n25123 & n25173 ) ;
  assign n25176 = ( n25174 & ~n25163 ) | ( n25174 & n25175 ) | ( ~n25163 & n25175 ) ;
  assign n25177 = ( n25116 & ~n25122 ) | ( n25116 & n25176 ) | ( ~n25122 & n25176 ) ;
  assign n25178 = ( n25122 & ~n25116 ) | ( n25122 & n25176 ) | ( ~n25116 & n25176 ) ;
  assign n25179 = ( n25177 & ~n25176 ) | ( n25177 & n25178 ) | ( ~n25176 & n25178 ) ;
  assign n25180 = n25120 | n25179 ;
  assign n25181 = ( n25120 & ~n25179 ) | ( n25120 & 1'b0 ) | ( ~n25179 & 1'b0 ) ;
  assign n25182 = ( n25180 & ~n25120 ) | ( n25180 & n25181 ) | ( ~n25120 & n25181 ) ;
  assign n25183 = ( n25116 & ~n25176 ) | ( n25116 & n25122 ) | ( ~n25176 & n25122 ) ;
  assign n25203 = ( n25098 & ~n25150 ) | ( n25098 & n25160 ) | ( ~n25150 & n25160 ) ;
  assign n25186 = n733 | n14540 ;
  assign n25187 = ( n548 & n616 ) | ( n548 & n25186 ) | ( n616 & n25186 ) ;
  assign n25188 = ( n548 & ~n25187 ) | ( n548 & 1'b0 ) | ( ~n25187 & 1'b0 ) ;
  assign n25189 = ( n20689 & ~n25188 ) | ( n20689 & n640 ) | ( ~n25188 & n640 ) ;
  assign n25190 = ( n640 & ~n25189 ) | ( n640 & 1'b0 ) | ( ~n25189 & 1'b0 ) ;
  assign n25191 = ( n485 & ~n785 ) | ( n485 & n25190 ) | ( ~n785 & n25190 ) ;
  assign n25192 = ~n485 & n25191 ;
  assign n25193 = ( n25147 & n25149 ) | ( n25147 & n25192 ) | ( n25149 & n25192 ) ;
  assign n25194 = ( n25147 & ~n25149 ) | ( n25147 & n25192 ) | ( ~n25149 & n25192 ) ;
  assign n25195 = ( n25149 & ~n25193 ) | ( n25149 & n25194 ) | ( ~n25193 & n25194 ) ;
  assign n25196 = n3644 | n21279 ;
  assign n25197 = ( n3652 & ~n20782 ) | ( n3652 & 1'b0 ) | ( ~n20782 & 1'b0 ) ;
  assign n25198 = n3657 &  n20777 ;
  assign n25199 = n25197 | n25198 ;
  assign n25200 = ~n3653 & n21271 ;
  assign n25201 = ( n3653 & ~n25199 ) | ( n3653 & n25200 ) | ( ~n25199 & n25200 ) ;
  assign n25202 = n25196 &  n25201 ;
  assign n25204 = ( n25195 & n25202 ) | ( n25195 & n25203 ) | ( n25202 & n25203 ) ;
  assign n25205 = ( n25195 & ~n25203 ) | ( n25195 & n25202 ) | ( ~n25203 & n25202 ) ;
  assign n25206 = ( n25203 & ~n25204 ) | ( n25203 & n25205 ) | ( ~n25204 & n25205 ) ;
  assign n25185 = ( n25123 & ~n25163 ) | ( n25123 & n25173 ) | ( ~n25163 & n25173 ) ;
  assign n25207 = ( n4478 & ~n22251 ) | ( n4478 & 1'b0 ) | ( ~n22251 & 1'b0 ) ;
  assign n25208 = ~n20747 & n22244 ;
  assign n25209 = n4482 | n22063 ;
  assign n25210 = ~n25208 & n25209 ;
  assign n25211 = ( n22251 & n25207 ) | ( n22251 & n25210 ) | ( n25207 & n25210 ) ;
  assign n25212 = ( n4430 & ~n21864 ) | ( n4430 & 1'b0 ) | ( ~n21864 & 1'b0 ) ;
  assign n25213 = ~n523 & n21475 ;
  assign n25214 = n3939 | n21675 ;
  assign n25215 = ~n25213 & n25214 ;
  assign n25216 = ( n21864 & n25212 ) | ( n21864 & n25215 ) | ( n25212 & n25215 ) ;
  assign n25217 = ~n601 & n21872 ;
  assign n25218 = ( n25216 & ~n25217 ) | ( n25216 & 1'b0 ) | ( ~n25217 & 1'b0 ) ;
  assign n25219 = x29 &  n25218 ;
  assign n25220 = x29 | n25218 ;
  assign n25221 = ~n25219 & n25220 ;
  assign n25222 = ( n25211 & ~x26 ) | ( n25211 & n25221 ) | ( ~x26 & n25221 ) ;
  assign n25223 = ( x26 & ~n25221 ) | ( x26 & n25211 ) | ( ~n25221 & n25211 ) ;
  assign n25224 = ( n25222 & ~n25211 ) | ( n25222 & n25223 ) | ( ~n25211 & n25223 ) ;
  assign n25229 = ( n25185 & n25206 ) | ( n25185 & n25224 ) | ( n25206 & n25224 ) ;
  assign n25228 = ( n25185 & ~n25206 ) | ( n25185 & n25224 ) | ( ~n25206 & n25224 ) ;
  assign n25230 = ( n25206 & ~n25229 ) | ( n25206 & n25228 ) | ( ~n25229 & n25228 ) ;
  assign n25184 = n25120 &  n25179 ;
  assign n25231 = ( n25183 & ~n25230 ) | ( n25183 & n25184 ) | ( ~n25230 & n25184 ) ;
  assign n25232 = ( n25183 & ~n25184 ) | ( n25183 & n25230 ) | ( ~n25184 & n25230 ) ;
  assign n25233 = ( n25231 & ~n25183 ) | ( n25231 & n25232 ) | ( ~n25183 & n25232 ) ;
  assign n25234 = ( n25183 & ~n25120 ) | ( n25183 & n25230 ) | ( ~n25120 & n25230 ) ;
  assign n25235 = ( n25179 & n25183 ) | ( n25179 & n25230 ) | ( n25183 & n25230 ) ;
  assign n25236 = ~n25234 & n25235 ;
  assign n25226 = n25206 &  n25224 ;
  assign n25225 = ~n25206 & n25224 ;
  assign n25227 = ( n25206 & ~n25226 ) | ( n25206 & n25225 ) | ( ~n25226 & n25225 ) ;
  assign n25237 = ( n25183 & ~n25227 ) | ( n25183 & n25185 ) | ( ~n25227 & n25185 ) ;
  assign n25238 = x26 | n25211 ;
  assign n25239 = x26 &  n25211 ;
  assign n25240 = ( n25238 & ~n25239 ) | ( n25238 & 1'b0 ) | ( ~n25239 & 1'b0 ) ;
  assign n25241 = ( n25221 & ~n25206 ) | ( n25221 & n25240 ) | ( ~n25206 & n25240 ) ;
  assign n25242 = ( n25149 & ~n25147 ) | ( n25149 & n25192 ) | ( ~n25147 & n25192 ) ;
  assign n25246 = ~n4430 & n22063 ;
  assign n25243 = n523 | n21675 ;
  assign n25244 = n3939 | n21864 ;
  assign n25245 = n25243 &  n25244 ;
  assign n25247 = ( n4430 & n25246 ) | ( n4430 & n25245 ) | ( n25246 & n25245 ) ;
  assign n25248 = n601 | n22071 ;
  assign n25249 = n25247 &  n25248 ;
  assign n25250 = ( n25202 & ~n25195 ) | ( n25202 & n25203 ) | ( ~n25195 & n25203 ) ;
  assign n25251 = ( n25249 & ~x29 ) | ( n25249 & n25250 ) | ( ~x29 & n25250 ) ;
  assign n25252 = ( x29 & ~n25249 ) | ( x29 & n25250 ) | ( ~n25249 & n25250 ) ;
  assign n25253 = ( n25251 & ~n25250 ) | ( n25251 & n25252 ) | ( ~n25250 & n25252 ) ;
  assign n25254 = n3644 | n21484 ;
  assign n25255 = n3652 &  n20777 ;
  assign n25256 = ( n3657 & ~n21271 ) | ( n3657 & 1'b0 ) | ( ~n21271 & 1'b0 ) ;
  assign n25257 = n25255 | n25256 ;
  assign n25258 = n3653 | n21475 ;
  assign n25259 = ( n25257 & ~n3653 ) | ( n25257 & n25258 ) | ( ~n3653 & n25258 ) ;
  assign n25260 = ( n25254 & ~n25259 ) | ( n25254 & 1'b0 ) | ( ~n25259 & 1'b0 ) ;
  assign n25262 = ( n25242 & n25253 ) | ( n25242 & n25260 ) | ( n25253 & n25260 ) ;
  assign n25261 = ( n25253 & ~n25242 ) | ( n25253 & n25260 ) | ( ~n25242 & n25260 ) ;
  assign n25263 = ( n25242 & ~n25262 ) | ( n25242 & n25261 ) | ( ~n25262 & n25261 ) ;
  assign n25269 = n20699 &  n22244 ;
  assign n25264 = n595 &  n699 ;
  assign n25265 = ~n237 & n25264 ;
  assign n25266 = x26 &  n25265 ;
  assign n25267 = x26 | n25265 ;
  assign n25268 = ~n25266 & n25267 ;
  assign n25270 = ( n25147 & ~n25269 ) | ( n25147 & n25268 ) | ( ~n25269 & n25268 ) ;
  assign n25271 = ( n25268 & ~n25147 ) | ( n25268 & n25269 ) | ( ~n25147 & n25269 ) ;
  assign n25272 = ( n25270 & ~n25268 ) | ( n25270 & n25271 ) | ( ~n25268 & n25271 ) ;
  assign n25273 = ( n25241 & n25263 ) | ( n25241 & n25272 ) | ( n25263 & n25272 ) ;
  assign n25274 = ( n25263 & ~n25241 ) | ( n25263 & n25272 ) | ( ~n25241 & n25272 ) ;
  assign n25275 = ( n25241 & ~n25273 ) | ( n25241 & n25274 ) | ( ~n25273 & n25274 ) ;
  assign n25276 = ( n25236 & n25237 ) | ( n25236 & n25275 ) | ( n25237 & n25275 ) ;
  assign n25277 = ( n25237 & ~n25236 ) | ( n25237 & n25275 ) | ( ~n25236 & n25275 ) ;
  assign n25278 = ( n25236 & ~n25276 ) | ( n25236 & n25277 ) | ( ~n25276 & n25277 ) ;
  assign y0 = ~n21292 ;
  assign y1 = ~n21495 ;
  assign y2 = ~n21695 ;
  assign y3 = ~n21883 ;
  assign y4 = ~n22082 ;
  assign y5 = ~n22264 ;
  assign y6 = ~n22446 ;
  assign y7 = n22620 ;
  assign y8 = n22820 ;
  assign y9 = n22971 ;
  assign y10 = n23148 ;
  assign y11 = n23309 ;
  assign y12 = n23488 ;
  assign y13 = ~n23619 ;
  assign y14 = n23752 ;
  assign y15 = n23886 ;
  assign y16 = ~n24010 ;
  assign y17 = n24123 ;
  assign y18 = n24242 ;
  assign y19 = ~n24350 ;
  assign y20 = ~n24450 ;
  assign y21 = ~n24556 ;
  assign y22 = n24649 ;
  assign y23 = n24738 ;
  assign y24 = n24822 ;
  assign y25 = ~n24907 ;
  assign y26 = ~n24981 ;
  assign y27 = ~n25053 ;
  assign y28 = n25121 ;
  assign y29 = n25182 ;
  assign y30 = n25233 ;
  assign y31 = ~n25278 ;
endmodule
