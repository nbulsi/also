module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 ;
  assign n196 = x85 | x86 ;
  assign n197 = x87 | x88 ;
  assign n198 = n196 | n197 ;
  assign n199 = x81 | x82 ;
  assign n200 = x83 | x84 ;
  assign n201 = n199 | n200 ;
  assign n202 = n198 | n201 ;
  assign n203 = x93 | x94 ;
  assign n204 = x95 | x96 ;
  assign n205 = n203 | n204 ;
  assign n206 = x89 | x90 ;
  assign n207 = x91 | x92 ;
  assign n208 = n206 | n207 ;
  assign n209 = n205 | n208 ;
  assign n210 = n202 | n209 ;
  assign n218 = x77 | x78 ;
  assign n219 = x79 | x80 ;
  assign n220 = n218 | n219 ;
  assign n221 = x73 | x74 ;
  assign n222 = x75 | x76 ;
  assign n223 = n221 | n222 ;
  assign n224 = n220 | n223 ;
  assign n211 = x69 | x70 ;
  assign n212 = x71 | x72 ;
  assign n213 = n211 | n212 ;
  assign n215 = x67 | x68 ;
  assign n214 = ( x64 & ~x66 ) | ( x64 & 1'b0 ) | ( ~x66 & 1'b0 ) ;
  assign n216 = ( n213 & ~n215 ) | ( n213 & n214 ) | ( ~n215 & n214 ) ;
  assign n217 = ~n213 & n216 ;
  assign n225 = ( n210 & ~n224 ) | ( n210 & n217 ) | ( ~n224 & n217 ) ;
  assign n226 = ~n210 & n225 ;
  assign n227 = x117 | x118 ;
  assign n228 = x119 | x120 ;
  assign n229 = n227 | n228 ;
  assign n230 = x113 | x114 ;
  assign n231 = x115 | x116 ;
  assign n232 = n230 | n231 ;
  assign n233 = n229 | n232 ;
  assign n234 = x125 | x126 ;
  assign n235 = x127 | n234 ;
  assign n236 = x121 | x122 ;
  assign n237 = x123 | x124 ;
  assign n238 = n236 | n237 ;
  assign n239 = n235 | n238 ;
  assign n240 = n233 | n239 ;
  assign n241 = x101 | x102 ;
  assign n242 = x103 | x104 ;
  assign n243 = n241 | n242 ;
  assign n244 = x97 | x98 ;
  assign n245 = x99 | x100 ;
  assign n246 = n244 | n245 ;
  assign n247 = n243 | n246 ;
  assign n248 = x109 | x110 ;
  assign n249 = x111 | x112 ;
  assign n250 = n248 | n249 ;
  assign n251 = x105 | x106 ;
  assign n252 = x107 | x108 ;
  assign n253 = n251 | n252 ;
  assign n254 = n250 | n253 ;
  assign n255 = n247 | n254 ;
  assign n256 = n240 | n255 ;
  assign n257 = ( n226 & ~n256 ) | ( n226 & 1'b0 ) | ( ~n256 & 1'b0 ) ;
  assign n130 = ~x63 & x64 ;
  assign n134 = x72 | x73 ;
  assign n135 = x74 | x75 ;
  assign n136 = n134 | n135 ;
  assign n137 = x68 | x69 ;
  assign n138 = x70 | x71 ;
  assign n139 = n137 | n138 ;
  assign n140 = n136 | n139 ;
  assign n141 = x80 | x81 ;
  assign n142 = x82 | x83 ;
  assign n143 = n141 | n142 ;
  assign n144 = x76 | x77 ;
  assign n145 = x78 | x79 ;
  assign n146 = n144 | n145 ;
  assign n147 = n143 | n146 ;
  assign n148 = n140 | n147 ;
  assign n131 = ( x64 & ~x65 ) | ( x64 & 1'b0 ) | ( ~x65 & 1'b0 ) ;
  assign n132 = x66 | x67 ;
  assign n133 = ( n131 & ~n132 ) | ( n131 & 1'b0 ) | ( ~n132 & 1'b0 ) ;
  assign n149 = ( n130 & ~n148 ) | ( n130 & n133 ) | ( ~n148 & n133 ) ;
  assign n150 = x124 | x125 ;
  assign n151 = x126 | x127 ;
  assign n152 = n150 | n151 ;
  assign n153 = x120 | x121 ;
  assign n154 = x122 | x123 ;
  assign n155 = n153 | n154 ;
  assign n156 = x116 | x117 ;
  assign n157 = x118 | x119 ;
  assign n158 = n156 | n157 ;
  assign n159 = n155 | n158 ;
  assign n160 = n152 | n159 ;
  assign n161 = x104 | x105 ;
  assign n162 = x106 | x107 ;
  assign n163 = n161 | n162 ;
  assign n164 = x100 | x101 ;
  assign n165 = x102 | x103 ;
  assign n166 = n164 | n165 ;
  assign n167 = n163 | n166 ;
  assign n168 = x112 | x113 ;
  assign n169 = x114 | x115 ;
  assign n170 = n168 | n169 ;
  assign n171 = x108 | x109 ;
  assign n172 = x110 | x111 ;
  assign n173 = n171 | n172 ;
  assign n174 = n170 | n173 ;
  assign n175 = n167 | n174 ;
  assign n176 = x88 | x89 ;
  assign n177 = x90 | x91 ;
  assign n178 = n176 | n177 ;
  assign n179 = x84 | x85 ;
  assign n180 = x86 | x87 ;
  assign n181 = n179 | n180 ;
  assign n182 = n178 | n181 ;
  assign n183 = x96 | x97 ;
  assign n184 = x98 | x99 ;
  assign n185 = n183 | n184 ;
  assign n186 = x92 | x93 ;
  assign n187 = x94 | x95 ;
  assign n188 = n186 | n187 ;
  assign n189 = n185 | n188 ;
  assign n190 = n182 | n189 ;
  assign n191 = ( n175 & ~n160 ) | ( n175 & n190 ) | ( ~n160 & n190 ) ;
  assign n192 = n160 | n191 ;
  assign n193 = n149 | n192 ;
  assign n194 = ( x63 & ~n193 ) | ( x63 & n192 ) | ( ~n193 & n192 ) ;
  assign n129 = ~x62 & x64 ;
  assign n195 = ( x65 & ~n194 ) | ( x65 & n129 ) | ( ~n194 & n129 ) ;
  assign n258 = n195 &  n257 ;
  assign n259 = ( x62 & ~n257 ) | ( x62 & n258 ) | ( ~n257 & n258 ) ;
  assign n260 = n143 | n181 ;
  assign n261 = n178 | n188 ;
  assign n262 = n260 | n261 ;
  assign n263 = n136 | n146 ;
  assign n264 = ( n129 & ~n132 ) | ( n129 & 1'b0 ) | ( ~n132 & 1'b0 ) ;
  assign n265 = ( n139 & ~n263 ) | ( n139 & n264 ) | ( ~n263 & n264 ) ;
  assign n266 = ~n139 & n265 ;
  assign n267 = ~n262 & n266 ;
  assign n268 = n158 | n170 ;
  assign n269 = n152 | n155 ;
  assign n270 = n268 | n269 ;
  assign n271 = n166 | n185 ;
  assign n272 = n163 | n173 ;
  assign n273 = n271 | n272 ;
  assign n274 = n270 | n273 ;
  assign n275 = ( n267 & ~n274 ) | ( n267 & 1'b0 ) | ( ~n274 & 1'b0 ) ;
  assign n276 = ~n195 & n275 ;
  assign n277 = n259 | n276 ;
  assign n302 = n213 | n215 ;
  assign n303 = n202 | n224 ;
  assign n304 = n302 | n303 ;
  assign n299 = ~x61 & x64 ;
  assign n305 = ( x65 & n239 ) | ( x65 & n299 ) | ( n239 & n299 ) ;
  assign n306 = n233 | n254 ;
  assign n307 = n209 | n247 ;
  assign n308 = n306 | n307 ;
  assign n309 = ( x65 & ~n308 ) | ( x65 & n299 ) | ( ~n308 & n299 ) ;
  assign n310 = ~n305 & n309 ;
  assign n311 = ~n304 & n310 ;
  assign n278 = n132 | n139 ;
  assign n279 = n263 | n278 ;
  assign n280 = ( x65 & n129 ) | ( x65 & n279 ) | ( n129 & n279 ) ;
  assign n281 = ( n262 & ~n270 ) | ( n262 & n273 ) | ( ~n270 & n273 ) ;
  assign n282 = n270 | n281 ;
  assign n283 = ( x65 & ~n282 ) | ( x65 & n129 ) | ( ~n282 & n129 ) ;
  assign n284 = ~n280 & n283 ;
  assign n285 = ~n194 & n284 ;
  assign n286 = ~n195 & n285 ;
  assign n287 = n260 | n263 ;
  assign n288 = n278 | n287 ;
  assign n289 = ( x65 & n129 ) | ( x65 & n269 ) | ( n129 & n269 ) ;
  assign n290 = n268 | n272 ;
  assign n291 = n261 | n271 ;
  assign n292 = n290 | n291 ;
  assign n293 = ( x65 & ~n292 ) | ( x65 & n129 ) | ( ~n292 & n129 ) ;
  assign n294 = ~n289 & n293 ;
  assign n295 = ~n288 & n294 ;
  assign n296 = n195 &  n295 ;
  assign n297 = ( n194 & ~n295 ) | ( n194 & n296 ) | ( ~n295 & n296 ) ;
  assign n298 = n286 | n297 ;
  assign n300 = ( x65 & ~n277 ) | ( x65 & n299 ) | ( ~n277 & n299 ) ;
  assign n301 = ( x66 & ~n298 ) | ( x66 & n300 ) | ( ~n298 & n300 ) ;
  assign n312 = n301 &  n311 ;
  assign n313 = ( n277 & ~n311 ) | ( n277 & n312 ) | ( ~n311 & n312 ) ;
  assign n314 = n224 | n302 ;
  assign n315 = ( x65 & n299 ) | ( x65 & n314 ) | ( n299 & n314 ) ;
  assign n316 = n210 | n255 ;
  assign n317 = n240 | n316 ;
  assign n318 = ( x65 & ~n317 ) | ( x65 & n299 ) | ( ~n317 & n299 ) ;
  assign n319 = ~n315 & n318 ;
  assign n320 = ( n259 & ~n276 ) | ( n259 & n319 ) | ( ~n276 & n319 ) ;
  assign n321 = ~n259 & n320 ;
  assign n322 = ~n301 & n321 ;
  assign n323 = n313 | n322 ;
  assign n324 = ( x64 & ~x67 ) | ( x64 & 1'b0 ) | ( ~x67 & 1'b0 ) ;
  assign n325 = ( n139 & ~n263 ) | ( n139 & n324 ) | ( ~n263 & n324 ) ;
  assign n326 = ~n139 & n325 ;
  assign n327 = ( n262 & ~n274 ) | ( n262 & n326 ) | ( ~n274 & n326 ) ;
  assign n328 = ~n262 & n327 ;
  assign n329 = n301 &  n328 ;
  assign n330 = ( x61 & ~n328 ) | ( x61 & n329 ) | ( ~n328 & n329 ) ;
  assign n331 = ~n215 & n299 ;
  assign n332 = ( n213 & ~n224 ) | ( n213 & n331 ) | ( ~n224 & n331 ) ;
  assign n333 = ~n213 & n332 ;
  assign n334 = ( n210 & ~n256 ) | ( n210 & n333 ) | ( ~n256 & n333 ) ;
  assign n335 = ~n210 & n334 ;
  assign n336 = ~n301 & n335 ;
  assign n337 = n330 | n336 ;
  assign n338 = ~x60 & x64 ;
  assign n339 = ( x65 & ~n337 ) | ( x65 & n338 ) | ( ~n337 & n338 ) ;
  assign n340 = ( x66 & ~n323 ) | ( x66 & n339 ) | ( ~n323 & n339 ) ;
  assign n355 = n148 | n190 ;
  assign n356 = n160 | n175 ;
  assign n357 = n355 | n356 ;
  assign n341 = ( n297 & ~n286 ) | ( n297 & n300 ) | ( ~n286 & n300 ) ;
  assign n342 = ~n297 & n341 ;
  assign n343 = ( x66 & ~n342 ) | ( x66 & n300 ) | ( ~n342 & n300 ) ;
  assign n344 = ( n256 & ~n210 ) | ( n256 & n314 ) | ( ~n210 & n314 ) ;
  assign n345 = n210 | n344 ;
  assign n346 = n301 | n345 ;
  assign n347 = n343 | n346 ;
  assign n348 = ( n298 & ~n347 ) | ( n298 & n346 ) | ( ~n347 & n346 ) ;
  assign n402 = ~x67 & n348 ;
  assign n403 = ( n340 & ~n357 ) | ( n340 & n402 ) | ( ~n357 & n402 ) ;
  assign n404 = ~n340 & n403 ;
  assign n349 = ( x67 & ~n348 ) | ( x67 & n340 ) | ( ~n348 & n340 ) ;
  assign n362 = n349 | n357 ;
  assign n405 = n348 &  n362 ;
  assign n406 = n404 | n405 ;
  assign n352 = n323 | x66 ;
  assign n350 = ( x66 & ~n322 ) | ( x66 & 1'b0 ) | ( ~n322 & 1'b0 ) ;
  assign n351 = ~n313 & n350 ;
  assign n353 = ( n352 & ~x66 ) | ( n352 & n351 ) | ( ~x66 & n351 ) ;
  assign n354 = n339 &  n353 ;
  assign n358 = ~n339 & n351 ;
  assign n359 = ( n339 & ~n357 ) | ( n339 & n358 ) | ( ~n357 & n358 ) ;
  assign n360 = ( n349 & ~n354 ) | ( n349 & n359 ) | ( ~n354 & n359 ) ;
  assign n361 = ~n349 & n360 ;
  assign n363 = ~x66 & n354 ;
  assign n364 = ( x66 & ~n362 ) | ( x66 & n363 ) | ( ~n362 & n363 ) ;
  assign n365 = ( n323 & ~n364 ) | ( n323 & 1'b0 ) | ( ~n364 & 1'b0 ) ;
  assign n366 = n361 | n365 ;
  assign n367 = n147 | n182 ;
  assign n368 = n140 | n367 ;
  assign n369 = n159 | n174 ;
  assign n370 = n167 | n189 ;
  assign n371 = n369 | n370 ;
  assign n372 = ( x65 & ~n371 ) | ( x65 & n338 ) | ( ~n371 & n338 ) ;
  assign n373 = ( x65 & n152 ) | ( x65 & n338 ) | ( n152 & n338 ) ;
  assign n374 = ( n372 & ~n373 ) | ( n372 & 1'b0 ) | ( ~n373 & 1'b0 ) ;
  assign n375 = ~n368 & n374 ;
  assign n376 = n349 &  n375 ;
  assign n377 = ( n337 & ~n375 ) | ( n337 & n376 ) | ( ~n375 & n376 ) ;
  assign n378 = ( x65 & n148 ) | ( x65 & n338 ) | ( n148 & n338 ) ;
  assign n379 = ( x65 & ~n192 ) | ( x65 & n338 ) | ( ~n192 & n338 ) ;
  assign n380 = ~n378 & n379 ;
  assign n381 = ( n330 & ~n336 ) | ( n330 & n380 ) | ( ~n336 & n380 ) ;
  assign n382 = ~n330 & n381 ;
  assign n383 = ~n349 & n382 ;
  assign n384 = n377 | n383 ;
  assign n386 = ( x64 & ~x68 ) | ( x64 & 1'b0 ) | ( ~x68 & 1'b0 ) ;
  assign n387 = ( n213 & ~n224 ) | ( n213 & n386 ) | ( ~n224 & n386 ) ;
  assign n388 = ~n213 & n387 ;
  assign n389 = ( n210 & ~n256 ) | ( n210 & n388 ) | ( ~n256 & n388 ) ;
  assign n390 = ~n210 & n389 ;
  assign n391 = n349 &  n390 ;
  assign n392 = ( x60 & ~n390 ) | ( x60 & n391 ) | ( ~n390 & n391 ) ;
  assign n393 = ~n139 & n338 ;
  assign n394 = ( n263 & ~n262 ) | ( n263 & n393 ) | ( ~n262 & n393 ) ;
  assign n395 = ~n263 & n394 ;
  assign n396 = ~n274 & n395 ;
  assign n397 = ~n349 & n396 ;
  assign n398 = n392 | n397 ;
  assign n385 = ~x59 & x64 ;
  assign n399 = ( x65 & ~n398 ) | ( x65 & n385 ) | ( ~n398 & n385 ) ;
  assign n400 = ( x66 & ~n384 ) | ( x66 & n399 ) | ( ~n384 & n399 ) ;
  assign n401 = ( x67 & ~n366 ) | ( x67 & n400 ) | ( ~n366 & n400 ) ;
  assign n407 = ( x68 & ~n406 ) | ( x68 & n401 ) | ( ~n406 & n401 ) ;
  assign n408 = ( x67 & ~n361 ) | ( x67 & 1'b0 ) | ( ~n361 & 1'b0 ) ;
  assign n409 = ~n365 & n408 ;
  assign n410 = n400 | n409 ;
  assign n411 = ~x67 & n366 ;
  assign n412 = ~x66 & n384 ;
  assign n413 = ( x66 & ~n383 ) | ( x66 & 1'b0 ) | ( ~n383 & 1'b0 ) ;
  assign n414 = ~n377 & n413 ;
  assign n415 = n399 | n414 ;
  assign n416 = ~n412 & n415 ;
  assign n417 = ( n409 & n411 ) | ( n409 & n416 ) | ( n411 & n416 ) ;
  assign n418 = n198 | n208 ;
  assign n419 = n205 | n246 ;
  assign n420 = n418 | n419 ;
  assign n421 = n213 | n223 ;
  assign n422 = n201 | n220 ;
  assign n423 = n421 | n422 ;
  assign n424 = n229 | n238 ;
  assign n425 = n235 | n424 ;
  assign n426 = n243 | n253 ;
  assign n427 = n232 | n250 ;
  assign n428 = n426 | n427 ;
  assign n429 = n425 | n428 ;
  assign n430 = ( n423 & ~n420 ) | ( n423 & n429 ) | ( ~n420 & n429 ) ;
  assign n431 = n420 | n430 ;
  assign n432 = ( n410 & n417 ) | ( n410 & n431 ) | ( n417 & n431 ) ;
  assign n433 = ( n410 & ~n432 ) | ( n410 & 1'b0 ) | ( ~n432 & 1'b0 ) ;
  assign n434 = ~n407 & n433 ;
  assign n435 = n407 | n431 ;
  assign n436 = ~x67 & n417 ;
  assign n437 = ( x67 & ~n435 ) | ( x67 & n436 ) | ( ~n435 & n436 ) ;
  assign n438 = ( n366 & ~n437 ) | ( n366 & 1'b0 ) | ( ~n437 & 1'b0 ) ;
  assign n439 = n434 | n438 ;
  assign n440 = n412 | n414 ;
  assign n441 = n399 &  n440 ;
  assign n442 = ( n415 & ~n431 ) | ( n415 & 1'b0 ) | ( ~n431 & 1'b0 ) ;
  assign n443 = ( n407 & ~n441 ) | ( n407 & n442 ) | ( ~n441 & n442 ) ;
  assign n444 = ~n407 & n443 ;
  assign n445 = ~x66 & n441 ;
  assign n446 = ( x66 & ~n435 ) | ( x66 & n445 ) | ( ~n435 & n445 ) ;
  assign n447 = ( n384 & ~n446 ) | ( n384 & 1'b0 ) | ( ~n446 & 1'b0 ) ;
  assign n448 = n444 | n447 ;
  assign n449 = n418 | n422 ;
  assign n450 = n421 | n449 ;
  assign n451 = n424 | n427 ;
  assign n452 = n419 | n426 ;
  assign n453 = n451 | n452 ;
  assign n454 = ( x65 & ~n453 ) | ( x65 & n385 ) | ( ~n453 & n385 ) ;
  assign n455 = ( x65 & n235 ) | ( x65 & n385 ) | ( n235 & n385 ) ;
  assign n456 = ( n454 & ~n455 ) | ( n454 & 1'b0 ) | ( ~n455 & 1'b0 ) ;
  assign n457 = ~n450 & n456 ;
  assign n458 = n407 &  n457 ;
  assign n459 = ( n398 & ~n457 ) | ( n398 & n458 ) | ( ~n457 & n458 ) ;
  assign n460 = ( x65 & n385 ) | ( x65 & n423 ) | ( n385 & n423 ) ;
  assign n461 = n420 | n428 ;
  assign n462 = n425 | n461 ;
  assign n463 = ( x65 & ~n462 ) | ( x65 & n385 ) | ( ~n462 & n385 ) ;
  assign n464 = ~n460 & n463 ;
  assign n465 = ( n392 & ~n397 ) | ( n392 & n464 ) | ( ~n397 & n464 ) ;
  assign n466 = ~n392 & n465 ;
  assign n467 = ~n407 & n466 ;
  assign n468 = n459 | n467 ;
  assign n469 = ( x64 & ~x69 ) | ( x64 & 1'b0 ) | ( ~x69 & 1'b0 ) ;
  assign n470 = ( n136 & ~n138 ) | ( n136 & n469 ) | ( ~n138 & n469 ) ;
  assign n471 = ~n136 & n470 ;
  assign n472 = ( n147 & ~n190 ) | ( n147 & n471 ) | ( ~n190 & n471 ) ;
  assign n473 = ~n147 & n472 ;
  assign n474 = ~n356 & n473 ;
  assign n475 = n407 &  n474 ;
  assign n476 = ( x59 & ~n474 ) | ( x59 & n475 ) | ( ~n474 & n475 ) ;
  assign n477 = ~n213 & n385 ;
  assign n478 = ( n210 & ~n224 ) | ( n210 & n477 ) | ( ~n224 & n477 ) ;
  assign n479 = ~n210 & n478 ;
  assign n480 = ~n256 & n479 ;
  assign n481 = ~n407 & n480 ;
  assign n482 = n476 | n481 ;
  assign n483 = ~x58 & x64 ;
  assign n484 = ( x65 & ~n482 ) | ( x65 & n483 ) | ( ~n482 & n483 ) ;
  assign n485 = ( x66 & ~n468 ) | ( x66 & n484 ) | ( ~n468 & n484 ) ;
  assign n486 = ( x67 & ~n448 ) | ( x67 & n485 ) | ( ~n448 & n485 ) ;
  assign n487 = ( x68 & ~n439 ) | ( x68 & n486 ) | ( ~n439 & n486 ) ;
  assign n490 = n406 | x68 ;
  assign n488 = ( x68 & ~n405 ) | ( x68 & 1'b0 ) | ( ~n405 & 1'b0 ) ;
  assign n489 = ~n404 & n488 ;
  assign n491 = ( n490 & ~x68 ) | ( n490 & n489 ) | ( ~x68 & n489 ) ;
  assign n492 = ~n411 & n491 ;
  assign n493 = n410 &  n492 ;
  assign n494 = n431 | n493 ;
  assign n495 = ~n401 & n489 ;
  assign n496 = ( n401 & ~n494 ) | ( n401 & n495 ) | ( ~n494 & n495 ) ;
  assign n497 = ~n407 & n496 ;
  assign n498 = ~x68 & n493 ;
  assign n499 = ( x68 & ~n435 ) | ( x68 & n498 ) | ( ~n435 & n498 ) ;
  assign n500 = ( n406 & ~n499 ) | ( n406 & 1'b0 ) | ( ~n499 & 1'b0 ) ;
  assign n501 = n497 | n500 ;
  assign n502 = x69 &  n501 ;
  assign n503 = x69 | n497 ;
  assign n504 = n500 | n503 ;
  assign n505 = ~n502 & n504 ;
  assign n506 = n136 | n138 ;
  assign n507 = ( n190 & ~n147 ) | ( n190 & n506 ) | ( ~n147 & n506 ) ;
  assign n508 = n147 | n507 ;
  assign n509 = n356 | n508 ;
  assign n510 = n505 | n509 ;
  assign n511 = n487 | n510 ;
  assign n512 = ~n431 & n501 ;
  assign n529 = ( n439 & ~n512 ) | ( n439 & 1'b0 ) | ( ~n512 & 1'b0 ) ;
  assign n530 = n511 &  n529 ;
  assign n513 = ( n511 & ~n512 ) | ( n511 & 1'b0 ) | ( ~n512 & 1'b0 ) ;
  assign n518 = x68 | n439 ;
  assign n519 = x68 &  n439 ;
  assign n520 = ( n518 & ~n519 ) | ( n518 & 1'b0 ) | ( ~n519 & 1'b0 ) ;
  assign n532 = ( n486 & n513 ) | ( n486 & n520 ) | ( n513 & n520 ) ;
  assign n531 = n486 | n520 ;
  assign n533 = ( n530 & ~n532 ) | ( n530 & n531 ) | ( ~n532 & n531 ) ;
  assign n521 = n431 &  n501 ;
  assign n522 = n511 &  n521 ;
  assign n524 = ( n487 & ~n512 ) | ( n487 & n505 ) | ( ~n512 & n505 ) ;
  assign n523 = n487 | n505 ;
  assign n525 = ( n522 & ~n524 ) | ( n522 & n523 ) | ( ~n524 & n523 ) ;
  assign n537 = ( n448 & ~n512 ) | ( n448 & 1'b0 ) | ( ~n512 & 1'b0 ) ;
  assign n538 = n511 &  n537 ;
  assign n526 = x67 | n448 ;
  assign n527 = x67 &  n448 ;
  assign n528 = ( n526 & ~n527 ) | ( n526 & 1'b0 ) | ( ~n527 & 1'b0 ) ;
  assign n540 = ( n485 & n513 ) | ( n485 & n528 ) | ( n513 & n528 ) ;
  assign n539 = n485 | n528 ;
  assign n541 = ( n538 & ~n540 ) | ( n538 & n539 ) | ( ~n540 & n539 ) ;
  assign n542 = ( n468 & ~n512 ) | ( n468 & 1'b0 ) | ( ~n512 & 1'b0 ) ;
  assign n543 = n511 &  n542 ;
  assign n534 = x66 | n468 ;
  assign n535 = x66 &  n468 ;
  assign n536 = ( n534 & ~n535 ) | ( n534 & 1'b0 ) | ( ~n535 & 1'b0 ) ;
  assign n544 = n484 &  n536 ;
  assign n545 = ( n484 & ~n513 ) | ( n484 & n536 ) | ( ~n513 & n536 ) ;
  assign n546 = ( n543 & ~n544 ) | ( n543 & n545 ) | ( ~n544 & n545 ) ;
  assign n547 = ( n482 & ~x65 ) | ( n482 & n483 ) | ( ~x65 & n483 ) ;
  assign n548 = ( n484 & ~n483 ) | ( n484 & n547 ) | ( ~n483 & n547 ) ;
  assign n549 = ~n513 & n548 ;
  assign n550 = ( n482 & ~n512 ) | ( n482 & 1'b0 ) | ( ~n512 & 1'b0 ) ;
  assign n551 = n511 &  n550 ;
  assign n552 = n549 | n551 ;
  assign n514 = ( x64 & ~n513 ) | ( x64 & 1'b0 ) | ( ~n513 & 1'b0 ) ;
  assign n515 = ( x58 & ~n514 ) | ( x58 & 1'b0 ) | ( ~n514 & 1'b0 ) ;
  assign n516 = ( n483 & ~n513 ) | ( n483 & 1'b0 ) | ( ~n513 & 1'b0 ) ;
  assign n517 = n515 | n516 ;
  assign n553 = ~x57 & x64 ;
  assign n554 = ( x65 & ~n517 ) | ( x65 & n553 ) | ( ~n517 & n553 ) ;
  assign n555 = ( x66 & ~n552 ) | ( x66 & n554 ) | ( ~n552 & n554 ) ;
  assign n556 = ( x67 & ~n546 ) | ( x67 & n555 ) | ( ~n546 & n555 ) ;
  assign n557 = ( x68 & ~n541 ) | ( x68 & n556 ) | ( ~n541 & n556 ) ;
  assign n558 = ( x69 & ~n533 ) | ( x69 & n557 ) | ( ~n533 & n557 ) ;
  assign n559 = ( x70 & ~n525 ) | ( x70 & n558 ) | ( ~n525 & n558 ) ;
  assign n560 = n212 | n223 ;
  assign n561 = ( n422 & ~n420 ) | ( n422 & n560 ) | ( ~n420 & n560 ) ;
  assign n562 = n420 | n561 ;
  assign n563 = n429 | n562 ;
  assign n564 = n559 | n563 ;
  assign n581 = n533 &  n564 ;
  assign n575 = x69 | n533 ;
  assign n576 = x69 &  n533 ;
  assign n577 = ( n575 & ~n576 ) | ( n575 & 1'b0 ) | ( ~n576 & 1'b0 ) ;
  assign n585 = ( n557 & n559 ) | ( n557 & n577 ) | ( n559 & n577 ) ;
  assign n586 = ( n557 & ~n563 ) | ( n557 & n577 ) | ( ~n563 & n577 ) ;
  assign n587 = ~n585 & n586 ;
  assign n588 = n581 | n587 ;
  assign n578 = x70 | n558 ;
  assign n579 = ( x70 & n558 ) | ( x70 & n563 ) | ( n558 & n563 ) ;
  assign n580 = ( n525 & ~n578 ) | ( n525 & n579 ) | ( ~n578 & n579 ) ;
  assign n589 = n541 &  n564 ;
  assign n582 = x68 | n541 ;
  assign n583 = x68 &  n541 ;
  assign n584 = ( n582 & ~n583 ) | ( n582 & 1'b0 ) | ( ~n583 & 1'b0 ) ;
  assign n593 = ( n556 & n559 ) | ( n556 & n584 ) | ( n559 & n584 ) ;
  assign n594 = ( n556 & ~n563 ) | ( n556 & n584 ) | ( ~n563 & n584 ) ;
  assign n595 = ~n593 & n594 ;
  assign n596 = n589 | n595 ;
  assign n597 = n546 &  n564 ;
  assign n590 = x67 | n546 ;
  assign n591 = x67 &  n546 ;
  assign n592 = ( n590 & ~n591 ) | ( n590 & 1'b0 ) | ( ~n591 & 1'b0 ) ;
  assign n601 = ( n555 & n559 ) | ( n555 & n592 ) | ( n559 & n592 ) ;
  assign n602 = ( n555 & ~n563 ) | ( n555 & n592 ) | ( ~n563 & n592 ) ;
  assign n603 = ~n601 & n602 ;
  assign n604 = n597 | n603 ;
  assign n605 = n552 &  n564 ;
  assign n598 = x66 | n552 ;
  assign n599 = x66 &  n552 ;
  assign n600 = ( n598 & ~n599 ) | ( n598 & 1'b0 ) | ( ~n599 & 1'b0 ) ;
  assign n606 = ( n554 & ~n559 ) | ( n554 & n600 ) | ( ~n559 & n600 ) ;
  assign n607 = ( n554 & n563 ) | ( n554 & n600 ) | ( n563 & n600 ) ;
  assign n608 = ( n606 & ~n607 ) | ( n606 & 1'b0 ) | ( ~n607 & 1'b0 ) ;
  assign n609 = n605 | n608 ;
  assign n565 = n517 &  n564 ;
  assign n566 = x65 &  n517 ;
  assign n567 = ( n515 & ~x65 ) | ( n515 & n516 ) | ( ~x65 & n516 ) ;
  assign n568 = x65 | n567 ;
  assign n569 = ( n553 & ~n566 ) | ( n553 & n568 ) | ( ~n566 & n568 ) ;
  assign n570 = ( x65 & n517 ) | ( x65 & n553 ) | ( n517 & n553 ) ;
  assign n571 = ( n563 & ~n566 ) | ( n563 & n570 ) | ( ~n566 & n570 ) ;
  assign n572 = ( n559 & n569 ) | ( n559 & n571 ) | ( n569 & n571 ) ;
  assign n573 = ( n569 & ~n572 ) | ( n569 & 1'b0 ) | ( ~n572 & 1'b0 ) ;
  assign n574 = n565 | n573 ;
  assign n610 = ( x64 & ~x71 ) | ( x64 & 1'b0 ) | ( ~x71 & 1'b0 ) ;
  assign n611 = ( n136 & ~n147 ) | ( n136 & n610 ) | ( ~n147 & n610 ) ;
  assign n612 = ~n136 & n611 ;
  assign n613 = ( n190 & ~n356 ) | ( n190 & n612 ) | ( ~n356 & n612 ) ;
  assign n614 = ~n190 & n613 ;
  assign n615 = n559 &  n614 ;
  assign n616 = ( x57 & ~n614 ) | ( x57 & n615 ) | ( ~n614 & n615 ) ;
  assign n617 = ~n212 & n553 ;
  assign n618 = ( n223 & ~n422 ) | ( n223 & n617 ) | ( ~n422 & n617 ) ;
  assign n619 = ~n223 & n618 ;
  assign n620 = ( n420 & ~n429 ) | ( n420 & n619 ) | ( ~n429 & n619 ) ;
  assign n621 = ~n420 & n620 ;
  assign n622 = ~n559 & n621 ;
  assign n623 = n616 | n622 ;
  assign n624 = ~x56 & x64 ;
  assign n625 = ( x65 & ~n623 ) | ( x65 & n624 ) | ( ~n623 & n624 ) ;
  assign n626 = ( x66 & ~n574 ) | ( x66 & n625 ) | ( ~n574 & n625 ) ;
  assign n627 = ( x67 & ~n609 ) | ( x67 & n626 ) | ( ~n609 & n626 ) ;
  assign n628 = ( x68 & ~n604 ) | ( x68 & n627 ) | ( ~n604 & n627 ) ;
  assign n629 = ( x69 & ~n596 ) | ( x69 & n628 ) | ( ~n596 & n628 ) ;
  assign n630 = ( x70 & ~n588 ) | ( x70 & n629 ) | ( ~n588 & n629 ) ;
  assign n631 = ( x71 & ~n580 ) | ( x71 & n630 ) | ( ~n580 & n630 ) ;
  assign n632 = n262 | n263 ;
  assign n633 = n274 | n632 ;
  assign n634 = n631 | n633 ;
  assign n684 = n588 &  n634 ;
  assign n688 = x70 | n588 ;
  assign n689 = x70 &  n588 ;
  assign n690 = ( n688 & ~n689 ) | ( n688 & 1'b0 ) | ( ~n689 & 1'b0 ) ;
  assign n691 = ( n629 & n631 ) | ( n629 & n690 ) | ( n631 & n690 ) ;
  assign n692 = ( n629 & ~n633 ) | ( n629 & n690 ) | ( ~n633 & n690 ) ;
  assign n693 = ~n691 & n692 ;
  assign n694 = n684 | n693 ;
  assign n695 = n596 &  n634 ;
  assign n685 = x69 | n596 ;
  assign n686 = x69 &  n596 ;
  assign n687 = ( n685 & ~n686 ) | ( n685 & 1'b0 ) | ( ~n686 & 1'b0 ) ;
  assign n699 = ( n628 & n631 ) | ( n628 & n687 ) | ( n631 & n687 ) ;
  assign n700 = ( n628 & ~n633 ) | ( n628 & n687 ) | ( ~n633 & n687 ) ;
  assign n701 = ~n699 & n700 ;
  assign n702 = n695 | n701 ;
  assign n703 = n604 &  n634 ;
  assign n696 = x68 | n604 ;
  assign n697 = x68 &  n604 ;
  assign n698 = ( n696 & ~n697 ) | ( n696 & 1'b0 ) | ( ~n697 & 1'b0 ) ;
  assign n704 = ( n627 & n631 ) | ( n627 & n698 ) | ( n631 & n698 ) ;
  assign n705 = ( n627 & ~n633 ) | ( n627 & n698 ) | ( ~n633 & n698 ) ;
  assign n706 = ~n704 & n705 ;
  assign n707 = n703 | n706 ;
  assign n673 = n609 &  n634 ;
  assign n674 = x67 | n609 ;
  assign n675 = x67 &  n609 ;
  assign n676 = ( n674 & ~n675 ) | ( n674 & 1'b0 ) | ( ~n675 & 1'b0 ) ;
  assign n677 = ( n626 & n631 ) | ( n626 & n676 ) | ( n631 & n676 ) ;
  assign n678 = ( n626 & ~n633 ) | ( n626 & n676 ) | ( ~n633 & n676 ) ;
  assign n679 = ~n677 & n678 ;
  assign n680 = n673 | n679 ;
  assign n635 = n574 &  n634 ;
  assign n640 = x66 | n574 ;
  assign n641 = x66 &  n574 ;
  assign n642 = ( n640 & ~n641 ) | ( n640 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n643 = ( n625 & n631 ) | ( n625 & n642 ) | ( n631 & n642 ) ;
  assign n644 = ( n625 & ~n633 ) | ( n625 & n642 ) | ( ~n633 & n642 ) ;
  assign n645 = ~n643 & n644 ;
  assign n646 = n635 | n645 ;
  assign n647 = n623 &  n634 ;
  assign n636 = x65 &  n623 ;
  assign n637 = x65 | n622 ;
  assign n638 = n616 | n637 ;
  assign n639 = ( n624 & ~n636 ) | ( n624 & n638 ) | ( ~n636 & n638 ) ;
  assign n648 = ( x65 & n623 ) | ( x65 & n624 ) | ( n623 & n624 ) ;
  assign n649 = ( n633 & ~n636 ) | ( n633 & n648 ) | ( ~n636 & n648 ) ;
  assign n650 = ( n631 & n639 ) | ( n631 & n649 ) | ( n639 & n649 ) ;
  assign n651 = ( n639 & ~n650 ) | ( n639 & 1'b0 ) | ( ~n650 & 1'b0 ) ;
  assign n652 = n647 | n651 ;
  assign n653 = ( x64 & ~x72 ) | ( x64 & 1'b0 ) | ( ~x72 & 1'b0 ) ;
  assign n654 = ( n223 & ~n422 ) | ( n223 & n653 ) | ( ~n422 & n653 ) ;
  assign n655 = ~n223 & n654 ;
  assign n656 = ( n420 & ~n429 ) | ( n420 & n655 ) | ( ~n429 & n655 ) ;
  assign n657 = ~n420 & n656 ;
  assign n658 = n631 &  n657 ;
  assign n659 = ( x56 & ~n657 ) | ( x56 & n658 ) | ( ~n657 & n658 ) ;
  assign n660 = ~n136 & n624 ;
  assign n661 = ( n147 & ~n190 ) | ( n147 & n660 ) | ( ~n190 & n660 ) ;
  assign n662 = ~n147 & n661 ;
  assign n663 = ~n356 & n662 ;
  assign n664 = ~n631 & n663 ;
  assign n665 = n659 | n664 ;
  assign n666 = ~x55 & x64 ;
  assign n667 = ( x65 & ~n665 ) | ( x65 & n666 ) | ( ~n665 & n666 ) ;
  assign n668 = ( x66 & ~n652 ) | ( x66 & n667 ) | ( ~n652 & n667 ) ;
  assign n672 = ( x67 & ~n646 ) | ( x67 & n668 ) | ( ~n646 & n668 ) ;
  assign n708 = ( x68 & ~n680 ) | ( x68 & n672 ) | ( ~n680 & n672 ) ;
  assign n709 = ( x69 & ~n707 ) | ( x69 & n708 ) | ( ~n707 & n708 ) ;
  assign n710 = ( x70 & ~n702 ) | ( x70 & n709 ) | ( ~n702 & n709 ) ;
  assign n711 = ( x71 & ~n694 ) | ( x71 & n710 ) | ( ~n694 & n710 ) ;
  assign n715 = n210 | n224 ;
  assign n716 = n256 | n715 ;
  assign n712 = x71 | n630 ;
  assign n713 = ( x71 & n630 ) | ( x71 & n633 ) | ( n630 & n633 ) ;
  assign n714 = ( n580 & ~n712 ) | ( n580 & n713 ) | ( ~n712 & n713 ) ;
  assign n718 = x72 &  n714 ;
  assign n717 = x72 | n714 ;
  assign n719 = ( n716 & ~n718 ) | ( n716 & n717 ) | ( ~n718 & n717 ) ;
  assign n720 = n711 | n719 ;
  assign n721 = ~n633 & n714 ;
  assign n741 = ( n694 & ~n721 ) | ( n694 & 1'b0 ) | ( ~n721 & 1'b0 ) ;
  assign n742 = n720 &  n741 ;
  assign n728 = x71 | n694 ;
  assign n729 = x71 &  n694 ;
  assign n730 = ( n728 & ~n729 ) | ( n728 & 1'b0 ) | ( ~n729 & 1'b0 ) ;
  assign n743 = n710 &  n730 ;
  assign n722 = ( n720 & ~n721 ) | ( n720 & 1'b0 ) | ( ~n721 & 1'b0 ) ;
  assign n744 = ( n710 & ~n722 ) | ( n710 & n730 ) | ( ~n722 & n730 ) ;
  assign n745 = ( n742 & ~n743 ) | ( n742 & n744 ) | ( ~n743 & n744 ) ;
  assign n731 = ( x72 & ~n714 ) | ( x72 & n711 ) | ( ~n714 & n711 ) ;
  assign n732 = ( n711 & ~x72 ) | ( n711 & n714 ) | ( ~x72 & n714 ) ;
  assign n733 = ( n731 & ~n711 ) | ( n731 & n732 ) | ( ~n711 & n732 ) ;
  assign n734 = ~n722 & n733 ;
  assign n735 = n580 &  n633 ;
  assign n736 = n720 &  n735 ;
  assign n737 = n734 | n736 ;
  assign n749 = ( n702 & ~n721 ) | ( n702 & 1'b0 ) | ( ~n721 & 1'b0 ) ;
  assign n750 = n720 &  n749 ;
  assign n738 = x70 | n702 ;
  assign n739 = x70 &  n702 ;
  assign n740 = ( n738 & ~n739 ) | ( n738 & 1'b0 ) | ( ~n739 & 1'b0 ) ;
  assign n751 = n709 &  n740 ;
  assign n752 = ( n709 & ~n722 ) | ( n709 & n740 ) | ( ~n722 & n740 ) ;
  assign n753 = ( n750 & ~n751 ) | ( n750 & n752 ) | ( ~n751 & n752 ) ;
  assign n754 = ( n707 & ~n721 ) | ( n707 & 1'b0 ) | ( ~n721 & 1'b0 ) ;
  assign n755 = n720 &  n754 ;
  assign n746 = x69 | n707 ;
  assign n747 = x69 &  n707 ;
  assign n748 = ( n746 & ~n747 ) | ( n746 & 1'b0 ) | ( ~n747 & 1'b0 ) ;
  assign n756 = n708 &  n748 ;
  assign n757 = ( n708 & ~n722 ) | ( n708 & n748 ) | ( ~n722 & n748 ) ;
  assign n758 = ( n755 & ~n756 ) | ( n755 & n757 ) | ( ~n756 & n757 ) ;
  assign n723 = ( n680 & ~n721 ) | ( n680 & 1'b0 ) | ( ~n721 & 1'b0 ) ;
  assign n724 = n720 &  n723 ;
  assign n681 = x68 | n680 ;
  assign n682 = x68 &  n680 ;
  assign n683 = ( n681 & ~n682 ) | ( n681 & 1'b0 ) | ( ~n682 & 1'b0 ) ;
  assign n726 = ( n672 & n683 ) | ( n672 & n722 ) | ( n683 & n722 ) ;
  assign n725 = n672 | n683 ;
  assign n727 = ( n724 & ~n726 ) | ( n724 & n725 ) | ( ~n726 & n725 ) ;
  assign n762 = ( n646 & ~n721 ) | ( n646 & 1'b0 ) | ( ~n721 & 1'b0 ) ;
  assign n763 = n720 &  n762 ;
  assign n669 = x67 | n646 ;
  assign n670 = x67 &  n646 ;
  assign n671 = ( n669 & ~n670 ) | ( n669 & 1'b0 ) | ( ~n670 & 1'b0 ) ;
  assign n765 = ( n668 & n671 ) | ( n668 & n722 ) | ( n671 & n722 ) ;
  assign n764 = n668 | n671 ;
  assign n766 = ( n763 & ~n765 ) | ( n763 & n764 ) | ( ~n765 & n764 ) ;
  assign n767 = ( n652 & ~n721 ) | ( n652 & 1'b0 ) | ( ~n721 & 1'b0 ) ;
  assign n768 = n720 &  n767 ;
  assign n759 = x66 | n652 ;
  assign n760 = x66 &  n652 ;
  assign n761 = ( n759 & ~n760 ) | ( n759 & 1'b0 ) | ( ~n760 & 1'b0 ) ;
  assign n770 = ( n667 & n722 ) | ( n667 & n761 ) | ( n722 & n761 ) ;
  assign n769 = n667 | n761 ;
  assign n771 = ( n768 & ~n770 ) | ( n768 & n769 ) | ( ~n770 & n769 ) ;
  assign n772 = ( n665 & ~x65 ) | ( n665 & n666 ) | ( ~x65 & n666 ) ;
  assign n773 = ( n667 & ~n666 ) | ( n667 & n772 ) | ( ~n666 & n772 ) ;
  assign n774 = ~n722 & n773 ;
  assign n775 = ( n665 & ~n721 ) | ( n665 & 1'b0 ) | ( ~n721 & 1'b0 ) ;
  assign n776 = n720 &  n775 ;
  assign n777 = n774 | n776 ;
  assign n778 = ( x64 & ~n722 ) | ( x64 & 1'b0 ) | ( ~n722 & 1'b0 ) ;
  assign n779 = ( x55 & ~n778 ) | ( x55 & 1'b0 ) | ( ~n778 & 1'b0 ) ;
  assign n780 = ( n666 & ~n722 ) | ( n666 & 1'b0 ) | ( ~n722 & 1'b0 ) ;
  assign n781 = n779 | n780 ;
  assign n782 = ~x54 & x64 ;
  assign n783 = ( x65 & ~n781 ) | ( x65 & n782 ) | ( ~n781 & n782 ) ;
  assign n784 = ( x66 & ~n777 ) | ( x66 & n783 ) | ( ~n777 & n783 ) ;
  assign n785 = ( x67 & ~n771 ) | ( x67 & n784 ) | ( ~n771 & n784 ) ;
  assign n786 = ( x68 & ~n766 ) | ( x68 & n785 ) | ( ~n766 & n785 ) ;
  assign n787 = ( x69 & ~n727 ) | ( x69 & n786 ) | ( ~n727 & n786 ) ;
  assign n788 = ( x70 & ~n758 ) | ( x70 & n787 ) | ( ~n758 & n787 ) ;
  assign n789 = ( x71 & ~n753 ) | ( x71 & n788 ) | ( ~n753 & n788 ) ;
  assign n790 = ( x72 & ~n745 ) | ( x72 & n789 ) | ( ~n745 & n789 ) ;
  assign n791 = ( x73 & ~n737 ) | ( x73 & n790 ) | ( ~n737 & n790 ) ;
  assign n792 = n135 | n146 ;
  assign n793 = ( n274 & ~n262 ) | ( n274 & n792 ) | ( ~n262 & n792 ) ;
  assign n794 = n262 | n793 ;
  assign n795 = n791 | n794 ;
  assign n813 = n745 &  n795 ;
  assign n807 = x72 | n745 ;
  assign n808 = x72 &  n745 ;
  assign n809 = ( n807 & ~n808 ) | ( n807 & 1'b0 ) | ( ~n808 & 1'b0 ) ;
  assign n817 = ( n789 & n791 ) | ( n789 & n809 ) | ( n791 & n809 ) ;
  assign n818 = ( n789 & ~n794 ) | ( n789 & n809 ) | ( ~n794 & n809 ) ;
  assign n819 = ~n817 & n818 ;
  assign n820 = n813 | n819 ;
  assign n810 = x73 | n790 ;
  assign n811 = ( x73 & n790 ) | ( x73 & n794 ) | ( n790 & n794 ) ;
  assign n812 = ( n737 & ~n810 ) | ( n737 & n811 ) | ( ~n810 & n811 ) ;
  assign n821 = n753 &  n795 ;
  assign n814 = x71 | n753 ;
  assign n815 = x71 &  n753 ;
  assign n816 = ( n814 & ~n815 ) | ( n814 & 1'b0 ) | ( ~n815 & 1'b0 ) ;
  assign n825 = ( n788 & n791 ) | ( n788 & n816 ) | ( n791 & n816 ) ;
  assign n826 = ( n788 & ~n794 ) | ( n788 & n816 ) | ( ~n794 & n816 ) ;
  assign n827 = ~n825 & n826 ;
  assign n828 = n821 | n827 ;
  assign n829 = n758 &  n795 ;
  assign n822 = x70 | n758 ;
  assign n823 = x70 &  n758 ;
  assign n824 = ( n822 & ~n823 ) | ( n822 & 1'b0 ) | ( ~n823 & 1'b0 ) ;
  assign n830 = ( n787 & n791 ) | ( n787 & n824 ) | ( n791 & n824 ) ;
  assign n831 = ( n787 & ~n794 ) | ( n787 & n824 ) | ( ~n794 & n824 ) ;
  assign n832 = ~n830 & n831 ;
  assign n833 = n829 | n832 ;
  assign n796 = n727 &  n795 ;
  assign n800 = x69 | n727 ;
  assign n801 = x69 &  n727 ;
  assign n802 = ( n800 & ~n801 ) | ( n800 & 1'b0 ) | ( ~n801 & 1'b0 ) ;
  assign n803 = ( n786 & n791 ) | ( n786 & n802 ) | ( n791 & n802 ) ;
  assign n804 = ( n786 & ~n794 ) | ( n786 & n802 ) | ( ~n794 & n802 ) ;
  assign n805 = ~n803 & n804 ;
  assign n806 = n796 | n805 ;
  assign n834 = n766 &  n795 ;
  assign n797 = x68 | n766 ;
  assign n798 = x68 &  n766 ;
  assign n799 = ( n797 & ~n798 ) | ( n797 & 1'b0 ) | ( ~n798 & 1'b0 ) ;
  assign n838 = ( n785 & n791 ) | ( n785 & n799 ) | ( n791 & n799 ) ;
  assign n839 = ( n785 & ~n794 ) | ( n785 & n799 ) | ( ~n794 & n799 ) ;
  assign n840 = ~n838 & n839 ;
  assign n841 = n834 | n840 ;
  assign n842 = n771 &  n795 ;
  assign n835 = x67 | n771 ;
  assign n836 = x67 &  n771 ;
  assign n837 = ( n835 & ~n836 ) | ( n835 & 1'b0 ) | ( ~n836 & 1'b0 ) ;
  assign n846 = ( n784 & n791 ) | ( n784 & n837 ) | ( n791 & n837 ) ;
  assign n847 = ( n784 & ~n794 ) | ( n784 & n837 ) | ( ~n794 & n837 ) ;
  assign n848 = ~n846 & n847 ;
  assign n849 = n842 | n848 ;
  assign n850 = n777 &  n795 ;
  assign n843 = x66 | n777 ;
  assign n844 = x66 &  n777 ;
  assign n845 = ( n843 & ~n844 ) | ( n843 & 1'b0 ) | ( ~n844 & 1'b0 ) ;
  assign n855 = ( n783 & n791 ) | ( n783 & n845 ) | ( n791 & n845 ) ;
  assign n856 = ( n783 & ~n794 ) | ( n783 & n845 ) | ( ~n794 & n845 ) ;
  assign n857 = ~n855 & n856 ;
  assign n858 = n850 | n857 ;
  assign n859 = n781 &  n795 ;
  assign n851 = x65 &  n781 ;
  assign n852 = ( n779 & ~x65 ) | ( n779 & n780 ) | ( ~x65 & n780 ) ;
  assign n853 = x65 | n852 ;
  assign n854 = ( n782 & ~n851 ) | ( n782 & n853 ) | ( ~n851 & n853 ) ;
  assign n860 = ( x65 & n781 ) | ( x65 & n782 ) | ( n781 & n782 ) ;
  assign n861 = ( n794 & ~n851 ) | ( n794 & n860 ) | ( ~n851 & n860 ) ;
  assign n862 = ( n791 & n854 ) | ( n791 & n861 ) | ( n854 & n861 ) ;
  assign n863 = ( n854 & ~n862 ) | ( n854 & 1'b0 ) | ( ~n862 & 1'b0 ) ;
  assign n864 = n859 | n863 ;
  assign n865 = ( x64 & ~x74 ) | ( x64 & 1'b0 ) | ( ~x74 & 1'b0 ) ;
  assign n866 = ( n220 & ~n222 ) | ( n220 & n865 ) | ( ~n222 & n865 ) ;
  assign n867 = ~n220 & n866 ;
  assign n868 = ( n210 & ~n256 ) | ( n210 & n867 ) | ( ~n256 & n867 ) ;
  assign n869 = ~n210 & n868 ;
  assign n870 = n791 &  n869 ;
  assign n871 = ( x54 & ~n869 ) | ( x54 & n870 ) | ( ~n869 & n870 ) ;
  assign n872 = ~n135 & n782 ;
  assign n873 = ( n146 & ~n262 ) | ( n146 & n872 ) | ( ~n262 & n872 ) ;
  assign n874 = ~n146 & n873 ;
  assign n875 = ~n274 & n874 ;
  assign n876 = ~n791 & n875 ;
  assign n877 = n871 | n876 ;
  assign n878 = ~x53 & x64 ;
  assign n879 = ( x65 & ~n877 ) | ( x65 & n878 ) | ( ~n877 & n878 ) ;
  assign n880 = ( x66 & ~n864 ) | ( x66 & n879 ) | ( ~n864 & n879 ) ;
  assign n881 = ( x67 & ~n858 ) | ( x67 & n880 ) | ( ~n858 & n880 ) ;
  assign n882 = ( x68 & ~n849 ) | ( x68 & n881 ) | ( ~n849 & n881 ) ;
  assign n883 = ( x69 & ~n841 ) | ( x69 & n882 ) | ( ~n841 & n882 ) ;
  assign n884 = ( x70 & ~n806 ) | ( x70 & n883 ) | ( ~n806 & n883 ) ;
  assign n885 = ( x71 & ~n833 ) | ( x71 & n884 ) | ( ~n833 & n884 ) ;
  assign n886 = ( x72 & ~n828 ) | ( x72 & n885 ) | ( ~n828 & n885 ) ;
  assign n887 = ( x73 & ~n820 ) | ( x73 & n886 ) | ( ~n820 & n886 ) ;
  assign n888 = ( x74 & ~n812 ) | ( x74 & n887 ) | ( ~n812 & n887 ) ;
  assign n889 = n220 | n222 ;
  assign n890 = ( n256 & ~n210 ) | ( n256 & n889 ) | ( ~n210 & n889 ) ;
  assign n891 = n210 | n890 ;
  assign n892 = n888 | n891 ;
  assign n977 = n820 &  n892 ;
  assign n981 = x73 | n820 ;
  assign n982 = x73 &  n820 ;
  assign n983 = ( n981 & ~n982 ) | ( n981 & 1'b0 ) | ( ~n982 & 1'b0 ) ;
  assign n984 = ( n886 & n888 ) | ( n886 & n983 ) | ( n888 & n983 ) ;
  assign n985 = ( n886 & ~n891 ) | ( n886 & n983 ) | ( ~n891 & n983 ) ;
  assign n986 = ~n984 & n985 ;
  assign n987 = n977 | n986 ;
  assign n988 = n828 &  n892 ;
  assign n978 = x72 | n828 ;
  assign n979 = x72 &  n828 ;
  assign n980 = ( n978 & ~n979 ) | ( n978 & 1'b0 ) | ( ~n979 & 1'b0 ) ;
  assign n989 = ( n885 & n888 ) | ( n885 & n980 ) | ( n888 & n980 ) ;
  assign n990 = ( n885 & ~n891 ) | ( n885 & n980 ) | ( ~n891 & n980 ) ;
  assign n991 = ~n989 & n990 ;
  assign n992 = n988 | n991 ;
  assign n966 = n833 &  n892 ;
  assign n967 = x71 | n833 ;
  assign n968 = x71 &  n833 ;
  assign n969 = ( n967 & ~n968 ) | ( n967 & 1'b0 ) | ( ~n968 & 1'b0 ) ;
  assign n970 = ( n884 & n888 ) | ( n884 & n969 ) | ( n888 & n969 ) ;
  assign n971 = ( n884 & ~n891 ) | ( n884 & n969 ) | ( ~n891 & n969 ) ;
  assign n972 = ~n970 & n971 ;
  assign n973 = n966 | n972 ;
  assign n893 = n806 &  n892 ;
  assign n897 = x70 | n806 ;
  assign n898 = x70 &  n806 ;
  assign n899 = ( n897 & ~n898 ) | ( n897 & 1'b0 ) | ( ~n898 & 1'b0 ) ;
  assign n900 = ( n883 & n888 ) | ( n883 & n899 ) | ( n888 & n899 ) ;
  assign n901 = ( n883 & ~n891 ) | ( n883 & n899 ) | ( ~n891 & n899 ) ;
  assign n902 = ~n900 & n901 ;
  assign n903 = n893 | n902 ;
  assign n904 = n841 &  n892 ;
  assign n894 = x69 | n841 ;
  assign n895 = x69 &  n841 ;
  assign n896 = ( n894 & ~n895 ) | ( n894 & 1'b0 ) | ( ~n895 & 1'b0 ) ;
  assign n908 = ( n882 & n888 ) | ( n882 & n896 ) | ( n888 & n896 ) ;
  assign n909 = ( n882 & ~n891 ) | ( n882 & n896 ) | ( ~n891 & n896 ) ;
  assign n910 = ~n908 & n909 ;
  assign n911 = n904 | n910 ;
  assign n912 = n849 &  n892 ;
  assign n905 = x68 | n849 ;
  assign n906 = x68 &  n849 ;
  assign n907 = ( n905 & ~n906 ) | ( n905 & 1'b0 ) | ( ~n906 & 1'b0 ) ;
  assign n916 = ( n881 & n888 ) | ( n881 & n907 ) | ( n888 & n907 ) ;
  assign n917 = ( n881 & ~n891 ) | ( n881 & n907 ) | ( ~n891 & n907 ) ;
  assign n918 = ~n916 & n917 ;
  assign n919 = n912 | n918 ;
  assign n920 = n858 &  n892 ;
  assign n913 = x67 | n858 ;
  assign n914 = x67 &  n858 ;
  assign n915 = ( n913 & ~n914 ) | ( n913 & 1'b0 ) | ( ~n914 & 1'b0 ) ;
  assign n924 = ( n880 & n888 ) | ( n880 & n915 ) | ( n888 & n915 ) ;
  assign n925 = ( n880 & ~n891 ) | ( n880 & n915 ) | ( ~n891 & n915 ) ;
  assign n926 = ~n924 & n925 ;
  assign n927 = n920 | n926 ;
  assign n928 = n864 &  n892 ;
  assign n921 = x66 | n864 ;
  assign n922 = x66 &  n864 ;
  assign n923 = ( n921 & ~n922 ) | ( n921 & 1'b0 ) | ( ~n922 & 1'b0 ) ;
  assign n933 = ( n879 & ~n888 ) | ( n879 & n923 ) | ( ~n888 & n923 ) ;
  assign n934 = ( n879 & n891 ) | ( n879 & n923 ) | ( n891 & n923 ) ;
  assign n935 = ( n933 & ~n934 ) | ( n933 & 1'b0 ) | ( ~n934 & 1'b0 ) ;
  assign n936 = n928 | n935 ;
  assign n937 = n877 &  n892 ;
  assign n929 = x65 &  n877 ;
  assign n930 = x65 | n876 ;
  assign n931 = n871 | n930 ;
  assign n932 = ( n878 & ~n929 ) | ( n878 & n931 ) | ( ~n929 & n931 ) ;
  assign n938 = ( x65 & n877 ) | ( x65 & n878 ) | ( n877 & n878 ) ;
  assign n939 = ( n891 & ~n929 ) | ( n891 & n938 ) | ( ~n929 & n938 ) ;
  assign n940 = ( n888 & n932 ) | ( n888 & n939 ) | ( n932 & n939 ) ;
  assign n941 = ( n932 & ~n940 ) | ( n932 & 1'b0 ) | ( ~n940 & 1'b0 ) ;
  assign n942 = n937 | n941 ;
  assign n943 = ( x64 & ~x75 ) | ( x64 & 1'b0 ) | ( ~x75 & 1'b0 ) ;
  assign n944 = ( n146 & ~n262 ) | ( n146 & n943 ) | ( ~n262 & n943 ) ;
  assign n945 = ~n146 & n944 ;
  assign n946 = ~n274 & n945 ;
  assign n947 = n888 &  n946 ;
  assign n948 = ( x53 & ~n946 ) | ( x53 & n947 ) | ( ~n946 & n947 ) ;
  assign n949 = ~n222 & n878 ;
  assign n950 = ( n210 & ~n220 ) | ( n210 & n949 ) | ( ~n220 & n949 ) ;
  assign n951 = ~n210 & n950 ;
  assign n952 = ~n256 & n951 ;
  assign n953 = ~n888 & n952 ;
  assign n954 = n948 | n953 ;
  assign n955 = ~x52 & x64 ;
  assign n956 = ( x65 & ~n954 ) | ( x65 & n955 ) | ( ~n954 & n955 ) ;
  assign n957 = ( x66 & ~n942 ) | ( x66 & n956 ) | ( ~n942 & n956 ) ;
  assign n958 = ( x67 & ~n936 ) | ( x67 & n957 ) | ( ~n936 & n957 ) ;
  assign n959 = ( x68 & ~n927 ) | ( x68 & n958 ) | ( ~n927 & n958 ) ;
  assign n960 = ( x69 & ~n919 ) | ( x69 & n959 ) | ( ~n919 & n959 ) ;
  assign n961 = ( x70 & ~n911 ) | ( x70 & n960 ) | ( ~n911 & n960 ) ;
  assign n965 = ( x71 & ~n903 ) | ( x71 & n961 ) | ( ~n903 & n961 ) ;
  assign n993 = ( x72 & ~n973 ) | ( x72 & n965 ) | ( ~n973 & n965 ) ;
  assign n994 = ( x73 & ~n992 ) | ( x73 & n993 ) | ( ~n992 & n993 ) ;
  assign n995 = ( x74 & ~n987 ) | ( x74 & n994 ) | ( ~n987 & n994 ) ;
  assign n999 = n147 | n190 ;
  assign n1000 = n356 | n999 ;
  assign n996 = x74 | n887 ;
  assign n997 = ( x74 & n887 ) | ( x74 & n891 ) | ( n887 & n891 ) ;
  assign n998 = ( n812 & ~n996 ) | ( n812 & n997 ) | ( ~n996 & n997 ) ;
  assign n1002 = x75 &  n998 ;
  assign n1001 = x75 | n998 ;
  assign n1003 = ( n1000 & ~n1002 ) | ( n1000 & n1001 ) | ( ~n1002 & n1001 ) ;
  assign n1004 = n995 | n1003 ;
  assign n1005 = ~n891 & n998 ;
  assign n1025 = ( n987 & ~n1005 ) | ( n987 & 1'b0 ) | ( ~n1005 & 1'b0 ) ;
  assign n1026 = n1004 &  n1025 ;
  assign n1012 = x74 | n987 ;
  assign n1013 = x74 &  n987 ;
  assign n1014 = ( n1012 & ~n1013 ) | ( n1012 & 1'b0 ) | ( ~n1013 & 1'b0 ) ;
  assign n1027 = n994 &  n1014 ;
  assign n1006 = ( n1004 & ~n1005 ) | ( n1004 & 1'b0 ) | ( ~n1005 & 1'b0 ) ;
  assign n1028 = ( n994 & ~n1006 ) | ( n994 & n1014 ) | ( ~n1006 & n1014 ) ;
  assign n1029 = ( n1026 & ~n1027 ) | ( n1026 & n1028 ) | ( ~n1027 & n1028 ) ;
  assign n1016 = ( x75 & n995 ) | ( x75 & n998 ) | ( n995 & n998 ) ;
  assign n1015 = ( x75 & ~n995 ) | ( x75 & n998 ) | ( ~n995 & n998 ) ;
  assign n1017 = ( n995 & ~n1016 ) | ( n995 & n1015 ) | ( ~n1016 & n1015 ) ;
  assign n1018 = ~n1006 & n1017 ;
  assign n1019 = n812 &  n891 ;
  assign n1020 = n1004 &  n1019 ;
  assign n1021 = n1018 | n1020 ;
  assign n1030 = ( n992 & ~n1005 ) | ( n992 & 1'b0 ) | ( ~n1005 & 1'b0 ) ;
  assign n1031 = n1004 &  n1030 ;
  assign n1022 = x73 | n992 ;
  assign n1023 = x73 &  n992 ;
  assign n1024 = ( n1022 & ~n1023 ) | ( n1022 & 1'b0 ) | ( ~n1023 & 1'b0 ) ;
  assign n1032 = n993 &  n1024 ;
  assign n1033 = ( n993 & ~n1006 ) | ( n993 & n1024 ) | ( ~n1006 & n1024 ) ;
  assign n1034 = ( n1031 & ~n1032 ) | ( n1031 & n1033 ) | ( ~n1032 & n1033 ) ;
  assign n1007 = ( n973 & ~n1005 ) | ( n973 & 1'b0 ) | ( ~n1005 & 1'b0 ) ;
  assign n1008 = n1004 &  n1007 ;
  assign n974 = x72 | n973 ;
  assign n975 = x72 &  n973 ;
  assign n976 = ( n974 & ~n975 ) | ( n974 & 1'b0 ) | ( ~n975 & 1'b0 ) ;
  assign n1009 = n965 &  n976 ;
  assign n1010 = ( n965 & ~n1006 ) | ( n965 & n976 ) | ( ~n1006 & n976 ) ;
  assign n1011 = ( n1008 & ~n1009 ) | ( n1008 & n1010 ) | ( ~n1009 & n1010 ) ;
  assign n1038 = ( n903 & ~n1005 ) | ( n903 & 1'b0 ) | ( ~n1005 & 1'b0 ) ;
  assign n1039 = n1004 &  n1038 ;
  assign n962 = x71 | n903 ;
  assign n963 = x71 &  n903 ;
  assign n964 = ( n962 & ~n963 ) | ( n962 & 1'b0 ) | ( ~n963 & 1'b0 ) ;
  assign n1041 = ( n961 & n964 ) | ( n961 & n1006 ) | ( n964 & n1006 ) ;
  assign n1040 = n961 | n964 ;
  assign n1042 = ( n1039 & ~n1041 ) | ( n1039 & n1040 ) | ( ~n1041 & n1040 ) ;
  assign n1046 = ( n911 & ~n1005 ) | ( n911 & 1'b0 ) | ( ~n1005 & 1'b0 ) ;
  assign n1047 = n1004 &  n1046 ;
  assign n1035 = x70 | n911 ;
  assign n1036 = x70 &  n911 ;
  assign n1037 = ( n1035 & ~n1036 ) | ( n1035 & 1'b0 ) | ( ~n1036 & 1'b0 ) ;
  assign n1048 = n960 &  n1037 ;
  assign n1049 = ( n960 & ~n1006 ) | ( n960 & n1037 ) | ( ~n1006 & n1037 ) ;
  assign n1050 = ( n1047 & ~n1048 ) | ( n1047 & n1049 ) | ( ~n1048 & n1049 ) ;
  assign n1054 = ( n919 & ~n1005 ) | ( n919 & 1'b0 ) | ( ~n1005 & 1'b0 ) ;
  assign n1055 = n1004 &  n1054 ;
  assign n1043 = x69 | n919 ;
  assign n1044 = x69 &  n919 ;
  assign n1045 = ( n1043 & ~n1044 ) | ( n1043 & 1'b0 ) | ( ~n1044 & 1'b0 ) ;
  assign n1057 = ( n959 & n1006 ) | ( n959 & n1045 ) | ( n1006 & n1045 ) ;
  assign n1056 = n959 | n1045 ;
  assign n1058 = ( n1055 & ~n1057 ) | ( n1055 & n1056 ) | ( ~n1057 & n1056 ) ;
  assign n1062 = ( n927 & ~n1005 ) | ( n927 & 1'b0 ) | ( ~n1005 & 1'b0 ) ;
  assign n1063 = n1004 &  n1062 ;
  assign n1051 = x68 | n927 ;
  assign n1052 = x68 &  n927 ;
  assign n1053 = ( n1051 & ~n1052 ) | ( n1051 & 1'b0 ) | ( ~n1052 & 1'b0 ) ;
  assign n1065 = ( n958 & n1006 ) | ( n958 & n1053 ) | ( n1006 & n1053 ) ;
  assign n1064 = n958 | n1053 ;
  assign n1066 = ( n1063 & ~n1065 ) | ( n1063 & n1064 ) | ( ~n1065 & n1064 ) ;
  assign n1070 = ( n936 & ~n1005 ) | ( n936 & 1'b0 ) | ( ~n1005 & 1'b0 ) ;
  assign n1071 = n1004 &  n1070 ;
  assign n1059 = x67 | n936 ;
  assign n1060 = x67 &  n936 ;
  assign n1061 = ( n1059 & ~n1060 ) | ( n1059 & 1'b0 ) | ( ~n1060 & 1'b0 ) ;
  assign n1073 = ( n957 & n1006 ) | ( n957 & n1061 ) | ( n1006 & n1061 ) ;
  assign n1072 = n957 | n1061 ;
  assign n1074 = ( n1071 & ~n1073 ) | ( n1071 & n1072 ) | ( ~n1073 & n1072 ) ;
  assign n1075 = ( n942 & ~n1005 ) | ( n942 & 1'b0 ) | ( ~n1005 & 1'b0 ) ;
  assign n1076 = n1004 &  n1075 ;
  assign n1067 = x66 | n942 ;
  assign n1068 = x66 &  n942 ;
  assign n1069 = ( n1067 & ~n1068 ) | ( n1067 & 1'b0 ) | ( ~n1068 & 1'b0 ) ;
  assign n1077 = n956 &  n1069 ;
  assign n1078 = ( n956 & ~n1006 ) | ( n956 & n1069 ) | ( ~n1006 & n1069 ) ;
  assign n1079 = ( n1076 & ~n1077 ) | ( n1076 & n1078 ) | ( ~n1077 & n1078 ) ;
  assign n1080 = ( n954 & ~x65 ) | ( n954 & n955 ) | ( ~x65 & n955 ) ;
  assign n1081 = ( n956 & ~n955 ) | ( n956 & n1080 ) | ( ~n955 & n1080 ) ;
  assign n1082 = ~n1006 & n1081 ;
  assign n1083 = ( n954 & ~n1005 ) | ( n954 & 1'b0 ) | ( ~n1005 & 1'b0 ) ;
  assign n1084 = n1004 &  n1083 ;
  assign n1085 = n1082 | n1084 ;
  assign n1086 = ( x64 & ~n1006 ) | ( x64 & 1'b0 ) | ( ~n1006 & 1'b0 ) ;
  assign n1087 = ( x52 & ~n1086 ) | ( x52 & 1'b0 ) | ( ~n1086 & 1'b0 ) ;
  assign n1088 = ( n955 & ~n1006 ) | ( n955 & 1'b0 ) | ( ~n1006 & 1'b0 ) ;
  assign n1089 = n1087 | n1088 ;
  assign n1090 = ~x51 & x64 ;
  assign n1091 = ( x65 & ~n1089 ) | ( x65 & n1090 ) | ( ~n1089 & n1090 ) ;
  assign n1092 = ( x66 & ~n1085 ) | ( x66 & n1091 ) | ( ~n1085 & n1091 ) ;
  assign n1093 = ( x67 & ~n1079 ) | ( x67 & n1092 ) | ( ~n1079 & n1092 ) ;
  assign n1094 = ( x68 & ~n1074 ) | ( x68 & n1093 ) | ( ~n1074 & n1093 ) ;
  assign n1095 = ( x69 & ~n1066 ) | ( x69 & n1094 ) | ( ~n1066 & n1094 ) ;
  assign n1096 = ( x70 & ~n1058 ) | ( x70 & n1095 ) | ( ~n1058 & n1095 ) ;
  assign n1097 = ( x71 & ~n1050 ) | ( x71 & n1096 ) | ( ~n1050 & n1096 ) ;
  assign n1098 = ( x72 & ~n1042 ) | ( x72 & n1097 ) | ( ~n1042 & n1097 ) ;
  assign n1099 = ( x73 & ~n1011 ) | ( x73 & n1098 ) | ( ~n1011 & n1098 ) ;
  assign n1100 = ( x74 & ~n1034 ) | ( x74 & n1099 ) | ( ~n1034 & n1099 ) ;
  assign n1101 = ( x75 & ~n1029 ) | ( x75 & n1100 ) | ( ~n1029 & n1100 ) ;
  assign n1102 = ( x76 & ~n1021 ) | ( x76 & n1101 ) | ( ~n1021 & n1101 ) ;
  assign n1103 = n420 | n422 ;
  assign n1104 = n429 | n1103 ;
  assign n1105 = n1102 | n1104 ;
  assign n1123 = n1029 &  n1105 ;
  assign n1117 = x75 | n1029 ;
  assign n1118 = x75 &  n1029 ;
  assign n1119 = ( n1117 & ~n1118 ) | ( n1117 & 1'b0 ) | ( ~n1118 & 1'b0 ) ;
  assign n1127 = ( n1100 & n1102 ) | ( n1100 & n1119 ) | ( n1102 & n1119 ) ;
  assign n1128 = ( n1100 & ~n1104 ) | ( n1100 & n1119 ) | ( ~n1104 & n1119 ) ;
  assign n1129 = ~n1127 & n1128 ;
  assign n1130 = n1123 | n1129 ;
  assign n1120 = x76 | n1101 ;
  assign n1121 = ( x76 & n1101 ) | ( x76 & n1104 ) | ( n1101 & n1104 ) ;
  assign n1122 = ( n1021 & ~n1120 ) | ( n1021 & n1121 ) | ( ~n1120 & n1121 ) ;
  assign n1131 = n1034 &  n1105 ;
  assign n1124 = x74 | n1034 ;
  assign n1125 = x74 &  n1034 ;
  assign n1126 = ( n1124 & ~n1125 ) | ( n1124 & 1'b0 ) | ( ~n1125 & 1'b0 ) ;
  assign n1132 = ( n1099 & n1102 ) | ( n1099 & n1126 ) | ( n1102 & n1126 ) ;
  assign n1133 = ( n1099 & ~n1104 ) | ( n1099 & n1126 ) | ( ~n1104 & n1126 ) ;
  assign n1134 = ~n1132 & n1133 ;
  assign n1135 = n1131 | n1134 ;
  assign n1106 = n1011 &  n1105 ;
  assign n1110 = x73 | n1011 ;
  assign n1111 = x73 &  n1011 ;
  assign n1112 = ( n1110 & ~n1111 ) | ( n1110 & 1'b0 ) | ( ~n1111 & 1'b0 ) ;
  assign n1113 = ( n1098 & n1102 ) | ( n1098 & n1112 ) | ( n1102 & n1112 ) ;
  assign n1114 = ( n1098 & ~n1104 ) | ( n1098 & n1112 ) | ( ~n1104 & n1112 ) ;
  assign n1115 = ~n1113 & n1114 ;
  assign n1116 = n1106 | n1115 ;
  assign n1136 = n1042 &  n1105 ;
  assign n1107 = x72 | n1042 ;
  assign n1108 = x72 &  n1042 ;
  assign n1109 = ( n1107 & ~n1108 ) | ( n1107 & 1'b0 ) | ( ~n1108 & 1'b0 ) ;
  assign n1140 = ( n1097 & n1102 ) | ( n1097 & n1109 ) | ( n1102 & n1109 ) ;
  assign n1141 = ( n1097 & ~n1104 ) | ( n1097 & n1109 ) | ( ~n1104 & n1109 ) ;
  assign n1142 = ~n1140 & n1141 ;
  assign n1143 = n1136 | n1142 ;
  assign n1144 = n1050 &  n1105 ;
  assign n1137 = x71 | n1050 ;
  assign n1138 = x71 &  n1050 ;
  assign n1139 = ( n1137 & ~n1138 ) | ( n1137 & 1'b0 ) | ( ~n1138 & 1'b0 ) ;
  assign n1148 = ( n1096 & n1102 ) | ( n1096 & n1139 ) | ( n1102 & n1139 ) ;
  assign n1149 = ( n1096 & ~n1104 ) | ( n1096 & n1139 ) | ( ~n1104 & n1139 ) ;
  assign n1150 = ~n1148 & n1149 ;
  assign n1151 = n1144 | n1150 ;
  assign n1152 = n1058 &  n1105 ;
  assign n1145 = x70 | n1058 ;
  assign n1146 = x70 &  n1058 ;
  assign n1147 = ( n1145 & ~n1146 ) | ( n1145 & 1'b0 ) | ( ~n1146 & 1'b0 ) ;
  assign n1156 = ( n1095 & n1102 ) | ( n1095 & n1147 ) | ( n1102 & n1147 ) ;
  assign n1157 = ( n1095 & ~n1104 ) | ( n1095 & n1147 ) | ( ~n1104 & n1147 ) ;
  assign n1158 = ~n1156 & n1157 ;
  assign n1159 = n1152 | n1158 ;
  assign n1160 = n1066 &  n1105 ;
  assign n1153 = x69 | n1066 ;
  assign n1154 = x69 &  n1066 ;
  assign n1155 = ( n1153 & ~n1154 ) | ( n1153 & 1'b0 ) | ( ~n1154 & 1'b0 ) ;
  assign n1164 = ( n1094 & n1102 ) | ( n1094 & n1155 ) | ( n1102 & n1155 ) ;
  assign n1165 = ( n1094 & ~n1104 ) | ( n1094 & n1155 ) | ( ~n1104 & n1155 ) ;
  assign n1166 = ~n1164 & n1165 ;
  assign n1167 = n1160 | n1166 ;
  assign n1168 = n1074 &  n1105 ;
  assign n1161 = x68 | n1074 ;
  assign n1162 = x68 &  n1074 ;
  assign n1163 = ( n1161 & ~n1162 ) | ( n1161 & 1'b0 ) | ( ~n1162 & 1'b0 ) ;
  assign n1172 = ( n1093 & n1102 ) | ( n1093 & n1163 ) | ( n1102 & n1163 ) ;
  assign n1173 = ( n1093 & ~n1104 ) | ( n1093 & n1163 ) | ( ~n1104 & n1163 ) ;
  assign n1174 = ~n1172 & n1173 ;
  assign n1175 = n1168 | n1174 ;
  assign n1176 = n1079 &  n1105 ;
  assign n1169 = x67 | n1079 ;
  assign n1170 = x67 &  n1079 ;
  assign n1171 = ( n1169 & ~n1170 ) | ( n1169 & 1'b0 ) | ( ~n1170 & 1'b0 ) ;
  assign n1180 = ( n1092 & n1102 ) | ( n1092 & n1171 ) | ( n1102 & n1171 ) ;
  assign n1181 = ( n1092 & ~n1104 ) | ( n1092 & n1171 ) | ( ~n1104 & n1171 ) ;
  assign n1182 = ~n1180 & n1181 ;
  assign n1183 = n1176 | n1182 ;
  assign n1184 = n1085 &  n1105 ;
  assign n1177 = x66 | n1085 ;
  assign n1178 = x66 &  n1085 ;
  assign n1179 = ( n1177 & ~n1178 ) | ( n1177 & 1'b0 ) | ( ~n1178 & 1'b0 ) ;
  assign n1189 = ( n1091 & ~n1102 ) | ( n1091 & n1179 ) | ( ~n1102 & n1179 ) ;
  assign n1190 = ( n1091 & n1104 ) | ( n1091 & n1179 ) | ( n1104 & n1179 ) ;
  assign n1191 = ( n1189 & ~n1190 ) | ( n1189 & 1'b0 ) | ( ~n1190 & 1'b0 ) ;
  assign n1192 = n1184 | n1191 ;
  assign n1193 = n1089 &  n1105 ;
  assign n1185 = x65 &  n1089 ;
  assign n1186 = ( n1087 & ~x65 ) | ( n1087 & n1088 ) | ( ~x65 & n1088 ) ;
  assign n1187 = x65 | n1186 ;
  assign n1188 = ( n1090 & ~n1185 ) | ( n1090 & n1187 ) | ( ~n1185 & n1187 ) ;
  assign n1194 = ( x65 & n1089 ) | ( x65 & n1090 ) | ( n1089 & n1090 ) ;
  assign n1195 = ( n1104 & ~n1185 ) | ( n1104 & n1194 ) | ( ~n1185 & n1194 ) ;
  assign n1196 = ( n1102 & n1188 ) | ( n1102 & n1195 ) | ( n1188 & n1195 ) ;
  assign n1197 = ( n1188 & ~n1196 ) | ( n1188 & 1'b0 ) | ( ~n1196 & 1'b0 ) ;
  assign n1198 = n1193 | n1197 ;
  assign n1199 = ( x64 & ~x77 ) | ( x64 & 1'b0 ) | ( ~x77 & 1'b0 ) ;
  assign n1200 = ( n143 & ~n145 ) | ( n143 & n1199 ) | ( ~n145 & n1199 ) ;
  assign n1201 = ~n143 & n1200 ;
  assign n1202 = ( n190 & ~n356 ) | ( n190 & n1201 ) | ( ~n356 & n1201 ) ;
  assign n1203 = ~n190 & n1202 ;
  assign n1204 = n1102 &  n1203 ;
  assign n1205 = ( x51 & ~n1203 ) | ( x51 & n1204 ) | ( ~n1203 & n1204 ) ;
  assign n1206 = ~n220 & n1090 ;
  assign n1207 = ( n210 & ~n256 ) | ( n210 & n1206 ) | ( ~n256 & n1206 ) ;
  assign n1208 = ~n210 & n1207 ;
  assign n1209 = ~n1102 & n1208 ;
  assign n1210 = n1205 | n1209 ;
  assign n1211 = ~x50 & x64 ;
  assign n1212 = ( x65 & ~n1210 ) | ( x65 & n1211 ) | ( ~n1210 & n1211 ) ;
  assign n1213 = ( x66 & ~n1198 ) | ( x66 & n1212 ) | ( ~n1198 & n1212 ) ;
  assign n1214 = ( x67 & ~n1192 ) | ( x67 & n1213 ) | ( ~n1192 & n1213 ) ;
  assign n1215 = ( x68 & ~n1183 ) | ( x68 & n1214 ) | ( ~n1183 & n1214 ) ;
  assign n1216 = ( x69 & ~n1175 ) | ( x69 & n1215 ) | ( ~n1175 & n1215 ) ;
  assign n1217 = ( x70 & ~n1167 ) | ( x70 & n1216 ) | ( ~n1167 & n1216 ) ;
  assign n1218 = ( x71 & ~n1159 ) | ( x71 & n1217 ) | ( ~n1159 & n1217 ) ;
  assign n1219 = ( x72 & ~n1151 ) | ( x72 & n1218 ) | ( ~n1151 & n1218 ) ;
  assign n1220 = ( x73 & ~n1143 ) | ( x73 & n1219 ) | ( ~n1143 & n1219 ) ;
  assign n1221 = ( x74 & ~n1116 ) | ( x74 & n1220 ) | ( ~n1116 & n1220 ) ;
  assign n1222 = ( x75 & ~n1135 ) | ( x75 & n1221 ) | ( ~n1135 & n1221 ) ;
  assign n1223 = ( x76 & ~n1130 ) | ( x76 & n1222 ) | ( ~n1130 & n1222 ) ;
  assign n1224 = ( x77 & ~n1122 ) | ( x77 & n1223 ) | ( ~n1122 & n1223 ) ;
  assign n1225 = n143 | n145 ;
  assign n1226 = ( n356 & ~n190 ) | ( n356 & n1225 ) | ( ~n190 & n1225 ) ;
  assign n1227 = n190 | n1226 ;
  assign n1228 = n1224 | n1227 ;
  assign n1350 = n1130 &  n1228 ;
  assign n1351 = x76 | n1130 ;
  assign n1352 = x76 &  n1130 ;
  assign n1353 = ( n1351 & ~n1352 ) | ( n1351 & 1'b0 ) | ( ~n1352 & 1'b0 ) ;
  assign n1354 = ( n1222 & n1224 ) | ( n1222 & n1353 ) | ( n1224 & n1353 ) ;
  assign n1355 = ( n1222 & ~n1227 ) | ( n1222 & n1353 ) | ( ~n1227 & n1353 ) ;
  assign n1356 = ~n1354 & n1355 ;
  assign n1357 = n1350 | n1356 ;
  assign n1339 = n1135 &  n1228 ;
  assign n1340 = x75 | n1135 ;
  assign n1341 = x75 &  n1135 ;
  assign n1342 = ( n1340 & ~n1341 ) | ( n1340 & 1'b0 ) | ( ~n1341 & 1'b0 ) ;
  assign n1343 = ( n1221 & n1224 ) | ( n1221 & n1342 ) | ( n1224 & n1342 ) ;
  assign n1344 = ( n1221 & ~n1227 ) | ( n1221 & n1342 ) | ( ~n1227 & n1342 ) ;
  assign n1345 = ~n1343 & n1344 ;
  assign n1346 = n1339 | n1345 ;
  assign n1229 = n1116 &  n1228 ;
  assign n1233 = x74 | n1116 ;
  assign n1234 = x74 &  n1116 ;
  assign n1235 = ( n1233 & ~n1234 ) | ( n1233 & 1'b0 ) | ( ~n1234 & 1'b0 ) ;
  assign n1236 = ( n1220 & n1224 ) | ( n1220 & n1235 ) | ( n1224 & n1235 ) ;
  assign n1237 = ( n1220 & ~n1227 ) | ( n1220 & n1235 ) | ( ~n1227 & n1235 ) ;
  assign n1238 = ~n1236 & n1237 ;
  assign n1239 = n1229 | n1238 ;
  assign n1240 = n1143 &  n1228 ;
  assign n1230 = x73 | n1143 ;
  assign n1231 = x73 &  n1143 ;
  assign n1232 = ( n1230 & ~n1231 ) | ( n1230 & 1'b0 ) | ( ~n1231 & 1'b0 ) ;
  assign n1244 = ( n1219 & n1224 ) | ( n1219 & n1232 ) | ( n1224 & n1232 ) ;
  assign n1245 = ( n1219 & ~n1227 ) | ( n1219 & n1232 ) | ( ~n1227 & n1232 ) ;
  assign n1246 = ~n1244 & n1245 ;
  assign n1247 = n1240 | n1246 ;
  assign n1248 = n1151 &  n1228 ;
  assign n1241 = x72 | n1151 ;
  assign n1242 = x72 &  n1151 ;
  assign n1243 = ( n1241 & ~n1242 ) | ( n1241 & 1'b0 ) | ( ~n1242 & 1'b0 ) ;
  assign n1252 = ( n1218 & n1224 ) | ( n1218 & n1243 ) | ( n1224 & n1243 ) ;
  assign n1253 = ( n1218 & ~n1227 ) | ( n1218 & n1243 ) | ( ~n1227 & n1243 ) ;
  assign n1254 = ~n1252 & n1253 ;
  assign n1255 = n1248 | n1254 ;
  assign n1256 = n1159 &  n1228 ;
  assign n1249 = x71 | n1159 ;
  assign n1250 = x71 &  n1159 ;
  assign n1251 = ( n1249 & ~n1250 ) | ( n1249 & 1'b0 ) | ( ~n1250 & 1'b0 ) ;
  assign n1260 = ( n1217 & n1224 ) | ( n1217 & n1251 ) | ( n1224 & n1251 ) ;
  assign n1261 = ( n1217 & ~n1227 ) | ( n1217 & n1251 ) | ( ~n1227 & n1251 ) ;
  assign n1262 = ~n1260 & n1261 ;
  assign n1263 = n1256 | n1262 ;
  assign n1264 = n1167 &  n1228 ;
  assign n1257 = x70 | n1167 ;
  assign n1258 = x70 &  n1167 ;
  assign n1259 = ( n1257 & ~n1258 ) | ( n1257 & 1'b0 ) | ( ~n1258 & 1'b0 ) ;
  assign n1268 = ( n1216 & n1224 ) | ( n1216 & n1259 ) | ( n1224 & n1259 ) ;
  assign n1269 = ( n1216 & ~n1227 ) | ( n1216 & n1259 ) | ( ~n1227 & n1259 ) ;
  assign n1270 = ~n1268 & n1269 ;
  assign n1271 = n1264 | n1270 ;
  assign n1272 = n1175 &  n1228 ;
  assign n1265 = x69 | n1175 ;
  assign n1266 = x69 &  n1175 ;
  assign n1267 = ( n1265 & ~n1266 ) | ( n1265 & 1'b0 ) | ( ~n1266 & 1'b0 ) ;
  assign n1276 = ( n1215 & n1224 ) | ( n1215 & n1267 ) | ( n1224 & n1267 ) ;
  assign n1277 = ( n1215 & ~n1227 ) | ( n1215 & n1267 ) | ( ~n1227 & n1267 ) ;
  assign n1278 = ~n1276 & n1277 ;
  assign n1279 = n1272 | n1278 ;
  assign n1280 = n1183 &  n1228 ;
  assign n1273 = x68 | n1183 ;
  assign n1274 = x68 &  n1183 ;
  assign n1275 = ( n1273 & ~n1274 ) | ( n1273 & 1'b0 ) | ( ~n1274 & 1'b0 ) ;
  assign n1284 = ( n1214 & n1224 ) | ( n1214 & n1275 ) | ( n1224 & n1275 ) ;
  assign n1285 = ( n1214 & ~n1227 ) | ( n1214 & n1275 ) | ( ~n1227 & n1275 ) ;
  assign n1286 = ~n1284 & n1285 ;
  assign n1287 = n1280 | n1286 ;
  assign n1288 = n1192 &  n1228 ;
  assign n1281 = x67 | n1192 ;
  assign n1282 = x67 &  n1192 ;
  assign n1283 = ( n1281 & ~n1282 ) | ( n1281 & 1'b0 ) | ( ~n1282 & 1'b0 ) ;
  assign n1292 = ( n1213 & n1224 ) | ( n1213 & n1283 ) | ( n1224 & n1283 ) ;
  assign n1293 = ( n1213 & ~n1227 ) | ( n1213 & n1283 ) | ( ~n1227 & n1283 ) ;
  assign n1294 = ~n1292 & n1293 ;
  assign n1295 = n1288 | n1294 ;
  assign n1296 = n1198 &  n1228 ;
  assign n1289 = x66 | n1198 ;
  assign n1290 = x66 &  n1198 ;
  assign n1291 = ( n1289 & ~n1290 ) | ( n1289 & 1'b0 ) | ( ~n1290 & 1'b0 ) ;
  assign n1301 = ( n1212 & ~n1224 ) | ( n1212 & n1291 ) | ( ~n1224 & n1291 ) ;
  assign n1302 = ( n1212 & n1227 ) | ( n1212 & n1291 ) | ( n1227 & n1291 ) ;
  assign n1303 = ( n1301 & ~n1302 ) | ( n1301 & 1'b0 ) | ( ~n1302 & 1'b0 ) ;
  assign n1304 = n1296 | n1303 ;
  assign n1305 = n1210 &  n1228 ;
  assign n1297 = x65 &  n1210 ;
  assign n1298 = x65 | n1209 ;
  assign n1299 = n1205 | n1298 ;
  assign n1300 = ( n1211 & ~n1297 ) | ( n1211 & n1299 ) | ( ~n1297 & n1299 ) ;
  assign n1306 = ( x65 & n1210 ) | ( x65 & n1211 ) | ( n1210 & n1211 ) ;
  assign n1307 = ( n1227 & ~n1297 ) | ( n1227 & n1306 ) | ( ~n1297 & n1306 ) ;
  assign n1308 = ( n1224 & n1300 ) | ( n1224 & n1307 ) | ( n1300 & n1307 ) ;
  assign n1309 = ( n1300 & ~n1308 ) | ( n1300 & 1'b0 ) | ( ~n1308 & 1'b0 ) ;
  assign n1310 = n1305 | n1309 ;
  assign n1311 = ( x64 & ~x78 ) | ( x64 & 1'b0 ) | ( ~x78 & 1'b0 ) ;
  assign n1312 = ( n201 & ~n219 ) | ( n201 & n1311 ) | ( ~n219 & n1311 ) ;
  assign n1313 = ~n201 & n1312 ;
  assign n1314 = ( n420 & ~n429 ) | ( n420 & n1313 ) | ( ~n429 & n1313 ) ;
  assign n1315 = ~n420 & n1314 ;
  assign n1316 = n1224 &  n1315 ;
  assign n1317 = ( x50 & ~n1315 ) | ( x50 & n1316 ) | ( ~n1315 & n1316 ) ;
  assign n1318 = ~n145 & n1211 ;
  assign n1319 = ( n143 & ~n190 ) | ( n143 & n1318 ) | ( ~n190 & n1318 ) ;
  assign n1320 = ~n143 & n1319 ;
  assign n1321 = ~n356 & n1320 ;
  assign n1322 = ~n1224 & n1321 ;
  assign n1323 = n1317 | n1322 ;
  assign n1324 = ~x49 & x64 ;
  assign n1325 = ( x65 & ~n1323 ) | ( x65 & n1324 ) | ( ~n1323 & n1324 ) ;
  assign n1326 = ( x66 & ~n1310 ) | ( x66 & n1325 ) | ( ~n1310 & n1325 ) ;
  assign n1327 = ( x67 & ~n1304 ) | ( x67 & n1326 ) | ( ~n1304 & n1326 ) ;
  assign n1328 = ( x68 & ~n1295 ) | ( x68 & n1327 ) | ( ~n1295 & n1327 ) ;
  assign n1329 = ( x69 & ~n1287 ) | ( x69 & n1328 ) | ( ~n1287 & n1328 ) ;
  assign n1330 = ( x70 & ~n1279 ) | ( x70 & n1329 ) | ( ~n1279 & n1329 ) ;
  assign n1331 = ( x71 & ~n1271 ) | ( x71 & n1330 ) | ( ~n1271 & n1330 ) ;
  assign n1332 = ( x72 & ~n1263 ) | ( x72 & n1331 ) | ( ~n1263 & n1331 ) ;
  assign n1333 = ( x73 & ~n1255 ) | ( x73 & n1332 ) | ( ~n1255 & n1332 ) ;
  assign n1334 = ( x74 & ~n1247 ) | ( x74 & n1333 ) | ( ~n1247 & n1333 ) ;
  assign n1338 = ( x75 & ~n1239 ) | ( x75 & n1334 ) | ( ~n1239 & n1334 ) ;
  assign n1358 = ( x76 & ~n1346 ) | ( x76 & n1338 ) | ( ~n1346 & n1338 ) ;
  assign n1359 = ( x77 & ~n1357 ) | ( x77 & n1358 ) | ( ~n1357 & n1358 ) ;
  assign n1363 = n201 | n219 ;
  assign n1364 = ( n429 & ~n420 ) | ( n429 & n1363 ) | ( ~n420 & n1363 ) ;
  assign n1365 = n420 | n1364 ;
  assign n1360 = x77 | n1223 ;
  assign n1361 = ( x77 & n1223 ) | ( x77 & n1227 ) | ( n1223 & n1227 ) ;
  assign n1362 = ( n1122 & ~n1360 ) | ( n1122 & n1361 ) | ( ~n1360 & n1361 ) ;
  assign n1367 = x78 &  n1362 ;
  assign n1366 = x78 | n1362 ;
  assign n1368 = ( n1365 & ~n1367 ) | ( n1365 & n1366 ) | ( ~n1367 & n1366 ) ;
  assign n1369 = n1359 | n1368 ;
  assign n1370 = ~n1227 & n1362 ;
  assign n1387 = ( n1357 & ~n1370 ) | ( n1357 & 1'b0 ) | ( ~n1370 & 1'b0 ) ;
  assign n1388 = n1369 &  n1387 ;
  assign n1377 = x77 | n1357 ;
  assign n1378 = x77 &  n1357 ;
  assign n1379 = ( n1377 & ~n1378 ) | ( n1377 & 1'b0 ) | ( ~n1378 & 1'b0 ) ;
  assign n1389 = n1358 &  n1379 ;
  assign n1371 = ( n1369 & ~n1370 ) | ( n1369 & 1'b0 ) | ( ~n1370 & 1'b0 ) ;
  assign n1390 = ( n1358 & ~n1371 ) | ( n1358 & n1379 ) | ( ~n1371 & n1379 ) ;
  assign n1391 = ( n1388 & ~n1389 ) | ( n1388 & n1390 ) | ( ~n1389 & n1390 ) ;
  assign n1381 = ( x78 & n1359 ) | ( x78 & n1362 ) | ( n1359 & n1362 ) ;
  assign n1380 = ( x78 & ~n1359 ) | ( x78 & n1362 ) | ( ~n1359 & n1362 ) ;
  assign n1382 = ( n1359 & ~n1381 ) | ( n1359 & n1380 ) | ( ~n1381 & n1380 ) ;
  assign n1383 = ~n1371 & n1382 ;
  assign n1384 = n1122 &  n1227 ;
  assign n1385 = n1369 &  n1384 ;
  assign n1386 = n1383 | n1385 ;
  assign n1372 = ( n1346 & ~n1370 ) | ( n1346 & 1'b0 ) | ( ~n1370 & 1'b0 ) ;
  assign n1373 = n1369 &  n1372 ;
  assign n1347 = x76 | n1346 ;
  assign n1348 = x76 &  n1346 ;
  assign n1349 = ( n1347 & ~n1348 ) | ( n1347 & 1'b0 ) | ( ~n1348 & 1'b0 ) ;
  assign n1374 = n1338 &  n1349 ;
  assign n1375 = ( n1338 & ~n1371 ) | ( n1338 & n1349 ) | ( ~n1371 & n1349 ) ;
  assign n1376 = ( n1373 & ~n1374 ) | ( n1373 & n1375 ) | ( ~n1374 & n1375 ) ;
  assign n1395 = ( n1239 & ~n1370 ) | ( n1239 & 1'b0 ) | ( ~n1370 & 1'b0 ) ;
  assign n1396 = n1369 &  n1395 ;
  assign n1335 = x75 | n1239 ;
  assign n1336 = x75 &  n1239 ;
  assign n1337 = ( n1335 & ~n1336 ) | ( n1335 & 1'b0 ) | ( ~n1336 & 1'b0 ) ;
  assign n1398 = ( n1334 & n1337 ) | ( n1334 & n1371 ) | ( n1337 & n1371 ) ;
  assign n1397 = n1334 | n1337 ;
  assign n1399 = ( n1396 & ~n1398 ) | ( n1396 & n1397 ) | ( ~n1398 & n1397 ) ;
  assign n1403 = ( n1247 & ~n1370 ) | ( n1247 & 1'b0 ) | ( ~n1370 & 1'b0 ) ;
  assign n1404 = n1369 &  n1403 ;
  assign n1392 = x74 | n1247 ;
  assign n1393 = x74 &  n1247 ;
  assign n1394 = ( n1392 & ~n1393 ) | ( n1392 & 1'b0 ) | ( ~n1393 & 1'b0 ) ;
  assign n1405 = n1333 &  n1394 ;
  assign n1406 = ( n1333 & ~n1371 ) | ( n1333 & n1394 ) | ( ~n1371 & n1394 ) ;
  assign n1407 = ( n1404 & ~n1405 ) | ( n1404 & n1406 ) | ( ~n1405 & n1406 ) ;
  assign n1411 = ( n1255 & ~n1370 ) | ( n1255 & 1'b0 ) | ( ~n1370 & 1'b0 ) ;
  assign n1412 = n1369 &  n1411 ;
  assign n1400 = x73 | n1255 ;
  assign n1401 = x73 &  n1255 ;
  assign n1402 = ( n1400 & ~n1401 ) | ( n1400 & 1'b0 ) | ( ~n1401 & 1'b0 ) ;
  assign n1413 = n1332 &  n1402 ;
  assign n1414 = ( n1332 & ~n1371 ) | ( n1332 & n1402 ) | ( ~n1371 & n1402 ) ;
  assign n1415 = ( n1412 & ~n1413 ) | ( n1412 & n1414 ) | ( ~n1413 & n1414 ) ;
  assign n1419 = ( n1263 & ~n1370 ) | ( n1263 & 1'b0 ) | ( ~n1370 & 1'b0 ) ;
  assign n1420 = n1369 &  n1419 ;
  assign n1408 = x72 | n1263 ;
  assign n1409 = x72 &  n1263 ;
  assign n1410 = ( n1408 & ~n1409 ) | ( n1408 & 1'b0 ) | ( ~n1409 & 1'b0 ) ;
  assign n1422 = ( n1331 & n1371 ) | ( n1331 & n1410 ) | ( n1371 & n1410 ) ;
  assign n1421 = n1331 | n1410 ;
  assign n1423 = ( n1420 & ~n1422 ) | ( n1420 & n1421 ) | ( ~n1422 & n1421 ) ;
  assign n1427 = ( n1271 & ~n1370 ) | ( n1271 & 1'b0 ) | ( ~n1370 & 1'b0 ) ;
  assign n1428 = n1369 &  n1427 ;
  assign n1416 = x71 | n1271 ;
  assign n1417 = x71 &  n1271 ;
  assign n1418 = ( n1416 & ~n1417 ) | ( n1416 & 1'b0 ) | ( ~n1417 & 1'b0 ) ;
  assign n1430 = ( n1330 & n1371 ) | ( n1330 & n1418 ) | ( n1371 & n1418 ) ;
  assign n1429 = n1330 | n1418 ;
  assign n1431 = ( n1428 & ~n1430 ) | ( n1428 & n1429 ) | ( ~n1430 & n1429 ) ;
  assign n1435 = ( n1279 & ~n1370 ) | ( n1279 & 1'b0 ) | ( ~n1370 & 1'b0 ) ;
  assign n1436 = n1369 &  n1435 ;
  assign n1424 = x70 | n1279 ;
  assign n1425 = x70 &  n1279 ;
  assign n1426 = ( n1424 & ~n1425 ) | ( n1424 & 1'b0 ) | ( ~n1425 & 1'b0 ) ;
  assign n1438 = ( n1329 & n1371 ) | ( n1329 & n1426 ) | ( n1371 & n1426 ) ;
  assign n1437 = n1329 | n1426 ;
  assign n1439 = ( n1436 & ~n1438 ) | ( n1436 & n1437 ) | ( ~n1438 & n1437 ) ;
  assign n1443 = ( n1287 & ~n1370 ) | ( n1287 & 1'b0 ) | ( ~n1370 & 1'b0 ) ;
  assign n1444 = n1369 &  n1443 ;
  assign n1432 = x69 | n1287 ;
  assign n1433 = x69 &  n1287 ;
  assign n1434 = ( n1432 & ~n1433 ) | ( n1432 & 1'b0 ) | ( ~n1433 & 1'b0 ) ;
  assign n1446 = ( n1328 & n1371 ) | ( n1328 & n1434 ) | ( n1371 & n1434 ) ;
  assign n1445 = n1328 | n1434 ;
  assign n1447 = ( n1444 & ~n1446 ) | ( n1444 & n1445 ) | ( ~n1446 & n1445 ) ;
  assign n1451 = ( n1295 & ~n1370 ) | ( n1295 & 1'b0 ) | ( ~n1370 & 1'b0 ) ;
  assign n1452 = n1369 &  n1451 ;
  assign n1440 = x68 | n1295 ;
  assign n1441 = x68 &  n1295 ;
  assign n1442 = ( n1440 & ~n1441 ) | ( n1440 & 1'b0 ) | ( ~n1441 & 1'b0 ) ;
  assign n1454 = ( n1327 & n1371 ) | ( n1327 & n1442 ) | ( n1371 & n1442 ) ;
  assign n1453 = n1327 | n1442 ;
  assign n1455 = ( n1452 & ~n1454 ) | ( n1452 & n1453 ) | ( ~n1454 & n1453 ) ;
  assign n1459 = ( n1304 & ~n1370 ) | ( n1304 & 1'b0 ) | ( ~n1370 & 1'b0 ) ;
  assign n1460 = n1369 &  n1459 ;
  assign n1448 = x67 | n1304 ;
  assign n1449 = x67 &  n1304 ;
  assign n1450 = ( n1448 & ~n1449 ) | ( n1448 & 1'b0 ) | ( ~n1449 & 1'b0 ) ;
  assign n1462 = ( n1326 & n1371 ) | ( n1326 & n1450 ) | ( n1371 & n1450 ) ;
  assign n1461 = n1326 | n1450 ;
  assign n1463 = ( n1460 & ~n1462 ) | ( n1460 & n1461 ) | ( ~n1462 & n1461 ) ;
  assign n1464 = ( n1310 & ~n1370 ) | ( n1310 & 1'b0 ) | ( ~n1370 & 1'b0 ) ;
  assign n1465 = n1369 &  n1464 ;
  assign n1456 = x66 | n1310 ;
  assign n1457 = x66 &  n1310 ;
  assign n1458 = ( n1456 & ~n1457 ) | ( n1456 & 1'b0 ) | ( ~n1457 & 1'b0 ) ;
  assign n1466 = n1325 &  n1458 ;
  assign n1467 = ( n1325 & ~n1371 ) | ( n1325 & n1458 ) | ( ~n1371 & n1458 ) ;
  assign n1468 = ( n1465 & ~n1466 ) | ( n1465 & n1467 ) | ( ~n1466 & n1467 ) ;
  assign n1469 = ( n1323 & ~x65 ) | ( n1323 & n1324 ) | ( ~x65 & n1324 ) ;
  assign n1470 = ( n1325 & ~n1324 ) | ( n1325 & n1469 ) | ( ~n1324 & n1469 ) ;
  assign n1471 = ~n1371 & n1470 ;
  assign n1472 = ( n1323 & ~n1370 ) | ( n1323 & 1'b0 ) | ( ~n1370 & 1'b0 ) ;
  assign n1473 = n1369 &  n1472 ;
  assign n1474 = n1471 | n1473 ;
  assign n1475 = ( x64 & ~n1371 ) | ( x64 & 1'b0 ) | ( ~n1371 & 1'b0 ) ;
  assign n1476 = ( x49 & ~n1475 ) | ( x49 & 1'b0 ) | ( ~n1475 & 1'b0 ) ;
  assign n1477 = ( n1324 & ~n1371 ) | ( n1324 & 1'b0 ) | ( ~n1371 & 1'b0 ) ;
  assign n1478 = n1476 | n1477 ;
  assign n1479 = ~x48 & x64 ;
  assign n1480 = ( x65 & ~n1478 ) | ( x65 & n1479 ) | ( ~n1478 & n1479 ) ;
  assign n1481 = ( x66 & ~n1474 ) | ( x66 & n1480 ) | ( ~n1474 & n1480 ) ;
  assign n1482 = ( x67 & ~n1468 ) | ( x67 & n1481 ) | ( ~n1468 & n1481 ) ;
  assign n1483 = ( x68 & ~n1463 ) | ( x68 & n1482 ) | ( ~n1463 & n1482 ) ;
  assign n1484 = ( x69 & ~n1455 ) | ( x69 & n1483 ) | ( ~n1455 & n1483 ) ;
  assign n1485 = ( x70 & ~n1447 ) | ( x70 & n1484 ) | ( ~n1447 & n1484 ) ;
  assign n1486 = ( x71 & ~n1439 ) | ( x71 & n1485 ) | ( ~n1439 & n1485 ) ;
  assign n1487 = ( x72 & ~n1431 ) | ( x72 & n1486 ) | ( ~n1431 & n1486 ) ;
  assign n1488 = ( x73 & ~n1423 ) | ( x73 & n1487 ) | ( ~n1423 & n1487 ) ;
  assign n1489 = ( x74 & ~n1415 ) | ( x74 & n1488 ) | ( ~n1415 & n1488 ) ;
  assign n1490 = ( x75 & ~n1407 ) | ( x75 & n1489 ) | ( ~n1407 & n1489 ) ;
  assign n1491 = ( x76 & ~n1399 ) | ( x76 & n1490 ) | ( ~n1399 & n1490 ) ;
  assign n1492 = ( x77 & ~n1376 ) | ( x77 & n1491 ) | ( ~n1376 & n1491 ) ;
  assign n1493 = ( x78 & ~n1391 ) | ( x78 & n1492 ) | ( ~n1391 & n1492 ) ;
  assign n1494 = ( x79 & ~n1386 ) | ( x79 & n1493 ) | ( ~n1386 & n1493 ) ;
  assign n1495 = n282 | n1494 ;
  assign n1513 = n1391 &  n1495 ;
  assign n1507 = x78 | n1391 ;
  assign n1508 = x78 &  n1391 ;
  assign n1509 = ( n1507 & ~n1508 ) | ( n1507 & 1'b0 ) | ( ~n1508 & 1'b0 ) ;
  assign n1514 = ( n282 & n1492 ) | ( n282 & n1509 ) | ( n1492 & n1509 ) ;
  assign n1515 = ( n1492 & ~n1494 ) | ( n1492 & n1509 ) | ( ~n1494 & n1509 ) ;
  assign n1516 = ~n1514 & n1515 ;
  assign n1517 = n1513 | n1516 ;
  assign n1511 = ( x79 & ~n282 ) | ( x79 & n1493 ) | ( ~n282 & n1493 ) ;
  assign n1510 = x79 &  n1493 ;
  assign n1512 = ( n1386 & ~n1511 ) | ( n1386 & n1510 ) | ( ~n1511 & n1510 ) ;
  assign n1496 = n1376 &  n1495 ;
  assign n1500 = x77 | n1376 ;
  assign n1501 = x77 &  n1376 ;
  assign n1502 = ( n1500 & ~n1501 ) | ( n1500 & 1'b0 ) | ( ~n1501 & 1'b0 ) ;
  assign n1503 = ( n282 & n1491 ) | ( n282 & n1502 ) | ( n1491 & n1502 ) ;
  assign n1504 = ( n1491 & ~n1494 ) | ( n1491 & n1502 ) | ( ~n1494 & n1502 ) ;
  assign n1505 = ~n1503 & n1504 ;
  assign n1506 = n1496 | n1505 ;
  assign n1518 = n1399 &  n1495 ;
  assign n1497 = x76 | n1399 ;
  assign n1498 = x76 &  n1399 ;
  assign n1499 = ( n1497 & ~n1498 ) | ( n1497 & 1'b0 ) | ( ~n1498 & 1'b0 ) ;
  assign n1522 = ( n282 & n1490 ) | ( n282 & n1499 ) | ( n1490 & n1499 ) ;
  assign n1523 = ( n1490 & ~n1494 ) | ( n1490 & n1499 ) | ( ~n1494 & n1499 ) ;
  assign n1524 = ~n1522 & n1523 ;
  assign n1525 = n1518 | n1524 ;
  assign n1526 = n1407 &  n1495 ;
  assign n1519 = x75 | n1407 ;
  assign n1520 = x75 &  n1407 ;
  assign n1521 = ( n1519 & ~n1520 ) | ( n1519 & 1'b0 ) | ( ~n1520 & 1'b0 ) ;
  assign n1530 = ( n282 & n1489 ) | ( n282 & n1521 ) | ( n1489 & n1521 ) ;
  assign n1531 = ( n1489 & ~n1494 ) | ( n1489 & n1521 ) | ( ~n1494 & n1521 ) ;
  assign n1532 = ~n1530 & n1531 ;
  assign n1533 = n1526 | n1532 ;
  assign n1534 = n1415 &  n1495 ;
  assign n1527 = x74 | n1415 ;
  assign n1528 = x74 &  n1415 ;
  assign n1529 = ( n1527 & ~n1528 ) | ( n1527 & 1'b0 ) | ( ~n1528 & 1'b0 ) ;
  assign n1538 = ( n282 & n1488 ) | ( n282 & n1529 ) | ( n1488 & n1529 ) ;
  assign n1539 = ( n1488 & ~n1494 ) | ( n1488 & n1529 ) | ( ~n1494 & n1529 ) ;
  assign n1540 = ~n1538 & n1539 ;
  assign n1541 = n1534 | n1540 ;
  assign n1542 = n1423 &  n1495 ;
  assign n1535 = x73 | n1423 ;
  assign n1536 = x73 &  n1423 ;
  assign n1537 = ( n1535 & ~n1536 ) | ( n1535 & 1'b0 ) | ( ~n1536 & 1'b0 ) ;
  assign n1546 = ( n282 & n1487 ) | ( n282 & n1537 ) | ( n1487 & n1537 ) ;
  assign n1547 = ( n1487 & ~n1494 ) | ( n1487 & n1537 ) | ( ~n1494 & n1537 ) ;
  assign n1548 = ~n1546 & n1547 ;
  assign n1549 = n1542 | n1548 ;
  assign n1550 = n1431 &  n1495 ;
  assign n1543 = x72 | n1431 ;
  assign n1544 = x72 &  n1431 ;
  assign n1545 = ( n1543 & ~n1544 ) | ( n1543 & 1'b0 ) | ( ~n1544 & 1'b0 ) ;
  assign n1554 = ( n282 & n1486 ) | ( n282 & n1545 ) | ( n1486 & n1545 ) ;
  assign n1555 = ( n1486 & ~n1494 ) | ( n1486 & n1545 ) | ( ~n1494 & n1545 ) ;
  assign n1556 = ~n1554 & n1555 ;
  assign n1557 = n1550 | n1556 ;
  assign n1558 = n1439 &  n1495 ;
  assign n1551 = x71 | n1439 ;
  assign n1552 = x71 &  n1439 ;
  assign n1553 = ( n1551 & ~n1552 ) | ( n1551 & 1'b0 ) | ( ~n1552 & 1'b0 ) ;
  assign n1562 = ( n282 & n1485 ) | ( n282 & n1553 ) | ( n1485 & n1553 ) ;
  assign n1563 = ( n1485 & ~n1494 ) | ( n1485 & n1553 ) | ( ~n1494 & n1553 ) ;
  assign n1564 = ~n1562 & n1563 ;
  assign n1565 = n1558 | n1564 ;
  assign n1566 = n1447 &  n1495 ;
  assign n1559 = x70 | n1447 ;
  assign n1560 = x70 &  n1447 ;
  assign n1561 = ( n1559 & ~n1560 ) | ( n1559 & 1'b0 ) | ( ~n1560 & 1'b0 ) ;
  assign n1570 = ( n282 & n1484 ) | ( n282 & n1561 ) | ( n1484 & n1561 ) ;
  assign n1571 = ( n1484 & ~n1494 ) | ( n1484 & n1561 ) | ( ~n1494 & n1561 ) ;
  assign n1572 = ~n1570 & n1571 ;
  assign n1573 = n1566 | n1572 ;
  assign n1574 = n1455 &  n1495 ;
  assign n1567 = x69 | n1455 ;
  assign n1568 = x69 &  n1455 ;
  assign n1569 = ( n1567 & ~n1568 ) | ( n1567 & 1'b0 ) | ( ~n1568 & 1'b0 ) ;
  assign n1578 = ( n282 & n1483 ) | ( n282 & n1569 ) | ( n1483 & n1569 ) ;
  assign n1579 = ( n1483 & ~n1494 ) | ( n1483 & n1569 ) | ( ~n1494 & n1569 ) ;
  assign n1580 = ~n1578 & n1579 ;
  assign n1581 = n1574 | n1580 ;
  assign n1582 = n1463 &  n1495 ;
  assign n1575 = x68 | n1463 ;
  assign n1576 = x68 &  n1463 ;
  assign n1577 = ( n1575 & ~n1576 ) | ( n1575 & 1'b0 ) | ( ~n1576 & 1'b0 ) ;
  assign n1586 = ( n282 & n1482 ) | ( n282 & n1577 ) | ( n1482 & n1577 ) ;
  assign n1587 = ( n1482 & ~n1494 ) | ( n1482 & n1577 ) | ( ~n1494 & n1577 ) ;
  assign n1588 = ~n1586 & n1587 ;
  assign n1589 = n1582 | n1588 ;
  assign n1590 = n1468 &  n1495 ;
  assign n1583 = x67 | n1468 ;
  assign n1584 = x67 &  n1468 ;
  assign n1585 = ( n1583 & ~n1584 ) | ( n1583 & 1'b0 ) | ( ~n1584 & 1'b0 ) ;
  assign n1594 = ( n282 & n1481 ) | ( n282 & n1585 ) | ( n1481 & n1585 ) ;
  assign n1595 = ( n1481 & ~n1494 ) | ( n1481 & n1585 ) | ( ~n1494 & n1585 ) ;
  assign n1596 = ~n1594 & n1595 ;
  assign n1597 = n1590 | n1596 ;
  assign n1598 = n1474 &  n1495 ;
  assign n1591 = x66 | n1474 ;
  assign n1592 = x66 &  n1474 ;
  assign n1593 = ( n1591 & ~n1592 ) | ( n1591 & 1'b0 ) | ( ~n1592 & 1'b0 ) ;
  assign n1599 = ( n1480 & ~n282 ) | ( n1480 & n1593 ) | ( ~n282 & n1593 ) ;
  assign n1600 = ( n1480 & n1494 ) | ( n1480 & n1593 ) | ( n1494 & n1593 ) ;
  assign n1601 = ( n1599 & ~n1600 ) | ( n1599 & 1'b0 ) | ( ~n1600 & 1'b0 ) ;
  assign n1602 = n1598 | n1601 ;
  assign n1603 = n1478 &  n1495 ;
  assign n1604 = ( x65 & ~x49 ) | ( x65 & n1475 ) | ( ~x49 & n1475 ) ;
  assign n1605 = ( x49 & ~n1475 ) | ( x49 & x65 ) | ( ~n1475 & x65 ) ;
  assign n1606 = ( n1604 & ~x65 ) | ( n1604 & n1605 ) | ( ~x65 & n1605 ) ;
  assign n1607 = ( n1479 & ~n1494 ) | ( n1479 & n1606 ) | ( ~n1494 & n1606 ) ;
  assign n1608 = ( n282 & n1479 ) | ( n282 & n1606 ) | ( n1479 & n1606 ) ;
  assign n1609 = ( n1607 & ~n1608 ) | ( n1607 & 1'b0 ) | ( ~n1608 & 1'b0 ) ;
  assign n1610 = n1603 | n1609 ;
  assign n1611 = ( x64 & ~x80 ) | ( x64 & 1'b0 ) | ( ~x80 & 1'b0 ) ;
  assign n1612 = ( n201 & ~n420 ) | ( n201 & n1611 ) | ( ~n420 & n1611 ) ;
  assign n1613 = ~n201 & n1612 ;
  assign n1614 = ~n429 & n1613 ;
  assign n1615 = n1494 &  n1614 ;
  assign n1616 = ( x48 & ~n1614 ) | ( x48 & n1615 ) | ( ~n1614 & n1615 ) ;
  assign n1617 = ~n143 & n1479 ;
  assign n1618 = ( n190 & ~n356 ) | ( n190 & n1617 ) | ( ~n356 & n1617 ) ;
  assign n1619 = ~n190 & n1618 ;
  assign n1620 = ~n1494 & n1619 ;
  assign n1621 = n1616 | n1620 ;
  assign n1622 = ~x47 & x64 ;
  assign n1623 = ( x65 & ~n1621 ) | ( x65 & n1622 ) | ( ~n1621 & n1622 ) ;
  assign n1624 = ( x66 & ~n1610 ) | ( x66 & n1623 ) | ( ~n1610 & n1623 ) ;
  assign n1625 = ( x67 & ~n1602 ) | ( x67 & n1624 ) | ( ~n1602 & n1624 ) ;
  assign n1626 = ( x68 & ~n1597 ) | ( x68 & n1625 ) | ( ~n1597 & n1625 ) ;
  assign n1627 = ( x69 & ~n1589 ) | ( x69 & n1626 ) | ( ~n1589 & n1626 ) ;
  assign n1628 = ( x70 & ~n1581 ) | ( x70 & n1627 ) | ( ~n1581 & n1627 ) ;
  assign n1629 = ( x71 & ~n1573 ) | ( x71 & n1628 ) | ( ~n1573 & n1628 ) ;
  assign n1630 = ( x72 & ~n1565 ) | ( x72 & n1629 ) | ( ~n1565 & n1629 ) ;
  assign n1631 = ( x73 & ~n1557 ) | ( x73 & n1630 ) | ( ~n1557 & n1630 ) ;
  assign n1632 = ( x74 & ~n1549 ) | ( x74 & n1631 ) | ( ~n1549 & n1631 ) ;
  assign n1633 = ( x75 & ~n1541 ) | ( x75 & n1632 ) | ( ~n1541 & n1632 ) ;
  assign n1634 = ( x76 & ~n1533 ) | ( x76 & n1633 ) | ( ~n1533 & n1633 ) ;
  assign n1635 = ( x77 & ~n1525 ) | ( x77 & n1634 ) | ( ~n1525 & n1634 ) ;
  assign n1636 = ( x78 & ~n1506 ) | ( x78 & n1635 ) | ( ~n1506 & n1635 ) ;
  assign n1637 = ( x79 & ~n1517 ) | ( x79 & n1636 ) | ( ~n1517 & n1636 ) ;
  assign n1638 = ( x80 & ~n1512 ) | ( x80 & n1637 ) | ( ~n1512 & n1637 ) ;
  assign n1639 = n317 | n1638 ;
  assign n1785 = n1517 &  n1639 ;
  assign n1786 = x79 | n1517 ;
  assign n1787 = x79 &  n1517 ;
  assign n1788 = ( n1786 & ~n1787 ) | ( n1786 & 1'b0 ) | ( ~n1787 & 1'b0 ) ;
  assign n1789 = ( n317 & n1636 ) | ( n317 & n1788 ) | ( n1636 & n1788 ) ;
  assign n1790 = ( n1636 & ~n1638 ) | ( n1636 & n1788 ) | ( ~n1638 & n1788 ) ;
  assign n1791 = ~n1789 & n1790 ;
  assign n1792 = n1785 | n1791 ;
  assign n1640 = n1506 &  n1639 ;
  assign n1644 = x78 | n1506 ;
  assign n1645 = x78 &  n1506 ;
  assign n1646 = ( n1644 & ~n1645 ) | ( n1644 & 1'b0 ) | ( ~n1645 & 1'b0 ) ;
  assign n1647 = ( n317 & n1635 ) | ( n317 & n1646 ) | ( n1635 & n1646 ) ;
  assign n1648 = ( n1635 & ~n1638 ) | ( n1635 & n1646 ) | ( ~n1638 & n1646 ) ;
  assign n1649 = ~n1647 & n1648 ;
  assign n1650 = n1640 | n1649 ;
  assign n1651 = n1525 &  n1639 ;
  assign n1641 = x77 | n1525 ;
  assign n1642 = x77 &  n1525 ;
  assign n1643 = ( n1641 & ~n1642 ) | ( n1641 & 1'b0 ) | ( ~n1642 & 1'b0 ) ;
  assign n1655 = ( n317 & n1634 ) | ( n317 & n1643 ) | ( n1634 & n1643 ) ;
  assign n1656 = ( n1634 & ~n1638 ) | ( n1634 & n1643 ) | ( ~n1638 & n1643 ) ;
  assign n1657 = ~n1655 & n1656 ;
  assign n1658 = n1651 | n1657 ;
  assign n1659 = n1533 &  n1639 ;
  assign n1652 = x76 | n1533 ;
  assign n1653 = x76 &  n1533 ;
  assign n1654 = ( n1652 & ~n1653 ) | ( n1652 & 1'b0 ) | ( ~n1653 & 1'b0 ) ;
  assign n1663 = ( n317 & n1633 ) | ( n317 & n1654 ) | ( n1633 & n1654 ) ;
  assign n1664 = ( n1633 & ~n1638 ) | ( n1633 & n1654 ) | ( ~n1638 & n1654 ) ;
  assign n1665 = ~n1663 & n1664 ;
  assign n1666 = n1659 | n1665 ;
  assign n1667 = n1541 &  n1639 ;
  assign n1660 = x75 | n1541 ;
  assign n1661 = x75 &  n1541 ;
  assign n1662 = ( n1660 & ~n1661 ) | ( n1660 & 1'b0 ) | ( ~n1661 & 1'b0 ) ;
  assign n1671 = ( n317 & n1632 ) | ( n317 & n1662 ) | ( n1632 & n1662 ) ;
  assign n1672 = ( n1632 & ~n1638 ) | ( n1632 & n1662 ) | ( ~n1638 & n1662 ) ;
  assign n1673 = ~n1671 & n1672 ;
  assign n1674 = n1667 | n1673 ;
  assign n1675 = n1549 &  n1639 ;
  assign n1668 = x74 | n1549 ;
  assign n1669 = x74 &  n1549 ;
  assign n1670 = ( n1668 & ~n1669 ) | ( n1668 & 1'b0 ) | ( ~n1669 & 1'b0 ) ;
  assign n1679 = ( n317 & n1631 ) | ( n317 & n1670 ) | ( n1631 & n1670 ) ;
  assign n1680 = ( n1631 & ~n1638 ) | ( n1631 & n1670 ) | ( ~n1638 & n1670 ) ;
  assign n1681 = ~n1679 & n1680 ;
  assign n1682 = n1675 | n1681 ;
  assign n1683 = n1557 &  n1639 ;
  assign n1676 = x73 | n1557 ;
  assign n1677 = x73 &  n1557 ;
  assign n1678 = ( n1676 & ~n1677 ) | ( n1676 & 1'b0 ) | ( ~n1677 & 1'b0 ) ;
  assign n1687 = ( n317 & n1630 ) | ( n317 & n1678 ) | ( n1630 & n1678 ) ;
  assign n1688 = ( n1630 & ~n1638 ) | ( n1630 & n1678 ) | ( ~n1638 & n1678 ) ;
  assign n1689 = ~n1687 & n1688 ;
  assign n1690 = n1683 | n1689 ;
  assign n1691 = n1565 &  n1639 ;
  assign n1684 = x72 | n1565 ;
  assign n1685 = x72 &  n1565 ;
  assign n1686 = ( n1684 & ~n1685 ) | ( n1684 & 1'b0 ) | ( ~n1685 & 1'b0 ) ;
  assign n1695 = ( n317 & n1629 ) | ( n317 & n1686 ) | ( n1629 & n1686 ) ;
  assign n1696 = ( n1629 & ~n1638 ) | ( n1629 & n1686 ) | ( ~n1638 & n1686 ) ;
  assign n1697 = ~n1695 & n1696 ;
  assign n1698 = n1691 | n1697 ;
  assign n1699 = n1573 &  n1639 ;
  assign n1692 = x71 | n1573 ;
  assign n1693 = x71 &  n1573 ;
  assign n1694 = ( n1692 & ~n1693 ) | ( n1692 & 1'b0 ) | ( ~n1693 & 1'b0 ) ;
  assign n1703 = ( n317 & n1628 ) | ( n317 & n1694 ) | ( n1628 & n1694 ) ;
  assign n1704 = ( n1628 & ~n1638 ) | ( n1628 & n1694 ) | ( ~n1638 & n1694 ) ;
  assign n1705 = ~n1703 & n1704 ;
  assign n1706 = n1699 | n1705 ;
  assign n1707 = n1581 &  n1639 ;
  assign n1700 = x70 | n1581 ;
  assign n1701 = x70 &  n1581 ;
  assign n1702 = ( n1700 & ~n1701 ) | ( n1700 & 1'b0 ) | ( ~n1701 & 1'b0 ) ;
  assign n1711 = ( n317 & n1627 ) | ( n317 & n1702 ) | ( n1627 & n1702 ) ;
  assign n1712 = ( n1627 & ~n1638 ) | ( n1627 & n1702 ) | ( ~n1638 & n1702 ) ;
  assign n1713 = ~n1711 & n1712 ;
  assign n1714 = n1707 | n1713 ;
  assign n1715 = n1589 &  n1639 ;
  assign n1708 = x69 | n1589 ;
  assign n1709 = x69 &  n1589 ;
  assign n1710 = ( n1708 & ~n1709 ) | ( n1708 & 1'b0 ) | ( ~n1709 & 1'b0 ) ;
  assign n1719 = ( n317 & n1626 ) | ( n317 & n1710 ) | ( n1626 & n1710 ) ;
  assign n1720 = ( n1626 & ~n1638 ) | ( n1626 & n1710 ) | ( ~n1638 & n1710 ) ;
  assign n1721 = ~n1719 & n1720 ;
  assign n1722 = n1715 | n1721 ;
  assign n1723 = n1597 &  n1639 ;
  assign n1716 = x68 | n1597 ;
  assign n1717 = x68 &  n1597 ;
  assign n1718 = ( n1716 & ~n1717 ) | ( n1716 & 1'b0 ) | ( ~n1717 & 1'b0 ) ;
  assign n1727 = ( n317 & n1625 ) | ( n317 & n1718 ) | ( n1625 & n1718 ) ;
  assign n1728 = ( n1625 & ~n1638 ) | ( n1625 & n1718 ) | ( ~n1638 & n1718 ) ;
  assign n1729 = ~n1727 & n1728 ;
  assign n1730 = n1723 | n1729 ;
  assign n1731 = n1602 &  n1639 ;
  assign n1724 = x67 | n1602 ;
  assign n1725 = x67 &  n1602 ;
  assign n1726 = ( n1724 & ~n1725 ) | ( n1724 & 1'b0 ) | ( ~n1725 & 1'b0 ) ;
  assign n1735 = ( n317 & n1624 ) | ( n317 & n1726 ) | ( n1624 & n1726 ) ;
  assign n1736 = ( n1624 & ~n1638 ) | ( n1624 & n1726 ) | ( ~n1638 & n1726 ) ;
  assign n1737 = ~n1735 & n1736 ;
  assign n1738 = n1731 | n1737 ;
  assign n1739 = n1610 &  n1639 ;
  assign n1732 = x66 | n1610 ;
  assign n1733 = x66 &  n1610 ;
  assign n1734 = ( n1732 & ~n1733 ) | ( n1732 & 1'b0 ) | ( ~n1733 & 1'b0 ) ;
  assign n1743 = ( n1623 & ~n317 ) | ( n1623 & n1734 ) | ( ~n317 & n1734 ) ;
  assign n1744 = ( n1623 & n1638 ) | ( n1623 & n1734 ) | ( n1638 & n1734 ) ;
  assign n1745 = ( n1743 & ~n1744 ) | ( n1743 & 1'b0 ) | ( ~n1744 & 1'b0 ) ;
  assign n1746 = n1739 | n1745 ;
  assign n1747 = n1621 &  n1639 ;
  assign n1740 = x65 &  n1621 ;
  assign n1741 = x65 | n1620 ;
  assign n1742 = n1616 | n1741 ;
  assign n1748 = ~n1740 & n1742 ;
  assign n1749 = ( n1622 & ~n1638 ) | ( n1622 & n1748 ) | ( ~n1638 & n1748 ) ;
  assign n1750 = ( n317 & n1622 ) | ( n317 & n1748 ) | ( n1622 & n1748 ) ;
  assign n1751 = ( n1749 & ~n1750 ) | ( n1749 & 1'b0 ) | ( ~n1750 & 1'b0 ) ;
  assign n1752 = n1747 | n1751 ;
  assign n1753 = ( x64 & ~x81 ) | ( x64 & 1'b0 ) | ( ~x81 & 1'b0 ) ;
  assign n1754 = ( n142 & ~n181 ) | ( n142 & n1753 ) | ( ~n181 & n1753 ) ;
  assign n1755 = ~n142 & n1754 ;
  assign n1756 = ( n273 & ~n261 ) | ( n273 & n1755 ) | ( ~n261 & n1755 ) ;
  assign n1757 = ~n273 & n1756 ;
  assign n1758 = ~n270 & n1757 ;
  assign n1759 = n1638 &  n1758 ;
  assign n1760 = ( x47 & ~n1758 ) | ( x47 & n1759 ) | ( ~n1758 & n1759 ) ;
  assign n1761 = ~n201 & n1622 ;
  assign n1762 = ( n420 & ~n429 ) | ( n420 & n1761 ) | ( ~n429 & n1761 ) ;
  assign n1763 = ~n420 & n1762 ;
  assign n1764 = ~n1638 & n1763 ;
  assign n1765 = n1760 | n1764 ;
  assign n1766 = ~x46 & x64 ;
  assign n1767 = ( x65 & ~n1765 ) | ( x65 & n1766 ) | ( ~n1765 & n1766 ) ;
  assign n1768 = ( x66 & ~n1752 ) | ( x66 & n1767 ) | ( ~n1752 & n1767 ) ;
  assign n1769 = ( x67 & ~n1746 ) | ( x67 & n1768 ) | ( ~n1746 & n1768 ) ;
  assign n1770 = ( x68 & ~n1738 ) | ( x68 & n1769 ) | ( ~n1738 & n1769 ) ;
  assign n1771 = ( x69 & ~n1730 ) | ( x69 & n1770 ) | ( ~n1730 & n1770 ) ;
  assign n1772 = ( x70 & ~n1722 ) | ( x70 & n1771 ) | ( ~n1722 & n1771 ) ;
  assign n1773 = ( x71 & ~n1714 ) | ( x71 & n1772 ) | ( ~n1714 & n1772 ) ;
  assign n1774 = ( x72 & ~n1706 ) | ( x72 & n1773 ) | ( ~n1706 & n1773 ) ;
  assign n1775 = ( x73 & ~n1698 ) | ( x73 & n1774 ) | ( ~n1698 & n1774 ) ;
  assign n1776 = ( x74 & ~n1690 ) | ( x74 & n1775 ) | ( ~n1690 & n1775 ) ;
  assign n1777 = ( x75 & ~n1682 ) | ( x75 & n1776 ) | ( ~n1682 & n1776 ) ;
  assign n1778 = ( x76 & ~n1674 ) | ( x76 & n1777 ) | ( ~n1674 & n1777 ) ;
  assign n1779 = ( x77 & ~n1666 ) | ( x77 & n1778 ) | ( ~n1666 & n1778 ) ;
  assign n1780 = ( x78 & ~n1658 ) | ( x78 & n1779 ) | ( ~n1658 & n1779 ) ;
  assign n1784 = ( x79 & ~n1650 ) | ( x79 & n1780 ) | ( ~n1650 & n1780 ) ;
  assign n1796 = ( x80 & ~n1792 ) | ( x80 & n1784 ) | ( ~n1792 & n1784 ) ;
  assign n1800 = n142 | n181 ;
  assign n1801 = ( n261 & ~n273 ) | ( n261 & n1800 ) | ( ~n273 & n1800 ) ;
  assign n1802 = n273 | n1801 ;
  assign n1803 = n270 | n1802 ;
  assign n1798 = ( x80 & ~n317 ) | ( x80 & n1637 ) | ( ~n317 & n1637 ) ;
  assign n1797 = x80 &  n1637 ;
  assign n1799 = ( n1512 & ~n1798 ) | ( n1512 & n1797 ) | ( ~n1798 & n1797 ) ;
  assign n1805 = x81 &  n1799 ;
  assign n1804 = x81 | n1799 ;
  assign n1806 = ( n1803 & ~n1805 ) | ( n1803 & n1804 ) | ( ~n1805 & n1804 ) ;
  assign n1807 = n1796 | n1806 ;
  assign n1808 = ~n317 & n1799 ;
  assign n1810 = ( n1792 & ~n1808 ) | ( n1792 & 1'b0 ) | ( ~n1808 & 1'b0 ) ;
  assign n1811 = n1807 &  n1810 ;
  assign n1793 = x80 | n1792 ;
  assign n1794 = x80 &  n1792 ;
  assign n1795 = ( n1793 & ~n1794 ) | ( n1793 & 1'b0 ) | ( ~n1794 & 1'b0 ) ;
  assign n1812 = n1784 &  n1795 ;
  assign n1809 = ( n1807 & ~n1808 ) | ( n1807 & 1'b0 ) | ( ~n1808 & 1'b0 ) ;
  assign n1813 = ( n1784 & ~n1809 ) | ( n1784 & n1795 ) | ( ~n1809 & n1795 ) ;
  assign n1814 = ( n1811 & ~n1812 ) | ( n1811 & n1813 ) | ( ~n1812 & n1813 ) ;
  assign n1816 = ( x81 & n1796 ) | ( x81 & n1799 ) | ( n1796 & n1799 ) ;
  assign n1815 = ( x81 & ~n1796 ) | ( x81 & n1799 ) | ( ~n1796 & n1799 ) ;
  assign n1817 = ( n1796 & ~n1816 ) | ( n1796 & n1815 ) | ( ~n1816 & n1815 ) ;
  assign n1818 = ~n1809 & n1817 ;
  assign n1819 = n317 &  n1512 ;
  assign n1820 = n1807 &  n1819 ;
  assign n1821 = n1818 | n1820 ;
  assign n1825 = ( n1650 & ~n1808 ) | ( n1650 & 1'b0 ) | ( ~n1808 & 1'b0 ) ;
  assign n1826 = n1807 &  n1825 ;
  assign n1781 = x79 | n1650 ;
  assign n1782 = x79 &  n1650 ;
  assign n1783 = ( n1781 & ~n1782 ) | ( n1781 & 1'b0 ) | ( ~n1782 & 1'b0 ) ;
  assign n1828 = ( n1780 & n1783 ) | ( n1780 & n1809 ) | ( n1783 & n1809 ) ;
  assign n1827 = n1780 | n1783 ;
  assign n1829 = ( n1826 & ~n1828 ) | ( n1826 & n1827 ) | ( ~n1828 & n1827 ) ;
  assign n1833 = ( n1658 & ~n1808 ) | ( n1658 & 1'b0 ) | ( ~n1808 & 1'b0 ) ;
  assign n1834 = n1807 &  n1833 ;
  assign n1822 = x78 | n1658 ;
  assign n1823 = x78 &  n1658 ;
  assign n1824 = ( n1822 & ~n1823 ) | ( n1822 & 1'b0 ) | ( ~n1823 & 1'b0 ) ;
  assign n1835 = n1779 &  n1824 ;
  assign n1836 = ( n1779 & ~n1809 ) | ( n1779 & n1824 ) | ( ~n1809 & n1824 ) ;
  assign n1837 = ( n1834 & ~n1835 ) | ( n1834 & n1836 ) | ( ~n1835 & n1836 ) ;
  assign n1841 = ( n1666 & ~n1808 ) | ( n1666 & 1'b0 ) | ( ~n1808 & 1'b0 ) ;
  assign n1842 = n1807 &  n1841 ;
  assign n1830 = x77 | n1666 ;
  assign n1831 = x77 &  n1666 ;
  assign n1832 = ( n1830 & ~n1831 ) | ( n1830 & 1'b0 ) | ( ~n1831 & 1'b0 ) ;
  assign n1843 = n1778 &  n1832 ;
  assign n1844 = ( n1778 & ~n1809 ) | ( n1778 & n1832 ) | ( ~n1809 & n1832 ) ;
  assign n1845 = ( n1842 & ~n1843 ) | ( n1842 & n1844 ) | ( ~n1843 & n1844 ) ;
  assign n1849 = ( n1674 & ~n1808 ) | ( n1674 & 1'b0 ) | ( ~n1808 & 1'b0 ) ;
  assign n1850 = n1807 &  n1849 ;
  assign n1838 = x76 | n1674 ;
  assign n1839 = x76 &  n1674 ;
  assign n1840 = ( n1838 & ~n1839 ) | ( n1838 & 1'b0 ) | ( ~n1839 & 1'b0 ) ;
  assign n1851 = n1777 &  n1840 ;
  assign n1852 = ( n1777 & ~n1809 ) | ( n1777 & n1840 ) | ( ~n1809 & n1840 ) ;
  assign n1853 = ( n1850 & ~n1851 ) | ( n1850 & n1852 ) | ( ~n1851 & n1852 ) ;
  assign n1857 = ( n1682 & ~n1808 ) | ( n1682 & 1'b0 ) | ( ~n1808 & 1'b0 ) ;
  assign n1858 = n1807 &  n1857 ;
  assign n1846 = x75 | n1682 ;
  assign n1847 = x75 &  n1682 ;
  assign n1848 = ( n1846 & ~n1847 ) | ( n1846 & 1'b0 ) | ( ~n1847 & 1'b0 ) ;
  assign n1860 = ( n1776 & n1809 ) | ( n1776 & n1848 ) | ( n1809 & n1848 ) ;
  assign n1859 = n1776 | n1848 ;
  assign n1861 = ( n1858 & ~n1860 ) | ( n1858 & n1859 ) | ( ~n1860 & n1859 ) ;
  assign n1865 = ( n1690 & ~n1808 ) | ( n1690 & 1'b0 ) | ( ~n1808 & 1'b0 ) ;
  assign n1866 = n1807 &  n1865 ;
  assign n1854 = x74 | n1690 ;
  assign n1855 = x74 &  n1690 ;
  assign n1856 = ( n1854 & ~n1855 ) | ( n1854 & 1'b0 ) | ( ~n1855 & 1'b0 ) ;
  assign n1868 = ( n1775 & n1809 ) | ( n1775 & n1856 ) | ( n1809 & n1856 ) ;
  assign n1867 = n1775 | n1856 ;
  assign n1869 = ( n1866 & ~n1868 ) | ( n1866 & n1867 ) | ( ~n1868 & n1867 ) ;
  assign n1873 = ( n1698 & ~n1808 ) | ( n1698 & 1'b0 ) | ( ~n1808 & 1'b0 ) ;
  assign n1874 = n1807 &  n1873 ;
  assign n1862 = x73 | n1698 ;
  assign n1863 = x73 &  n1698 ;
  assign n1864 = ( n1862 & ~n1863 ) | ( n1862 & 1'b0 ) | ( ~n1863 & 1'b0 ) ;
  assign n1876 = ( n1774 & n1809 ) | ( n1774 & n1864 ) | ( n1809 & n1864 ) ;
  assign n1875 = n1774 | n1864 ;
  assign n1877 = ( n1874 & ~n1876 ) | ( n1874 & n1875 ) | ( ~n1876 & n1875 ) ;
  assign n1881 = ( n1706 & ~n1808 ) | ( n1706 & 1'b0 ) | ( ~n1808 & 1'b0 ) ;
  assign n1882 = n1807 &  n1881 ;
  assign n1870 = x72 | n1706 ;
  assign n1871 = x72 &  n1706 ;
  assign n1872 = ( n1870 & ~n1871 ) | ( n1870 & 1'b0 ) | ( ~n1871 & 1'b0 ) ;
  assign n1884 = ( n1773 & n1809 ) | ( n1773 & n1872 ) | ( n1809 & n1872 ) ;
  assign n1883 = n1773 | n1872 ;
  assign n1885 = ( n1882 & ~n1884 ) | ( n1882 & n1883 ) | ( ~n1884 & n1883 ) ;
  assign n1889 = ( n1714 & ~n1808 ) | ( n1714 & 1'b0 ) | ( ~n1808 & 1'b0 ) ;
  assign n1890 = n1807 &  n1889 ;
  assign n1878 = x71 | n1714 ;
  assign n1879 = x71 &  n1714 ;
  assign n1880 = ( n1878 & ~n1879 ) | ( n1878 & 1'b0 ) | ( ~n1879 & 1'b0 ) ;
  assign n1892 = ( n1772 & n1809 ) | ( n1772 & n1880 ) | ( n1809 & n1880 ) ;
  assign n1891 = n1772 | n1880 ;
  assign n1893 = ( n1890 & ~n1892 ) | ( n1890 & n1891 ) | ( ~n1892 & n1891 ) ;
  assign n1897 = ( n1722 & ~n1808 ) | ( n1722 & 1'b0 ) | ( ~n1808 & 1'b0 ) ;
  assign n1898 = n1807 &  n1897 ;
  assign n1886 = x70 | n1722 ;
  assign n1887 = x70 &  n1722 ;
  assign n1888 = ( n1886 & ~n1887 ) | ( n1886 & 1'b0 ) | ( ~n1887 & 1'b0 ) ;
  assign n1900 = ( n1771 & n1809 ) | ( n1771 & n1888 ) | ( n1809 & n1888 ) ;
  assign n1899 = n1771 | n1888 ;
  assign n1901 = ( n1898 & ~n1900 ) | ( n1898 & n1899 ) | ( ~n1900 & n1899 ) ;
  assign n1905 = ( n1730 & ~n1808 ) | ( n1730 & 1'b0 ) | ( ~n1808 & 1'b0 ) ;
  assign n1906 = n1807 &  n1905 ;
  assign n1894 = x69 | n1730 ;
  assign n1895 = x69 &  n1730 ;
  assign n1896 = ( n1894 & ~n1895 ) | ( n1894 & 1'b0 ) | ( ~n1895 & 1'b0 ) ;
  assign n1908 = ( n1770 & n1809 ) | ( n1770 & n1896 ) | ( n1809 & n1896 ) ;
  assign n1907 = n1770 | n1896 ;
  assign n1909 = ( n1906 & ~n1908 ) | ( n1906 & n1907 ) | ( ~n1908 & n1907 ) ;
  assign n1913 = ( n1738 & ~n1808 ) | ( n1738 & 1'b0 ) | ( ~n1808 & 1'b0 ) ;
  assign n1914 = n1807 &  n1913 ;
  assign n1902 = x68 | n1738 ;
  assign n1903 = x68 &  n1738 ;
  assign n1904 = ( n1902 & ~n1903 ) | ( n1902 & 1'b0 ) | ( ~n1903 & 1'b0 ) ;
  assign n1916 = ( n1769 & n1809 ) | ( n1769 & n1904 ) | ( n1809 & n1904 ) ;
  assign n1915 = n1769 | n1904 ;
  assign n1917 = ( n1914 & ~n1916 ) | ( n1914 & n1915 ) | ( ~n1916 & n1915 ) ;
  assign n1921 = ( n1746 & ~n1808 ) | ( n1746 & 1'b0 ) | ( ~n1808 & 1'b0 ) ;
  assign n1922 = n1807 &  n1921 ;
  assign n1910 = x67 | n1746 ;
  assign n1911 = x67 &  n1746 ;
  assign n1912 = ( n1910 & ~n1911 ) | ( n1910 & 1'b0 ) | ( ~n1911 & 1'b0 ) ;
  assign n1924 = ( n1768 & n1809 ) | ( n1768 & n1912 ) | ( n1809 & n1912 ) ;
  assign n1923 = n1768 | n1912 ;
  assign n1925 = ( n1922 & ~n1924 ) | ( n1922 & n1923 ) | ( ~n1924 & n1923 ) ;
  assign n1926 = ( n1752 & ~n1808 ) | ( n1752 & 1'b0 ) | ( ~n1808 & 1'b0 ) ;
  assign n1927 = n1807 &  n1926 ;
  assign n1918 = x66 | n1752 ;
  assign n1919 = x66 &  n1752 ;
  assign n1920 = ( n1918 & ~n1919 ) | ( n1918 & 1'b0 ) | ( ~n1919 & 1'b0 ) ;
  assign n1928 = n1767 &  n1920 ;
  assign n1929 = ( n1767 & ~n1809 ) | ( n1767 & n1920 ) | ( ~n1809 & n1920 ) ;
  assign n1930 = ( n1927 & ~n1928 ) | ( n1927 & n1929 ) | ( ~n1928 & n1929 ) ;
  assign n1931 = ( n1765 & ~x65 ) | ( n1765 & n1766 ) | ( ~x65 & n1766 ) ;
  assign n1932 = ( n1767 & ~n1766 ) | ( n1767 & n1931 ) | ( ~n1766 & n1931 ) ;
  assign n1933 = ~n1809 & n1932 ;
  assign n1934 = ( n1765 & ~n1808 ) | ( n1765 & 1'b0 ) | ( ~n1808 & 1'b0 ) ;
  assign n1935 = n1807 &  n1934 ;
  assign n1936 = n1933 | n1935 ;
  assign n1937 = ( x64 & ~n1809 ) | ( x64 & 1'b0 ) | ( ~n1809 & 1'b0 ) ;
  assign n1938 = ( x46 & ~n1937 ) | ( x46 & 1'b0 ) | ( ~n1937 & 1'b0 ) ;
  assign n1939 = ( n1766 & ~n1809 ) | ( n1766 & 1'b0 ) | ( ~n1809 & 1'b0 ) ;
  assign n1940 = n1938 | n1939 ;
  assign n1941 = ~x45 & x64 ;
  assign n1942 = ( x65 & ~n1940 ) | ( x65 & n1941 ) | ( ~n1940 & n1941 ) ;
  assign n1943 = ( x66 & ~n1936 ) | ( x66 & n1942 ) | ( ~n1936 & n1942 ) ;
  assign n1944 = ( x67 & ~n1930 ) | ( x67 & n1943 ) | ( ~n1930 & n1943 ) ;
  assign n1945 = ( x68 & ~n1925 ) | ( x68 & n1944 ) | ( ~n1925 & n1944 ) ;
  assign n1946 = ( x69 & ~n1917 ) | ( x69 & n1945 ) | ( ~n1917 & n1945 ) ;
  assign n1947 = ( x70 & ~n1909 ) | ( x70 & n1946 ) | ( ~n1909 & n1946 ) ;
  assign n1948 = ( x71 & ~n1901 ) | ( x71 & n1947 ) | ( ~n1901 & n1947 ) ;
  assign n1949 = ( x72 & ~n1893 ) | ( x72 & n1948 ) | ( ~n1893 & n1948 ) ;
  assign n1950 = ( x73 & ~n1885 ) | ( x73 & n1949 ) | ( ~n1885 & n1949 ) ;
  assign n1951 = ( x74 & ~n1877 ) | ( x74 & n1950 ) | ( ~n1877 & n1950 ) ;
  assign n1952 = ( x75 & ~n1869 ) | ( x75 & n1951 ) | ( ~n1869 & n1951 ) ;
  assign n1953 = ( x76 & ~n1861 ) | ( x76 & n1952 ) | ( ~n1861 & n1952 ) ;
  assign n1954 = ( x77 & ~n1853 ) | ( x77 & n1953 ) | ( ~n1853 & n1953 ) ;
  assign n1955 = ( x78 & ~n1845 ) | ( x78 & n1954 ) | ( ~n1845 & n1954 ) ;
  assign n1956 = ( x79 & ~n1837 ) | ( x79 & n1955 ) | ( ~n1837 & n1955 ) ;
  assign n1957 = ( x80 & ~n1829 ) | ( x80 & n1956 ) | ( ~n1829 & n1956 ) ;
  assign n1958 = ( x81 & ~n1814 ) | ( x81 & n1957 ) | ( ~n1814 & n1957 ) ;
  assign n1959 = ( x82 & ~n1821 ) | ( x82 & n1958 ) | ( ~n1821 & n1958 ) ;
  assign n1960 = n198 | n200 ;
  assign n1961 = ( n255 & ~n209 ) | ( n255 & n1960 ) | ( ~n209 & n1960 ) ;
  assign n1962 = n209 | n1961 ;
  assign n1963 = n240 | n1962 ;
  assign n1964 = n1959 | n1963 ;
  assign n1965 = n1814 &  n1964 ;
  assign n1969 = x81 | n1814 ;
  assign n1970 = x81 &  n1814 ;
  assign n1971 = ( n1969 & ~n1970 ) | ( n1969 & 1'b0 ) | ( ~n1970 & 1'b0 ) ;
  assign n1972 = ( n1957 & n1959 ) | ( n1957 & n1971 ) | ( n1959 & n1971 ) ;
  assign n1973 = ( n1957 & ~n1963 ) | ( n1957 & n1971 ) | ( ~n1963 & n1971 ) ;
  assign n1974 = ~n1972 & n1973 ;
  assign n1975 = n1965 | n1974 ;
  assign n1976 = x82 | n1958 ;
  assign n1977 = ( x82 & n1958 ) | ( x82 & n1963 ) | ( n1958 & n1963 ) ;
  assign n1978 = ( n1821 & ~n1976 ) | ( n1821 & n1977 ) | ( ~n1976 & n1977 ) ;
  assign n1979 = n1829 &  n1964 ;
  assign n1966 = x80 | n1829 ;
  assign n1967 = x80 &  n1829 ;
  assign n1968 = ( n1966 & ~n1967 ) | ( n1966 & 1'b0 ) | ( ~n1967 & 1'b0 ) ;
  assign n1983 = ( n1956 & n1959 ) | ( n1956 & n1968 ) | ( n1959 & n1968 ) ;
  assign n1984 = ( n1956 & ~n1963 ) | ( n1956 & n1968 ) | ( ~n1963 & n1968 ) ;
  assign n1985 = ~n1983 & n1984 ;
  assign n1986 = n1979 | n1985 ;
  assign n1987 = n1837 &  n1964 ;
  assign n1980 = x79 | n1837 ;
  assign n1981 = x79 &  n1837 ;
  assign n1982 = ( n1980 & ~n1981 ) | ( n1980 & 1'b0 ) | ( ~n1981 & 1'b0 ) ;
  assign n1991 = ( n1955 & n1959 ) | ( n1955 & n1982 ) | ( n1959 & n1982 ) ;
  assign n1992 = ( n1955 & ~n1963 ) | ( n1955 & n1982 ) | ( ~n1963 & n1982 ) ;
  assign n1993 = ~n1991 & n1992 ;
  assign n1994 = n1987 | n1993 ;
  assign n1995 = n1845 &  n1964 ;
  assign n1988 = x78 | n1845 ;
  assign n1989 = x78 &  n1845 ;
  assign n1990 = ( n1988 & ~n1989 ) | ( n1988 & 1'b0 ) | ( ~n1989 & 1'b0 ) ;
  assign n1999 = ( n1954 & n1959 ) | ( n1954 & n1990 ) | ( n1959 & n1990 ) ;
  assign n2000 = ( n1954 & ~n1963 ) | ( n1954 & n1990 ) | ( ~n1963 & n1990 ) ;
  assign n2001 = ~n1999 & n2000 ;
  assign n2002 = n1995 | n2001 ;
  assign n2003 = n1853 &  n1964 ;
  assign n1996 = x77 | n1853 ;
  assign n1997 = x77 &  n1853 ;
  assign n1998 = ( n1996 & ~n1997 ) | ( n1996 & 1'b0 ) | ( ~n1997 & 1'b0 ) ;
  assign n2007 = ( n1953 & n1959 ) | ( n1953 & n1998 ) | ( n1959 & n1998 ) ;
  assign n2008 = ( n1953 & ~n1963 ) | ( n1953 & n1998 ) | ( ~n1963 & n1998 ) ;
  assign n2009 = ~n2007 & n2008 ;
  assign n2010 = n2003 | n2009 ;
  assign n2011 = n1861 &  n1964 ;
  assign n2004 = x76 | n1861 ;
  assign n2005 = x76 &  n1861 ;
  assign n2006 = ( n2004 & ~n2005 ) | ( n2004 & 1'b0 ) | ( ~n2005 & 1'b0 ) ;
  assign n2015 = ( n1952 & n1959 ) | ( n1952 & n2006 ) | ( n1959 & n2006 ) ;
  assign n2016 = ( n1952 & ~n1963 ) | ( n1952 & n2006 ) | ( ~n1963 & n2006 ) ;
  assign n2017 = ~n2015 & n2016 ;
  assign n2018 = n2011 | n2017 ;
  assign n2019 = n1869 &  n1964 ;
  assign n2012 = x75 | n1869 ;
  assign n2013 = x75 &  n1869 ;
  assign n2014 = ( n2012 & ~n2013 ) | ( n2012 & 1'b0 ) | ( ~n2013 & 1'b0 ) ;
  assign n2023 = ( n1951 & n1959 ) | ( n1951 & n2014 ) | ( n1959 & n2014 ) ;
  assign n2024 = ( n1951 & ~n1963 ) | ( n1951 & n2014 ) | ( ~n1963 & n2014 ) ;
  assign n2025 = ~n2023 & n2024 ;
  assign n2026 = n2019 | n2025 ;
  assign n2027 = n1877 &  n1964 ;
  assign n2020 = x74 | n1877 ;
  assign n2021 = x74 &  n1877 ;
  assign n2022 = ( n2020 & ~n2021 ) | ( n2020 & 1'b0 ) | ( ~n2021 & 1'b0 ) ;
  assign n2031 = ( n1950 & n1959 ) | ( n1950 & n2022 ) | ( n1959 & n2022 ) ;
  assign n2032 = ( n1950 & ~n1963 ) | ( n1950 & n2022 ) | ( ~n1963 & n2022 ) ;
  assign n2033 = ~n2031 & n2032 ;
  assign n2034 = n2027 | n2033 ;
  assign n2035 = n1885 &  n1964 ;
  assign n2028 = x73 | n1885 ;
  assign n2029 = x73 &  n1885 ;
  assign n2030 = ( n2028 & ~n2029 ) | ( n2028 & 1'b0 ) | ( ~n2029 & 1'b0 ) ;
  assign n2039 = ( n1949 & n1959 ) | ( n1949 & n2030 ) | ( n1959 & n2030 ) ;
  assign n2040 = ( n1949 & ~n1963 ) | ( n1949 & n2030 ) | ( ~n1963 & n2030 ) ;
  assign n2041 = ~n2039 & n2040 ;
  assign n2042 = n2035 | n2041 ;
  assign n2043 = n1893 &  n1964 ;
  assign n2036 = x72 | n1893 ;
  assign n2037 = x72 &  n1893 ;
  assign n2038 = ( n2036 & ~n2037 ) | ( n2036 & 1'b0 ) | ( ~n2037 & 1'b0 ) ;
  assign n2047 = ( n1948 & n1959 ) | ( n1948 & n2038 ) | ( n1959 & n2038 ) ;
  assign n2048 = ( n1948 & ~n1963 ) | ( n1948 & n2038 ) | ( ~n1963 & n2038 ) ;
  assign n2049 = ~n2047 & n2048 ;
  assign n2050 = n2043 | n2049 ;
  assign n2051 = n1901 &  n1964 ;
  assign n2044 = x71 | n1901 ;
  assign n2045 = x71 &  n1901 ;
  assign n2046 = ( n2044 & ~n2045 ) | ( n2044 & 1'b0 ) | ( ~n2045 & 1'b0 ) ;
  assign n2055 = ( n1947 & n1959 ) | ( n1947 & n2046 ) | ( n1959 & n2046 ) ;
  assign n2056 = ( n1947 & ~n1963 ) | ( n1947 & n2046 ) | ( ~n1963 & n2046 ) ;
  assign n2057 = ~n2055 & n2056 ;
  assign n2058 = n2051 | n2057 ;
  assign n2059 = n1909 &  n1964 ;
  assign n2052 = x70 | n1909 ;
  assign n2053 = x70 &  n1909 ;
  assign n2054 = ( n2052 & ~n2053 ) | ( n2052 & 1'b0 ) | ( ~n2053 & 1'b0 ) ;
  assign n2063 = ( n1946 & n1959 ) | ( n1946 & n2054 ) | ( n1959 & n2054 ) ;
  assign n2064 = ( n1946 & ~n1963 ) | ( n1946 & n2054 ) | ( ~n1963 & n2054 ) ;
  assign n2065 = ~n2063 & n2064 ;
  assign n2066 = n2059 | n2065 ;
  assign n2067 = n1917 &  n1964 ;
  assign n2060 = x69 | n1917 ;
  assign n2061 = x69 &  n1917 ;
  assign n2062 = ( n2060 & ~n2061 ) | ( n2060 & 1'b0 ) | ( ~n2061 & 1'b0 ) ;
  assign n2071 = ( n1945 & n1959 ) | ( n1945 & n2062 ) | ( n1959 & n2062 ) ;
  assign n2072 = ( n1945 & ~n1963 ) | ( n1945 & n2062 ) | ( ~n1963 & n2062 ) ;
  assign n2073 = ~n2071 & n2072 ;
  assign n2074 = n2067 | n2073 ;
  assign n2075 = n1925 &  n1964 ;
  assign n2068 = x68 | n1925 ;
  assign n2069 = x68 &  n1925 ;
  assign n2070 = ( n2068 & ~n2069 ) | ( n2068 & 1'b0 ) | ( ~n2069 & 1'b0 ) ;
  assign n2079 = ( n1944 & n1959 ) | ( n1944 & n2070 ) | ( n1959 & n2070 ) ;
  assign n2080 = ( n1944 & ~n1963 ) | ( n1944 & n2070 ) | ( ~n1963 & n2070 ) ;
  assign n2081 = ~n2079 & n2080 ;
  assign n2082 = n2075 | n2081 ;
  assign n2083 = n1930 &  n1964 ;
  assign n2076 = x67 | n1930 ;
  assign n2077 = x67 &  n1930 ;
  assign n2078 = ( n2076 & ~n2077 ) | ( n2076 & 1'b0 ) | ( ~n2077 & 1'b0 ) ;
  assign n2087 = ( n1943 & n1959 ) | ( n1943 & n2078 ) | ( n1959 & n2078 ) ;
  assign n2088 = ( n1943 & ~n1963 ) | ( n1943 & n2078 ) | ( ~n1963 & n2078 ) ;
  assign n2089 = ~n2087 & n2088 ;
  assign n2090 = n2083 | n2089 ;
  assign n2091 = n1936 &  n1964 ;
  assign n2084 = x66 | n1936 ;
  assign n2085 = x66 &  n1936 ;
  assign n2086 = ( n2084 & ~n2085 ) | ( n2084 & 1'b0 ) | ( ~n2085 & 1'b0 ) ;
  assign n2096 = ( n1942 & ~n1959 ) | ( n1942 & n2086 ) | ( ~n1959 & n2086 ) ;
  assign n2097 = ( n1942 & n1963 ) | ( n1942 & n2086 ) | ( n1963 & n2086 ) ;
  assign n2098 = ( n2096 & ~n2097 ) | ( n2096 & 1'b0 ) | ( ~n2097 & 1'b0 ) ;
  assign n2099 = n2091 | n2098 ;
  assign n2100 = n1940 &  n1964 ;
  assign n2092 = x65 &  n1940 ;
  assign n2093 = ( n1938 & ~x65 ) | ( n1938 & n1939 ) | ( ~x65 & n1939 ) ;
  assign n2094 = x65 | n2093 ;
  assign n2095 = ( n1941 & ~n2092 ) | ( n1941 & n2094 ) | ( ~n2092 & n2094 ) ;
  assign n2101 = ( x65 & n1940 ) | ( x65 & n1941 ) | ( n1940 & n1941 ) ;
  assign n2102 = ( n1963 & ~n2092 ) | ( n1963 & n2101 ) | ( ~n2092 & n2101 ) ;
  assign n2103 = ( n1959 & n2095 ) | ( n1959 & n2102 ) | ( n2095 & n2102 ) ;
  assign n2104 = ( n2095 & ~n2103 ) | ( n2095 & 1'b0 ) | ( ~n2103 & 1'b0 ) ;
  assign n2105 = n2100 | n2104 ;
  assign n2106 = ( x64 & ~x83 ) | ( x64 & 1'b0 ) | ( ~x83 & 1'b0 ) ;
  assign n2107 = ( n181 & ~n261 ) | ( n181 & n2106 ) | ( ~n261 & n2106 ) ;
  assign n2108 = ~n181 & n2107 ;
  assign n2109 = ( n270 & ~n273 ) | ( n270 & n2108 ) | ( ~n273 & n2108 ) ;
  assign n2110 = ~n270 & n2109 ;
  assign n2111 = n1959 &  n2110 ;
  assign n2112 = ( x45 & ~n2110 ) | ( x45 & n2111 ) | ( ~n2110 & n2111 ) ;
  assign n2113 = ~n200 & n1941 ;
  assign n2114 = ( n198 & ~n209 ) | ( n198 & n2113 ) | ( ~n209 & n2113 ) ;
  assign n2115 = ~n198 & n2114 ;
  assign n2116 = ( n240 & ~n255 ) | ( n240 & n2115 ) | ( ~n255 & n2115 ) ;
  assign n2117 = ~n240 & n2116 ;
  assign n2118 = ~n1959 & n2117 ;
  assign n2119 = n2112 | n2118 ;
  assign n2120 = ~x44 & x64 ;
  assign n2121 = ( x65 & ~n2119 ) | ( x65 & n2120 ) | ( ~n2119 & n2120 ) ;
  assign n2122 = ( x66 & ~n2105 ) | ( x66 & n2121 ) | ( ~n2105 & n2121 ) ;
  assign n2123 = ( x67 & ~n2099 ) | ( x67 & n2122 ) | ( ~n2099 & n2122 ) ;
  assign n2124 = ( x68 & ~n2090 ) | ( x68 & n2123 ) | ( ~n2090 & n2123 ) ;
  assign n2125 = ( x69 & ~n2082 ) | ( x69 & n2124 ) | ( ~n2082 & n2124 ) ;
  assign n2126 = ( x70 & ~n2074 ) | ( x70 & n2125 ) | ( ~n2074 & n2125 ) ;
  assign n2127 = ( x71 & ~n2066 ) | ( x71 & n2126 ) | ( ~n2066 & n2126 ) ;
  assign n2128 = ( x72 & ~n2058 ) | ( x72 & n2127 ) | ( ~n2058 & n2127 ) ;
  assign n2129 = ( x73 & ~n2050 ) | ( x73 & n2128 ) | ( ~n2050 & n2128 ) ;
  assign n2130 = ( x74 & ~n2042 ) | ( x74 & n2129 ) | ( ~n2042 & n2129 ) ;
  assign n2131 = ( x75 & ~n2034 ) | ( x75 & n2130 ) | ( ~n2034 & n2130 ) ;
  assign n2132 = ( x76 & ~n2026 ) | ( x76 & n2131 ) | ( ~n2026 & n2131 ) ;
  assign n2133 = ( x77 & ~n2018 ) | ( x77 & n2132 ) | ( ~n2018 & n2132 ) ;
  assign n2134 = ( x78 & ~n2010 ) | ( x78 & n2133 ) | ( ~n2010 & n2133 ) ;
  assign n2135 = ( x79 & ~n2002 ) | ( x79 & n2134 ) | ( ~n2002 & n2134 ) ;
  assign n2136 = ( x80 & ~n1994 ) | ( x80 & n2135 ) | ( ~n1994 & n2135 ) ;
  assign n2137 = ( x81 & ~n1986 ) | ( x81 & n2136 ) | ( ~n1986 & n2136 ) ;
  assign n2138 = ( x82 & ~n1975 ) | ( x82 & n2137 ) | ( ~n1975 & n2137 ) ;
  assign n2139 = ( x83 & ~n1978 ) | ( x83 & n2138 ) | ( ~n1978 & n2138 ) ;
  assign n2140 = n192 | n2139 ;
  assign n2141 = n1975 &  n2140 ;
  assign n2145 = x82 | n1975 ;
  assign n2146 = x82 &  n1975 ;
  assign n2147 = ( n2145 & ~n2146 ) | ( n2145 & 1'b0 ) | ( ~n2146 & 1'b0 ) ;
  assign n2148 = ( n192 & n2137 ) | ( n192 & n2147 ) | ( n2137 & n2147 ) ;
  assign n2149 = ( n2137 & ~n2139 ) | ( n2137 & n2147 ) | ( ~n2139 & n2147 ) ;
  assign n2150 = ~n2148 & n2149 ;
  assign n2151 = n2141 | n2150 ;
  assign n2152 = n1986 &  n2140 ;
  assign n2142 = x81 | n1986 ;
  assign n2143 = x81 &  n1986 ;
  assign n2144 = ( n2142 & ~n2143 ) | ( n2142 & 1'b0 ) | ( ~n2143 & 1'b0 ) ;
  assign n2156 = ( n192 & n2136 ) | ( n192 & n2144 ) | ( n2136 & n2144 ) ;
  assign n2157 = ( n2136 & ~n2139 ) | ( n2136 & n2144 ) | ( ~n2139 & n2144 ) ;
  assign n2158 = ~n2156 & n2157 ;
  assign n2159 = n2152 | n2158 ;
  assign n2160 = n1994 &  n2140 ;
  assign n2153 = x80 | n1994 ;
  assign n2154 = x80 &  n1994 ;
  assign n2155 = ( n2153 & ~n2154 ) | ( n2153 & 1'b0 ) | ( ~n2154 & 1'b0 ) ;
  assign n2164 = ( n192 & n2135 ) | ( n192 & n2155 ) | ( n2135 & n2155 ) ;
  assign n2165 = ( n2135 & ~n2139 ) | ( n2135 & n2155 ) | ( ~n2139 & n2155 ) ;
  assign n2166 = ~n2164 & n2165 ;
  assign n2167 = n2160 | n2166 ;
  assign n2168 = n2002 &  n2140 ;
  assign n2161 = x79 | n2002 ;
  assign n2162 = x79 &  n2002 ;
  assign n2163 = ( n2161 & ~n2162 ) | ( n2161 & 1'b0 ) | ( ~n2162 & 1'b0 ) ;
  assign n2172 = ( n192 & n2134 ) | ( n192 & n2163 ) | ( n2134 & n2163 ) ;
  assign n2173 = ( n2134 & ~n2139 ) | ( n2134 & n2163 ) | ( ~n2139 & n2163 ) ;
  assign n2174 = ~n2172 & n2173 ;
  assign n2175 = n2168 | n2174 ;
  assign n2176 = n2010 &  n2140 ;
  assign n2169 = x78 | n2010 ;
  assign n2170 = x78 &  n2010 ;
  assign n2171 = ( n2169 & ~n2170 ) | ( n2169 & 1'b0 ) | ( ~n2170 & 1'b0 ) ;
  assign n2180 = ( n192 & n2133 ) | ( n192 & n2171 ) | ( n2133 & n2171 ) ;
  assign n2181 = ( n2133 & ~n2139 ) | ( n2133 & n2171 ) | ( ~n2139 & n2171 ) ;
  assign n2182 = ~n2180 & n2181 ;
  assign n2183 = n2176 | n2182 ;
  assign n2184 = n2018 &  n2140 ;
  assign n2177 = x77 | n2018 ;
  assign n2178 = x77 &  n2018 ;
  assign n2179 = ( n2177 & ~n2178 ) | ( n2177 & 1'b0 ) | ( ~n2178 & 1'b0 ) ;
  assign n2188 = ( n192 & n2132 ) | ( n192 & n2179 ) | ( n2132 & n2179 ) ;
  assign n2189 = ( n2132 & ~n2139 ) | ( n2132 & n2179 ) | ( ~n2139 & n2179 ) ;
  assign n2190 = ~n2188 & n2189 ;
  assign n2191 = n2184 | n2190 ;
  assign n2192 = n2026 &  n2140 ;
  assign n2185 = x76 | n2026 ;
  assign n2186 = x76 &  n2026 ;
  assign n2187 = ( n2185 & ~n2186 ) | ( n2185 & 1'b0 ) | ( ~n2186 & 1'b0 ) ;
  assign n2196 = ( n192 & n2131 ) | ( n192 & n2187 ) | ( n2131 & n2187 ) ;
  assign n2197 = ( n2131 & ~n2139 ) | ( n2131 & n2187 ) | ( ~n2139 & n2187 ) ;
  assign n2198 = ~n2196 & n2197 ;
  assign n2199 = n2192 | n2198 ;
  assign n2200 = n2034 &  n2140 ;
  assign n2193 = x75 | n2034 ;
  assign n2194 = x75 &  n2034 ;
  assign n2195 = ( n2193 & ~n2194 ) | ( n2193 & 1'b0 ) | ( ~n2194 & 1'b0 ) ;
  assign n2204 = ( n192 & n2130 ) | ( n192 & n2195 ) | ( n2130 & n2195 ) ;
  assign n2205 = ( n2130 & ~n2139 ) | ( n2130 & n2195 ) | ( ~n2139 & n2195 ) ;
  assign n2206 = ~n2204 & n2205 ;
  assign n2207 = n2200 | n2206 ;
  assign n2208 = n2042 &  n2140 ;
  assign n2201 = x74 | n2042 ;
  assign n2202 = x74 &  n2042 ;
  assign n2203 = ( n2201 & ~n2202 ) | ( n2201 & 1'b0 ) | ( ~n2202 & 1'b0 ) ;
  assign n2212 = ( n192 & n2129 ) | ( n192 & n2203 ) | ( n2129 & n2203 ) ;
  assign n2213 = ( n2129 & ~n2139 ) | ( n2129 & n2203 ) | ( ~n2139 & n2203 ) ;
  assign n2214 = ~n2212 & n2213 ;
  assign n2215 = n2208 | n2214 ;
  assign n2216 = n2050 &  n2140 ;
  assign n2209 = x73 | n2050 ;
  assign n2210 = x73 &  n2050 ;
  assign n2211 = ( n2209 & ~n2210 ) | ( n2209 & 1'b0 ) | ( ~n2210 & 1'b0 ) ;
  assign n2220 = ( n192 & n2128 ) | ( n192 & n2211 ) | ( n2128 & n2211 ) ;
  assign n2221 = ( n2128 & ~n2139 ) | ( n2128 & n2211 ) | ( ~n2139 & n2211 ) ;
  assign n2222 = ~n2220 & n2221 ;
  assign n2223 = n2216 | n2222 ;
  assign n2224 = n2058 &  n2140 ;
  assign n2217 = x72 | n2058 ;
  assign n2218 = x72 &  n2058 ;
  assign n2219 = ( n2217 & ~n2218 ) | ( n2217 & 1'b0 ) | ( ~n2218 & 1'b0 ) ;
  assign n2228 = ( n192 & n2127 ) | ( n192 & n2219 ) | ( n2127 & n2219 ) ;
  assign n2229 = ( n2127 & ~n2139 ) | ( n2127 & n2219 ) | ( ~n2139 & n2219 ) ;
  assign n2230 = ~n2228 & n2229 ;
  assign n2231 = n2224 | n2230 ;
  assign n2232 = n2066 &  n2140 ;
  assign n2225 = x71 | n2066 ;
  assign n2226 = x71 &  n2066 ;
  assign n2227 = ( n2225 & ~n2226 ) | ( n2225 & 1'b0 ) | ( ~n2226 & 1'b0 ) ;
  assign n2236 = ( n192 & n2126 ) | ( n192 & n2227 ) | ( n2126 & n2227 ) ;
  assign n2237 = ( n2126 & ~n2139 ) | ( n2126 & n2227 ) | ( ~n2139 & n2227 ) ;
  assign n2238 = ~n2236 & n2237 ;
  assign n2239 = n2232 | n2238 ;
  assign n2240 = n2074 &  n2140 ;
  assign n2233 = x70 | n2074 ;
  assign n2234 = x70 &  n2074 ;
  assign n2235 = ( n2233 & ~n2234 ) | ( n2233 & 1'b0 ) | ( ~n2234 & 1'b0 ) ;
  assign n2244 = ( n192 & n2125 ) | ( n192 & n2235 ) | ( n2125 & n2235 ) ;
  assign n2245 = ( n2125 & ~n2139 ) | ( n2125 & n2235 ) | ( ~n2139 & n2235 ) ;
  assign n2246 = ~n2244 & n2245 ;
  assign n2247 = n2240 | n2246 ;
  assign n2248 = n2082 &  n2140 ;
  assign n2241 = x69 | n2082 ;
  assign n2242 = x69 &  n2082 ;
  assign n2243 = ( n2241 & ~n2242 ) | ( n2241 & 1'b0 ) | ( ~n2242 & 1'b0 ) ;
  assign n2252 = ( n192 & n2124 ) | ( n192 & n2243 ) | ( n2124 & n2243 ) ;
  assign n2253 = ( n2124 & ~n2139 ) | ( n2124 & n2243 ) | ( ~n2139 & n2243 ) ;
  assign n2254 = ~n2252 & n2253 ;
  assign n2255 = n2248 | n2254 ;
  assign n2256 = n2090 &  n2140 ;
  assign n2249 = x68 | n2090 ;
  assign n2250 = x68 &  n2090 ;
  assign n2251 = ( n2249 & ~n2250 ) | ( n2249 & 1'b0 ) | ( ~n2250 & 1'b0 ) ;
  assign n2260 = ( n192 & n2123 ) | ( n192 & n2251 ) | ( n2123 & n2251 ) ;
  assign n2261 = ( n2123 & ~n2139 ) | ( n2123 & n2251 ) | ( ~n2139 & n2251 ) ;
  assign n2262 = ~n2260 & n2261 ;
  assign n2263 = n2256 | n2262 ;
  assign n2264 = n2099 &  n2140 ;
  assign n2257 = x67 | n2099 ;
  assign n2258 = x67 &  n2099 ;
  assign n2259 = ( n2257 & ~n2258 ) | ( n2257 & 1'b0 ) | ( ~n2258 & 1'b0 ) ;
  assign n2268 = ( n192 & n2122 ) | ( n192 & n2259 ) | ( n2122 & n2259 ) ;
  assign n2269 = ( n2122 & ~n2139 ) | ( n2122 & n2259 ) | ( ~n2139 & n2259 ) ;
  assign n2270 = ~n2268 & n2269 ;
  assign n2271 = n2264 | n2270 ;
  assign n2272 = n2105 &  n2140 ;
  assign n2265 = x66 | n2105 ;
  assign n2266 = x66 &  n2105 ;
  assign n2267 = ( n2265 & ~n2266 ) | ( n2265 & 1'b0 ) | ( ~n2266 & 1'b0 ) ;
  assign n2276 = ( n2121 & ~n192 ) | ( n2121 & n2267 ) | ( ~n192 & n2267 ) ;
  assign n2277 = ( n2121 & n2139 ) | ( n2121 & n2267 ) | ( n2139 & n2267 ) ;
  assign n2278 = ( n2276 & ~n2277 ) | ( n2276 & 1'b0 ) | ( ~n2277 & 1'b0 ) ;
  assign n2279 = n2272 | n2278 ;
  assign n2280 = n2119 &  n2140 ;
  assign n2273 = x65 &  n2119 ;
  assign n2274 = x65 | n2118 ;
  assign n2275 = n2112 | n2274 ;
  assign n2281 = ~n2273 & n2275 ;
  assign n2282 = ( n2120 & ~n2139 ) | ( n2120 & n2281 ) | ( ~n2139 & n2281 ) ;
  assign n2283 = ( n192 & n2120 ) | ( n192 & n2281 ) | ( n2120 & n2281 ) ;
  assign n2284 = ( n2282 & ~n2283 ) | ( n2282 & 1'b0 ) | ( ~n2283 & 1'b0 ) ;
  assign n2285 = n2280 | n2284 ;
  assign n2286 = ( x64 & ~x84 ) | ( x64 & 1'b0 ) | ( ~x84 & 1'b0 ) ;
  assign n2287 = ( n198 & ~n209 ) | ( n198 & n2286 ) | ( ~n209 & n2286 ) ;
  assign n2288 = ~n198 & n2287 ;
  assign n2289 = ( n240 & ~n255 ) | ( n240 & n2288 ) | ( ~n255 & n2288 ) ;
  assign n2290 = ~n240 & n2289 ;
  assign n2291 = n2139 &  n2290 ;
  assign n2292 = ( x44 & ~n2290 ) | ( x44 & n2291 ) | ( ~n2290 & n2291 ) ;
  assign n2293 = ~n181 & n2120 ;
  assign n2294 = ( n273 & ~n261 ) | ( n273 & n2293 ) | ( ~n261 & n2293 ) ;
  assign n2295 = ~n273 & n2294 ;
  assign n2296 = ~n270 & n2295 ;
  assign n2297 = ~n2139 & n2296 ;
  assign n2298 = n2292 | n2297 ;
  assign n2299 = ~x43 & x64 ;
  assign n2300 = ( x65 & ~n2298 ) | ( x65 & n2299 ) | ( ~n2298 & n2299 ) ;
  assign n2301 = ( x66 & ~n2285 ) | ( x66 & n2300 ) | ( ~n2285 & n2300 ) ;
  assign n2302 = ( x67 & ~n2279 ) | ( x67 & n2301 ) | ( ~n2279 & n2301 ) ;
  assign n2303 = ( x68 & ~n2271 ) | ( x68 & n2302 ) | ( ~n2271 & n2302 ) ;
  assign n2304 = ( x69 & ~n2263 ) | ( x69 & n2303 ) | ( ~n2263 & n2303 ) ;
  assign n2305 = ( x70 & ~n2255 ) | ( x70 & n2304 ) | ( ~n2255 & n2304 ) ;
  assign n2306 = ( x71 & ~n2247 ) | ( x71 & n2305 ) | ( ~n2247 & n2305 ) ;
  assign n2307 = ( x72 & ~n2239 ) | ( x72 & n2306 ) | ( ~n2239 & n2306 ) ;
  assign n2308 = ( x73 & ~n2231 ) | ( x73 & n2307 ) | ( ~n2231 & n2307 ) ;
  assign n2309 = ( x74 & ~n2223 ) | ( x74 & n2308 ) | ( ~n2223 & n2308 ) ;
  assign n2310 = ( x75 & ~n2215 ) | ( x75 & n2309 ) | ( ~n2215 & n2309 ) ;
  assign n2311 = ( x76 & ~n2207 ) | ( x76 & n2310 ) | ( ~n2207 & n2310 ) ;
  assign n2312 = ( x77 & ~n2199 ) | ( x77 & n2311 ) | ( ~n2199 & n2311 ) ;
  assign n2313 = ( x78 & ~n2191 ) | ( x78 & n2312 ) | ( ~n2191 & n2312 ) ;
  assign n2314 = ( x79 & ~n2183 ) | ( x79 & n2313 ) | ( ~n2183 & n2313 ) ;
  assign n2315 = ( x80 & ~n2175 ) | ( x80 & n2314 ) | ( ~n2175 & n2314 ) ;
  assign n2316 = ( x81 & ~n2167 ) | ( x81 & n2315 ) | ( ~n2167 & n2315 ) ;
  assign n2317 = ( x82 & ~n2159 ) | ( x82 & n2316 ) | ( ~n2159 & n2316 ) ;
  assign n2318 = ( x83 & ~n2151 ) | ( x83 & n2317 ) | ( ~n2151 & n2317 ) ;
  assign n2319 = n1978 &  n2140 ;
  assign n2320 = ( n192 & n1978 ) | ( n192 & n2138 ) | ( n1978 & n2138 ) ;
  assign n2321 = ( x83 & ~n2320 ) | ( x83 & n1978 ) | ( ~n2320 & n1978 ) ;
  assign n2322 = ~x83 & n2321 ;
  assign n2323 = n2319 | n2322 ;
  assign n2324 = ~x84 & n2323 ;
  assign n2325 = ( x84 & ~n2319 ) | ( x84 & 1'b0 ) | ( ~n2319 & 1'b0 ) ;
  assign n2326 = ~n2322 & n2325 ;
  assign n2327 = n462 | n2326 ;
  assign n2328 = n2324 | n2327 ;
  assign n2329 = n2318 | n2328 ;
  assign n2330 = ~n192 & n2323 ;
  assign n2344 = ( n2151 & ~n2330 ) | ( n2151 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2345 = n2329 &  n2344 ;
  assign n2332 = x83 | n2151 ;
  assign n2333 = x83 &  n2151 ;
  assign n2334 = ( n2332 & ~n2333 ) | ( n2332 & 1'b0 ) | ( ~n2333 & 1'b0 ) ;
  assign n2346 = n2317 &  n2334 ;
  assign n2331 = ( n2329 & ~n2330 ) | ( n2329 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2347 = ( n2317 & ~n2331 ) | ( n2317 & n2334 ) | ( ~n2331 & n2334 ) ;
  assign n2348 = ( n2345 & ~n2346 ) | ( n2345 & n2347 ) | ( ~n2346 & n2347 ) ;
  assign n2336 = n192 &  n1978 ;
  assign n2337 = n2329 &  n2336 ;
  assign n2335 = n2324 | n2326 ;
  assign n2339 = ( n2318 & n2331 ) | ( n2318 & n2335 ) | ( n2331 & n2335 ) ;
  assign n2338 = n2318 | n2335 ;
  assign n2340 = ( n2337 & ~n2339 ) | ( n2337 & n2338 ) | ( ~n2339 & n2338 ) ;
  assign n2352 = ( n2159 & ~n2330 ) | ( n2159 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2353 = n2329 &  n2352 ;
  assign n2341 = x82 | n2159 ;
  assign n2342 = x82 &  n2159 ;
  assign n2343 = ( n2341 & ~n2342 ) | ( n2341 & 1'b0 ) | ( ~n2342 & 1'b0 ) ;
  assign n2354 = n2316 &  n2343 ;
  assign n2355 = ( n2316 & ~n2331 ) | ( n2316 & n2343 ) | ( ~n2331 & n2343 ) ;
  assign n2356 = ( n2353 & ~n2354 ) | ( n2353 & n2355 ) | ( ~n2354 & n2355 ) ;
  assign n2360 = ( n2167 & ~n2330 ) | ( n2167 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2361 = n2329 &  n2360 ;
  assign n2349 = x81 | n2167 ;
  assign n2350 = x81 &  n2167 ;
  assign n2351 = ( n2349 & ~n2350 ) | ( n2349 & 1'b0 ) | ( ~n2350 & 1'b0 ) ;
  assign n2362 = n2315 &  n2351 ;
  assign n2363 = ( n2315 & ~n2331 ) | ( n2315 & n2351 ) | ( ~n2331 & n2351 ) ;
  assign n2364 = ( n2361 & ~n2362 ) | ( n2361 & n2363 ) | ( ~n2362 & n2363 ) ;
  assign n2368 = ( n2175 & ~n2330 ) | ( n2175 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2369 = n2329 &  n2368 ;
  assign n2357 = x80 | n2175 ;
  assign n2358 = x80 &  n2175 ;
  assign n2359 = ( n2357 & ~n2358 ) | ( n2357 & 1'b0 ) | ( ~n2358 & 1'b0 ) ;
  assign n2370 = n2314 &  n2359 ;
  assign n2371 = ( n2314 & ~n2331 ) | ( n2314 & n2359 ) | ( ~n2331 & n2359 ) ;
  assign n2372 = ( n2369 & ~n2370 ) | ( n2369 & n2371 ) | ( ~n2370 & n2371 ) ;
  assign n2376 = ( n2183 & ~n2330 ) | ( n2183 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2377 = n2329 &  n2376 ;
  assign n2365 = x79 | n2183 ;
  assign n2366 = x79 &  n2183 ;
  assign n2367 = ( n2365 & ~n2366 ) | ( n2365 & 1'b0 ) | ( ~n2366 & 1'b0 ) ;
  assign n2378 = n2313 &  n2367 ;
  assign n2379 = ( n2313 & ~n2331 ) | ( n2313 & n2367 ) | ( ~n2331 & n2367 ) ;
  assign n2380 = ( n2377 & ~n2378 ) | ( n2377 & n2379 ) | ( ~n2378 & n2379 ) ;
  assign n2384 = ( n2191 & ~n2330 ) | ( n2191 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2385 = n2329 &  n2384 ;
  assign n2373 = x78 | n2191 ;
  assign n2374 = x78 &  n2191 ;
  assign n2375 = ( n2373 & ~n2374 ) | ( n2373 & 1'b0 ) | ( ~n2374 & 1'b0 ) ;
  assign n2387 = ( n2312 & n2331 ) | ( n2312 & n2375 ) | ( n2331 & n2375 ) ;
  assign n2386 = n2312 | n2375 ;
  assign n2388 = ( n2385 & ~n2387 ) | ( n2385 & n2386 ) | ( ~n2387 & n2386 ) ;
  assign n2392 = ( n2199 & ~n2330 ) | ( n2199 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2393 = n2329 &  n2392 ;
  assign n2381 = x77 | n2199 ;
  assign n2382 = x77 &  n2199 ;
  assign n2383 = ( n2381 & ~n2382 ) | ( n2381 & 1'b0 ) | ( ~n2382 & 1'b0 ) ;
  assign n2395 = ( n2311 & n2331 ) | ( n2311 & n2383 ) | ( n2331 & n2383 ) ;
  assign n2394 = n2311 | n2383 ;
  assign n2396 = ( n2393 & ~n2395 ) | ( n2393 & n2394 ) | ( ~n2395 & n2394 ) ;
  assign n2400 = ( n2207 & ~n2330 ) | ( n2207 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2401 = n2329 &  n2400 ;
  assign n2389 = x76 | n2207 ;
  assign n2390 = x76 &  n2207 ;
  assign n2391 = ( n2389 & ~n2390 ) | ( n2389 & 1'b0 ) | ( ~n2390 & 1'b0 ) ;
  assign n2403 = ( n2310 & n2331 ) | ( n2310 & n2391 ) | ( n2331 & n2391 ) ;
  assign n2402 = n2310 | n2391 ;
  assign n2404 = ( n2401 & ~n2403 ) | ( n2401 & n2402 ) | ( ~n2403 & n2402 ) ;
  assign n2408 = ( n2215 & ~n2330 ) | ( n2215 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2409 = n2329 &  n2408 ;
  assign n2397 = x75 | n2215 ;
  assign n2398 = x75 &  n2215 ;
  assign n2399 = ( n2397 & ~n2398 ) | ( n2397 & 1'b0 ) | ( ~n2398 & 1'b0 ) ;
  assign n2411 = ( n2309 & n2331 ) | ( n2309 & n2399 ) | ( n2331 & n2399 ) ;
  assign n2410 = n2309 | n2399 ;
  assign n2412 = ( n2409 & ~n2411 ) | ( n2409 & n2410 ) | ( ~n2411 & n2410 ) ;
  assign n2416 = ( n2223 & ~n2330 ) | ( n2223 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2417 = n2329 &  n2416 ;
  assign n2405 = x74 | n2223 ;
  assign n2406 = x74 &  n2223 ;
  assign n2407 = ( n2405 & ~n2406 ) | ( n2405 & 1'b0 ) | ( ~n2406 & 1'b0 ) ;
  assign n2419 = ( n2308 & n2331 ) | ( n2308 & n2407 ) | ( n2331 & n2407 ) ;
  assign n2418 = n2308 | n2407 ;
  assign n2420 = ( n2417 & ~n2419 ) | ( n2417 & n2418 ) | ( ~n2419 & n2418 ) ;
  assign n2424 = ( n2231 & ~n2330 ) | ( n2231 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2425 = n2329 &  n2424 ;
  assign n2413 = x73 | n2231 ;
  assign n2414 = x73 &  n2231 ;
  assign n2415 = ( n2413 & ~n2414 ) | ( n2413 & 1'b0 ) | ( ~n2414 & 1'b0 ) ;
  assign n2427 = ( n2307 & n2331 ) | ( n2307 & n2415 ) | ( n2331 & n2415 ) ;
  assign n2426 = n2307 | n2415 ;
  assign n2428 = ( n2425 & ~n2427 ) | ( n2425 & n2426 ) | ( ~n2427 & n2426 ) ;
  assign n2432 = ( n2239 & ~n2330 ) | ( n2239 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2433 = n2329 &  n2432 ;
  assign n2421 = x72 | n2239 ;
  assign n2422 = x72 &  n2239 ;
  assign n2423 = ( n2421 & ~n2422 ) | ( n2421 & 1'b0 ) | ( ~n2422 & 1'b0 ) ;
  assign n2435 = ( n2306 & n2331 ) | ( n2306 & n2423 ) | ( n2331 & n2423 ) ;
  assign n2434 = n2306 | n2423 ;
  assign n2436 = ( n2433 & ~n2435 ) | ( n2433 & n2434 ) | ( ~n2435 & n2434 ) ;
  assign n2440 = ( n2247 & ~n2330 ) | ( n2247 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2441 = n2329 &  n2440 ;
  assign n2429 = x71 | n2247 ;
  assign n2430 = x71 &  n2247 ;
  assign n2431 = ( n2429 & ~n2430 ) | ( n2429 & 1'b0 ) | ( ~n2430 & 1'b0 ) ;
  assign n2443 = ( n2305 & n2331 ) | ( n2305 & n2431 ) | ( n2331 & n2431 ) ;
  assign n2442 = n2305 | n2431 ;
  assign n2444 = ( n2441 & ~n2443 ) | ( n2441 & n2442 ) | ( ~n2443 & n2442 ) ;
  assign n2448 = ( n2255 & ~n2330 ) | ( n2255 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2449 = n2329 &  n2448 ;
  assign n2437 = x70 | n2255 ;
  assign n2438 = x70 &  n2255 ;
  assign n2439 = ( n2437 & ~n2438 ) | ( n2437 & 1'b0 ) | ( ~n2438 & 1'b0 ) ;
  assign n2451 = ( n2304 & n2331 ) | ( n2304 & n2439 ) | ( n2331 & n2439 ) ;
  assign n2450 = n2304 | n2439 ;
  assign n2452 = ( n2449 & ~n2451 ) | ( n2449 & n2450 ) | ( ~n2451 & n2450 ) ;
  assign n2456 = ( n2263 & ~n2330 ) | ( n2263 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2457 = n2329 &  n2456 ;
  assign n2445 = x69 | n2263 ;
  assign n2446 = x69 &  n2263 ;
  assign n2447 = ( n2445 & ~n2446 ) | ( n2445 & 1'b0 ) | ( ~n2446 & 1'b0 ) ;
  assign n2459 = ( n2303 & n2331 ) | ( n2303 & n2447 ) | ( n2331 & n2447 ) ;
  assign n2458 = n2303 | n2447 ;
  assign n2460 = ( n2457 & ~n2459 ) | ( n2457 & n2458 ) | ( ~n2459 & n2458 ) ;
  assign n2464 = ( n2271 & ~n2330 ) | ( n2271 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2465 = n2329 &  n2464 ;
  assign n2453 = x68 | n2271 ;
  assign n2454 = x68 &  n2271 ;
  assign n2455 = ( n2453 & ~n2454 ) | ( n2453 & 1'b0 ) | ( ~n2454 & 1'b0 ) ;
  assign n2467 = ( n2302 & n2331 ) | ( n2302 & n2455 ) | ( n2331 & n2455 ) ;
  assign n2466 = n2302 | n2455 ;
  assign n2468 = ( n2465 & ~n2467 ) | ( n2465 & n2466 ) | ( ~n2467 & n2466 ) ;
  assign n2472 = ( n2279 & ~n2330 ) | ( n2279 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2473 = n2329 &  n2472 ;
  assign n2461 = x67 | n2279 ;
  assign n2462 = x67 &  n2279 ;
  assign n2463 = ( n2461 & ~n2462 ) | ( n2461 & 1'b0 ) | ( ~n2462 & 1'b0 ) ;
  assign n2475 = ( n2301 & n2331 ) | ( n2301 & n2463 ) | ( n2331 & n2463 ) ;
  assign n2474 = n2301 | n2463 ;
  assign n2476 = ( n2473 & ~n2475 ) | ( n2473 & n2474 ) | ( ~n2475 & n2474 ) ;
  assign n2477 = ( n2285 & ~n2330 ) | ( n2285 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2478 = n2329 &  n2477 ;
  assign n2469 = x66 | n2285 ;
  assign n2470 = x66 &  n2285 ;
  assign n2471 = ( n2469 & ~n2470 ) | ( n2469 & 1'b0 ) | ( ~n2470 & 1'b0 ) ;
  assign n2479 = n2300 &  n2471 ;
  assign n2480 = ( n2300 & ~n2331 ) | ( n2300 & n2471 ) | ( ~n2331 & n2471 ) ;
  assign n2481 = ( n2478 & ~n2479 ) | ( n2478 & n2480 ) | ( ~n2479 & n2480 ) ;
  assign n2482 = ( n2298 & ~x65 ) | ( n2298 & n2299 ) | ( ~x65 & n2299 ) ;
  assign n2483 = ( n2300 & ~n2299 ) | ( n2300 & n2482 ) | ( ~n2299 & n2482 ) ;
  assign n2484 = ~n2331 & n2483 ;
  assign n2485 = ( n2298 & ~n2330 ) | ( n2298 & 1'b0 ) | ( ~n2330 & 1'b0 ) ;
  assign n2486 = n2329 &  n2485 ;
  assign n2487 = n2484 | n2486 ;
  assign n2488 = ( x64 & ~n2331 ) | ( x64 & 1'b0 ) | ( ~n2331 & 1'b0 ) ;
  assign n2489 = ( x43 & ~n2488 ) | ( x43 & 1'b0 ) | ( ~n2488 & 1'b0 ) ;
  assign n2490 = ( n2299 & ~n2331 ) | ( n2299 & 1'b0 ) | ( ~n2331 & 1'b0 ) ;
  assign n2491 = n2489 | n2490 ;
  assign n2492 = ~x42 & x64 ;
  assign n2493 = ( x65 & ~n2491 ) | ( x65 & n2492 ) | ( ~n2491 & n2492 ) ;
  assign n2494 = ( x66 & ~n2487 ) | ( x66 & n2493 ) | ( ~n2487 & n2493 ) ;
  assign n2495 = ( x67 & ~n2481 ) | ( x67 & n2494 ) | ( ~n2481 & n2494 ) ;
  assign n2496 = ( x68 & ~n2476 ) | ( x68 & n2495 ) | ( ~n2476 & n2495 ) ;
  assign n2497 = ( x69 & ~n2468 ) | ( x69 & n2496 ) | ( ~n2468 & n2496 ) ;
  assign n2498 = ( x70 & ~n2460 ) | ( x70 & n2497 ) | ( ~n2460 & n2497 ) ;
  assign n2499 = ( x71 & ~n2452 ) | ( x71 & n2498 ) | ( ~n2452 & n2498 ) ;
  assign n2500 = ( x72 & ~n2444 ) | ( x72 & n2499 ) | ( ~n2444 & n2499 ) ;
  assign n2501 = ( x73 & ~n2436 ) | ( x73 & n2500 ) | ( ~n2436 & n2500 ) ;
  assign n2502 = ( x74 & ~n2428 ) | ( x74 & n2501 ) | ( ~n2428 & n2501 ) ;
  assign n2503 = ( x75 & ~n2420 ) | ( x75 & n2502 ) | ( ~n2420 & n2502 ) ;
  assign n2504 = ( x76 & ~n2412 ) | ( x76 & n2503 ) | ( ~n2412 & n2503 ) ;
  assign n2505 = ( x77 & ~n2404 ) | ( x77 & n2504 ) | ( ~n2404 & n2504 ) ;
  assign n2506 = ( x78 & ~n2396 ) | ( x78 & n2505 ) | ( ~n2396 & n2505 ) ;
  assign n2507 = ( x79 & ~n2388 ) | ( x79 & n2506 ) | ( ~n2388 & n2506 ) ;
  assign n2508 = ( x80 & ~n2380 ) | ( x80 & n2507 ) | ( ~n2380 & n2507 ) ;
  assign n2509 = ( x81 & ~n2372 ) | ( x81 & n2508 ) | ( ~n2372 & n2508 ) ;
  assign n2510 = ( x82 & ~n2364 ) | ( x82 & n2509 ) | ( ~n2364 & n2509 ) ;
  assign n2511 = ( x83 & ~n2356 ) | ( x83 & n2510 ) | ( ~n2356 & n2510 ) ;
  assign n2512 = ( x84 & ~n2348 ) | ( x84 & n2511 ) | ( ~n2348 & n2511 ) ;
  assign n2513 = ( x85 & ~n2340 ) | ( x85 & n2512 ) | ( ~n2340 & n2512 ) ;
  assign n2514 = n178 | n180 ;
  assign n2515 = ( n189 & ~n175 ) | ( n189 & n2514 ) | ( ~n175 & n2514 ) ;
  assign n2516 = n175 | n2515 ;
  assign n2517 = n160 | n2516 ;
  assign n2518 = n2513 | n2517 ;
  assign n2525 = n2348 &  n2518 ;
  assign n2519 = x84 | n2348 ;
  assign n2520 = x84 &  n2348 ;
  assign n2521 = ( n2519 & ~n2520 ) | ( n2519 & 1'b0 ) | ( ~n2520 & 1'b0 ) ;
  assign n2529 = ( n2511 & n2513 ) | ( n2511 & n2521 ) | ( n2513 & n2521 ) ;
  assign n2530 = ( n2511 & ~n2517 ) | ( n2511 & n2521 ) | ( ~n2517 & n2521 ) ;
  assign n2531 = ~n2529 & n2530 ;
  assign n2532 = n2525 | n2531 ;
  assign n2522 = x85 | n2512 ;
  assign n2523 = ( x85 & n2512 ) | ( x85 & n2517 ) | ( n2512 & n2517 ) ;
  assign n2524 = ( n2340 & ~n2522 ) | ( n2340 & n2523 ) | ( ~n2522 & n2523 ) ;
  assign n2533 = n2356 &  n2518 ;
  assign n2526 = x83 | n2356 ;
  assign n2527 = x83 &  n2356 ;
  assign n2528 = ( n2526 & ~n2527 ) | ( n2526 & 1'b0 ) | ( ~n2527 & 1'b0 ) ;
  assign n2537 = ( n2510 & n2513 ) | ( n2510 & n2528 ) | ( n2513 & n2528 ) ;
  assign n2538 = ( n2510 & ~n2517 ) | ( n2510 & n2528 ) | ( ~n2517 & n2528 ) ;
  assign n2539 = ~n2537 & n2538 ;
  assign n2540 = n2533 | n2539 ;
  assign n2541 = n2364 &  n2518 ;
  assign n2534 = x82 | n2364 ;
  assign n2535 = x82 &  n2364 ;
  assign n2536 = ( n2534 & ~n2535 ) | ( n2534 & 1'b0 ) | ( ~n2535 & 1'b0 ) ;
  assign n2545 = ( n2509 & n2513 ) | ( n2509 & n2536 ) | ( n2513 & n2536 ) ;
  assign n2546 = ( n2509 & ~n2517 ) | ( n2509 & n2536 ) | ( ~n2517 & n2536 ) ;
  assign n2547 = ~n2545 & n2546 ;
  assign n2548 = n2541 | n2547 ;
  assign n2549 = n2372 &  n2518 ;
  assign n2542 = x81 | n2372 ;
  assign n2543 = x81 &  n2372 ;
  assign n2544 = ( n2542 & ~n2543 ) | ( n2542 & 1'b0 ) | ( ~n2543 & 1'b0 ) ;
  assign n2553 = ( n2508 & n2513 ) | ( n2508 & n2544 ) | ( n2513 & n2544 ) ;
  assign n2554 = ( n2508 & ~n2517 ) | ( n2508 & n2544 ) | ( ~n2517 & n2544 ) ;
  assign n2555 = ~n2553 & n2554 ;
  assign n2556 = n2549 | n2555 ;
  assign n2557 = n2380 &  n2518 ;
  assign n2550 = x80 | n2380 ;
  assign n2551 = x80 &  n2380 ;
  assign n2552 = ( n2550 & ~n2551 ) | ( n2550 & 1'b0 ) | ( ~n2551 & 1'b0 ) ;
  assign n2561 = ( n2507 & n2513 ) | ( n2507 & n2552 ) | ( n2513 & n2552 ) ;
  assign n2562 = ( n2507 & ~n2517 ) | ( n2507 & n2552 ) | ( ~n2517 & n2552 ) ;
  assign n2563 = ~n2561 & n2562 ;
  assign n2564 = n2557 | n2563 ;
  assign n2565 = n2388 &  n2518 ;
  assign n2558 = x79 | n2388 ;
  assign n2559 = x79 &  n2388 ;
  assign n2560 = ( n2558 & ~n2559 ) | ( n2558 & 1'b0 ) | ( ~n2559 & 1'b0 ) ;
  assign n2569 = ( n2506 & n2513 ) | ( n2506 & n2560 ) | ( n2513 & n2560 ) ;
  assign n2570 = ( n2506 & ~n2517 ) | ( n2506 & n2560 ) | ( ~n2517 & n2560 ) ;
  assign n2571 = ~n2569 & n2570 ;
  assign n2572 = n2565 | n2571 ;
  assign n2573 = n2396 &  n2518 ;
  assign n2566 = x78 | n2396 ;
  assign n2567 = x78 &  n2396 ;
  assign n2568 = ( n2566 & ~n2567 ) | ( n2566 & 1'b0 ) | ( ~n2567 & 1'b0 ) ;
  assign n2577 = ( n2505 & n2513 ) | ( n2505 & n2568 ) | ( n2513 & n2568 ) ;
  assign n2578 = ( n2505 & ~n2517 ) | ( n2505 & n2568 ) | ( ~n2517 & n2568 ) ;
  assign n2579 = ~n2577 & n2578 ;
  assign n2580 = n2573 | n2579 ;
  assign n2581 = n2404 &  n2518 ;
  assign n2574 = x77 | n2404 ;
  assign n2575 = x77 &  n2404 ;
  assign n2576 = ( n2574 & ~n2575 ) | ( n2574 & 1'b0 ) | ( ~n2575 & 1'b0 ) ;
  assign n2585 = ( n2504 & n2513 ) | ( n2504 & n2576 ) | ( n2513 & n2576 ) ;
  assign n2586 = ( n2504 & ~n2517 ) | ( n2504 & n2576 ) | ( ~n2517 & n2576 ) ;
  assign n2587 = ~n2585 & n2586 ;
  assign n2588 = n2581 | n2587 ;
  assign n2589 = n2412 &  n2518 ;
  assign n2582 = x76 | n2412 ;
  assign n2583 = x76 &  n2412 ;
  assign n2584 = ( n2582 & ~n2583 ) | ( n2582 & 1'b0 ) | ( ~n2583 & 1'b0 ) ;
  assign n2593 = ( n2503 & n2513 ) | ( n2503 & n2584 ) | ( n2513 & n2584 ) ;
  assign n2594 = ( n2503 & ~n2517 ) | ( n2503 & n2584 ) | ( ~n2517 & n2584 ) ;
  assign n2595 = ~n2593 & n2594 ;
  assign n2596 = n2589 | n2595 ;
  assign n2597 = n2420 &  n2518 ;
  assign n2590 = x75 | n2420 ;
  assign n2591 = x75 &  n2420 ;
  assign n2592 = ( n2590 & ~n2591 ) | ( n2590 & 1'b0 ) | ( ~n2591 & 1'b0 ) ;
  assign n2601 = ( n2502 & n2513 ) | ( n2502 & n2592 ) | ( n2513 & n2592 ) ;
  assign n2602 = ( n2502 & ~n2517 ) | ( n2502 & n2592 ) | ( ~n2517 & n2592 ) ;
  assign n2603 = ~n2601 & n2602 ;
  assign n2604 = n2597 | n2603 ;
  assign n2605 = n2428 &  n2518 ;
  assign n2598 = x74 | n2428 ;
  assign n2599 = x74 &  n2428 ;
  assign n2600 = ( n2598 & ~n2599 ) | ( n2598 & 1'b0 ) | ( ~n2599 & 1'b0 ) ;
  assign n2609 = ( n2501 & n2513 ) | ( n2501 & n2600 ) | ( n2513 & n2600 ) ;
  assign n2610 = ( n2501 & ~n2517 ) | ( n2501 & n2600 ) | ( ~n2517 & n2600 ) ;
  assign n2611 = ~n2609 & n2610 ;
  assign n2612 = n2605 | n2611 ;
  assign n2613 = n2436 &  n2518 ;
  assign n2606 = x73 | n2436 ;
  assign n2607 = x73 &  n2436 ;
  assign n2608 = ( n2606 & ~n2607 ) | ( n2606 & 1'b0 ) | ( ~n2607 & 1'b0 ) ;
  assign n2617 = ( n2500 & n2513 ) | ( n2500 & n2608 ) | ( n2513 & n2608 ) ;
  assign n2618 = ( n2500 & ~n2517 ) | ( n2500 & n2608 ) | ( ~n2517 & n2608 ) ;
  assign n2619 = ~n2617 & n2618 ;
  assign n2620 = n2613 | n2619 ;
  assign n2621 = n2444 &  n2518 ;
  assign n2614 = x72 | n2444 ;
  assign n2615 = x72 &  n2444 ;
  assign n2616 = ( n2614 & ~n2615 ) | ( n2614 & 1'b0 ) | ( ~n2615 & 1'b0 ) ;
  assign n2625 = ( n2499 & n2513 ) | ( n2499 & n2616 ) | ( n2513 & n2616 ) ;
  assign n2626 = ( n2499 & ~n2517 ) | ( n2499 & n2616 ) | ( ~n2517 & n2616 ) ;
  assign n2627 = ~n2625 & n2626 ;
  assign n2628 = n2621 | n2627 ;
  assign n2629 = n2452 &  n2518 ;
  assign n2622 = x71 | n2452 ;
  assign n2623 = x71 &  n2452 ;
  assign n2624 = ( n2622 & ~n2623 ) | ( n2622 & 1'b0 ) | ( ~n2623 & 1'b0 ) ;
  assign n2633 = ( n2498 & n2513 ) | ( n2498 & n2624 ) | ( n2513 & n2624 ) ;
  assign n2634 = ( n2498 & ~n2517 ) | ( n2498 & n2624 ) | ( ~n2517 & n2624 ) ;
  assign n2635 = ~n2633 & n2634 ;
  assign n2636 = n2629 | n2635 ;
  assign n2637 = n2460 &  n2518 ;
  assign n2630 = x70 | n2460 ;
  assign n2631 = x70 &  n2460 ;
  assign n2632 = ( n2630 & ~n2631 ) | ( n2630 & 1'b0 ) | ( ~n2631 & 1'b0 ) ;
  assign n2641 = ( n2497 & n2513 ) | ( n2497 & n2632 ) | ( n2513 & n2632 ) ;
  assign n2642 = ( n2497 & ~n2517 ) | ( n2497 & n2632 ) | ( ~n2517 & n2632 ) ;
  assign n2643 = ~n2641 & n2642 ;
  assign n2644 = n2637 | n2643 ;
  assign n2645 = n2468 &  n2518 ;
  assign n2638 = x69 | n2468 ;
  assign n2639 = x69 &  n2468 ;
  assign n2640 = ( n2638 & ~n2639 ) | ( n2638 & 1'b0 ) | ( ~n2639 & 1'b0 ) ;
  assign n2649 = ( n2496 & n2513 ) | ( n2496 & n2640 ) | ( n2513 & n2640 ) ;
  assign n2650 = ( n2496 & ~n2517 ) | ( n2496 & n2640 ) | ( ~n2517 & n2640 ) ;
  assign n2651 = ~n2649 & n2650 ;
  assign n2652 = n2645 | n2651 ;
  assign n2653 = n2476 &  n2518 ;
  assign n2646 = x68 | n2476 ;
  assign n2647 = x68 &  n2476 ;
  assign n2648 = ( n2646 & ~n2647 ) | ( n2646 & 1'b0 ) | ( ~n2647 & 1'b0 ) ;
  assign n2657 = ( n2495 & n2513 ) | ( n2495 & n2648 ) | ( n2513 & n2648 ) ;
  assign n2658 = ( n2495 & ~n2517 ) | ( n2495 & n2648 ) | ( ~n2517 & n2648 ) ;
  assign n2659 = ~n2657 & n2658 ;
  assign n2660 = n2653 | n2659 ;
  assign n2661 = n2481 &  n2518 ;
  assign n2654 = x67 | n2481 ;
  assign n2655 = x67 &  n2481 ;
  assign n2656 = ( n2654 & ~n2655 ) | ( n2654 & 1'b0 ) | ( ~n2655 & 1'b0 ) ;
  assign n2665 = ( n2494 & n2513 ) | ( n2494 & n2656 ) | ( n2513 & n2656 ) ;
  assign n2666 = ( n2494 & ~n2517 ) | ( n2494 & n2656 ) | ( ~n2517 & n2656 ) ;
  assign n2667 = ~n2665 & n2666 ;
  assign n2668 = n2661 | n2667 ;
  assign n2669 = n2487 &  n2518 ;
  assign n2662 = x66 | n2487 ;
  assign n2663 = x66 &  n2487 ;
  assign n2664 = ( n2662 & ~n2663 ) | ( n2662 & 1'b0 ) | ( ~n2663 & 1'b0 ) ;
  assign n2674 = ( n2493 & ~n2513 ) | ( n2493 & n2664 ) | ( ~n2513 & n2664 ) ;
  assign n2675 = ( n2493 & n2517 ) | ( n2493 & n2664 ) | ( n2517 & n2664 ) ;
  assign n2676 = ( n2674 & ~n2675 ) | ( n2674 & 1'b0 ) | ( ~n2675 & 1'b0 ) ;
  assign n2677 = n2669 | n2676 ;
  assign n2678 = n2491 &  n2518 ;
  assign n2670 = x65 &  n2491 ;
  assign n2671 = ( n2489 & ~x65 ) | ( n2489 & n2490 ) | ( ~x65 & n2490 ) ;
  assign n2672 = x65 | n2671 ;
  assign n2673 = ( n2492 & ~n2670 ) | ( n2492 & n2672 ) | ( ~n2670 & n2672 ) ;
  assign n2679 = ( x65 & n2491 ) | ( x65 & n2492 ) | ( n2491 & n2492 ) ;
  assign n2680 = ( n2517 & ~n2670 ) | ( n2517 & n2679 ) | ( ~n2670 & n2679 ) ;
  assign n2681 = ( n2513 & n2673 ) | ( n2513 & n2680 ) | ( n2673 & n2680 ) ;
  assign n2682 = ( n2673 & ~n2681 ) | ( n2673 & 1'b0 ) | ( ~n2681 & 1'b0 ) ;
  assign n2683 = n2678 | n2682 ;
  assign n2684 = ( x64 & ~x86 ) | ( x64 & 1'b0 ) | ( ~x86 & 1'b0 ) ;
  assign n2685 = ( n197 & ~n208 ) | ( n197 & n2684 ) | ( ~n208 & n2684 ) ;
  assign n2686 = ~n197 & n2685 ;
  assign n2687 = ( n419 & ~n428 ) | ( n419 & n2686 ) | ( ~n428 & n2686 ) ;
  assign n2688 = ~n419 & n2687 ;
  assign n2689 = ~n425 & n2688 ;
  assign n2690 = n2513 &  n2689 ;
  assign n2691 = ( x42 & ~n2689 ) | ( x42 & n2690 ) | ( ~n2689 & n2690 ) ;
  assign n2692 = ~n180 & n2492 ;
  assign n2693 = ( n178 & ~n189 ) | ( n178 & n2692 ) | ( ~n189 & n2692 ) ;
  assign n2694 = ~n178 & n2693 ;
  assign n2695 = ( n160 & ~n175 ) | ( n160 & n2694 ) | ( ~n175 & n2694 ) ;
  assign n2696 = ~n160 & n2695 ;
  assign n2697 = ~n2513 & n2696 ;
  assign n2698 = n2691 | n2697 ;
  assign n2699 = ~x41 & x64 ;
  assign n2700 = ( x65 & ~n2698 ) | ( x65 & n2699 ) | ( ~n2698 & n2699 ) ;
  assign n2701 = ( x66 & ~n2683 ) | ( x66 & n2700 ) | ( ~n2683 & n2700 ) ;
  assign n2702 = ( x67 & ~n2677 ) | ( x67 & n2701 ) | ( ~n2677 & n2701 ) ;
  assign n2703 = ( x68 & ~n2668 ) | ( x68 & n2702 ) | ( ~n2668 & n2702 ) ;
  assign n2704 = ( x69 & ~n2660 ) | ( x69 & n2703 ) | ( ~n2660 & n2703 ) ;
  assign n2705 = ( x70 & ~n2652 ) | ( x70 & n2704 ) | ( ~n2652 & n2704 ) ;
  assign n2706 = ( x71 & ~n2644 ) | ( x71 & n2705 ) | ( ~n2644 & n2705 ) ;
  assign n2707 = ( x72 & ~n2636 ) | ( x72 & n2706 ) | ( ~n2636 & n2706 ) ;
  assign n2708 = ( x73 & ~n2628 ) | ( x73 & n2707 ) | ( ~n2628 & n2707 ) ;
  assign n2709 = ( x74 & ~n2620 ) | ( x74 & n2708 ) | ( ~n2620 & n2708 ) ;
  assign n2710 = ( x75 & ~n2612 ) | ( x75 & n2709 ) | ( ~n2612 & n2709 ) ;
  assign n2711 = ( x76 & ~n2604 ) | ( x76 & n2710 ) | ( ~n2604 & n2710 ) ;
  assign n2712 = ( x77 & ~n2596 ) | ( x77 & n2711 ) | ( ~n2596 & n2711 ) ;
  assign n2713 = ( x78 & ~n2588 ) | ( x78 & n2712 ) | ( ~n2588 & n2712 ) ;
  assign n2714 = ( x79 & ~n2580 ) | ( x79 & n2713 ) | ( ~n2580 & n2713 ) ;
  assign n2715 = ( x80 & ~n2572 ) | ( x80 & n2714 ) | ( ~n2572 & n2714 ) ;
  assign n2716 = ( x81 & ~n2564 ) | ( x81 & n2715 ) | ( ~n2564 & n2715 ) ;
  assign n2717 = ( x82 & ~n2556 ) | ( x82 & n2716 ) | ( ~n2556 & n2716 ) ;
  assign n2718 = ( x83 & ~n2548 ) | ( x83 & n2717 ) | ( ~n2548 & n2717 ) ;
  assign n2719 = ( x84 & ~n2540 ) | ( x84 & n2718 ) | ( ~n2540 & n2718 ) ;
  assign n2720 = ( x85 & ~n2532 ) | ( x85 & n2719 ) | ( ~n2532 & n2719 ) ;
  assign n2721 = ( x86 & ~n2524 ) | ( x86 & n2720 ) | ( ~n2524 & n2720 ) ;
  assign n2738 = n197 | n208 ;
  assign n2739 = ( n428 & ~n419 ) | ( n428 & n2738 ) | ( ~n419 & n2738 ) ;
  assign n2740 = n419 | n2739 ;
  assign n2741 = n425 | n2740 ;
  assign n2742 = n2721 | n2741 ;
  assign n2756 = n2532 &  n2742 ;
  assign n2760 = x85 | n2532 ;
  assign n2761 = x85 &  n2532 ;
  assign n2762 = ( n2760 & ~n2761 ) | ( n2760 & 1'b0 ) | ( ~n2761 & 1'b0 ) ;
  assign n2763 = ( n2719 & n2721 ) | ( n2719 & n2762 ) | ( n2721 & n2762 ) ;
  assign n2764 = ( n2719 & ~n2741 ) | ( n2719 & n2762 ) | ( ~n2741 & n2762 ) ;
  assign n2765 = ~n2763 & n2764 ;
  assign n2766 = n2756 | n2765 ;
  assign n2767 = n2540 &  n2742 ;
  assign n2757 = x84 | n2540 ;
  assign n2758 = x84 &  n2540 ;
  assign n2759 = ( n2757 & ~n2758 ) | ( n2757 & 1'b0 ) | ( ~n2758 & 1'b0 ) ;
  assign n2771 = ( n2718 & n2721 ) | ( n2718 & n2759 ) | ( n2721 & n2759 ) ;
  assign n2772 = ( n2718 & ~n2741 ) | ( n2718 & n2759 ) | ( ~n2741 & n2759 ) ;
  assign n2773 = ~n2771 & n2772 ;
  assign n2774 = n2767 | n2773 ;
  assign n2775 = n2548 &  n2742 ;
  assign n2768 = x83 | n2548 ;
  assign n2769 = x83 &  n2548 ;
  assign n2770 = ( n2768 & ~n2769 ) | ( n2768 & 1'b0 ) | ( ~n2769 & 1'b0 ) ;
  assign n2779 = ( n2717 & n2721 ) | ( n2717 & n2770 ) | ( n2721 & n2770 ) ;
  assign n2780 = ( n2717 & ~n2741 ) | ( n2717 & n2770 ) | ( ~n2741 & n2770 ) ;
  assign n2781 = ~n2779 & n2780 ;
  assign n2782 = n2775 | n2781 ;
  assign n2783 = n2556 &  n2742 ;
  assign n2776 = x82 | n2556 ;
  assign n2777 = x82 &  n2556 ;
  assign n2778 = ( n2776 & ~n2777 ) | ( n2776 & 1'b0 ) | ( ~n2777 & 1'b0 ) ;
  assign n2787 = ( n2716 & n2721 ) | ( n2716 & n2778 ) | ( n2721 & n2778 ) ;
  assign n2788 = ( n2716 & ~n2741 ) | ( n2716 & n2778 ) | ( ~n2741 & n2778 ) ;
  assign n2789 = ~n2787 & n2788 ;
  assign n2790 = n2783 | n2789 ;
  assign n2791 = n2564 &  n2742 ;
  assign n2784 = x81 | n2564 ;
  assign n2785 = x81 &  n2564 ;
  assign n2786 = ( n2784 & ~n2785 ) | ( n2784 & 1'b0 ) | ( ~n2785 & 1'b0 ) ;
  assign n2795 = ( n2715 & n2721 ) | ( n2715 & n2786 ) | ( n2721 & n2786 ) ;
  assign n2796 = ( n2715 & ~n2741 ) | ( n2715 & n2786 ) | ( ~n2741 & n2786 ) ;
  assign n2797 = ~n2795 & n2796 ;
  assign n2798 = n2791 | n2797 ;
  assign n2799 = n2572 &  n2742 ;
  assign n2792 = x80 | n2572 ;
  assign n2793 = x80 &  n2572 ;
  assign n2794 = ( n2792 & ~n2793 ) | ( n2792 & 1'b0 ) | ( ~n2793 & 1'b0 ) ;
  assign n2803 = ( n2714 & n2721 ) | ( n2714 & n2794 ) | ( n2721 & n2794 ) ;
  assign n2804 = ( n2714 & ~n2741 ) | ( n2714 & n2794 ) | ( ~n2741 & n2794 ) ;
  assign n2805 = ~n2803 & n2804 ;
  assign n2806 = n2799 | n2805 ;
  assign n2807 = n2580 &  n2742 ;
  assign n2800 = x79 | n2580 ;
  assign n2801 = x79 &  n2580 ;
  assign n2802 = ( n2800 & ~n2801 ) | ( n2800 & 1'b0 ) | ( ~n2801 & 1'b0 ) ;
  assign n2811 = ( n2713 & n2721 ) | ( n2713 & n2802 ) | ( n2721 & n2802 ) ;
  assign n2812 = ( n2713 & ~n2741 ) | ( n2713 & n2802 ) | ( ~n2741 & n2802 ) ;
  assign n2813 = ~n2811 & n2812 ;
  assign n2814 = n2807 | n2813 ;
  assign n2815 = n2588 &  n2742 ;
  assign n2808 = x78 | n2588 ;
  assign n2809 = x78 &  n2588 ;
  assign n2810 = ( n2808 & ~n2809 ) | ( n2808 & 1'b0 ) | ( ~n2809 & 1'b0 ) ;
  assign n2819 = ( n2712 & n2721 ) | ( n2712 & n2810 ) | ( n2721 & n2810 ) ;
  assign n2820 = ( n2712 & ~n2741 ) | ( n2712 & n2810 ) | ( ~n2741 & n2810 ) ;
  assign n2821 = ~n2819 & n2820 ;
  assign n2822 = n2815 | n2821 ;
  assign n2823 = n2596 &  n2742 ;
  assign n2816 = x77 | n2596 ;
  assign n2817 = x77 &  n2596 ;
  assign n2818 = ( n2816 & ~n2817 ) | ( n2816 & 1'b0 ) | ( ~n2817 & 1'b0 ) ;
  assign n2827 = ( n2711 & n2721 ) | ( n2711 & n2818 ) | ( n2721 & n2818 ) ;
  assign n2828 = ( n2711 & ~n2741 ) | ( n2711 & n2818 ) | ( ~n2741 & n2818 ) ;
  assign n2829 = ~n2827 & n2828 ;
  assign n2830 = n2823 | n2829 ;
  assign n2831 = n2604 &  n2742 ;
  assign n2824 = x76 | n2604 ;
  assign n2825 = x76 &  n2604 ;
  assign n2826 = ( n2824 & ~n2825 ) | ( n2824 & 1'b0 ) | ( ~n2825 & 1'b0 ) ;
  assign n2835 = ( n2710 & n2721 ) | ( n2710 & n2826 ) | ( n2721 & n2826 ) ;
  assign n2836 = ( n2710 & ~n2741 ) | ( n2710 & n2826 ) | ( ~n2741 & n2826 ) ;
  assign n2837 = ~n2835 & n2836 ;
  assign n2838 = n2831 | n2837 ;
  assign n2839 = n2612 &  n2742 ;
  assign n2832 = x75 | n2612 ;
  assign n2833 = x75 &  n2612 ;
  assign n2834 = ( n2832 & ~n2833 ) | ( n2832 & 1'b0 ) | ( ~n2833 & 1'b0 ) ;
  assign n2843 = ( n2709 & n2721 ) | ( n2709 & n2834 ) | ( n2721 & n2834 ) ;
  assign n2844 = ( n2709 & ~n2741 ) | ( n2709 & n2834 ) | ( ~n2741 & n2834 ) ;
  assign n2845 = ~n2843 & n2844 ;
  assign n2846 = n2839 | n2845 ;
  assign n2847 = n2620 &  n2742 ;
  assign n2840 = x74 | n2620 ;
  assign n2841 = x74 &  n2620 ;
  assign n2842 = ( n2840 & ~n2841 ) | ( n2840 & 1'b0 ) | ( ~n2841 & 1'b0 ) ;
  assign n2851 = ( n2708 & n2721 ) | ( n2708 & n2842 ) | ( n2721 & n2842 ) ;
  assign n2852 = ( n2708 & ~n2741 ) | ( n2708 & n2842 ) | ( ~n2741 & n2842 ) ;
  assign n2853 = ~n2851 & n2852 ;
  assign n2854 = n2847 | n2853 ;
  assign n2855 = n2628 &  n2742 ;
  assign n2848 = x73 | n2628 ;
  assign n2849 = x73 &  n2628 ;
  assign n2850 = ( n2848 & ~n2849 ) | ( n2848 & 1'b0 ) | ( ~n2849 & 1'b0 ) ;
  assign n2859 = ( n2707 & n2721 ) | ( n2707 & n2850 ) | ( n2721 & n2850 ) ;
  assign n2860 = ( n2707 & ~n2741 ) | ( n2707 & n2850 ) | ( ~n2741 & n2850 ) ;
  assign n2861 = ~n2859 & n2860 ;
  assign n2862 = n2855 | n2861 ;
  assign n2863 = n2636 &  n2742 ;
  assign n2856 = x72 | n2636 ;
  assign n2857 = x72 &  n2636 ;
  assign n2858 = ( n2856 & ~n2857 ) | ( n2856 & 1'b0 ) | ( ~n2857 & 1'b0 ) ;
  assign n2867 = ( n2706 & n2721 ) | ( n2706 & n2858 ) | ( n2721 & n2858 ) ;
  assign n2868 = ( n2706 & ~n2741 ) | ( n2706 & n2858 ) | ( ~n2741 & n2858 ) ;
  assign n2869 = ~n2867 & n2868 ;
  assign n2870 = n2863 | n2869 ;
  assign n2871 = n2644 &  n2742 ;
  assign n2864 = x71 | n2644 ;
  assign n2865 = x71 &  n2644 ;
  assign n2866 = ( n2864 & ~n2865 ) | ( n2864 & 1'b0 ) | ( ~n2865 & 1'b0 ) ;
  assign n2875 = ( n2705 & n2721 ) | ( n2705 & n2866 ) | ( n2721 & n2866 ) ;
  assign n2876 = ( n2705 & ~n2741 ) | ( n2705 & n2866 ) | ( ~n2741 & n2866 ) ;
  assign n2877 = ~n2875 & n2876 ;
  assign n2878 = n2871 | n2877 ;
  assign n2879 = n2652 &  n2742 ;
  assign n2872 = x70 | n2652 ;
  assign n2873 = x70 &  n2652 ;
  assign n2874 = ( n2872 & ~n2873 ) | ( n2872 & 1'b0 ) | ( ~n2873 & 1'b0 ) ;
  assign n2883 = ( n2704 & n2721 ) | ( n2704 & n2874 ) | ( n2721 & n2874 ) ;
  assign n2884 = ( n2704 & ~n2741 ) | ( n2704 & n2874 ) | ( ~n2741 & n2874 ) ;
  assign n2885 = ~n2883 & n2884 ;
  assign n2886 = n2879 | n2885 ;
  assign n2887 = n2660 &  n2742 ;
  assign n2880 = x69 | n2660 ;
  assign n2881 = x69 &  n2660 ;
  assign n2882 = ( n2880 & ~n2881 ) | ( n2880 & 1'b0 ) | ( ~n2881 & 1'b0 ) ;
  assign n2891 = ( n2703 & n2721 ) | ( n2703 & n2882 ) | ( n2721 & n2882 ) ;
  assign n2892 = ( n2703 & ~n2741 ) | ( n2703 & n2882 ) | ( ~n2741 & n2882 ) ;
  assign n2893 = ~n2891 & n2892 ;
  assign n2894 = n2887 | n2893 ;
  assign n2895 = n2668 &  n2742 ;
  assign n2888 = x68 | n2668 ;
  assign n2889 = x68 &  n2668 ;
  assign n2890 = ( n2888 & ~n2889 ) | ( n2888 & 1'b0 ) | ( ~n2889 & 1'b0 ) ;
  assign n2899 = ( n2702 & n2721 ) | ( n2702 & n2890 ) | ( n2721 & n2890 ) ;
  assign n2900 = ( n2702 & ~n2741 ) | ( n2702 & n2890 ) | ( ~n2741 & n2890 ) ;
  assign n2901 = ~n2899 & n2900 ;
  assign n2902 = n2895 | n2901 ;
  assign n2903 = n2677 &  n2742 ;
  assign n2896 = x67 | n2677 ;
  assign n2897 = x67 &  n2677 ;
  assign n2898 = ( n2896 & ~n2897 ) | ( n2896 & 1'b0 ) | ( ~n2897 & 1'b0 ) ;
  assign n2907 = ( n2701 & n2721 ) | ( n2701 & n2898 ) | ( n2721 & n2898 ) ;
  assign n2908 = ( n2701 & ~n2741 ) | ( n2701 & n2898 ) | ( ~n2741 & n2898 ) ;
  assign n2909 = ~n2907 & n2908 ;
  assign n2910 = n2903 | n2909 ;
  assign n2911 = n2683 &  n2742 ;
  assign n2904 = x66 | n2683 ;
  assign n2905 = x66 &  n2683 ;
  assign n2906 = ( n2904 & ~n2905 ) | ( n2904 & 1'b0 ) | ( ~n2905 & 1'b0 ) ;
  assign n2912 = ( n2700 & ~n2721 ) | ( n2700 & n2906 ) | ( ~n2721 & n2906 ) ;
  assign n2913 = ( n2700 & n2741 ) | ( n2700 & n2906 ) | ( n2741 & n2906 ) ;
  assign n2914 = ( n2912 & ~n2913 ) | ( n2912 & 1'b0 ) | ( ~n2913 & 1'b0 ) ;
  assign n2915 = n2911 | n2914 ;
  assign n2743 = n2698 &  n2742 ;
  assign n2744 = x65 &  n2698 ;
  assign n2745 = x65 | n2697 ;
  assign n2746 = n2691 | n2745 ;
  assign n2747 = ( n2699 & ~n2744 ) | ( n2699 & n2746 ) | ( ~n2744 & n2746 ) ;
  assign n2748 = ( x65 & n2698 ) | ( x65 & n2699 ) | ( n2698 & n2699 ) ;
  assign n2749 = ( n2741 & ~n2744 ) | ( n2741 & n2748 ) | ( ~n2744 & n2748 ) ;
  assign n2750 = ( n2721 & n2747 ) | ( n2721 & n2749 ) | ( n2747 & n2749 ) ;
  assign n2751 = ( n2747 & ~n2750 ) | ( n2747 & 1'b0 ) | ( ~n2750 & 1'b0 ) ;
  assign n2752 = n2743 | n2751 ;
  assign n2722 = ( x64 & ~x87 ) | ( x64 & 1'b0 ) | ( ~x87 & 1'b0 ) ;
  assign n2723 = ( n178 & ~n189 ) | ( n178 & n2722 ) | ( ~n189 & n2722 ) ;
  assign n2724 = ~n178 & n2723 ;
  assign n2725 = ( n160 & ~n175 ) | ( n160 & n2724 ) | ( ~n175 & n2724 ) ;
  assign n2726 = ~n160 & n2725 ;
  assign n2727 = n2721 &  n2726 ;
  assign n2728 = ( x41 & ~n2726 ) | ( x41 & n2727 ) | ( ~n2726 & n2727 ) ;
  assign n2729 = ~n197 & n2699 ;
  assign n2730 = ( n208 & ~n419 ) | ( n208 & n2729 ) | ( ~n419 & n2729 ) ;
  assign n2731 = ~n208 & n2730 ;
  assign n2732 = ( n425 & ~n428 ) | ( n425 & n2731 ) | ( ~n428 & n2731 ) ;
  assign n2733 = ~n425 & n2732 ;
  assign n2734 = ~n2721 & n2733 ;
  assign n2735 = n2728 | n2734 ;
  assign n2736 = ~x40 & x64 ;
  assign n2737 = ( x65 & ~n2735 ) | ( x65 & n2736 ) | ( ~n2735 & n2736 ) ;
  assign n2916 = ( x66 & ~n2752 ) | ( x66 & n2737 ) | ( ~n2752 & n2737 ) ;
  assign n2917 = ( x67 & ~n2915 ) | ( x67 & n2916 ) | ( ~n2915 & n2916 ) ;
  assign n2918 = ( x68 & ~n2910 ) | ( x68 & n2917 ) | ( ~n2910 & n2917 ) ;
  assign n2919 = ( x69 & ~n2902 ) | ( x69 & n2918 ) | ( ~n2902 & n2918 ) ;
  assign n2920 = ( x70 & ~n2894 ) | ( x70 & n2919 ) | ( ~n2894 & n2919 ) ;
  assign n2921 = ( x71 & ~n2886 ) | ( x71 & n2920 ) | ( ~n2886 & n2920 ) ;
  assign n2922 = ( x72 & ~n2878 ) | ( x72 & n2921 ) | ( ~n2878 & n2921 ) ;
  assign n2923 = ( x73 & ~n2870 ) | ( x73 & n2922 ) | ( ~n2870 & n2922 ) ;
  assign n2924 = ( x74 & ~n2862 ) | ( x74 & n2923 ) | ( ~n2862 & n2923 ) ;
  assign n2925 = ( x75 & ~n2854 ) | ( x75 & n2924 ) | ( ~n2854 & n2924 ) ;
  assign n2926 = ( x76 & ~n2846 ) | ( x76 & n2925 ) | ( ~n2846 & n2925 ) ;
  assign n2927 = ( x77 & ~n2838 ) | ( x77 & n2926 ) | ( ~n2838 & n2926 ) ;
  assign n2928 = ( x78 & ~n2830 ) | ( x78 & n2927 ) | ( ~n2830 & n2927 ) ;
  assign n2929 = ( x79 & ~n2822 ) | ( x79 & n2928 ) | ( ~n2822 & n2928 ) ;
  assign n2930 = ( x80 & ~n2814 ) | ( x80 & n2929 ) | ( ~n2814 & n2929 ) ;
  assign n2931 = ( x81 & ~n2806 ) | ( x81 & n2930 ) | ( ~n2806 & n2930 ) ;
  assign n2932 = ( x82 & ~n2798 ) | ( x82 & n2931 ) | ( ~n2798 & n2931 ) ;
  assign n2933 = ( x83 & ~n2790 ) | ( x83 & n2932 ) | ( ~n2790 & n2932 ) ;
  assign n2934 = ( x84 & ~n2782 ) | ( x84 & n2933 ) | ( ~n2782 & n2933 ) ;
  assign n2935 = ( x85 & ~n2774 ) | ( x85 & n2934 ) | ( ~n2774 & n2934 ) ;
  assign n2936 = ( x86 & ~n2766 ) | ( x86 & n2935 ) | ( ~n2766 & n2935 ) ;
  assign n2940 = n261 | n273 ;
  assign n2941 = n270 | n2940 ;
  assign n2937 = x86 | n2720 ;
  assign n2938 = ( x86 & n2720 ) | ( x86 & n2741 ) | ( n2720 & n2741 ) ;
  assign n2939 = ( n2524 & ~n2937 ) | ( n2524 & n2938 ) | ( ~n2937 & n2938 ) ;
  assign n2943 = x87 &  n2939 ;
  assign n2942 = x87 | n2939 ;
  assign n2944 = ( n2941 & ~n2943 ) | ( n2941 & n2942 ) | ( ~n2943 & n2942 ) ;
  assign n2945 = n2936 | n2944 ;
  assign n2946 = ~n2939 |  n2741 ;
  assign n2966 = n2766 &  n2946 ;
  assign n2967 = n2945 &  n2966 ;
  assign n2953 = x86 | n2766 ;
  assign n2954 = x86 &  n2766 ;
  assign n2955 = ( n2953 & ~n2954 ) | ( n2953 & 1'b0 ) | ( ~n2954 & 1'b0 ) ;
  assign n2968 = n2935 &  n2955 ;
  assign n2947 = n2945 &  n2946 ;
  assign n2969 = ( n2935 & ~n2947 ) | ( n2935 & n2955 ) | ( ~n2947 & n2955 ) ;
  assign n2970 = ( n2967 & ~n2968 ) | ( n2967 & n2969 ) | ( ~n2968 & n2969 ) ;
  assign n2957 = ( x87 & n2936 ) | ( x87 & n2939 ) | ( n2936 & n2939 ) ;
  assign n2956 = ( x87 & ~n2936 ) | ( x87 & n2939 ) | ( ~n2936 & n2939 ) ;
  assign n2958 = ( n2936 & ~n2957 ) | ( n2936 & n2956 ) | ( ~n2957 & n2956 ) ;
  assign n2959 = ~n2947 & n2958 ;
  assign n2960 = n2524 &  n2741 ;
  assign n2961 = n2945 &  n2960 ;
  assign n2962 = n2959 | n2961 ;
  assign n2974 = n2774 &  n2946 ;
  assign n2975 = n2945 &  n2974 ;
  assign n2963 = x85 | n2774 ;
  assign n2964 = x85 &  n2774 ;
  assign n2965 = ( n2963 & ~n2964 ) | ( n2963 & 1'b0 ) | ( ~n2964 & 1'b0 ) ;
  assign n2976 = n2934 &  n2965 ;
  assign n2977 = ( n2934 & ~n2947 ) | ( n2934 & n2965 ) | ( ~n2947 & n2965 ) ;
  assign n2978 = ( n2975 & ~n2976 ) | ( n2975 & n2977 ) | ( ~n2976 & n2977 ) ;
  assign n2982 = n2782 &  n2946 ;
  assign n2983 = n2945 &  n2982 ;
  assign n2971 = x84 | n2782 ;
  assign n2972 = x84 &  n2782 ;
  assign n2973 = ( n2971 & ~n2972 ) | ( n2971 & 1'b0 ) | ( ~n2972 & 1'b0 ) ;
  assign n2984 = n2933 &  n2973 ;
  assign n2985 = ( n2933 & ~n2947 ) | ( n2933 & n2973 ) | ( ~n2947 & n2973 ) ;
  assign n2986 = ( n2983 & ~n2984 ) | ( n2983 & n2985 ) | ( ~n2984 & n2985 ) ;
  assign n2990 = n2790 &  n2946 ;
  assign n2991 = n2945 &  n2990 ;
  assign n2979 = x83 | n2790 ;
  assign n2980 = x83 &  n2790 ;
  assign n2981 = ( n2979 & ~n2980 ) | ( n2979 & 1'b0 ) | ( ~n2980 & 1'b0 ) ;
  assign n2992 = n2932 &  n2981 ;
  assign n2993 = ( n2932 & ~n2947 ) | ( n2932 & n2981 ) | ( ~n2947 & n2981 ) ;
  assign n2994 = ( n2991 & ~n2992 ) | ( n2991 & n2993 ) | ( ~n2992 & n2993 ) ;
  assign n2998 = n2798 &  n2946 ;
  assign n2999 = n2945 &  n2998 ;
  assign n2987 = x82 | n2798 ;
  assign n2988 = x82 &  n2798 ;
  assign n2989 = ( n2987 & ~n2988 ) | ( n2987 & 1'b0 ) | ( ~n2988 & 1'b0 ) ;
  assign n3000 = n2931 &  n2989 ;
  assign n3001 = ( n2931 & ~n2947 ) | ( n2931 & n2989 ) | ( ~n2947 & n2989 ) ;
  assign n3002 = ( n2999 & ~n3000 ) | ( n2999 & n3001 ) | ( ~n3000 & n3001 ) ;
  assign n3006 = n2806 &  n2946 ;
  assign n3007 = n2945 &  n3006 ;
  assign n2995 = x81 | n2806 ;
  assign n2996 = x81 &  n2806 ;
  assign n2997 = ( n2995 & ~n2996 ) | ( n2995 & 1'b0 ) | ( ~n2996 & 1'b0 ) ;
  assign n3009 = ( n2930 & n2947 ) | ( n2930 & n2997 ) | ( n2947 & n2997 ) ;
  assign n3008 = n2930 | n2997 ;
  assign n3010 = ( n3007 & ~n3009 ) | ( n3007 & n3008 ) | ( ~n3009 & n3008 ) ;
  assign n3014 = n2814 &  n2946 ;
  assign n3015 = n2945 &  n3014 ;
  assign n3003 = x80 | n2814 ;
  assign n3004 = x80 &  n2814 ;
  assign n3005 = ( n3003 & ~n3004 ) | ( n3003 & 1'b0 ) | ( ~n3004 & 1'b0 ) ;
  assign n3017 = ( n2929 & n2947 ) | ( n2929 & n3005 ) | ( n2947 & n3005 ) ;
  assign n3016 = n2929 | n3005 ;
  assign n3018 = ( n3015 & ~n3017 ) | ( n3015 & n3016 ) | ( ~n3017 & n3016 ) ;
  assign n3022 = n2822 &  n2946 ;
  assign n3023 = n2945 &  n3022 ;
  assign n3011 = x79 | n2822 ;
  assign n3012 = x79 &  n2822 ;
  assign n3013 = ( n3011 & ~n3012 ) | ( n3011 & 1'b0 ) | ( ~n3012 & 1'b0 ) ;
  assign n3025 = ( n2928 & n2947 ) | ( n2928 & n3013 ) | ( n2947 & n3013 ) ;
  assign n3024 = n2928 | n3013 ;
  assign n3026 = ( n3023 & ~n3025 ) | ( n3023 & n3024 ) | ( ~n3025 & n3024 ) ;
  assign n3030 = n2830 &  n2946 ;
  assign n3031 = n2945 &  n3030 ;
  assign n3019 = x78 | n2830 ;
  assign n3020 = x78 &  n2830 ;
  assign n3021 = ( n3019 & ~n3020 ) | ( n3019 & 1'b0 ) | ( ~n3020 & 1'b0 ) ;
  assign n3033 = ( n2927 & n2947 ) | ( n2927 & n3021 ) | ( n2947 & n3021 ) ;
  assign n3032 = n2927 | n3021 ;
  assign n3034 = ( n3031 & ~n3033 ) | ( n3031 & n3032 ) | ( ~n3033 & n3032 ) ;
  assign n3038 = n2838 &  n2946 ;
  assign n3039 = n2945 &  n3038 ;
  assign n3027 = x77 | n2838 ;
  assign n3028 = x77 &  n2838 ;
  assign n3029 = ( n3027 & ~n3028 ) | ( n3027 & 1'b0 ) | ( ~n3028 & 1'b0 ) ;
  assign n3041 = ( n2926 & n2947 ) | ( n2926 & n3029 ) | ( n2947 & n3029 ) ;
  assign n3040 = n2926 | n3029 ;
  assign n3042 = ( n3039 & ~n3041 ) | ( n3039 & n3040 ) | ( ~n3041 & n3040 ) ;
  assign n3046 = n2846 &  n2946 ;
  assign n3047 = n2945 &  n3046 ;
  assign n3035 = x76 | n2846 ;
  assign n3036 = x76 &  n2846 ;
  assign n3037 = ( n3035 & ~n3036 ) | ( n3035 & 1'b0 ) | ( ~n3036 & 1'b0 ) ;
  assign n3049 = ( n2925 & n2947 ) | ( n2925 & n3037 ) | ( n2947 & n3037 ) ;
  assign n3048 = n2925 | n3037 ;
  assign n3050 = ( n3047 & ~n3049 ) | ( n3047 & n3048 ) | ( ~n3049 & n3048 ) ;
  assign n3054 = n2854 &  n2946 ;
  assign n3055 = n2945 &  n3054 ;
  assign n3043 = x75 | n2854 ;
  assign n3044 = x75 &  n2854 ;
  assign n3045 = ( n3043 & ~n3044 ) | ( n3043 & 1'b0 ) | ( ~n3044 & 1'b0 ) ;
  assign n3057 = ( n2924 & n2947 ) | ( n2924 & n3045 ) | ( n2947 & n3045 ) ;
  assign n3056 = n2924 | n3045 ;
  assign n3058 = ( n3055 & ~n3057 ) | ( n3055 & n3056 ) | ( ~n3057 & n3056 ) ;
  assign n3062 = n2862 &  n2946 ;
  assign n3063 = n2945 &  n3062 ;
  assign n3051 = x74 | n2862 ;
  assign n3052 = x74 &  n2862 ;
  assign n3053 = ( n3051 & ~n3052 ) | ( n3051 & 1'b0 ) | ( ~n3052 & 1'b0 ) ;
  assign n3065 = ( n2923 & n2947 ) | ( n2923 & n3053 ) | ( n2947 & n3053 ) ;
  assign n3064 = n2923 | n3053 ;
  assign n3066 = ( n3063 & ~n3065 ) | ( n3063 & n3064 ) | ( ~n3065 & n3064 ) ;
  assign n3070 = n2870 &  n2946 ;
  assign n3071 = n2945 &  n3070 ;
  assign n3059 = x73 | n2870 ;
  assign n3060 = x73 &  n2870 ;
  assign n3061 = ( n3059 & ~n3060 ) | ( n3059 & 1'b0 ) | ( ~n3060 & 1'b0 ) ;
  assign n3073 = ( n2922 & n2947 ) | ( n2922 & n3061 ) | ( n2947 & n3061 ) ;
  assign n3072 = n2922 | n3061 ;
  assign n3074 = ( n3071 & ~n3073 ) | ( n3071 & n3072 ) | ( ~n3073 & n3072 ) ;
  assign n3078 = n2878 &  n2946 ;
  assign n3079 = n2945 &  n3078 ;
  assign n3067 = x72 | n2878 ;
  assign n3068 = x72 &  n2878 ;
  assign n3069 = ( n3067 & ~n3068 ) | ( n3067 & 1'b0 ) | ( ~n3068 & 1'b0 ) ;
  assign n3081 = ( n2921 & n2947 ) | ( n2921 & n3069 ) | ( n2947 & n3069 ) ;
  assign n3080 = n2921 | n3069 ;
  assign n3082 = ( n3079 & ~n3081 ) | ( n3079 & n3080 ) | ( ~n3081 & n3080 ) ;
  assign n3086 = n2886 &  n2946 ;
  assign n3087 = n2945 &  n3086 ;
  assign n3075 = x71 | n2886 ;
  assign n3076 = x71 &  n2886 ;
  assign n3077 = ( n3075 & ~n3076 ) | ( n3075 & 1'b0 ) | ( ~n3076 & 1'b0 ) ;
  assign n3089 = ( n2920 & n2947 ) | ( n2920 & n3077 ) | ( n2947 & n3077 ) ;
  assign n3088 = n2920 | n3077 ;
  assign n3090 = ( n3087 & ~n3089 ) | ( n3087 & n3088 ) | ( ~n3089 & n3088 ) ;
  assign n3094 = n2894 &  n2946 ;
  assign n3095 = n2945 &  n3094 ;
  assign n3083 = x70 | n2894 ;
  assign n3084 = x70 &  n2894 ;
  assign n3085 = ( n3083 & ~n3084 ) | ( n3083 & 1'b0 ) | ( ~n3084 & 1'b0 ) ;
  assign n3097 = ( n2919 & n2947 ) | ( n2919 & n3085 ) | ( n2947 & n3085 ) ;
  assign n3096 = n2919 | n3085 ;
  assign n3098 = ( n3095 & ~n3097 ) | ( n3095 & n3096 ) | ( ~n3097 & n3096 ) ;
  assign n3102 = n2902 &  n2946 ;
  assign n3103 = n2945 &  n3102 ;
  assign n3091 = x69 | n2902 ;
  assign n3092 = x69 &  n2902 ;
  assign n3093 = ( n3091 & ~n3092 ) | ( n3091 & 1'b0 ) | ( ~n3092 & 1'b0 ) ;
  assign n3105 = ( n2918 & n2947 ) | ( n2918 & n3093 ) | ( n2947 & n3093 ) ;
  assign n3104 = n2918 | n3093 ;
  assign n3106 = ( n3103 & ~n3105 ) | ( n3103 & n3104 ) | ( ~n3105 & n3104 ) ;
  assign n3110 = n2910 &  n2946 ;
  assign n3111 = n2945 &  n3110 ;
  assign n3099 = x68 | n2910 ;
  assign n3100 = x68 &  n2910 ;
  assign n3101 = ( n3099 & ~n3100 ) | ( n3099 & 1'b0 ) | ( ~n3100 & 1'b0 ) ;
  assign n3113 = ( n2917 & n2947 ) | ( n2917 & n3101 ) | ( n2947 & n3101 ) ;
  assign n3112 = n2917 | n3101 ;
  assign n3114 = ( n3111 & ~n3113 ) | ( n3111 & n3112 ) | ( ~n3113 & n3112 ) ;
  assign n3115 = n2915 &  n2946 ;
  assign n3116 = n2945 &  n3115 ;
  assign n3107 = x67 | n2915 ;
  assign n3108 = x67 &  n2915 ;
  assign n3109 = ( n3107 & ~n3108 ) | ( n3107 & 1'b0 ) | ( ~n3108 & 1'b0 ) ;
  assign n3118 = ( n2916 & n2947 ) | ( n2916 & n3109 ) | ( n2947 & n3109 ) ;
  assign n3117 = n2916 | n3109 ;
  assign n3119 = ( n3116 & ~n3118 ) | ( n3116 & n3117 ) | ( ~n3118 & n3117 ) ;
  assign n2948 = n2752 &  n2946 ;
  assign n2949 = n2945 &  n2948 ;
  assign n2753 = x66 | n2752 ;
  assign n2754 = x66 &  n2752 ;
  assign n2755 = ( n2753 & ~n2754 ) | ( n2753 & 1'b0 ) | ( ~n2754 & 1'b0 ) ;
  assign n2951 = ( n2737 & n2755 ) | ( n2737 & n2947 ) | ( n2755 & n2947 ) ;
  assign n2950 = n2737 | n2755 ;
  assign n2952 = ( n2949 & ~n2951 ) | ( n2949 & n2950 ) | ( ~n2951 & n2950 ) ;
  assign n3120 = ( n2735 & ~x65 ) | ( n2735 & n2736 ) | ( ~x65 & n2736 ) ;
  assign n3121 = ( n2737 & ~n2736 ) | ( n2737 & n3120 ) | ( ~n2736 & n3120 ) ;
  assign n3122 = ~n2947 & n3121 ;
  assign n3123 = n2735 &  n2946 ;
  assign n3124 = n2945 &  n3123 ;
  assign n3125 = n3122 | n3124 ;
  assign n3126 = ( x64 & ~n2947 ) | ( x64 & 1'b0 ) | ( ~n2947 & 1'b0 ) ;
  assign n3127 = ( x40 & ~n3126 ) | ( x40 & 1'b0 ) | ( ~n3126 & 1'b0 ) ;
  assign n3128 = ( n2736 & ~n2947 ) | ( n2736 & 1'b0 ) | ( ~n2947 & 1'b0 ) ;
  assign n3129 = n3127 | n3128 ;
  assign n3130 = ~x39 & x64 ;
  assign n3131 = ( x65 & ~n3129 ) | ( x65 & n3130 ) | ( ~n3129 & n3130 ) ;
  assign n3132 = ( x66 & ~n3125 ) | ( x66 & n3131 ) | ( ~n3125 & n3131 ) ;
  assign n3133 = ( x67 & ~n2952 ) | ( x67 & n3132 ) | ( ~n2952 & n3132 ) ;
  assign n3134 = ( x68 & ~n3119 ) | ( x68 & n3133 ) | ( ~n3119 & n3133 ) ;
  assign n3135 = ( x69 & ~n3114 ) | ( x69 & n3134 ) | ( ~n3114 & n3134 ) ;
  assign n3136 = ( x70 & ~n3106 ) | ( x70 & n3135 ) | ( ~n3106 & n3135 ) ;
  assign n3137 = ( x71 & ~n3098 ) | ( x71 & n3136 ) | ( ~n3098 & n3136 ) ;
  assign n3138 = ( x72 & ~n3090 ) | ( x72 & n3137 ) | ( ~n3090 & n3137 ) ;
  assign n3139 = ( x73 & ~n3082 ) | ( x73 & n3138 ) | ( ~n3082 & n3138 ) ;
  assign n3140 = ( x74 & ~n3074 ) | ( x74 & n3139 ) | ( ~n3074 & n3139 ) ;
  assign n3141 = ( x75 & ~n3066 ) | ( x75 & n3140 ) | ( ~n3066 & n3140 ) ;
  assign n3142 = ( x76 & ~n3058 ) | ( x76 & n3141 ) | ( ~n3058 & n3141 ) ;
  assign n3143 = ( x77 & ~n3050 ) | ( x77 & n3142 ) | ( ~n3050 & n3142 ) ;
  assign n3144 = ( x78 & ~n3042 ) | ( x78 & n3143 ) | ( ~n3042 & n3143 ) ;
  assign n3145 = ( x79 & ~n3034 ) | ( x79 & n3144 ) | ( ~n3034 & n3144 ) ;
  assign n3146 = ( x80 & ~n3026 ) | ( x80 & n3145 ) | ( ~n3026 & n3145 ) ;
  assign n3147 = ( x81 & ~n3018 ) | ( x81 & n3146 ) | ( ~n3018 & n3146 ) ;
  assign n3148 = ( x82 & ~n3010 ) | ( x82 & n3147 ) | ( ~n3010 & n3147 ) ;
  assign n3149 = ( x83 & ~n3002 ) | ( x83 & n3148 ) | ( ~n3002 & n3148 ) ;
  assign n3150 = ( x84 & ~n2994 ) | ( x84 & n3149 ) | ( ~n2994 & n3149 ) ;
  assign n3151 = ( x85 & ~n2986 ) | ( x85 & n3150 ) | ( ~n2986 & n3150 ) ;
  assign n3152 = ( x86 & ~n2978 ) | ( x86 & n3151 ) | ( ~n2978 & n3151 ) ;
  assign n3153 = ( x87 & ~n2970 ) | ( x87 & n3152 ) | ( ~n2970 & n3152 ) ;
  assign n3154 = ( x88 & ~n2962 ) | ( x88 & n3153 ) | ( ~n2962 & n3153 ) ;
  assign n3155 = n209 | n255 ;
  assign n3156 = n240 | n3155 ;
  assign n3157 = n3154 | n3156 ;
  assign n3175 = n2970 &  n3157 ;
  assign n3169 = x87 | n2970 ;
  assign n3170 = x87 &  n2970 ;
  assign n3171 = ( n3169 & ~n3170 ) | ( n3169 & 1'b0 ) | ( ~n3170 & 1'b0 ) ;
  assign n3179 = ( n3152 & n3154 ) | ( n3152 & n3171 ) | ( n3154 & n3171 ) ;
  assign n3180 = ( n3152 & ~n3156 ) | ( n3152 & n3171 ) | ( ~n3156 & n3171 ) ;
  assign n3181 = ~n3179 & n3180 ;
  assign n3182 = n3175 | n3181 ;
  assign n3172 = x88 | n3153 ;
  assign n3173 = ( x88 & n3153 ) | ( x88 & n3156 ) | ( n3153 & n3156 ) ;
  assign n3174 = ( n2962 & ~n3172 ) | ( n2962 & n3173 ) | ( ~n3172 & n3173 ) ;
  assign n3183 = n2978 &  n3157 ;
  assign n3176 = x86 | n2978 ;
  assign n3177 = x86 &  n2978 ;
  assign n3178 = ( n3176 & ~n3177 ) | ( n3176 & 1'b0 ) | ( ~n3177 & 1'b0 ) ;
  assign n3187 = ( n3151 & n3154 ) | ( n3151 & n3178 ) | ( n3154 & n3178 ) ;
  assign n3188 = ( n3151 & ~n3156 ) | ( n3151 & n3178 ) | ( ~n3156 & n3178 ) ;
  assign n3189 = ~n3187 & n3188 ;
  assign n3190 = n3183 | n3189 ;
  assign n3191 = n2986 &  n3157 ;
  assign n3184 = x85 | n2986 ;
  assign n3185 = x85 &  n2986 ;
  assign n3186 = ( n3184 & ~n3185 ) | ( n3184 & 1'b0 ) | ( ~n3185 & 1'b0 ) ;
  assign n3195 = ( n3150 & n3154 ) | ( n3150 & n3186 ) | ( n3154 & n3186 ) ;
  assign n3196 = ( n3150 & ~n3156 ) | ( n3150 & n3186 ) | ( ~n3156 & n3186 ) ;
  assign n3197 = ~n3195 & n3196 ;
  assign n3198 = n3191 | n3197 ;
  assign n3199 = n2994 &  n3157 ;
  assign n3192 = x84 | n2994 ;
  assign n3193 = x84 &  n2994 ;
  assign n3194 = ( n3192 & ~n3193 ) | ( n3192 & 1'b0 ) | ( ~n3193 & 1'b0 ) ;
  assign n3203 = ( n3149 & n3154 ) | ( n3149 & n3194 ) | ( n3154 & n3194 ) ;
  assign n3204 = ( n3149 & ~n3156 ) | ( n3149 & n3194 ) | ( ~n3156 & n3194 ) ;
  assign n3205 = ~n3203 & n3204 ;
  assign n3206 = n3199 | n3205 ;
  assign n3207 = n3002 &  n3157 ;
  assign n3200 = x83 | n3002 ;
  assign n3201 = x83 &  n3002 ;
  assign n3202 = ( n3200 & ~n3201 ) | ( n3200 & 1'b0 ) | ( ~n3201 & 1'b0 ) ;
  assign n3211 = ( n3148 & n3154 ) | ( n3148 & n3202 ) | ( n3154 & n3202 ) ;
  assign n3212 = ( n3148 & ~n3156 ) | ( n3148 & n3202 ) | ( ~n3156 & n3202 ) ;
  assign n3213 = ~n3211 & n3212 ;
  assign n3214 = n3207 | n3213 ;
  assign n3215 = n3010 &  n3157 ;
  assign n3208 = x82 | n3010 ;
  assign n3209 = x82 &  n3010 ;
  assign n3210 = ( n3208 & ~n3209 ) | ( n3208 & 1'b0 ) | ( ~n3209 & 1'b0 ) ;
  assign n3219 = ( n3147 & n3154 ) | ( n3147 & n3210 ) | ( n3154 & n3210 ) ;
  assign n3220 = ( n3147 & ~n3156 ) | ( n3147 & n3210 ) | ( ~n3156 & n3210 ) ;
  assign n3221 = ~n3219 & n3220 ;
  assign n3222 = n3215 | n3221 ;
  assign n3223 = n3018 &  n3157 ;
  assign n3216 = x81 | n3018 ;
  assign n3217 = x81 &  n3018 ;
  assign n3218 = ( n3216 & ~n3217 ) | ( n3216 & 1'b0 ) | ( ~n3217 & 1'b0 ) ;
  assign n3227 = ( n3146 & n3154 ) | ( n3146 & n3218 ) | ( n3154 & n3218 ) ;
  assign n3228 = ( n3146 & ~n3156 ) | ( n3146 & n3218 ) | ( ~n3156 & n3218 ) ;
  assign n3229 = ~n3227 & n3228 ;
  assign n3230 = n3223 | n3229 ;
  assign n3231 = n3026 &  n3157 ;
  assign n3224 = x80 | n3026 ;
  assign n3225 = x80 &  n3026 ;
  assign n3226 = ( n3224 & ~n3225 ) | ( n3224 & 1'b0 ) | ( ~n3225 & 1'b0 ) ;
  assign n3235 = ( n3145 & n3154 ) | ( n3145 & n3226 ) | ( n3154 & n3226 ) ;
  assign n3236 = ( n3145 & ~n3156 ) | ( n3145 & n3226 ) | ( ~n3156 & n3226 ) ;
  assign n3237 = ~n3235 & n3236 ;
  assign n3238 = n3231 | n3237 ;
  assign n3239 = n3034 &  n3157 ;
  assign n3232 = x79 | n3034 ;
  assign n3233 = x79 &  n3034 ;
  assign n3234 = ( n3232 & ~n3233 ) | ( n3232 & 1'b0 ) | ( ~n3233 & 1'b0 ) ;
  assign n3243 = ( n3144 & n3154 ) | ( n3144 & n3234 ) | ( n3154 & n3234 ) ;
  assign n3244 = ( n3144 & ~n3156 ) | ( n3144 & n3234 ) | ( ~n3156 & n3234 ) ;
  assign n3245 = ~n3243 & n3244 ;
  assign n3246 = n3239 | n3245 ;
  assign n3247 = n3042 &  n3157 ;
  assign n3240 = x78 | n3042 ;
  assign n3241 = x78 &  n3042 ;
  assign n3242 = ( n3240 & ~n3241 ) | ( n3240 & 1'b0 ) | ( ~n3241 & 1'b0 ) ;
  assign n3251 = ( n3143 & n3154 ) | ( n3143 & n3242 ) | ( n3154 & n3242 ) ;
  assign n3252 = ( n3143 & ~n3156 ) | ( n3143 & n3242 ) | ( ~n3156 & n3242 ) ;
  assign n3253 = ~n3251 & n3252 ;
  assign n3254 = n3247 | n3253 ;
  assign n3255 = n3050 &  n3157 ;
  assign n3248 = x77 | n3050 ;
  assign n3249 = x77 &  n3050 ;
  assign n3250 = ( n3248 & ~n3249 ) | ( n3248 & 1'b0 ) | ( ~n3249 & 1'b0 ) ;
  assign n3259 = ( n3142 & n3154 ) | ( n3142 & n3250 ) | ( n3154 & n3250 ) ;
  assign n3260 = ( n3142 & ~n3156 ) | ( n3142 & n3250 ) | ( ~n3156 & n3250 ) ;
  assign n3261 = ~n3259 & n3260 ;
  assign n3262 = n3255 | n3261 ;
  assign n3263 = n3058 &  n3157 ;
  assign n3256 = x76 | n3058 ;
  assign n3257 = x76 &  n3058 ;
  assign n3258 = ( n3256 & ~n3257 ) | ( n3256 & 1'b0 ) | ( ~n3257 & 1'b0 ) ;
  assign n3267 = ( n3141 & n3154 ) | ( n3141 & n3258 ) | ( n3154 & n3258 ) ;
  assign n3268 = ( n3141 & ~n3156 ) | ( n3141 & n3258 ) | ( ~n3156 & n3258 ) ;
  assign n3269 = ~n3267 & n3268 ;
  assign n3270 = n3263 | n3269 ;
  assign n3271 = n3066 &  n3157 ;
  assign n3264 = x75 | n3066 ;
  assign n3265 = x75 &  n3066 ;
  assign n3266 = ( n3264 & ~n3265 ) | ( n3264 & 1'b0 ) | ( ~n3265 & 1'b0 ) ;
  assign n3275 = ( n3140 & n3154 ) | ( n3140 & n3266 ) | ( n3154 & n3266 ) ;
  assign n3276 = ( n3140 & ~n3156 ) | ( n3140 & n3266 ) | ( ~n3156 & n3266 ) ;
  assign n3277 = ~n3275 & n3276 ;
  assign n3278 = n3271 | n3277 ;
  assign n3279 = n3074 &  n3157 ;
  assign n3272 = x74 | n3074 ;
  assign n3273 = x74 &  n3074 ;
  assign n3274 = ( n3272 & ~n3273 ) | ( n3272 & 1'b0 ) | ( ~n3273 & 1'b0 ) ;
  assign n3283 = ( n3139 & n3154 ) | ( n3139 & n3274 ) | ( n3154 & n3274 ) ;
  assign n3284 = ( n3139 & ~n3156 ) | ( n3139 & n3274 ) | ( ~n3156 & n3274 ) ;
  assign n3285 = ~n3283 & n3284 ;
  assign n3286 = n3279 | n3285 ;
  assign n3287 = n3082 &  n3157 ;
  assign n3280 = x73 | n3082 ;
  assign n3281 = x73 &  n3082 ;
  assign n3282 = ( n3280 & ~n3281 ) | ( n3280 & 1'b0 ) | ( ~n3281 & 1'b0 ) ;
  assign n3291 = ( n3138 & n3154 ) | ( n3138 & n3282 ) | ( n3154 & n3282 ) ;
  assign n3292 = ( n3138 & ~n3156 ) | ( n3138 & n3282 ) | ( ~n3156 & n3282 ) ;
  assign n3293 = ~n3291 & n3292 ;
  assign n3294 = n3287 | n3293 ;
  assign n3295 = n3090 &  n3157 ;
  assign n3288 = x72 | n3090 ;
  assign n3289 = x72 &  n3090 ;
  assign n3290 = ( n3288 & ~n3289 ) | ( n3288 & 1'b0 ) | ( ~n3289 & 1'b0 ) ;
  assign n3299 = ( n3137 & n3154 ) | ( n3137 & n3290 ) | ( n3154 & n3290 ) ;
  assign n3300 = ( n3137 & ~n3156 ) | ( n3137 & n3290 ) | ( ~n3156 & n3290 ) ;
  assign n3301 = ~n3299 & n3300 ;
  assign n3302 = n3295 | n3301 ;
  assign n3303 = n3098 &  n3157 ;
  assign n3296 = x71 | n3098 ;
  assign n3297 = x71 &  n3098 ;
  assign n3298 = ( n3296 & ~n3297 ) | ( n3296 & 1'b0 ) | ( ~n3297 & 1'b0 ) ;
  assign n3307 = ( n3136 & n3154 ) | ( n3136 & n3298 ) | ( n3154 & n3298 ) ;
  assign n3308 = ( n3136 & ~n3156 ) | ( n3136 & n3298 ) | ( ~n3156 & n3298 ) ;
  assign n3309 = ~n3307 & n3308 ;
  assign n3310 = n3303 | n3309 ;
  assign n3311 = n3106 &  n3157 ;
  assign n3304 = x70 | n3106 ;
  assign n3305 = x70 &  n3106 ;
  assign n3306 = ( n3304 & ~n3305 ) | ( n3304 & 1'b0 ) | ( ~n3305 & 1'b0 ) ;
  assign n3315 = ( n3135 & n3154 ) | ( n3135 & n3306 ) | ( n3154 & n3306 ) ;
  assign n3316 = ( n3135 & ~n3156 ) | ( n3135 & n3306 ) | ( ~n3156 & n3306 ) ;
  assign n3317 = ~n3315 & n3316 ;
  assign n3318 = n3311 | n3317 ;
  assign n3319 = n3114 &  n3157 ;
  assign n3312 = x69 | n3114 ;
  assign n3313 = x69 &  n3114 ;
  assign n3314 = ( n3312 & ~n3313 ) | ( n3312 & 1'b0 ) | ( ~n3313 & 1'b0 ) ;
  assign n3323 = ( n3134 & n3154 ) | ( n3134 & n3314 ) | ( n3154 & n3314 ) ;
  assign n3324 = ( n3134 & ~n3156 ) | ( n3134 & n3314 ) | ( ~n3156 & n3314 ) ;
  assign n3325 = ~n3323 & n3324 ;
  assign n3326 = n3319 | n3325 ;
  assign n3327 = n3119 &  n3157 ;
  assign n3320 = x68 | n3119 ;
  assign n3321 = x68 &  n3119 ;
  assign n3322 = ( n3320 & ~n3321 ) | ( n3320 & 1'b0 ) | ( ~n3321 & 1'b0 ) ;
  assign n3328 = ( n3133 & n3154 ) | ( n3133 & n3322 ) | ( n3154 & n3322 ) ;
  assign n3329 = ( n3133 & ~n3156 ) | ( n3133 & n3322 ) | ( ~n3156 & n3322 ) ;
  assign n3330 = ~n3328 & n3329 ;
  assign n3331 = n3327 | n3330 ;
  assign n3158 = n2952 &  n3157 ;
  assign n3162 = x67 | n2952 ;
  assign n3163 = x67 &  n2952 ;
  assign n3164 = ( n3162 & ~n3163 ) | ( n3162 & 1'b0 ) | ( ~n3163 & 1'b0 ) ;
  assign n3165 = ( n3132 & n3154 ) | ( n3132 & n3164 ) | ( n3154 & n3164 ) ;
  assign n3166 = ( n3132 & ~n3156 ) | ( n3132 & n3164 ) | ( ~n3156 & n3164 ) ;
  assign n3167 = ~n3165 & n3166 ;
  assign n3168 = n3158 | n3167 ;
  assign n3332 = n3125 &  n3157 ;
  assign n3159 = x66 | n3125 ;
  assign n3160 = x66 &  n3125 ;
  assign n3161 = ( n3159 & ~n3160 ) | ( n3159 & 1'b0 ) | ( ~n3160 & 1'b0 ) ;
  assign n3337 = ( n3131 & ~n3154 ) | ( n3131 & n3161 ) | ( ~n3154 & n3161 ) ;
  assign n3338 = ( n3131 & n3156 ) | ( n3131 & n3161 ) | ( n3156 & n3161 ) ;
  assign n3339 = ( n3337 & ~n3338 ) | ( n3337 & 1'b0 ) | ( ~n3338 & 1'b0 ) ;
  assign n3340 = n3332 | n3339 ;
  assign n3341 = n3129 &  n3157 ;
  assign n3333 = x65 &  n3129 ;
  assign n3334 = ( n3127 & ~x65 ) | ( n3127 & n3128 ) | ( ~x65 & n3128 ) ;
  assign n3335 = x65 | n3334 ;
  assign n3336 = ( n3130 & ~n3333 ) | ( n3130 & n3335 ) | ( ~n3333 & n3335 ) ;
  assign n3342 = ( x65 & n3129 ) | ( x65 & n3130 ) | ( n3129 & n3130 ) ;
  assign n3343 = ( n3156 & ~n3333 ) | ( n3156 & n3342 ) | ( ~n3333 & n3342 ) ;
  assign n3344 = ( n3154 & n3336 ) | ( n3154 & n3343 ) | ( n3336 & n3343 ) ;
  assign n3345 = ( n3336 & ~n3344 ) | ( n3336 & 1'b0 ) | ( ~n3344 & 1'b0 ) ;
  assign n3346 = n3341 | n3345 ;
  assign n3347 = ( x64 & ~x89 ) | ( x64 & 1'b0 ) | ( ~x89 & 1'b0 ) ;
  assign n3348 = ( n177 & ~n188 ) | ( n177 & n3347 ) | ( ~n188 & n3347 ) ;
  assign n3349 = ~n177 & n3348 ;
  assign n3350 = ( n270 & ~n273 ) | ( n270 & n3349 ) | ( ~n273 & n3349 ) ;
  assign n3351 = ~n270 & n3350 ;
  assign n3352 = n3154 &  n3351 ;
  assign n3353 = ( x39 & ~n3351 ) | ( x39 & n3352 ) | ( ~n3351 & n3352 ) ;
  assign n3354 = ~n208 & n3130 ;
  assign n3355 = ( n419 & ~n428 ) | ( n419 & n3354 ) | ( ~n428 & n3354 ) ;
  assign n3356 = ~n419 & n3355 ;
  assign n3357 = ~n425 & n3356 ;
  assign n3358 = ~n3154 & n3357 ;
  assign n3359 = n3353 | n3358 ;
  assign n3360 = ~x38 & x64 ;
  assign n3361 = ( x65 & ~n3359 ) | ( x65 & n3360 ) | ( ~n3359 & n3360 ) ;
  assign n3362 = ( x66 & ~n3346 ) | ( x66 & n3361 ) | ( ~n3346 & n3361 ) ;
  assign n3363 = ( x67 & ~n3340 ) | ( x67 & n3362 ) | ( ~n3340 & n3362 ) ;
  assign n3364 = ( x68 & ~n3168 ) | ( x68 & n3363 ) | ( ~n3168 & n3363 ) ;
  assign n3365 = ( x69 & ~n3331 ) | ( x69 & n3364 ) | ( ~n3331 & n3364 ) ;
  assign n3366 = ( x70 & ~n3326 ) | ( x70 & n3365 ) | ( ~n3326 & n3365 ) ;
  assign n3367 = ( x71 & ~n3318 ) | ( x71 & n3366 ) | ( ~n3318 & n3366 ) ;
  assign n3368 = ( x72 & ~n3310 ) | ( x72 & n3367 ) | ( ~n3310 & n3367 ) ;
  assign n3369 = ( x73 & ~n3302 ) | ( x73 & n3368 ) | ( ~n3302 & n3368 ) ;
  assign n3370 = ( x74 & ~n3294 ) | ( x74 & n3369 ) | ( ~n3294 & n3369 ) ;
  assign n3371 = ( x75 & ~n3286 ) | ( x75 & n3370 ) | ( ~n3286 & n3370 ) ;
  assign n3372 = ( x76 & ~n3278 ) | ( x76 & n3371 ) | ( ~n3278 & n3371 ) ;
  assign n3373 = ( x77 & ~n3270 ) | ( x77 & n3372 ) | ( ~n3270 & n3372 ) ;
  assign n3374 = ( x78 & ~n3262 ) | ( x78 & n3373 ) | ( ~n3262 & n3373 ) ;
  assign n3375 = ( x79 & ~n3254 ) | ( x79 & n3374 ) | ( ~n3254 & n3374 ) ;
  assign n3376 = ( x80 & ~n3246 ) | ( x80 & n3375 ) | ( ~n3246 & n3375 ) ;
  assign n3377 = ( x81 & ~n3238 ) | ( x81 & n3376 ) | ( ~n3238 & n3376 ) ;
  assign n3378 = ( x82 & ~n3230 ) | ( x82 & n3377 ) | ( ~n3230 & n3377 ) ;
  assign n3379 = ( x83 & ~n3222 ) | ( x83 & n3378 ) | ( ~n3222 & n3378 ) ;
  assign n3380 = ( x84 & ~n3214 ) | ( x84 & n3379 ) | ( ~n3214 & n3379 ) ;
  assign n3381 = ( x85 & ~n3206 ) | ( x85 & n3380 ) | ( ~n3206 & n3380 ) ;
  assign n3382 = ( x86 & ~n3198 ) | ( x86 & n3381 ) | ( ~n3198 & n3381 ) ;
  assign n3383 = ( x87 & ~n3190 ) | ( x87 & n3382 ) | ( ~n3190 & n3382 ) ;
  assign n3384 = ( x88 & ~n3182 ) | ( x88 & n3383 ) | ( ~n3182 & n3383 ) ;
  assign n3385 = ( x89 & ~n3174 ) | ( x89 & n3384 ) | ( ~n3174 & n3384 ) ;
  assign n3386 = n177 | n188 ;
  assign n3387 = ( n273 & ~n270 ) | ( n273 & n3386 ) | ( ~n270 & n3386 ) ;
  assign n3388 = n270 | n3387 ;
  assign n3389 = n3385 | n3388 ;
  assign n3457 = n3182 &  n3389 ;
  assign n3461 = x88 | n3182 ;
  assign n3462 = x88 &  n3182 ;
  assign n3463 = ( n3461 & ~n3462 ) | ( n3461 & 1'b0 ) | ( ~n3462 & 1'b0 ) ;
  assign n3464 = ( n3383 & n3385 ) | ( n3383 & n3463 ) | ( n3385 & n3463 ) ;
  assign n3465 = ( n3383 & ~n3388 ) | ( n3383 & n3463 ) | ( ~n3388 & n3463 ) ;
  assign n3466 = ~n3464 & n3465 ;
  assign n3467 = n3457 | n3466 ;
  assign n3468 = n3190 &  n3389 ;
  assign n3458 = x87 | n3190 ;
  assign n3459 = x87 &  n3190 ;
  assign n3460 = ( n3458 & ~n3459 ) | ( n3458 & 1'b0 ) | ( ~n3459 & 1'b0 ) ;
  assign n3472 = ( n3382 & n3385 ) | ( n3382 & n3460 ) | ( n3385 & n3460 ) ;
  assign n3473 = ( n3382 & ~n3388 ) | ( n3382 & n3460 ) | ( ~n3388 & n3460 ) ;
  assign n3474 = ~n3472 & n3473 ;
  assign n3475 = n3468 | n3474 ;
  assign n3476 = n3198 &  n3389 ;
  assign n3469 = x86 | n3198 ;
  assign n3470 = x86 &  n3198 ;
  assign n3471 = ( n3469 & ~n3470 ) | ( n3469 & 1'b0 ) | ( ~n3470 & 1'b0 ) ;
  assign n3480 = ( n3381 & n3385 ) | ( n3381 & n3471 ) | ( n3385 & n3471 ) ;
  assign n3481 = ( n3381 & ~n3388 ) | ( n3381 & n3471 ) | ( ~n3388 & n3471 ) ;
  assign n3482 = ~n3480 & n3481 ;
  assign n3483 = n3476 | n3482 ;
  assign n3484 = n3206 &  n3389 ;
  assign n3477 = x85 | n3206 ;
  assign n3478 = x85 &  n3206 ;
  assign n3479 = ( n3477 & ~n3478 ) | ( n3477 & 1'b0 ) | ( ~n3478 & 1'b0 ) ;
  assign n3488 = ( n3380 & n3385 ) | ( n3380 & n3479 ) | ( n3385 & n3479 ) ;
  assign n3489 = ( n3380 & ~n3388 ) | ( n3380 & n3479 ) | ( ~n3388 & n3479 ) ;
  assign n3490 = ~n3488 & n3489 ;
  assign n3491 = n3484 | n3490 ;
  assign n3492 = n3214 &  n3389 ;
  assign n3485 = x84 | n3214 ;
  assign n3486 = x84 &  n3214 ;
  assign n3487 = ( n3485 & ~n3486 ) | ( n3485 & 1'b0 ) | ( ~n3486 & 1'b0 ) ;
  assign n3496 = ( n3379 & n3385 ) | ( n3379 & n3487 ) | ( n3385 & n3487 ) ;
  assign n3497 = ( n3379 & ~n3388 ) | ( n3379 & n3487 ) | ( ~n3388 & n3487 ) ;
  assign n3498 = ~n3496 & n3497 ;
  assign n3499 = n3492 | n3498 ;
  assign n3500 = n3222 &  n3389 ;
  assign n3493 = x83 | n3222 ;
  assign n3494 = x83 &  n3222 ;
  assign n3495 = ( n3493 & ~n3494 ) | ( n3493 & 1'b0 ) | ( ~n3494 & 1'b0 ) ;
  assign n3504 = ( n3378 & n3385 ) | ( n3378 & n3495 ) | ( n3385 & n3495 ) ;
  assign n3505 = ( n3378 & ~n3388 ) | ( n3378 & n3495 ) | ( ~n3388 & n3495 ) ;
  assign n3506 = ~n3504 & n3505 ;
  assign n3507 = n3500 | n3506 ;
  assign n3508 = n3230 &  n3389 ;
  assign n3501 = x82 | n3230 ;
  assign n3502 = x82 &  n3230 ;
  assign n3503 = ( n3501 & ~n3502 ) | ( n3501 & 1'b0 ) | ( ~n3502 & 1'b0 ) ;
  assign n3512 = ( n3377 & n3385 ) | ( n3377 & n3503 ) | ( n3385 & n3503 ) ;
  assign n3513 = ( n3377 & ~n3388 ) | ( n3377 & n3503 ) | ( ~n3388 & n3503 ) ;
  assign n3514 = ~n3512 & n3513 ;
  assign n3515 = n3508 | n3514 ;
  assign n3516 = n3238 &  n3389 ;
  assign n3509 = x81 | n3238 ;
  assign n3510 = x81 &  n3238 ;
  assign n3511 = ( n3509 & ~n3510 ) | ( n3509 & 1'b0 ) | ( ~n3510 & 1'b0 ) ;
  assign n3520 = ( n3376 & n3385 ) | ( n3376 & n3511 ) | ( n3385 & n3511 ) ;
  assign n3521 = ( n3376 & ~n3388 ) | ( n3376 & n3511 ) | ( ~n3388 & n3511 ) ;
  assign n3522 = ~n3520 & n3521 ;
  assign n3523 = n3516 | n3522 ;
  assign n3524 = n3246 &  n3389 ;
  assign n3517 = x80 | n3246 ;
  assign n3518 = x80 &  n3246 ;
  assign n3519 = ( n3517 & ~n3518 ) | ( n3517 & 1'b0 ) | ( ~n3518 & 1'b0 ) ;
  assign n3528 = ( n3375 & n3385 ) | ( n3375 & n3519 ) | ( n3385 & n3519 ) ;
  assign n3529 = ( n3375 & ~n3388 ) | ( n3375 & n3519 ) | ( ~n3388 & n3519 ) ;
  assign n3530 = ~n3528 & n3529 ;
  assign n3531 = n3524 | n3530 ;
  assign n3532 = n3254 &  n3389 ;
  assign n3525 = x79 | n3254 ;
  assign n3526 = x79 &  n3254 ;
  assign n3527 = ( n3525 & ~n3526 ) | ( n3525 & 1'b0 ) | ( ~n3526 & 1'b0 ) ;
  assign n3536 = ( n3374 & n3385 ) | ( n3374 & n3527 ) | ( n3385 & n3527 ) ;
  assign n3537 = ( n3374 & ~n3388 ) | ( n3374 & n3527 ) | ( ~n3388 & n3527 ) ;
  assign n3538 = ~n3536 & n3537 ;
  assign n3539 = n3532 | n3538 ;
  assign n3540 = n3262 &  n3389 ;
  assign n3533 = x78 | n3262 ;
  assign n3534 = x78 &  n3262 ;
  assign n3535 = ( n3533 & ~n3534 ) | ( n3533 & 1'b0 ) | ( ~n3534 & 1'b0 ) ;
  assign n3544 = ( n3373 & n3385 ) | ( n3373 & n3535 ) | ( n3385 & n3535 ) ;
  assign n3545 = ( n3373 & ~n3388 ) | ( n3373 & n3535 ) | ( ~n3388 & n3535 ) ;
  assign n3546 = ~n3544 & n3545 ;
  assign n3547 = n3540 | n3546 ;
  assign n3548 = n3270 &  n3389 ;
  assign n3541 = x77 | n3270 ;
  assign n3542 = x77 &  n3270 ;
  assign n3543 = ( n3541 & ~n3542 ) | ( n3541 & 1'b0 ) | ( ~n3542 & 1'b0 ) ;
  assign n3552 = ( n3372 & n3385 ) | ( n3372 & n3543 ) | ( n3385 & n3543 ) ;
  assign n3553 = ( n3372 & ~n3388 ) | ( n3372 & n3543 ) | ( ~n3388 & n3543 ) ;
  assign n3554 = ~n3552 & n3553 ;
  assign n3555 = n3548 | n3554 ;
  assign n3556 = n3278 &  n3389 ;
  assign n3549 = x76 | n3278 ;
  assign n3550 = x76 &  n3278 ;
  assign n3551 = ( n3549 & ~n3550 ) | ( n3549 & 1'b0 ) | ( ~n3550 & 1'b0 ) ;
  assign n3560 = ( n3371 & n3385 ) | ( n3371 & n3551 ) | ( n3385 & n3551 ) ;
  assign n3561 = ( n3371 & ~n3388 ) | ( n3371 & n3551 ) | ( ~n3388 & n3551 ) ;
  assign n3562 = ~n3560 & n3561 ;
  assign n3563 = n3556 | n3562 ;
  assign n3564 = n3286 &  n3389 ;
  assign n3557 = x75 | n3286 ;
  assign n3558 = x75 &  n3286 ;
  assign n3559 = ( n3557 & ~n3558 ) | ( n3557 & 1'b0 ) | ( ~n3558 & 1'b0 ) ;
  assign n3568 = ( n3370 & n3385 ) | ( n3370 & n3559 ) | ( n3385 & n3559 ) ;
  assign n3569 = ( n3370 & ~n3388 ) | ( n3370 & n3559 ) | ( ~n3388 & n3559 ) ;
  assign n3570 = ~n3568 & n3569 ;
  assign n3571 = n3564 | n3570 ;
  assign n3572 = n3294 &  n3389 ;
  assign n3565 = x74 | n3294 ;
  assign n3566 = x74 &  n3294 ;
  assign n3567 = ( n3565 & ~n3566 ) | ( n3565 & 1'b0 ) | ( ~n3566 & 1'b0 ) ;
  assign n3576 = ( n3369 & n3385 ) | ( n3369 & n3567 ) | ( n3385 & n3567 ) ;
  assign n3577 = ( n3369 & ~n3388 ) | ( n3369 & n3567 ) | ( ~n3388 & n3567 ) ;
  assign n3578 = ~n3576 & n3577 ;
  assign n3579 = n3572 | n3578 ;
  assign n3580 = n3302 &  n3389 ;
  assign n3573 = x73 | n3302 ;
  assign n3574 = x73 &  n3302 ;
  assign n3575 = ( n3573 & ~n3574 ) | ( n3573 & 1'b0 ) | ( ~n3574 & 1'b0 ) ;
  assign n3584 = ( n3368 & n3385 ) | ( n3368 & n3575 ) | ( n3385 & n3575 ) ;
  assign n3585 = ( n3368 & ~n3388 ) | ( n3368 & n3575 ) | ( ~n3388 & n3575 ) ;
  assign n3586 = ~n3584 & n3585 ;
  assign n3587 = n3580 | n3586 ;
  assign n3588 = n3310 &  n3389 ;
  assign n3581 = x72 | n3310 ;
  assign n3582 = x72 &  n3310 ;
  assign n3583 = ( n3581 & ~n3582 ) | ( n3581 & 1'b0 ) | ( ~n3582 & 1'b0 ) ;
  assign n3592 = ( n3367 & n3385 ) | ( n3367 & n3583 ) | ( n3385 & n3583 ) ;
  assign n3593 = ( n3367 & ~n3388 ) | ( n3367 & n3583 ) | ( ~n3388 & n3583 ) ;
  assign n3594 = ~n3592 & n3593 ;
  assign n3595 = n3588 | n3594 ;
  assign n3596 = n3318 &  n3389 ;
  assign n3589 = x71 | n3318 ;
  assign n3590 = x71 &  n3318 ;
  assign n3591 = ( n3589 & ~n3590 ) | ( n3589 & 1'b0 ) | ( ~n3590 & 1'b0 ) ;
  assign n3600 = ( n3366 & n3385 ) | ( n3366 & n3591 ) | ( n3385 & n3591 ) ;
  assign n3601 = ( n3366 & ~n3388 ) | ( n3366 & n3591 ) | ( ~n3388 & n3591 ) ;
  assign n3602 = ~n3600 & n3601 ;
  assign n3603 = n3596 | n3602 ;
  assign n3604 = n3326 &  n3389 ;
  assign n3597 = x70 | n3326 ;
  assign n3598 = x70 &  n3326 ;
  assign n3599 = ( n3597 & ~n3598 ) | ( n3597 & 1'b0 ) | ( ~n3598 & 1'b0 ) ;
  assign n3605 = ( n3365 & n3385 ) | ( n3365 & n3599 ) | ( n3385 & n3599 ) ;
  assign n3606 = ( n3365 & ~n3388 ) | ( n3365 & n3599 ) | ( ~n3388 & n3599 ) ;
  assign n3607 = ~n3605 & n3606 ;
  assign n3608 = n3604 | n3607 ;
  assign n3446 = n3331 &  n3389 ;
  assign n3447 = x69 | n3331 ;
  assign n3448 = x69 &  n3331 ;
  assign n3449 = ( n3447 & ~n3448 ) | ( n3447 & 1'b0 ) | ( ~n3448 & 1'b0 ) ;
  assign n3450 = ( n3364 & n3385 ) | ( n3364 & n3449 ) | ( n3385 & n3449 ) ;
  assign n3451 = ( n3364 & ~n3388 ) | ( n3364 & n3449 ) | ( ~n3388 & n3449 ) ;
  assign n3452 = ~n3450 & n3451 ;
  assign n3453 = n3446 | n3452 ;
  assign n3390 = n3168 &  n3389 ;
  assign n3394 = x68 | n3168 ;
  assign n3395 = x68 &  n3168 ;
  assign n3396 = ( n3394 & ~n3395 ) | ( n3394 & 1'b0 ) | ( ~n3395 & 1'b0 ) ;
  assign n3397 = ( n3363 & n3385 ) | ( n3363 & n3396 ) | ( n3385 & n3396 ) ;
  assign n3398 = ( n3363 & ~n3388 ) | ( n3363 & n3396 ) | ( ~n3388 & n3396 ) ;
  assign n3399 = ~n3397 & n3398 ;
  assign n3400 = n3390 | n3399 ;
  assign n3401 = n3340 &  n3389 ;
  assign n3391 = x67 | n3340 ;
  assign n3392 = x67 &  n3340 ;
  assign n3393 = ( n3391 & ~n3392 ) | ( n3391 & 1'b0 ) | ( ~n3392 & 1'b0 ) ;
  assign n3405 = ( n3362 & n3385 ) | ( n3362 & n3393 ) | ( n3385 & n3393 ) ;
  assign n3406 = ( n3362 & ~n3388 ) | ( n3362 & n3393 ) | ( ~n3388 & n3393 ) ;
  assign n3407 = ~n3405 & n3406 ;
  assign n3408 = n3401 | n3407 ;
  assign n3409 = n3346 &  n3389 ;
  assign n3402 = x66 | n3346 ;
  assign n3403 = x66 &  n3346 ;
  assign n3404 = ( n3402 & ~n3403 ) | ( n3402 & 1'b0 ) | ( ~n3403 & 1'b0 ) ;
  assign n3414 = ( n3361 & ~n3385 ) | ( n3361 & n3404 ) | ( ~n3385 & n3404 ) ;
  assign n3415 = ( n3361 & n3388 ) | ( n3361 & n3404 ) | ( n3388 & n3404 ) ;
  assign n3416 = ( n3414 & ~n3415 ) | ( n3414 & 1'b0 ) | ( ~n3415 & 1'b0 ) ;
  assign n3417 = n3409 | n3416 ;
  assign n3418 = n3359 &  n3389 ;
  assign n3410 = x65 &  n3359 ;
  assign n3411 = x65 | n3358 ;
  assign n3412 = n3353 | n3411 ;
  assign n3413 = ( n3360 & ~n3410 ) | ( n3360 & n3412 ) | ( ~n3410 & n3412 ) ;
  assign n3419 = ( x65 & n3359 ) | ( x65 & n3360 ) | ( n3359 & n3360 ) ;
  assign n3420 = ( n3388 & ~n3410 ) | ( n3388 & n3419 ) | ( ~n3410 & n3419 ) ;
  assign n3421 = ( n3385 & n3413 ) | ( n3385 & n3420 ) | ( n3413 & n3420 ) ;
  assign n3422 = ( n3413 & ~n3421 ) | ( n3413 & 1'b0 ) | ( ~n3421 & 1'b0 ) ;
  assign n3423 = n3418 | n3422 ;
  assign n3424 = ( x64 & ~x90 ) | ( x64 & 1'b0 ) | ( ~x90 & 1'b0 ) ;
  assign n3425 = ( n205 & ~n207 ) | ( n205 & n3424 ) | ( ~n207 & n3424 ) ;
  assign n3426 = ~n205 & n3425 ;
  assign n3427 = ( n240 & ~n255 ) | ( n240 & n3426 ) | ( ~n255 & n3426 ) ;
  assign n3428 = ~n240 & n3427 ;
  assign n3429 = n3385 &  n3428 ;
  assign n3430 = ( x38 & ~n3428 ) | ( x38 & n3429 ) | ( ~n3428 & n3429 ) ;
  assign n3431 = ~n177 & n3360 ;
  assign n3432 = ( n188 & ~n273 ) | ( n188 & n3431 ) | ( ~n273 & n3431 ) ;
  assign n3433 = ~n188 & n3432 ;
  assign n3434 = ~n270 & n3433 ;
  assign n3435 = ~n3385 & n3434 ;
  assign n3436 = n3430 | n3435 ;
  assign n3437 = ~x37 & x64 ;
  assign n3438 = ( x65 & ~n3436 ) | ( x65 & n3437 ) | ( ~n3436 & n3437 ) ;
  assign n3439 = ( x66 & ~n3423 ) | ( x66 & n3438 ) | ( ~n3423 & n3438 ) ;
  assign n3440 = ( x67 & ~n3417 ) | ( x67 & n3439 ) | ( ~n3417 & n3439 ) ;
  assign n3441 = ( x68 & ~n3408 ) | ( x68 & n3440 ) | ( ~n3408 & n3440 ) ;
  assign n3445 = ( x69 & ~n3400 ) | ( x69 & n3441 ) | ( ~n3400 & n3441 ) ;
  assign n3609 = ( x70 & ~n3453 ) | ( x70 & n3445 ) | ( ~n3453 & n3445 ) ;
  assign n3610 = ( x71 & ~n3608 ) | ( x71 & n3609 ) | ( ~n3608 & n3609 ) ;
  assign n3611 = ( x72 & ~n3603 ) | ( x72 & n3610 ) | ( ~n3603 & n3610 ) ;
  assign n3612 = ( x73 & ~n3595 ) | ( x73 & n3611 ) | ( ~n3595 & n3611 ) ;
  assign n3613 = ( x74 & ~n3587 ) | ( x74 & n3612 ) | ( ~n3587 & n3612 ) ;
  assign n3614 = ( x75 & ~n3579 ) | ( x75 & n3613 ) | ( ~n3579 & n3613 ) ;
  assign n3615 = ( x76 & ~n3571 ) | ( x76 & n3614 ) | ( ~n3571 & n3614 ) ;
  assign n3616 = ( x77 & ~n3563 ) | ( x77 & n3615 ) | ( ~n3563 & n3615 ) ;
  assign n3617 = ( x78 & ~n3555 ) | ( x78 & n3616 ) | ( ~n3555 & n3616 ) ;
  assign n3618 = ( x79 & ~n3547 ) | ( x79 & n3617 ) | ( ~n3547 & n3617 ) ;
  assign n3619 = ( x80 & ~n3539 ) | ( x80 & n3618 ) | ( ~n3539 & n3618 ) ;
  assign n3620 = ( x81 & ~n3531 ) | ( x81 & n3619 ) | ( ~n3531 & n3619 ) ;
  assign n3621 = ( x82 & ~n3523 ) | ( x82 & n3620 ) | ( ~n3523 & n3620 ) ;
  assign n3622 = ( x83 & ~n3515 ) | ( x83 & n3621 ) | ( ~n3515 & n3621 ) ;
  assign n3623 = ( x84 & ~n3507 ) | ( x84 & n3622 ) | ( ~n3507 & n3622 ) ;
  assign n3624 = ( x85 & ~n3499 ) | ( x85 & n3623 ) | ( ~n3499 & n3623 ) ;
  assign n3625 = ( x86 & ~n3491 ) | ( x86 & n3624 ) | ( ~n3491 & n3624 ) ;
  assign n3626 = ( x87 & ~n3483 ) | ( x87 & n3625 ) | ( ~n3483 & n3625 ) ;
  assign n3627 = ( x88 & ~n3475 ) | ( x88 & n3626 ) | ( ~n3475 & n3626 ) ;
  assign n3628 = ( x89 & ~n3467 ) | ( x89 & n3627 ) | ( ~n3467 & n3627 ) ;
  assign n3632 = n205 | n207 ;
  assign n3633 = ( n255 & ~n240 ) | ( n255 & n3632 ) | ( ~n240 & n3632 ) ;
  assign n3634 = n240 | n3633 ;
  assign n3629 = x89 | n3384 ;
  assign n3630 = ( x89 & n3384 ) | ( x89 & n3388 ) | ( n3384 & n3388 ) ;
  assign n3631 = ( n3174 & ~n3629 ) | ( n3174 & n3630 ) | ( ~n3629 & n3630 ) ;
  assign n3636 = x90 &  n3631 ;
  assign n3635 = x90 | n3631 ;
  assign n3637 = ( n3634 & ~n3636 ) | ( n3634 & n3635 ) | ( ~n3636 & n3635 ) ;
  assign n3638 = n3628 | n3637 ;
  assign n3639 = ~n3631 |  n3388 ;
  assign n3659 = n3467 &  n3639 ;
  assign n3660 = n3638 &  n3659 ;
  assign n3646 = x89 | n3467 ;
  assign n3647 = x89 &  n3467 ;
  assign n3648 = ( n3646 & ~n3647 ) | ( n3646 & 1'b0 ) | ( ~n3647 & 1'b0 ) ;
  assign n3661 = n3627 &  n3648 ;
  assign n3640 = n3638 &  n3639 ;
  assign n3662 = ( n3627 & ~n3640 ) | ( n3627 & n3648 ) | ( ~n3640 & n3648 ) ;
  assign n3663 = ( n3660 & ~n3661 ) | ( n3660 & n3662 ) | ( ~n3661 & n3662 ) ;
  assign n3650 = ( x90 & n3628 ) | ( x90 & n3631 ) | ( n3628 & n3631 ) ;
  assign n3649 = ( x90 & ~n3628 ) | ( x90 & n3631 ) | ( ~n3628 & n3631 ) ;
  assign n3651 = ( n3628 & ~n3650 ) | ( n3628 & n3649 ) | ( ~n3650 & n3649 ) ;
  assign n3652 = ~n3640 & n3651 ;
  assign n3653 = n3174 &  n3388 ;
  assign n3654 = n3638 &  n3653 ;
  assign n3655 = n3652 | n3654 ;
  assign n3667 = n3475 &  n3639 ;
  assign n3668 = n3638 &  n3667 ;
  assign n3656 = x88 | n3475 ;
  assign n3657 = x88 &  n3475 ;
  assign n3658 = ( n3656 & ~n3657 ) | ( n3656 & 1'b0 ) | ( ~n3657 & 1'b0 ) ;
  assign n3669 = n3626 &  n3658 ;
  assign n3670 = ( n3626 & ~n3640 ) | ( n3626 & n3658 ) | ( ~n3640 & n3658 ) ;
  assign n3671 = ( n3668 & ~n3669 ) | ( n3668 & n3670 ) | ( ~n3669 & n3670 ) ;
  assign n3675 = n3483 &  n3639 ;
  assign n3676 = n3638 &  n3675 ;
  assign n3664 = x87 | n3483 ;
  assign n3665 = x87 &  n3483 ;
  assign n3666 = ( n3664 & ~n3665 ) | ( n3664 & 1'b0 ) | ( ~n3665 & 1'b0 ) ;
  assign n3677 = n3625 &  n3666 ;
  assign n3678 = ( n3625 & ~n3640 ) | ( n3625 & n3666 ) | ( ~n3640 & n3666 ) ;
  assign n3679 = ( n3676 & ~n3677 ) | ( n3676 & n3678 ) | ( ~n3677 & n3678 ) ;
  assign n3683 = n3491 &  n3639 ;
  assign n3684 = n3638 &  n3683 ;
  assign n3672 = x86 | n3491 ;
  assign n3673 = x86 &  n3491 ;
  assign n3674 = ( n3672 & ~n3673 ) | ( n3672 & 1'b0 ) | ( ~n3673 & 1'b0 ) ;
  assign n3685 = n3624 &  n3674 ;
  assign n3686 = ( n3624 & ~n3640 ) | ( n3624 & n3674 ) | ( ~n3640 & n3674 ) ;
  assign n3687 = ( n3684 & ~n3685 ) | ( n3684 & n3686 ) | ( ~n3685 & n3686 ) ;
  assign n3691 = n3499 &  n3639 ;
  assign n3692 = n3638 &  n3691 ;
  assign n3680 = x85 | n3499 ;
  assign n3681 = x85 &  n3499 ;
  assign n3682 = ( n3680 & ~n3681 ) | ( n3680 & 1'b0 ) | ( ~n3681 & 1'b0 ) ;
  assign n3693 = n3623 &  n3682 ;
  assign n3694 = ( n3623 & ~n3640 ) | ( n3623 & n3682 ) | ( ~n3640 & n3682 ) ;
  assign n3695 = ( n3692 & ~n3693 ) | ( n3692 & n3694 ) | ( ~n3693 & n3694 ) ;
  assign n3699 = n3507 &  n3639 ;
  assign n3700 = n3638 &  n3699 ;
  assign n3688 = x84 | n3507 ;
  assign n3689 = x84 &  n3507 ;
  assign n3690 = ( n3688 & ~n3689 ) | ( n3688 & 1'b0 ) | ( ~n3689 & 1'b0 ) ;
  assign n3702 = ( n3622 & n3640 ) | ( n3622 & n3690 ) | ( n3640 & n3690 ) ;
  assign n3701 = n3622 | n3690 ;
  assign n3703 = ( n3700 & ~n3702 ) | ( n3700 & n3701 ) | ( ~n3702 & n3701 ) ;
  assign n3707 = n3515 &  n3639 ;
  assign n3708 = n3638 &  n3707 ;
  assign n3696 = x83 | n3515 ;
  assign n3697 = x83 &  n3515 ;
  assign n3698 = ( n3696 & ~n3697 ) | ( n3696 & 1'b0 ) | ( ~n3697 & 1'b0 ) ;
  assign n3710 = ( n3621 & n3640 ) | ( n3621 & n3698 ) | ( n3640 & n3698 ) ;
  assign n3709 = n3621 | n3698 ;
  assign n3711 = ( n3708 & ~n3710 ) | ( n3708 & n3709 ) | ( ~n3710 & n3709 ) ;
  assign n3715 = n3523 &  n3639 ;
  assign n3716 = n3638 &  n3715 ;
  assign n3704 = x82 | n3523 ;
  assign n3705 = x82 &  n3523 ;
  assign n3706 = ( n3704 & ~n3705 ) | ( n3704 & 1'b0 ) | ( ~n3705 & 1'b0 ) ;
  assign n3718 = ( n3620 & n3640 ) | ( n3620 & n3706 ) | ( n3640 & n3706 ) ;
  assign n3717 = n3620 | n3706 ;
  assign n3719 = ( n3716 & ~n3718 ) | ( n3716 & n3717 ) | ( ~n3718 & n3717 ) ;
  assign n3723 = n3531 &  n3639 ;
  assign n3724 = n3638 &  n3723 ;
  assign n3712 = x81 | n3531 ;
  assign n3713 = x81 &  n3531 ;
  assign n3714 = ( n3712 & ~n3713 ) | ( n3712 & 1'b0 ) | ( ~n3713 & 1'b0 ) ;
  assign n3726 = ( n3619 & n3640 ) | ( n3619 & n3714 ) | ( n3640 & n3714 ) ;
  assign n3725 = n3619 | n3714 ;
  assign n3727 = ( n3724 & ~n3726 ) | ( n3724 & n3725 ) | ( ~n3726 & n3725 ) ;
  assign n3731 = n3539 &  n3639 ;
  assign n3732 = n3638 &  n3731 ;
  assign n3720 = x80 | n3539 ;
  assign n3721 = x80 &  n3539 ;
  assign n3722 = ( n3720 & ~n3721 ) | ( n3720 & 1'b0 ) | ( ~n3721 & 1'b0 ) ;
  assign n3734 = ( n3618 & n3640 ) | ( n3618 & n3722 ) | ( n3640 & n3722 ) ;
  assign n3733 = n3618 | n3722 ;
  assign n3735 = ( n3732 & ~n3734 ) | ( n3732 & n3733 ) | ( ~n3734 & n3733 ) ;
  assign n3739 = n3547 &  n3639 ;
  assign n3740 = n3638 &  n3739 ;
  assign n3728 = x79 | n3547 ;
  assign n3729 = x79 &  n3547 ;
  assign n3730 = ( n3728 & ~n3729 ) | ( n3728 & 1'b0 ) | ( ~n3729 & 1'b0 ) ;
  assign n3742 = ( n3617 & n3640 ) | ( n3617 & n3730 ) | ( n3640 & n3730 ) ;
  assign n3741 = n3617 | n3730 ;
  assign n3743 = ( n3740 & ~n3742 ) | ( n3740 & n3741 ) | ( ~n3742 & n3741 ) ;
  assign n3747 = n3555 &  n3639 ;
  assign n3748 = n3638 &  n3747 ;
  assign n3736 = x78 | n3555 ;
  assign n3737 = x78 &  n3555 ;
  assign n3738 = ( n3736 & ~n3737 ) | ( n3736 & 1'b0 ) | ( ~n3737 & 1'b0 ) ;
  assign n3750 = ( n3616 & n3640 ) | ( n3616 & n3738 ) | ( n3640 & n3738 ) ;
  assign n3749 = n3616 | n3738 ;
  assign n3751 = ( n3748 & ~n3750 ) | ( n3748 & n3749 ) | ( ~n3750 & n3749 ) ;
  assign n3755 = n3563 &  n3639 ;
  assign n3756 = n3638 &  n3755 ;
  assign n3744 = x77 | n3563 ;
  assign n3745 = x77 &  n3563 ;
  assign n3746 = ( n3744 & ~n3745 ) | ( n3744 & 1'b0 ) | ( ~n3745 & 1'b0 ) ;
  assign n3758 = ( n3615 & n3640 ) | ( n3615 & n3746 ) | ( n3640 & n3746 ) ;
  assign n3757 = n3615 | n3746 ;
  assign n3759 = ( n3756 & ~n3758 ) | ( n3756 & n3757 ) | ( ~n3758 & n3757 ) ;
  assign n3763 = n3571 &  n3639 ;
  assign n3764 = n3638 &  n3763 ;
  assign n3752 = x76 | n3571 ;
  assign n3753 = x76 &  n3571 ;
  assign n3754 = ( n3752 & ~n3753 ) | ( n3752 & 1'b0 ) | ( ~n3753 & 1'b0 ) ;
  assign n3766 = ( n3614 & n3640 ) | ( n3614 & n3754 ) | ( n3640 & n3754 ) ;
  assign n3765 = n3614 | n3754 ;
  assign n3767 = ( n3764 & ~n3766 ) | ( n3764 & n3765 ) | ( ~n3766 & n3765 ) ;
  assign n3771 = n3579 &  n3639 ;
  assign n3772 = n3638 &  n3771 ;
  assign n3760 = x75 | n3579 ;
  assign n3761 = x75 &  n3579 ;
  assign n3762 = ( n3760 & ~n3761 ) | ( n3760 & 1'b0 ) | ( ~n3761 & 1'b0 ) ;
  assign n3774 = ( n3613 & n3640 ) | ( n3613 & n3762 ) | ( n3640 & n3762 ) ;
  assign n3773 = n3613 | n3762 ;
  assign n3775 = ( n3772 & ~n3774 ) | ( n3772 & n3773 ) | ( ~n3774 & n3773 ) ;
  assign n3779 = n3587 &  n3639 ;
  assign n3780 = n3638 &  n3779 ;
  assign n3768 = x74 | n3587 ;
  assign n3769 = x74 &  n3587 ;
  assign n3770 = ( n3768 & ~n3769 ) | ( n3768 & 1'b0 ) | ( ~n3769 & 1'b0 ) ;
  assign n3782 = ( n3612 & n3640 ) | ( n3612 & n3770 ) | ( n3640 & n3770 ) ;
  assign n3781 = n3612 | n3770 ;
  assign n3783 = ( n3780 & ~n3782 ) | ( n3780 & n3781 ) | ( ~n3782 & n3781 ) ;
  assign n3787 = n3595 &  n3639 ;
  assign n3788 = n3638 &  n3787 ;
  assign n3776 = x73 | n3595 ;
  assign n3777 = x73 &  n3595 ;
  assign n3778 = ( n3776 & ~n3777 ) | ( n3776 & 1'b0 ) | ( ~n3777 & 1'b0 ) ;
  assign n3790 = ( n3611 & n3640 ) | ( n3611 & n3778 ) | ( n3640 & n3778 ) ;
  assign n3789 = n3611 | n3778 ;
  assign n3791 = ( n3788 & ~n3790 ) | ( n3788 & n3789 ) | ( ~n3790 & n3789 ) ;
  assign n3795 = n3603 &  n3639 ;
  assign n3796 = n3638 &  n3795 ;
  assign n3784 = x72 | n3603 ;
  assign n3785 = x72 &  n3603 ;
  assign n3786 = ( n3784 & ~n3785 ) | ( n3784 & 1'b0 ) | ( ~n3785 & 1'b0 ) ;
  assign n3798 = ( n3610 & n3640 ) | ( n3610 & n3786 ) | ( n3640 & n3786 ) ;
  assign n3797 = n3610 | n3786 ;
  assign n3799 = ( n3796 & ~n3798 ) | ( n3796 & n3797 ) | ( ~n3798 & n3797 ) ;
  assign n3800 = n3608 &  n3639 ;
  assign n3801 = n3638 &  n3800 ;
  assign n3792 = x71 | n3608 ;
  assign n3793 = x71 &  n3608 ;
  assign n3794 = ( n3792 & ~n3793 ) | ( n3792 & 1'b0 ) | ( ~n3793 & 1'b0 ) ;
  assign n3803 = ( n3609 & n3640 ) | ( n3609 & n3794 ) | ( n3640 & n3794 ) ;
  assign n3802 = n3609 | n3794 ;
  assign n3804 = ( n3801 & ~n3803 ) | ( n3801 & n3802 ) | ( ~n3803 & n3802 ) ;
  assign n3641 = n3453 &  n3639 ;
  assign n3642 = n3638 &  n3641 ;
  assign n3454 = x70 | n3453 ;
  assign n3455 = x70 &  n3453 ;
  assign n3456 = ( n3454 & ~n3455 ) | ( n3454 & 1'b0 ) | ( ~n3455 & 1'b0 ) ;
  assign n3644 = ( n3445 & n3456 ) | ( n3445 & n3640 ) | ( n3456 & n3640 ) ;
  assign n3643 = n3445 | n3456 ;
  assign n3645 = ( n3642 & ~n3644 ) | ( n3642 & n3643 ) | ( ~n3644 & n3643 ) ;
  assign n3808 = n3400 &  n3639 ;
  assign n3809 = n3638 &  n3808 ;
  assign n3442 = x69 | n3400 ;
  assign n3443 = x69 &  n3400 ;
  assign n3444 = ( n3442 & ~n3443 ) | ( n3442 & 1'b0 ) | ( ~n3443 & 1'b0 ) ;
  assign n3810 = n3441 &  n3444 ;
  assign n3811 = ( n3441 & ~n3640 ) | ( n3441 & n3444 ) | ( ~n3640 & n3444 ) ;
  assign n3812 = ( n3809 & ~n3810 ) | ( n3809 & n3811 ) | ( ~n3810 & n3811 ) ;
  assign n3816 = n3408 &  n3639 ;
  assign n3817 = n3638 &  n3816 ;
  assign n3805 = x68 | n3408 ;
  assign n3806 = x68 &  n3408 ;
  assign n3807 = ( n3805 & ~n3806 ) | ( n3805 & 1'b0 ) | ( ~n3806 & 1'b0 ) ;
  assign n3819 = ( n3440 & n3640 ) | ( n3440 & n3807 ) | ( n3640 & n3807 ) ;
  assign n3818 = n3440 | n3807 ;
  assign n3820 = ( n3817 & ~n3819 ) | ( n3817 & n3818 ) | ( ~n3819 & n3818 ) ;
  assign n3824 = n3417 &  n3639 ;
  assign n3825 = n3638 &  n3824 ;
  assign n3813 = x67 | n3417 ;
  assign n3814 = x67 &  n3417 ;
  assign n3815 = ( n3813 & ~n3814 ) | ( n3813 & 1'b0 ) | ( ~n3814 & 1'b0 ) ;
  assign n3827 = ( n3439 & n3640 ) | ( n3439 & n3815 ) | ( n3640 & n3815 ) ;
  assign n3826 = n3439 | n3815 ;
  assign n3828 = ( n3825 & ~n3827 ) | ( n3825 & n3826 ) | ( ~n3827 & n3826 ) ;
  assign n3829 = n3423 &  n3639 ;
  assign n3830 = n3638 &  n3829 ;
  assign n3821 = x66 | n3423 ;
  assign n3822 = x66 &  n3423 ;
  assign n3823 = ( n3821 & ~n3822 ) | ( n3821 & 1'b0 ) | ( ~n3822 & 1'b0 ) ;
  assign n3831 = n3438 &  n3823 ;
  assign n3832 = ( n3438 & ~n3640 ) | ( n3438 & n3823 ) | ( ~n3640 & n3823 ) ;
  assign n3833 = ( n3830 & ~n3831 ) | ( n3830 & n3832 ) | ( ~n3831 & n3832 ) ;
  assign n3834 = ( n3436 & ~x65 ) | ( n3436 & n3437 ) | ( ~x65 & n3437 ) ;
  assign n3835 = ( n3438 & ~n3437 ) | ( n3438 & n3834 ) | ( ~n3437 & n3834 ) ;
  assign n3836 = ~n3640 & n3835 ;
  assign n3837 = n3436 &  n3639 ;
  assign n3838 = n3638 &  n3837 ;
  assign n3839 = n3836 | n3838 ;
  assign n3840 = ( x64 & ~n3640 ) | ( x64 & 1'b0 ) | ( ~n3640 & 1'b0 ) ;
  assign n3841 = ( x37 & ~n3840 ) | ( x37 & 1'b0 ) | ( ~n3840 & 1'b0 ) ;
  assign n3842 = ( n3437 & ~n3640 ) | ( n3437 & 1'b0 ) | ( ~n3640 & 1'b0 ) ;
  assign n3843 = n3841 | n3842 ;
  assign n3844 = ~x36 & x64 ;
  assign n3845 = ( x65 & ~n3843 ) | ( x65 & n3844 ) | ( ~n3843 & n3844 ) ;
  assign n3846 = ( x66 & ~n3839 ) | ( x66 & n3845 ) | ( ~n3839 & n3845 ) ;
  assign n3847 = ( x67 & ~n3833 ) | ( x67 & n3846 ) | ( ~n3833 & n3846 ) ;
  assign n3848 = ( x68 & ~n3828 ) | ( x68 & n3847 ) | ( ~n3828 & n3847 ) ;
  assign n3849 = ( x69 & ~n3820 ) | ( x69 & n3848 ) | ( ~n3820 & n3848 ) ;
  assign n3850 = ( x70 & ~n3812 ) | ( x70 & n3849 ) | ( ~n3812 & n3849 ) ;
  assign n3851 = ( x71 & ~n3645 ) | ( x71 & n3850 ) | ( ~n3645 & n3850 ) ;
  assign n3852 = ( x72 & ~n3804 ) | ( x72 & n3851 ) | ( ~n3804 & n3851 ) ;
  assign n3853 = ( x73 & ~n3799 ) | ( x73 & n3852 ) | ( ~n3799 & n3852 ) ;
  assign n3854 = ( x74 & ~n3791 ) | ( x74 & n3853 ) | ( ~n3791 & n3853 ) ;
  assign n3855 = ( x75 & ~n3783 ) | ( x75 & n3854 ) | ( ~n3783 & n3854 ) ;
  assign n3856 = ( x76 & ~n3775 ) | ( x76 & n3855 ) | ( ~n3775 & n3855 ) ;
  assign n3857 = ( x77 & ~n3767 ) | ( x77 & n3856 ) | ( ~n3767 & n3856 ) ;
  assign n3858 = ( x78 & ~n3759 ) | ( x78 & n3857 ) | ( ~n3759 & n3857 ) ;
  assign n3859 = ( x79 & ~n3751 ) | ( x79 & n3858 ) | ( ~n3751 & n3858 ) ;
  assign n3860 = ( x80 & ~n3743 ) | ( x80 & n3859 ) | ( ~n3743 & n3859 ) ;
  assign n3861 = ( x81 & ~n3735 ) | ( x81 & n3860 ) | ( ~n3735 & n3860 ) ;
  assign n3862 = ( x82 & ~n3727 ) | ( x82 & n3861 ) | ( ~n3727 & n3861 ) ;
  assign n3863 = ( x83 & ~n3719 ) | ( x83 & n3862 ) | ( ~n3719 & n3862 ) ;
  assign n3864 = ( x84 & ~n3711 ) | ( x84 & n3863 ) | ( ~n3711 & n3863 ) ;
  assign n3865 = ( x85 & ~n3703 ) | ( x85 & n3864 ) | ( ~n3703 & n3864 ) ;
  assign n3866 = ( x86 & ~n3695 ) | ( x86 & n3865 ) | ( ~n3695 & n3865 ) ;
  assign n3867 = ( x87 & ~n3687 ) | ( x87 & n3866 ) | ( ~n3687 & n3866 ) ;
  assign n3868 = ( x88 & ~n3679 ) | ( x88 & n3867 ) | ( ~n3679 & n3867 ) ;
  assign n3869 = ( x89 & ~n3671 ) | ( x89 & n3868 ) | ( ~n3671 & n3868 ) ;
  assign n3870 = ( x90 & ~n3663 ) | ( x90 & n3869 ) | ( ~n3663 & n3869 ) ;
  assign n3871 = ( x91 & ~n3655 ) | ( x91 & n3870 ) | ( ~n3655 & n3870 ) ;
  assign n3872 = n175 | n189 ;
  assign n3873 = n160 | n3872 ;
  assign n3874 = n3871 | n3873 ;
  assign n3892 = n3663 &  n3874 ;
  assign n3886 = x90 | n3663 ;
  assign n3887 = x90 &  n3663 ;
  assign n3888 = ( n3886 & ~n3887 ) | ( n3886 & 1'b0 ) | ( ~n3887 & 1'b0 ) ;
  assign n3896 = ( n3869 & n3871 ) | ( n3869 & n3888 ) | ( n3871 & n3888 ) ;
  assign n3897 = ( n3869 & ~n3873 ) | ( n3869 & n3888 ) | ( ~n3873 & n3888 ) ;
  assign n3898 = ~n3896 & n3897 ;
  assign n3899 = n3892 | n3898 ;
  assign n3889 = x91 | n3870 ;
  assign n3890 = ( x91 & n3870 ) | ( x91 & n3873 ) | ( n3870 & n3873 ) ;
  assign n3891 = ( n3655 & ~n3889 ) | ( n3655 & n3890 ) | ( ~n3889 & n3890 ) ;
  assign n3900 = n3671 &  n3874 ;
  assign n3893 = x89 | n3671 ;
  assign n3894 = x89 &  n3671 ;
  assign n3895 = ( n3893 & ~n3894 ) | ( n3893 & 1'b0 ) | ( ~n3894 & 1'b0 ) ;
  assign n3904 = ( n3868 & n3871 ) | ( n3868 & n3895 ) | ( n3871 & n3895 ) ;
  assign n3905 = ( n3868 & ~n3873 ) | ( n3868 & n3895 ) | ( ~n3873 & n3895 ) ;
  assign n3906 = ~n3904 & n3905 ;
  assign n3907 = n3900 | n3906 ;
  assign n3908 = n3679 &  n3874 ;
  assign n3901 = x88 | n3679 ;
  assign n3902 = x88 &  n3679 ;
  assign n3903 = ( n3901 & ~n3902 ) | ( n3901 & 1'b0 ) | ( ~n3902 & 1'b0 ) ;
  assign n3912 = ( n3867 & n3871 ) | ( n3867 & n3903 ) | ( n3871 & n3903 ) ;
  assign n3913 = ( n3867 & ~n3873 ) | ( n3867 & n3903 ) | ( ~n3873 & n3903 ) ;
  assign n3914 = ~n3912 & n3913 ;
  assign n3915 = n3908 | n3914 ;
  assign n3916 = n3687 &  n3874 ;
  assign n3909 = x87 | n3687 ;
  assign n3910 = x87 &  n3687 ;
  assign n3911 = ( n3909 & ~n3910 ) | ( n3909 & 1'b0 ) | ( ~n3910 & 1'b0 ) ;
  assign n3920 = ( n3866 & n3871 ) | ( n3866 & n3911 ) | ( n3871 & n3911 ) ;
  assign n3921 = ( n3866 & ~n3873 ) | ( n3866 & n3911 ) | ( ~n3873 & n3911 ) ;
  assign n3922 = ~n3920 & n3921 ;
  assign n3923 = n3916 | n3922 ;
  assign n3924 = n3695 &  n3874 ;
  assign n3917 = x86 | n3695 ;
  assign n3918 = x86 &  n3695 ;
  assign n3919 = ( n3917 & ~n3918 ) | ( n3917 & 1'b0 ) | ( ~n3918 & 1'b0 ) ;
  assign n3928 = ( n3865 & n3871 ) | ( n3865 & n3919 ) | ( n3871 & n3919 ) ;
  assign n3929 = ( n3865 & ~n3873 ) | ( n3865 & n3919 ) | ( ~n3873 & n3919 ) ;
  assign n3930 = ~n3928 & n3929 ;
  assign n3931 = n3924 | n3930 ;
  assign n3932 = n3703 &  n3874 ;
  assign n3925 = x85 | n3703 ;
  assign n3926 = x85 &  n3703 ;
  assign n3927 = ( n3925 & ~n3926 ) | ( n3925 & 1'b0 ) | ( ~n3926 & 1'b0 ) ;
  assign n3936 = ( n3864 & n3871 ) | ( n3864 & n3927 ) | ( n3871 & n3927 ) ;
  assign n3937 = ( n3864 & ~n3873 ) | ( n3864 & n3927 ) | ( ~n3873 & n3927 ) ;
  assign n3938 = ~n3936 & n3937 ;
  assign n3939 = n3932 | n3938 ;
  assign n3940 = n3711 &  n3874 ;
  assign n3933 = x84 | n3711 ;
  assign n3934 = x84 &  n3711 ;
  assign n3935 = ( n3933 & ~n3934 ) | ( n3933 & 1'b0 ) | ( ~n3934 & 1'b0 ) ;
  assign n3944 = ( n3863 & n3871 ) | ( n3863 & n3935 ) | ( n3871 & n3935 ) ;
  assign n3945 = ( n3863 & ~n3873 ) | ( n3863 & n3935 ) | ( ~n3873 & n3935 ) ;
  assign n3946 = ~n3944 & n3945 ;
  assign n3947 = n3940 | n3946 ;
  assign n3948 = n3719 &  n3874 ;
  assign n3941 = x83 | n3719 ;
  assign n3942 = x83 &  n3719 ;
  assign n3943 = ( n3941 & ~n3942 ) | ( n3941 & 1'b0 ) | ( ~n3942 & 1'b0 ) ;
  assign n3952 = ( n3862 & n3871 ) | ( n3862 & n3943 ) | ( n3871 & n3943 ) ;
  assign n3953 = ( n3862 & ~n3873 ) | ( n3862 & n3943 ) | ( ~n3873 & n3943 ) ;
  assign n3954 = ~n3952 & n3953 ;
  assign n3955 = n3948 | n3954 ;
  assign n3956 = n3727 &  n3874 ;
  assign n3949 = x82 | n3727 ;
  assign n3950 = x82 &  n3727 ;
  assign n3951 = ( n3949 & ~n3950 ) | ( n3949 & 1'b0 ) | ( ~n3950 & 1'b0 ) ;
  assign n3960 = ( n3861 & n3871 ) | ( n3861 & n3951 ) | ( n3871 & n3951 ) ;
  assign n3961 = ( n3861 & ~n3873 ) | ( n3861 & n3951 ) | ( ~n3873 & n3951 ) ;
  assign n3962 = ~n3960 & n3961 ;
  assign n3963 = n3956 | n3962 ;
  assign n3964 = n3735 &  n3874 ;
  assign n3957 = x81 | n3735 ;
  assign n3958 = x81 &  n3735 ;
  assign n3959 = ( n3957 & ~n3958 ) | ( n3957 & 1'b0 ) | ( ~n3958 & 1'b0 ) ;
  assign n3968 = ( n3860 & n3871 ) | ( n3860 & n3959 ) | ( n3871 & n3959 ) ;
  assign n3969 = ( n3860 & ~n3873 ) | ( n3860 & n3959 ) | ( ~n3873 & n3959 ) ;
  assign n3970 = ~n3968 & n3969 ;
  assign n3971 = n3964 | n3970 ;
  assign n3972 = n3743 &  n3874 ;
  assign n3965 = x80 | n3743 ;
  assign n3966 = x80 &  n3743 ;
  assign n3967 = ( n3965 & ~n3966 ) | ( n3965 & 1'b0 ) | ( ~n3966 & 1'b0 ) ;
  assign n3976 = ( n3859 & n3871 ) | ( n3859 & n3967 ) | ( n3871 & n3967 ) ;
  assign n3977 = ( n3859 & ~n3873 ) | ( n3859 & n3967 ) | ( ~n3873 & n3967 ) ;
  assign n3978 = ~n3976 & n3977 ;
  assign n3979 = n3972 | n3978 ;
  assign n3980 = n3751 &  n3874 ;
  assign n3973 = x79 | n3751 ;
  assign n3974 = x79 &  n3751 ;
  assign n3975 = ( n3973 & ~n3974 ) | ( n3973 & 1'b0 ) | ( ~n3974 & 1'b0 ) ;
  assign n3984 = ( n3858 & n3871 ) | ( n3858 & n3975 ) | ( n3871 & n3975 ) ;
  assign n3985 = ( n3858 & ~n3873 ) | ( n3858 & n3975 ) | ( ~n3873 & n3975 ) ;
  assign n3986 = ~n3984 & n3985 ;
  assign n3987 = n3980 | n3986 ;
  assign n3988 = n3759 &  n3874 ;
  assign n3981 = x78 | n3759 ;
  assign n3982 = x78 &  n3759 ;
  assign n3983 = ( n3981 & ~n3982 ) | ( n3981 & 1'b0 ) | ( ~n3982 & 1'b0 ) ;
  assign n3992 = ( n3857 & n3871 ) | ( n3857 & n3983 ) | ( n3871 & n3983 ) ;
  assign n3993 = ( n3857 & ~n3873 ) | ( n3857 & n3983 ) | ( ~n3873 & n3983 ) ;
  assign n3994 = ~n3992 & n3993 ;
  assign n3995 = n3988 | n3994 ;
  assign n3996 = n3767 &  n3874 ;
  assign n3989 = x77 | n3767 ;
  assign n3990 = x77 &  n3767 ;
  assign n3991 = ( n3989 & ~n3990 ) | ( n3989 & 1'b0 ) | ( ~n3990 & 1'b0 ) ;
  assign n4000 = ( n3856 & n3871 ) | ( n3856 & n3991 ) | ( n3871 & n3991 ) ;
  assign n4001 = ( n3856 & ~n3873 ) | ( n3856 & n3991 ) | ( ~n3873 & n3991 ) ;
  assign n4002 = ~n4000 & n4001 ;
  assign n4003 = n3996 | n4002 ;
  assign n4004 = n3775 &  n3874 ;
  assign n3997 = x76 | n3775 ;
  assign n3998 = x76 &  n3775 ;
  assign n3999 = ( n3997 & ~n3998 ) | ( n3997 & 1'b0 ) | ( ~n3998 & 1'b0 ) ;
  assign n4008 = ( n3855 & n3871 ) | ( n3855 & n3999 ) | ( n3871 & n3999 ) ;
  assign n4009 = ( n3855 & ~n3873 ) | ( n3855 & n3999 ) | ( ~n3873 & n3999 ) ;
  assign n4010 = ~n4008 & n4009 ;
  assign n4011 = n4004 | n4010 ;
  assign n4012 = n3783 &  n3874 ;
  assign n4005 = x75 | n3783 ;
  assign n4006 = x75 &  n3783 ;
  assign n4007 = ( n4005 & ~n4006 ) | ( n4005 & 1'b0 ) | ( ~n4006 & 1'b0 ) ;
  assign n4016 = ( n3854 & n3871 ) | ( n3854 & n4007 ) | ( n3871 & n4007 ) ;
  assign n4017 = ( n3854 & ~n3873 ) | ( n3854 & n4007 ) | ( ~n3873 & n4007 ) ;
  assign n4018 = ~n4016 & n4017 ;
  assign n4019 = n4012 | n4018 ;
  assign n4020 = n3791 &  n3874 ;
  assign n4013 = x74 | n3791 ;
  assign n4014 = x74 &  n3791 ;
  assign n4015 = ( n4013 & ~n4014 ) | ( n4013 & 1'b0 ) | ( ~n4014 & 1'b0 ) ;
  assign n4024 = ( n3853 & n3871 ) | ( n3853 & n4015 ) | ( n3871 & n4015 ) ;
  assign n4025 = ( n3853 & ~n3873 ) | ( n3853 & n4015 ) | ( ~n3873 & n4015 ) ;
  assign n4026 = ~n4024 & n4025 ;
  assign n4027 = n4020 | n4026 ;
  assign n4028 = n3799 &  n3874 ;
  assign n4021 = x73 | n3799 ;
  assign n4022 = x73 &  n3799 ;
  assign n4023 = ( n4021 & ~n4022 ) | ( n4021 & 1'b0 ) | ( ~n4022 & 1'b0 ) ;
  assign n4032 = ( n3852 & n3871 ) | ( n3852 & n4023 ) | ( n3871 & n4023 ) ;
  assign n4033 = ( n3852 & ~n3873 ) | ( n3852 & n4023 ) | ( ~n3873 & n4023 ) ;
  assign n4034 = ~n4032 & n4033 ;
  assign n4035 = n4028 | n4034 ;
  assign n4036 = n3804 &  n3874 ;
  assign n4029 = x72 | n3804 ;
  assign n4030 = x72 &  n3804 ;
  assign n4031 = ( n4029 & ~n4030 ) | ( n4029 & 1'b0 ) | ( ~n4030 & 1'b0 ) ;
  assign n4037 = ( n3851 & n3871 ) | ( n3851 & n4031 ) | ( n3871 & n4031 ) ;
  assign n4038 = ( n3851 & ~n3873 ) | ( n3851 & n4031 ) | ( ~n3873 & n4031 ) ;
  assign n4039 = ~n4037 & n4038 ;
  assign n4040 = n4036 | n4039 ;
  assign n3875 = n3645 &  n3874 ;
  assign n3879 = x71 | n3645 ;
  assign n3880 = x71 &  n3645 ;
  assign n3881 = ( n3879 & ~n3880 ) | ( n3879 & 1'b0 ) | ( ~n3880 & 1'b0 ) ;
  assign n3882 = ( n3850 & n3871 ) | ( n3850 & n3881 ) | ( n3871 & n3881 ) ;
  assign n3883 = ( n3850 & ~n3873 ) | ( n3850 & n3881 ) | ( ~n3873 & n3881 ) ;
  assign n3884 = ~n3882 & n3883 ;
  assign n3885 = n3875 | n3884 ;
  assign n4041 = n3812 &  n3874 ;
  assign n3876 = x70 | n3812 ;
  assign n3877 = x70 &  n3812 ;
  assign n3878 = ( n3876 & ~n3877 ) | ( n3876 & 1'b0 ) | ( ~n3877 & 1'b0 ) ;
  assign n4045 = ( n3849 & n3871 ) | ( n3849 & n3878 ) | ( n3871 & n3878 ) ;
  assign n4046 = ( n3849 & ~n3873 ) | ( n3849 & n3878 ) | ( ~n3873 & n3878 ) ;
  assign n4047 = ~n4045 & n4046 ;
  assign n4048 = n4041 | n4047 ;
  assign n4049 = n3820 &  n3874 ;
  assign n4042 = x69 | n3820 ;
  assign n4043 = x69 &  n3820 ;
  assign n4044 = ( n4042 & ~n4043 ) | ( n4042 & 1'b0 ) | ( ~n4043 & 1'b0 ) ;
  assign n4053 = ( n3848 & n3871 ) | ( n3848 & n4044 ) | ( n3871 & n4044 ) ;
  assign n4054 = ( n3848 & ~n3873 ) | ( n3848 & n4044 ) | ( ~n3873 & n4044 ) ;
  assign n4055 = ~n4053 & n4054 ;
  assign n4056 = n4049 | n4055 ;
  assign n4057 = n3828 &  n3874 ;
  assign n4050 = x68 | n3828 ;
  assign n4051 = x68 &  n3828 ;
  assign n4052 = ( n4050 & ~n4051 ) | ( n4050 & 1'b0 ) | ( ~n4051 & 1'b0 ) ;
  assign n4061 = ( n3847 & n3871 ) | ( n3847 & n4052 ) | ( n3871 & n4052 ) ;
  assign n4062 = ( n3847 & ~n3873 ) | ( n3847 & n4052 ) | ( ~n3873 & n4052 ) ;
  assign n4063 = ~n4061 & n4062 ;
  assign n4064 = n4057 | n4063 ;
  assign n4065 = n3833 &  n3874 ;
  assign n4058 = x67 | n3833 ;
  assign n4059 = x67 &  n3833 ;
  assign n4060 = ( n4058 & ~n4059 ) | ( n4058 & 1'b0 ) | ( ~n4059 & 1'b0 ) ;
  assign n4069 = ( n3846 & n3871 ) | ( n3846 & n4060 ) | ( n3871 & n4060 ) ;
  assign n4070 = ( n3846 & ~n3873 ) | ( n3846 & n4060 ) | ( ~n3873 & n4060 ) ;
  assign n4071 = ~n4069 & n4070 ;
  assign n4072 = n4065 | n4071 ;
  assign n4073 = n3839 &  n3874 ;
  assign n4066 = x66 | n3839 ;
  assign n4067 = x66 &  n3839 ;
  assign n4068 = ( n4066 & ~n4067 ) | ( n4066 & 1'b0 ) | ( ~n4067 & 1'b0 ) ;
  assign n4078 = ( n3845 & ~n3871 ) | ( n3845 & n4068 ) | ( ~n3871 & n4068 ) ;
  assign n4079 = ( n3845 & n3873 ) | ( n3845 & n4068 ) | ( n3873 & n4068 ) ;
  assign n4080 = ( n4078 & ~n4079 ) | ( n4078 & 1'b0 ) | ( ~n4079 & 1'b0 ) ;
  assign n4081 = n4073 | n4080 ;
  assign n4082 = n3843 &  n3874 ;
  assign n4074 = x65 &  n3843 ;
  assign n4075 = ( n3841 & ~x65 ) | ( n3841 & n3842 ) | ( ~x65 & n3842 ) ;
  assign n4076 = x65 | n4075 ;
  assign n4077 = ( n3844 & ~n4074 ) | ( n3844 & n4076 ) | ( ~n4074 & n4076 ) ;
  assign n4083 = ( x65 & n3843 ) | ( x65 & n3844 ) | ( n3843 & n3844 ) ;
  assign n4084 = ( n3873 & ~n4074 ) | ( n3873 & n4083 ) | ( ~n4074 & n4083 ) ;
  assign n4085 = ( n3871 & n4077 ) | ( n3871 & n4084 ) | ( n4077 & n4084 ) ;
  assign n4086 = ( n4077 & ~n4085 ) | ( n4077 & 1'b0 ) | ( ~n4085 & 1'b0 ) ;
  assign n4087 = n4082 | n4086 ;
  assign n4088 = ( x64 & ~x92 ) | ( x64 & 1'b0 ) | ( ~x92 & 1'b0 ) ;
  assign n4089 = ( n205 & ~n255 ) | ( n205 & n4088 ) | ( ~n255 & n4088 ) ;
  assign n4090 = ~n205 & n4089 ;
  assign n4091 = ~n240 & n4090 ;
  assign n4092 = n3871 &  n4091 ;
  assign n4093 = ( x36 & ~n4091 ) | ( x36 & n4092 ) | ( ~n4091 & n4092 ) ;
  assign n4094 = ~n188 & n3844 ;
  assign n4095 = ( n270 & ~n273 ) | ( n270 & n4094 ) | ( ~n273 & n4094 ) ;
  assign n4096 = ~n270 & n4095 ;
  assign n4097 = ~n3871 & n4096 ;
  assign n4098 = n4093 | n4097 ;
  assign n4099 = ~x35 & x64 ;
  assign n4100 = ( x65 & ~n4098 ) | ( x65 & n4099 ) | ( ~n4098 & n4099 ) ;
  assign n4101 = ( x66 & ~n4087 ) | ( x66 & n4100 ) | ( ~n4087 & n4100 ) ;
  assign n4102 = ( x67 & ~n4081 ) | ( x67 & n4101 ) | ( ~n4081 & n4101 ) ;
  assign n4103 = ( x68 & ~n4072 ) | ( x68 & n4102 ) | ( ~n4072 & n4102 ) ;
  assign n4104 = ( x69 & ~n4064 ) | ( x69 & n4103 ) | ( ~n4064 & n4103 ) ;
  assign n4105 = ( x70 & ~n4056 ) | ( x70 & n4104 ) | ( ~n4056 & n4104 ) ;
  assign n4106 = ( x71 & ~n4048 ) | ( x71 & n4105 ) | ( ~n4048 & n4105 ) ;
  assign n4107 = ( x72 & ~n3885 ) | ( x72 & n4106 ) | ( ~n3885 & n4106 ) ;
  assign n4108 = ( x73 & ~n4040 ) | ( x73 & n4107 ) | ( ~n4040 & n4107 ) ;
  assign n4109 = ( x74 & ~n4035 ) | ( x74 & n4108 ) | ( ~n4035 & n4108 ) ;
  assign n4110 = ( x75 & ~n4027 ) | ( x75 & n4109 ) | ( ~n4027 & n4109 ) ;
  assign n4111 = ( x76 & ~n4019 ) | ( x76 & n4110 ) | ( ~n4019 & n4110 ) ;
  assign n4112 = ( x77 & ~n4011 ) | ( x77 & n4111 ) | ( ~n4011 & n4111 ) ;
  assign n4113 = ( x78 & ~n4003 ) | ( x78 & n4112 ) | ( ~n4003 & n4112 ) ;
  assign n4114 = ( x79 & ~n3995 ) | ( x79 & n4113 ) | ( ~n3995 & n4113 ) ;
  assign n4115 = ( x80 & ~n3987 ) | ( x80 & n4114 ) | ( ~n3987 & n4114 ) ;
  assign n4116 = ( x81 & ~n3979 ) | ( x81 & n4115 ) | ( ~n3979 & n4115 ) ;
  assign n4117 = ( x82 & ~n3971 ) | ( x82 & n4116 ) | ( ~n3971 & n4116 ) ;
  assign n4118 = ( x83 & ~n3963 ) | ( x83 & n4117 ) | ( ~n3963 & n4117 ) ;
  assign n4119 = ( x84 & ~n3955 ) | ( x84 & n4118 ) | ( ~n3955 & n4118 ) ;
  assign n4120 = ( x85 & ~n3947 ) | ( x85 & n4119 ) | ( ~n3947 & n4119 ) ;
  assign n4121 = ( x86 & ~n3939 ) | ( x86 & n4120 ) | ( ~n3939 & n4120 ) ;
  assign n4122 = ( x87 & ~n3931 ) | ( x87 & n4121 ) | ( ~n3931 & n4121 ) ;
  assign n4123 = ( x88 & ~n3923 ) | ( x88 & n4122 ) | ( ~n3923 & n4122 ) ;
  assign n4124 = ( x89 & ~n3915 ) | ( x89 & n4123 ) | ( ~n3915 & n4123 ) ;
  assign n4125 = ( x90 & ~n3907 ) | ( x90 & n4124 ) | ( ~n3907 & n4124 ) ;
  assign n4126 = ( x91 & ~n3899 ) | ( x91 & n4125 ) | ( ~n3899 & n4125 ) ;
  assign n4127 = ( x92 & ~n3891 ) | ( x92 & n4126 ) | ( ~n3891 & n4126 ) ;
  assign n4128 = n419 | n428 ;
  assign n4129 = n425 | n4128 ;
  assign n4130 = n4127 | n4129 ;
  assign n4233 = n3899 &  n4130 ;
  assign n4237 = x91 | n3899 ;
  assign n4238 = x91 &  n3899 ;
  assign n4239 = ( n4237 & ~n4238 ) | ( n4237 & 1'b0 ) | ( ~n4238 & 1'b0 ) ;
  assign n4240 = ( n4125 & n4127 ) | ( n4125 & n4239 ) | ( n4127 & n4239 ) ;
  assign n4241 = ( n4125 & ~n4129 ) | ( n4125 & n4239 ) | ( ~n4129 & n4239 ) ;
  assign n4242 = ~n4240 & n4241 ;
  assign n4243 = n4233 | n4242 ;
  assign n4244 = n3907 &  n4130 ;
  assign n4234 = x90 | n3907 ;
  assign n4235 = x90 &  n3907 ;
  assign n4236 = ( n4234 & ~n4235 ) | ( n4234 & 1'b0 ) | ( ~n4235 & 1'b0 ) ;
  assign n4248 = ( n4124 & n4127 ) | ( n4124 & n4236 ) | ( n4127 & n4236 ) ;
  assign n4249 = ( n4124 & ~n4129 ) | ( n4124 & n4236 ) | ( ~n4129 & n4236 ) ;
  assign n4250 = ~n4248 & n4249 ;
  assign n4251 = n4244 | n4250 ;
  assign n4252 = n3915 &  n4130 ;
  assign n4245 = x89 | n3915 ;
  assign n4246 = x89 &  n3915 ;
  assign n4247 = ( n4245 & ~n4246 ) | ( n4245 & 1'b0 ) | ( ~n4246 & 1'b0 ) ;
  assign n4256 = ( n4123 & n4127 ) | ( n4123 & n4247 ) | ( n4127 & n4247 ) ;
  assign n4257 = ( n4123 & ~n4129 ) | ( n4123 & n4247 ) | ( ~n4129 & n4247 ) ;
  assign n4258 = ~n4256 & n4257 ;
  assign n4259 = n4252 | n4258 ;
  assign n4260 = n3923 &  n4130 ;
  assign n4253 = x88 | n3923 ;
  assign n4254 = x88 &  n3923 ;
  assign n4255 = ( n4253 & ~n4254 ) | ( n4253 & 1'b0 ) | ( ~n4254 & 1'b0 ) ;
  assign n4264 = ( n4122 & n4127 ) | ( n4122 & n4255 ) | ( n4127 & n4255 ) ;
  assign n4265 = ( n4122 & ~n4129 ) | ( n4122 & n4255 ) | ( ~n4129 & n4255 ) ;
  assign n4266 = ~n4264 & n4265 ;
  assign n4267 = n4260 | n4266 ;
  assign n4268 = n3931 &  n4130 ;
  assign n4261 = x87 | n3931 ;
  assign n4262 = x87 &  n3931 ;
  assign n4263 = ( n4261 & ~n4262 ) | ( n4261 & 1'b0 ) | ( ~n4262 & 1'b0 ) ;
  assign n4272 = ( n4121 & n4127 ) | ( n4121 & n4263 ) | ( n4127 & n4263 ) ;
  assign n4273 = ( n4121 & ~n4129 ) | ( n4121 & n4263 ) | ( ~n4129 & n4263 ) ;
  assign n4274 = ~n4272 & n4273 ;
  assign n4275 = n4268 | n4274 ;
  assign n4276 = n3939 &  n4130 ;
  assign n4269 = x86 | n3939 ;
  assign n4270 = x86 &  n3939 ;
  assign n4271 = ( n4269 & ~n4270 ) | ( n4269 & 1'b0 ) | ( ~n4270 & 1'b0 ) ;
  assign n4280 = ( n4120 & n4127 ) | ( n4120 & n4271 ) | ( n4127 & n4271 ) ;
  assign n4281 = ( n4120 & ~n4129 ) | ( n4120 & n4271 ) | ( ~n4129 & n4271 ) ;
  assign n4282 = ~n4280 & n4281 ;
  assign n4283 = n4276 | n4282 ;
  assign n4284 = n3947 &  n4130 ;
  assign n4277 = x85 | n3947 ;
  assign n4278 = x85 &  n3947 ;
  assign n4279 = ( n4277 & ~n4278 ) | ( n4277 & 1'b0 ) | ( ~n4278 & 1'b0 ) ;
  assign n4288 = ( n4119 & n4127 ) | ( n4119 & n4279 ) | ( n4127 & n4279 ) ;
  assign n4289 = ( n4119 & ~n4129 ) | ( n4119 & n4279 ) | ( ~n4129 & n4279 ) ;
  assign n4290 = ~n4288 & n4289 ;
  assign n4291 = n4284 | n4290 ;
  assign n4292 = n3955 &  n4130 ;
  assign n4285 = x84 | n3955 ;
  assign n4286 = x84 &  n3955 ;
  assign n4287 = ( n4285 & ~n4286 ) | ( n4285 & 1'b0 ) | ( ~n4286 & 1'b0 ) ;
  assign n4296 = ( n4118 & n4127 ) | ( n4118 & n4287 ) | ( n4127 & n4287 ) ;
  assign n4297 = ( n4118 & ~n4129 ) | ( n4118 & n4287 ) | ( ~n4129 & n4287 ) ;
  assign n4298 = ~n4296 & n4297 ;
  assign n4299 = n4292 | n4298 ;
  assign n4300 = n3963 &  n4130 ;
  assign n4293 = x83 | n3963 ;
  assign n4294 = x83 &  n3963 ;
  assign n4295 = ( n4293 & ~n4294 ) | ( n4293 & 1'b0 ) | ( ~n4294 & 1'b0 ) ;
  assign n4304 = ( n4117 & n4127 ) | ( n4117 & n4295 ) | ( n4127 & n4295 ) ;
  assign n4305 = ( n4117 & ~n4129 ) | ( n4117 & n4295 ) | ( ~n4129 & n4295 ) ;
  assign n4306 = ~n4304 & n4305 ;
  assign n4307 = n4300 | n4306 ;
  assign n4308 = n3971 &  n4130 ;
  assign n4301 = x82 | n3971 ;
  assign n4302 = x82 &  n3971 ;
  assign n4303 = ( n4301 & ~n4302 ) | ( n4301 & 1'b0 ) | ( ~n4302 & 1'b0 ) ;
  assign n4312 = ( n4116 & n4127 ) | ( n4116 & n4303 ) | ( n4127 & n4303 ) ;
  assign n4313 = ( n4116 & ~n4129 ) | ( n4116 & n4303 ) | ( ~n4129 & n4303 ) ;
  assign n4314 = ~n4312 & n4313 ;
  assign n4315 = n4308 | n4314 ;
  assign n4316 = n3979 &  n4130 ;
  assign n4309 = x81 | n3979 ;
  assign n4310 = x81 &  n3979 ;
  assign n4311 = ( n4309 & ~n4310 ) | ( n4309 & 1'b0 ) | ( ~n4310 & 1'b0 ) ;
  assign n4320 = ( n4115 & n4127 ) | ( n4115 & n4311 ) | ( n4127 & n4311 ) ;
  assign n4321 = ( n4115 & ~n4129 ) | ( n4115 & n4311 ) | ( ~n4129 & n4311 ) ;
  assign n4322 = ~n4320 & n4321 ;
  assign n4323 = n4316 | n4322 ;
  assign n4324 = n3987 &  n4130 ;
  assign n4317 = x80 | n3987 ;
  assign n4318 = x80 &  n3987 ;
  assign n4319 = ( n4317 & ~n4318 ) | ( n4317 & 1'b0 ) | ( ~n4318 & 1'b0 ) ;
  assign n4328 = ( n4114 & n4127 ) | ( n4114 & n4319 ) | ( n4127 & n4319 ) ;
  assign n4329 = ( n4114 & ~n4129 ) | ( n4114 & n4319 ) | ( ~n4129 & n4319 ) ;
  assign n4330 = ~n4328 & n4329 ;
  assign n4331 = n4324 | n4330 ;
  assign n4332 = n3995 &  n4130 ;
  assign n4325 = x79 | n3995 ;
  assign n4326 = x79 &  n3995 ;
  assign n4327 = ( n4325 & ~n4326 ) | ( n4325 & 1'b0 ) | ( ~n4326 & 1'b0 ) ;
  assign n4336 = ( n4113 & n4127 ) | ( n4113 & n4327 ) | ( n4127 & n4327 ) ;
  assign n4337 = ( n4113 & ~n4129 ) | ( n4113 & n4327 ) | ( ~n4129 & n4327 ) ;
  assign n4338 = ~n4336 & n4337 ;
  assign n4339 = n4332 | n4338 ;
  assign n4340 = n4003 &  n4130 ;
  assign n4333 = x78 | n4003 ;
  assign n4334 = x78 &  n4003 ;
  assign n4335 = ( n4333 & ~n4334 ) | ( n4333 & 1'b0 ) | ( ~n4334 & 1'b0 ) ;
  assign n4344 = ( n4112 & n4127 ) | ( n4112 & n4335 ) | ( n4127 & n4335 ) ;
  assign n4345 = ( n4112 & ~n4129 ) | ( n4112 & n4335 ) | ( ~n4129 & n4335 ) ;
  assign n4346 = ~n4344 & n4345 ;
  assign n4347 = n4340 | n4346 ;
  assign n4348 = n4011 &  n4130 ;
  assign n4341 = x77 | n4011 ;
  assign n4342 = x77 &  n4011 ;
  assign n4343 = ( n4341 & ~n4342 ) | ( n4341 & 1'b0 ) | ( ~n4342 & 1'b0 ) ;
  assign n4352 = ( n4111 & n4127 ) | ( n4111 & n4343 ) | ( n4127 & n4343 ) ;
  assign n4353 = ( n4111 & ~n4129 ) | ( n4111 & n4343 ) | ( ~n4129 & n4343 ) ;
  assign n4354 = ~n4352 & n4353 ;
  assign n4355 = n4348 | n4354 ;
  assign n4356 = n4019 &  n4130 ;
  assign n4349 = x76 | n4019 ;
  assign n4350 = x76 &  n4019 ;
  assign n4351 = ( n4349 & ~n4350 ) | ( n4349 & 1'b0 ) | ( ~n4350 & 1'b0 ) ;
  assign n4360 = ( n4110 & n4127 ) | ( n4110 & n4351 ) | ( n4127 & n4351 ) ;
  assign n4361 = ( n4110 & ~n4129 ) | ( n4110 & n4351 ) | ( ~n4129 & n4351 ) ;
  assign n4362 = ~n4360 & n4361 ;
  assign n4363 = n4356 | n4362 ;
  assign n4364 = n4027 &  n4130 ;
  assign n4357 = x75 | n4027 ;
  assign n4358 = x75 &  n4027 ;
  assign n4359 = ( n4357 & ~n4358 ) | ( n4357 & 1'b0 ) | ( ~n4358 & 1'b0 ) ;
  assign n4368 = ( n4109 & n4127 ) | ( n4109 & n4359 ) | ( n4127 & n4359 ) ;
  assign n4369 = ( n4109 & ~n4129 ) | ( n4109 & n4359 ) | ( ~n4129 & n4359 ) ;
  assign n4370 = ~n4368 & n4369 ;
  assign n4371 = n4364 | n4370 ;
  assign n4372 = n4035 &  n4130 ;
  assign n4365 = x74 | n4035 ;
  assign n4366 = x74 &  n4035 ;
  assign n4367 = ( n4365 & ~n4366 ) | ( n4365 & 1'b0 ) | ( ~n4366 & 1'b0 ) ;
  assign n4373 = ( n4108 & n4127 ) | ( n4108 & n4367 ) | ( n4127 & n4367 ) ;
  assign n4374 = ( n4108 & ~n4129 ) | ( n4108 & n4367 ) | ( ~n4129 & n4367 ) ;
  assign n4375 = ~n4373 & n4374 ;
  assign n4376 = n4372 | n4375 ;
  assign n4222 = n4040 &  n4130 ;
  assign n4223 = x73 | n4040 ;
  assign n4224 = x73 &  n4040 ;
  assign n4225 = ( n4223 & ~n4224 ) | ( n4223 & 1'b0 ) | ( ~n4224 & 1'b0 ) ;
  assign n4226 = ( n4107 & n4127 ) | ( n4107 & n4225 ) | ( n4127 & n4225 ) ;
  assign n4227 = ( n4107 & ~n4129 ) | ( n4107 & n4225 ) | ( ~n4129 & n4225 ) ;
  assign n4228 = ~n4226 & n4227 ;
  assign n4229 = n4222 | n4228 ;
  assign n4131 = n3885 &  n4130 ;
  assign n4135 = x72 | n3885 ;
  assign n4136 = x72 &  n3885 ;
  assign n4137 = ( n4135 & ~n4136 ) | ( n4135 & 1'b0 ) | ( ~n4136 & 1'b0 ) ;
  assign n4138 = ( n4106 & n4127 ) | ( n4106 & n4137 ) | ( n4127 & n4137 ) ;
  assign n4139 = ( n4106 & ~n4129 ) | ( n4106 & n4137 ) | ( ~n4129 & n4137 ) ;
  assign n4140 = ~n4138 & n4139 ;
  assign n4141 = n4131 | n4140 ;
  assign n4142 = n4048 &  n4130 ;
  assign n4132 = x71 | n4048 ;
  assign n4133 = x71 &  n4048 ;
  assign n4134 = ( n4132 & ~n4133 ) | ( n4132 & 1'b0 ) | ( ~n4133 & 1'b0 ) ;
  assign n4146 = ( n4105 & n4127 ) | ( n4105 & n4134 ) | ( n4127 & n4134 ) ;
  assign n4147 = ( n4105 & ~n4129 ) | ( n4105 & n4134 ) | ( ~n4129 & n4134 ) ;
  assign n4148 = ~n4146 & n4147 ;
  assign n4149 = n4142 | n4148 ;
  assign n4150 = n4056 &  n4130 ;
  assign n4143 = x70 | n4056 ;
  assign n4144 = x70 &  n4056 ;
  assign n4145 = ( n4143 & ~n4144 ) | ( n4143 & 1'b0 ) | ( ~n4144 & 1'b0 ) ;
  assign n4154 = ( n4104 & n4127 ) | ( n4104 & n4145 ) | ( n4127 & n4145 ) ;
  assign n4155 = ( n4104 & ~n4129 ) | ( n4104 & n4145 ) | ( ~n4129 & n4145 ) ;
  assign n4156 = ~n4154 & n4155 ;
  assign n4157 = n4150 | n4156 ;
  assign n4158 = n4064 &  n4130 ;
  assign n4151 = x69 | n4064 ;
  assign n4152 = x69 &  n4064 ;
  assign n4153 = ( n4151 & ~n4152 ) | ( n4151 & 1'b0 ) | ( ~n4152 & 1'b0 ) ;
  assign n4162 = ( n4103 & n4127 ) | ( n4103 & n4153 ) | ( n4127 & n4153 ) ;
  assign n4163 = ( n4103 & ~n4129 ) | ( n4103 & n4153 ) | ( ~n4129 & n4153 ) ;
  assign n4164 = ~n4162 & n4163 ;
  assign n4165 = n4158 | n4164 ;
  assign n4166 = n4072 &  n4130 ;
  assign n4159 = x68 | n4072 ;
  assign n4160 = x68 &  n4072 ;
  assign n4161 = ( n4159 & ~n4160 ) | ( n4159 & 1'b0 ) | ( ~n4160 & 1'b0 ) ;
  assign n4170 = ( n4102 & n4127 ) | ( n4102 & n4161 ) | ( n4127 & n4161 ) ;
  assign n4171 = ( n4102 & ~n4129 ) | ( n4102 & n4161 ) | ( ~n4129 & n4161 ) ;
  assign n4172 = ~n4170 & n4171 ;
  assign n4173 = n4166 | n4172 ;
  assign n4174 = n4081 &  n4130 ;
  assign n4167 = x67 | n4081 ;
  assign n4168 = x67 &  n4081 ;
  assign n4169 = ( n4167 & ~n4168 ) | ( n4167 & 1'b0 ) | ( ~n4168 & 1'b0 ) ;
  assign n4178 = ( n4101 & n4127 ) | ( n4101 & n4169 ) | ( n4127 & n4169 ) ;
  assign n4179 = ( n4101 & ~n4129 ) | ( n4101 & n4169 ) | ( ~n4129 & n4169 ) ;
  assign n4180 = ~n4178 & n4179 ;
  assign n4181 = n4174 | n4180 ;
  assign n4182 = n4087 &  n4130 ;
  assign n4175 = x66 | n4087 ;
  assign n4176 = x66 &  n4087 ;
  assign n4177 = ( n4175 & ~n4176 ) | ( n4175 & 1'b0 ) | ( ~n4176 & 1'b0 ) ;
  assign n4187 = ( n4100 & ~n4127 ) | ( n4100 & n4177 ) | ( ~n4127 & n4177 ) ;
  assign n4188 = ( n4100 & n4129 ) | ( n4100 & n4177 ) | ( n4129 & n4177 ) ;
  assign n4189 = ( n4187 & ~n4188 ) | ( n4187 & 1'b0 ) | ( ~n4188 & 1'b0 ) ;
  assign n4190 = n4182 | n4189 ;
  assign n4191 = n4098 &  n4130 ;
  assign n4183 = x65 &  n4098 ;
  assign n4184 = x65 | n4097 ;
  assign n4185 = n4093 | n4184 ;
  assign n4186 = ( n4099 & ~n4183 ) | ( n4099 & n4185 ) | ( ~n4183 & n4185 ) ;
  assign n4192 = ( x65 & n4098 ) | ( x65 & n4099 ) | ( n4098 & n4099 ) ;
  assign n4193 = ( n4129 & ~n4183 ) | ( n4129 & n4192 ) | ( ~n4183 & n4192 ) ;
  assign n4194 = ( n4127 & n4186 ) | ( n4127 & n4193 ) | ( n4186 & n4193 ) ;
  assign n4195 = ( n4186 & ~n4194 ) | ( n4186 & 1'b0 ) | ( ~n4194 & 1'b0 ) ;
  assign n4196 = n4191 | n4195 ;
  assign n4197 = ( x64 & ~x93 ) | ( x64 & 1'b0 ) | ( ~x93 & 1'b0 ) ;
  assign n4198 = ( n185 & ~n187 ) | ( n185 & n4197 ) | ( ~n187 & n4197 ) ;
  assign n4199 = ~n185 & n4198 ;
  assign n4200 = ( n160 & ~n175 ) | ( n160 & n4199 ) | ( ~n175 & n4199 ) ;
  assign n4201 = ~n160 & n4200 ;
  assign n4202 = n4127 &  n4201 ;
  assign n4203 = ( x35 & ~n4201 ) | ( x35 & n4202 ) | ( ~n4201 & n4202 ) ;
  assign n4204 = ~n205 & n4099 ;
  assign n4205 = ( n240 & ~n255 ) | ( n240 & n4204 ) | ( ~n255 & n4204 ) ;
  assign n4206 = ~n240 & n4205 ;
  assign n4207 = ~n4127 & n4206 ;
  assign n4208 = n4203 | n4207 ;
  assign n4209 = ~x34 & x64 ;
  assign n4210 = ( x65 & ~n4208 ) | ( x65 & n4209 ) | ( ~n4208 & n4209 ) ;
  assign n4211 = ( x66 & ~n4196 ) | ( x66 & n4210 ) | ( ~n4196 & n4210 ) ;
  assign n4212 = ( x67 & ~n4190 ) | ( x67 & n4211 ) | ( ~n4190 & n4211 ) ;
  assign n4213 = ( x68 & ~n4181 ) | ( x68 & n4212 ) | ( ~n4181 & n4212 ) ;
  assign n4214 = ( x69 & ~n4173 ) | ( x69 & n4213 ) | ( ~n4173 & n4213 ) ;
  assign n4215 = ( x70 & ~n4165 ) | ( x70 & n4214 ) | ( ~n4165 & n4214 ) ;
  assign n4216 = ( x71 & ~n4157 ) | ( x71 & n4215 ) | ( ~n4157 & n4215 ) ;
  assign n4217 = ( x72 & ~n4149 ) | ( x72 & n4216 ) | ( ~n4149 & n4216 ) ;
  assign n4221 = ( x73 & ~n4141 ) | ( x73 & n4217 ) | ( ~n4141 & n4217 ) ;
  assign n4377 = ( x74 & ~n4229 ) | ( x74 & n4221 ) | ( ~n4229 & n4221 ) ;
  assign n4378 = ( x75 & ~n4376 ) | ( x75 & n4377 ) | ( ~n4376 & n4377 ) ;
  assign n4379 = ( x76 & ~n4371 ) | ( x76 & n4378 ) | ( ~n4371 & n4378 ) ;
  assign n4380 = ( x77 & ~n4363 ) | ( x77 & n4379 ) | ( ~n4363 & n4379 ) ;
  assign n4381 = ( x78 & ~n4355 ) | ( x78 & n4380 ) | ( ~n4355 & n4380 ) ;
  assign n4382 = ( x79 & ~n4347 ) | ( x79 & n4381 ) | ( ~n4347 & n4381 ) ;
  assign n4383 = ( x80 & ~n4339 ) | ( x80 & n4382 ) | ( ~n4339 & n4382 ) ;
  assign n4384 = ( x81 & ~n4331 ) | ( x81 & n4383 ) | ( ~n4331 & n4383 ) ;
  assign n4385 = ( x82 & ~n4323 ) | ( x82 & n4384 ) | ( ~n4323 & n4384 ) ;
  assign n4386 = ( x83 & ~n4315 ) | ( x83 & n4385 ) | ( ~n4315 & n4385 ) ;
  assign n4387 = ( x84 & ~n4307 ) | ( x84 & n4386 ) | ( ~n4307 & n4386 ) ;
  assign n4388 = ( x85 & ~n4299 ) | ( x85 & n4387 ) | ( ~n4299 & n4387 ) ;
  assign n4389 = ( x86 & ~n4291 ) | ( x86 & n4388 ) | ( ~n4291 & n4388 ) ;
  assign n4390 = ( x87 & ~n4283 ) | ( x87 & n4389 ) | ( ~n4283 & n4389 ) ;
  assign n4391 = ( x88 & ~n4275 ) | ( x88 & n4390 ) | ( ~n4275 & n4390 ) ;
  assign n4392 = ( x89 & ~n4267 ) | ( x89 & n4391 ) | ( ~n4267 & n4391 ) ;
  assign n4393 = ( x90 & ~n4259 ) | ( x90 & n4392 ) | ( ~n4259 & n4392 ) ;
  assign n4394 = ( x91 & ~n4251 ) | ( x91 & n4393 ) | ( ~n4251 & n4393 ) ;
  assign n4395 = ( x92 & ~n4243 ) | ( x92 & n4394 ) | ( ~n4243 & n4394 ) ;
  assign n4399 = n185 | n187 ;
  assign n4400 = ( n175 & ~n160 ) | ( n175 & n4399 ) | ( ~n160 & n4399 ) ;
  assign n4401 = n160 | n4400 ;
  assign n4396 = x92 | n4126 ;
  assign n4397 = ( x92 & n4126 ) | ( x92 & n4129 ) | ( n4126 & n4129 ) ;
  assign n4398 = ( n3891 & ~n4396 ) | ( n3891 & n4397 ) | ( ~n4396 & n4397 ) ;
  assign n4403 = x93 &  n4398 ;
  assign n4402 = x93 | n4398 ;
  assign n4404 = ( n4401 & ~n4403 ) | ( n4401 & n4402 ) | ( ~n4403 & n4402 ) ;
  assign n4405 = n4395 | n4404 ;
  assign n4406 = ~n4398 |  n4129 ;
  assign n4426 = n4243 &  n4406 ;
  assign n4427 = n4405 &  n4426 ;
  assign n4413 = x92 | n4243 ;
  assign n4414 = x92 &  n4243 ;
  assign n4415 = ( n4413 & ~n4414 ) | ( n4413 & 1'b0 ) | ( ~n4414 & 1'b0 ) ;
  assign n4428 = n4394 &  n4415 ;
  assign n4407 = n4405 &  n4406 ;
  assign n4429 = ( n4394 & ~n4407 ) | ( n4394 & n4415 ) | ( ~n4407 & n4415 ) ;
  assign n4430 = ( n4427 & ~n4428 ) | ( n4427 & n4429 ) | ( ~n4428 & n4429 ) ;
  assign n4417 = ( x93 & n4395 ) | ( x93 & n4398 ) | ( n4395 & n4398 ) ;
  assign n4416 = ( x93 & ~n4395 ) | ( x93 & n4398 ) | ( ~n4395 & n4398 ) ;
  assign n4418 = ( n4395 & ~n4417 ) | ( n4395 & n4416 ) | ( ~n4417 & n4416 ) ;
  assign n4419 = ~n4407 & n4418 ;
  assign n4420 = n3891 &  n4129 ;
  assign n4421 = n4405 &  n4420 ;
  assign n4422 = n4419 | n4421 ;
  assign n4434 = n4251 &  n4406 ;
  assign n4435 = n4405 &  n4434 ;
  assign n4423 = x91 | n4251 ;
  assign n4424 = x91 &  n4251 ;
  assign n4425 = ( n4423 & ~n4424 ) | ( n4423 & 1'b0 ) | ( ~n4424 & 1'b0 ) ;
  assign n4436 = n4393 &  n4425 ;
  assign n4437 = ( n4393 & ~n4407 ) | ( n4393 & n4425 ) | ( ~n4407 & n4425 ) ;
  assign n4438 = ( n4435 & ~n4436 ) | ( n4435 & n4437 ) | ( ~n4436 & n4437 ) ;
  assign n4442 = n4259 &  n4406 ;
  assign n4443 = n4405 &  n4442 ;
  assign n4431 = x90 | n4259 ;
  assign n4432 = x90 &  n4259 ;
  assign n4433 = ( n4431 & ~n4432 ) | ( n4431 & 1'b0 ) | ( ~n4432 & 1'b0 ) ;
  assign n4444 = n4392 &  n4433 ;
  assign n4445 = ( n4392 & ~n4407 ) | ( n4392 & n4433 ) | ( ~n4407 & n4433 ) ;
  assign n4446 = ( n4443 & ~n4444 ) | ( n4443 & n4445 ) | ( ~n4444 & n4445 ) ;
  assign n4450 = n4267 &  n4406 ;
  assign n4451 = n4405 &  n4450 ;
  assign n4439 = x89 | n4267 ;
  assign n4440 = x89 &  n4267 ;
  assign n4441 = ( n4439 & ~n4440 ) | ( n4439 & 1'b0 ) | ( ~n4440 & 1'b0 ) ;
  assign n4452 = n4391 &  n4441 ;
  assign n4453 = ( n4391 & ~n4407 ) | ( n4391 & n4441 ) | ( ~n4407 & n4441 ) ;
  assign n4454 = ( n4451 & ~n4452 ) | ( n4451 & n4453 ) | ( ~n4452 & n4453 ) ;
  assign n4458 = n4275 &  n4406 ;
  assign n4459 = n4405 &  n4458 ;
  assign n4447 = x88 | n4275 ;
  assign n4448 = x88 &  n4275 ;
  assign n4449 = ( n4447 & ~n4448 ) | ( n4447 & 1'b0 ) | ( ~n4448 & 1'b0 ) ;
  assign n4460 = n4390 &  n4449 ;
  assign n4461 = ( n4390 & ~n4407 ) | ( n4390 & n4449 ) | ( ~n4407 & n4449 ) ;
  assign n4462 = ( n4459 & ~n4460 ) | ( n4459 & n4461 ) | ( ~n4460 & n4461 ) ;
  assign n4466 = n4283 &  n4406 ;
  assign n4467 = n4405 &  n4466 ;
  assign n4455 = x87 | n4283 ;
  assign n4456 = x87 &  n4283 ;
  assign n4457 = ( n4455 & ~n4456 ) | ( n4455 & 1'b0 ) | ( ~n4456 & 1'b0 ) ;
  assign n4469 = ( n4389 & n4407 ) | ( n4389 & n4457 ) | ( n4407 & n4457 ) ;
  assign n4468 = n4389 | n4457 ;
  assign n4470 = ( n4467 & ~n4469 ) | ( n4467 & n4468 ) | ( ~n4469 & n4468 ) ;
  assign n4474 = n4291 &  n4406 ;
  assign n4475 = n4405 &  n4474 ;
  assign n4463 = x86 | n4291 ;
  assign n4464 = x86 &  n4291 ;
  assign n4465 = ( n4463 & ~n4464 ) | ( n4463 & 1'b0 ) | ( ~n4464 & 1'b0 ) ;
  assign n4477 = ( n4388 & n4407 ) | ( n4388 & n4465 ) | ( n4407 & n4465 ) ;
  assign n4476 = n4388 | n4465 ;
  assign n4478 = ( n4475 & ~n4477 ) | ( n4475 & n4476 ) | ( ~n4477 & n4476 ) ;
  assign n4482 = n4299 &  n4406 ;
  assign n4483 = n4405 &  n4482 ;
  assign n4471 = x85 | n4299 ;
  assign n4472 = x85 &  n4299 ;
  assign n4473 = ( n4471 & ~n4472 ) | ( n4471 & 1'b0 ) | ( ~n4472 & 1'b0 ) ;
  assign n4485 = ( n4387 & n4407 ) | ( n4387 & n4473 ) | ( n4407 & n4473 ) ;
  assign n4484 = n4387 | n4473 ;
  assign n4486 = ( n4483 & ~n4485 ) | ( n4483 & n4484 ) | ( ~n4485 & n4484 ) ;
  assign n4490 = n4307 &  n4406 ;
  assign n4491 = n4405 &  n4490 ;
  assign n4479 = x84 | n4307 ;
  assign n4480 = x84 &  n4307 ;
  assign n4481 = ( n4479 & ~n4480 ) | ( n4479 & 1'b0 ) | ( ~n4480 & 1'b0 ) ;
  assign n4493 = ( n4386 & n4407 ) | ( n4386 & n4481 ) | ( n4407 & n4481 ) ;
  assign n4492 = n4386 | n4481 ;
  assign n4494 = ( n4491 & ~n4493 ) | ( n4491 & n4492 ) | ( ~n4493 & n4492 ) ;
  assign n4498 = n4315 &  n4406 ;
  assign n4499 = n4405 &  n4498 ;
  assign n4487 = x83 | n4315 ;
  assign n4488 = x83 &  n4315 ;
  assign n4489 = ( n4487 & ~n4488 ) | ( n4487 & 1'b0 ) | ( ~n4488 & 1'b0 ) ;
  assign n4501 = ( n4385 & n4407 ) | ( n4385 & n4489 ) | ( n4407 & n4489 ) ;
  assign n4500 = n4385 | n4489 ;
  assign n4502 = ( n4499 & ~n4501 ) | ( n4499 & n4500 ) | ( ~n4501 & n4500 ) ;
  assign n4506 = n4323 &  n4406 ;
  assign n4507 = n4405 &  n4506 ;
  assign n4495 = x82 | n4323 ;
  assign n4496 = x82 &  n4323 ;
  assign n4497 = ( n4495 & ~n4496 ) | ( n4495 & 1'b0 ) | ( ~n4496 & 1'b0 ) ;
  assign n4509 = ( n4384 & n4407 ) | ( n4384 & n4497 ) | ( n4407 & n4497 ) ;
  assign n4508 = n4384 | n4497 ;
  assign n4510 = ( n4507 & ~n4509 ) | ( n4507 & n4508 ) | ( ~n4509 & n4508 ) ;
  assign n4514 = n4331 &  n4406 ;
  assign n4515 = n4405 &  n4514 ;
  assign n4503 = x81 | n4331 ;
  assign n4504 = x81 &  n4331 ;
  assign n4505 = ( n4503 & ~n4504 ) | ( n4503 & 1'b0 ) | ( ~n4504 & 1'b0 ) ;
  assign n4517 = ( n4383 & n4407 ) | ( n4383 & n4505 ) | ( n4407 & n4505 ) ;
  assign n4516 = n4383 | n4505 ;
  assign n4518 = ( n4515 & ~n4517 ) | ( n4515 & n4516 ) | ( ~n4517 & n4516 ) ;
  assign n4522 = n4339 &  n4406 ;
  assign n4523 = n4405 &  n4522 ;
  assign n4511 = x80 | n4339 ;
  assign n4512 = x80 &  n4339 ;
  assign n4513 = ( n4511 & ~n4512 ) | ( n4511 & 1'b0 ) | ( ~n4512 & 1'b0 ) ;
  assign n4525 = ( n4382 & n4407 ) | ( n4382 & n4513 ) | ( n4407 & n4513 ) ;
  assign n4524 = n4382 | n4513 ;
  assign n4526 = ( n4523 & ~n4525 ) | ( n4523 & n4524 ) | ( ~n4525 & n4524 ) ;
  assign n4530 = n4347 &  n4406 ;
  assign n4531 = n4405 &  n4530 ;
  assign n4519 = x79 | n4347 ;
  assign n4520 = x79 &  n4347 ;
  assign n4521 = ( n4519 & ~n4520 ) | ( n4519 & 1'b0 ) | ( ~n4520 & 1'b0 ) ;
  assign n4533 = ( n4381 & n4407 ) | ( n4381 & n4521 ) | ( n4407 & n4521 ) ;
  assign n4532 = n4381 | n4521 ;
  assign n4534 = ( n4531 & ~n4533 ) | ( n4531 & n4532 ) | ( ~n4533 & n4532 ) ;
  assign n4538 = n4355 &  n4406 ;
  assign n4539 = n4405 &  n4538 ;
  assign n4527 = x78 | n4355 ;
  assign n4528 = x78 &  n4355 ;
  assign n4529 = ( n4527 & ~n4528 ) | ( n4527 & 1'b0 ) | ( ~n4528 & 1'b0 ) ;
  assign n4541 = ( n4380 & n4407 ) | ( n4380 & n4529 ) | ( n4407 & n4529 ) ;
  assign n4540 = n4380 | n4529 ;
  assign n4542 = ( n4539 & ~n4541 ) | ( n4539 & n4540 ) | ( ~n4541 & n4540 ) ;
  assign n4546 = n4363 &  n4406 ;
  assign n4547 = n4405 &  n4546 ;
  assign n4535 = x77 | n4363 ;
  assign n4536 = x77 &  n4363 ;
  assign n4537 = ( n4535 & ~n4536 ) | ( n4535 & 1'b0 ) | ( ~n4536 & 1'b0 ) ;
  assign n4549 = ( n4379 & n4407 ) | ( n4379 & n4537 ) | ( n4407 & n4537 ) ;
  assign n4548 = n4379 | n4537 ;
  assign n4550 = ( n4547 & ~n4549 ) | ( n4547 & n4548 ) | ( ~n4549 & n4548 ) ;
  assign n4554 = n4371 &  n4406 ;
  assign n4555 = n4405 &  n4554 ;
  assign n4543 = x76 | n4371 ;
  assign n4544 = x76 &  n4371 ;
  assign n4545 = ( n4543 & ~n4544 ) | ( n4543 & 1'b0 ) | ( ~n4544 & 1'b0 ) ;
  assign n4557 = ( n4378 & n4407 ) | ( n4378 & n4545 ) | ( n4407 & n4545 ) ;
  assign n4556 = n4378 | n4545 ;
  assign n4558 = ( n4555 & ~n4557 ) | ( n4555 & n4556 ) | ( ~n4557 & n4556 ) ;
  assign n4559 = n4376 &  n4406 ;
  assign n4560 = n4405 &  n4559 ;
  assign n4551 = x75 | n4376 ;
  assign n4552 = x75 &  n4376 ;
  assign n4553 = ( n4551 & ~n4552 ) | ( n4551 & 1'b0 ) | ( ~n4552 & 1'b0 ) ;
  assign n4562 = ( n4377 & n4407 ) | ( n4377 & n4553 ) | ( n4407 & n4553 ) ;
  assign n4561 = n4377 | n4553 ;
  assign n4563 = ( n4560 & ~n4562 ) | ( n4560 & n4561 ) | ( ~n4562 & n4561 ) ;
  assign n4408 = n4229 &  n4406 ;
  assign n4409 = n4405 &  n4408 ;
  assign n4230 = x74 | n4229 ;
  assign n4231 = x74 &  n4229 ;
  assign n4232 = ( n4230 & ~n4231 ) | ( n4230 & 1'b0 ) | ( ~n4231 & 1'b0 ) ;
  assign n4411 = ( n4221 & n4232 ) | ( n4221 & n4407 ) | ( n4232 & n4407 ) ;
  assign n4410 = n4221 | n4232 ;
  assign n4412 = ( n4409 & ~n4411 ) | ( n4409 & n4410 ) | ( ~n4411 & n4410 ) ;
  assign n4567 = n4141 &  n4406 ;
  assign n4568 = n4405 &  n4567 ;
  assign n4218 = x73 | n4141 ;
  assign n4219 = x73 &  n4141 ;
  assign n4220 = ( n4218 & ~n4219 ) | ( n4218 & 1'b0 ) | ( ~n4219 & 1'b0 ) ;
  assign n4569 = n4217 &  n4220 ;
  assign n4570 = ( n4217 & ~n4407 ) | ( n4217 & n4220 ) | ( ~n4407 & n4220 ) ;
  assign n4571 = ( n4568 & ~n4569 ) | ( n4568 & n4570 ) | ( ~n4569 & n4570 ) ;
  assign n4575 = n4149 &  n4406 ;
  assign n4576 = n4405 &  n4575 ;
  assign n4564 = x72 | n4149 ;
  assign n4565 = x72 &  n4149 ;
  assign n4566 = ( n4564 & ~n4565 ) | ( n4564 & 1'b0 ) | ( ~n4565 & 1'b0 ) ;
  assign n4578 = ( n4216 & n4407 ) | ( n4216 & n4566 ) | ( n4407 & n4566 ) ;
  assign n4577 = n4216 | n4566 ;
  assign n4579 = ( n4576 & ~n4578 ) | ( n4576 & n4577 ) | ( ~n4578 & n4577 ) ;
  assign n4583 = n4157 &  n4406 ;
  assign n4584 = n4405 &  n4583 ;
  assign n4572 = x71 | n4157 ;
  assign n4573 = x71 &  n4157 ;
  assign n4574 = ( n4572 & ~n4573 ) | ( n4572 & 1'b0 ) | ( ~n4573 & 1'b0 ) ;
  assign n4586 = ( n4215 & n4407 ) | ( n4215 & n4574 ) | ( n4407 & n4574 ) ;
  assign n4585 = n4215 | n4574 ;
  assign n4587 = ( n4584 & ~n4586 ) | ( n4584 & n4585 ) | ( ~n4586 & n4585 ) ;
  assign n4591 = n4165 &  n4406 ;
  assign n4592 = n4405 &  n4591 ;
  assign n4580 = x70 | n4165 ;
  assign n4581 = x70 &  n4165 ;
  assign n4582 = ( n4580 & ~n4581 ) | ( n4580 & 1'b0 ) | ( ~n4581 & 1'b0 ) ;
  assign n4594 = ( n4214 & n4407 ) | ( n4214 & n4582 ) | ( n4407 & n4582 ) ;
  assign n4593 = n4214 | n4582 ;
  assign n4595 = ( n4592 & ~n4594 ) | ( n4592 & n4593 ) | ( ~n4594 & n4593 ) ;
  assign n4599 = n4173 &  n4406 ;
  assign n4600 = n4405 &  n4599 ;
  assign n4588 = x69 | n4173 ;
  assign n4589 = x69 &  n4173 ;
  assign n4590 = ( n4588 & ~n4589 ) | ( n4588 & 1'b0 ) | ( ~n4589 & 1'b0 ) ;
  assign n4602 = ( n4213 & n4407 ) | ( n4213 & n4590 ) | ( n4407 & n4590 ) ;
  assign n4601 = n4213 | n4590 ;
  assign n4603 = ( n4600 & ~n4602 ) | ( n4600 & n4601 ) | ( ~n4602 & n4601 ) ;
  assign n4607 = n4181 &  n4406 ;
  assign n4608 = n4405 &  n4607 ;
  assign n4596 = x68 | n4181 ;
  assign n4597 = x68 &  n4181 ;
  assign n4598 = ( n4596 & ~n4597 ) | ( n4596 & 1'b0 ) | ( ~n4597 & 1'b0 ) ;
  assign n4610 = ( n4212 & n4407 ) | ( n4212 & n4598 ) | ( n4407 & n4598 ) ;
  assign n4609 = n4212 | n4598 ;
  assign n4611 = ( n4608 & ~n4610 ) | ( n4608 & n4609 ) | ( ~n4610 & n4609 ) ;
  assign n4615 = n4190 &  n4406 ;
  assign n4616 = n4405 &  n4615 ;
  assign n4604 = x67 | n4190 ;
  assign n4605 = x67 &  n4190 ;
  assign n4606 = ( n4604 & ~n4605 ) | ( n4604 & 1'b0 ) | ( ~n4605 & 1'b0 ) ;
  assign n4618 = ( n4211 & n4407 ) | ( n4211 & n4606 ) | ( n4407 & n4606 ) ;
  assign n4617 = n4211 | n4606 ;
  assign n4619 = ( n4616 & ~n4618 ) | ( n4616 & n4617 ) | ( ~n4618 & n4617 ) ;
  assign n4620 = n4196 &  n4406 ;
  assign n4621 = n4405 &  n4620 ;
  assign n4612 = x66 | n4196 ;
  assign n4613 = x66 &  n4196 ;
  assign n4614 = ( n4612 & ~n4613 ) | ( n4612 & 1'b0 ) | ( ~n4613 & 1'b0 ) ;
  assign n4622 = n4210 &  n4614 ;
  assign n4623 = ( n4210 & ~n4407 ) | ( n4210 & n4614 ) | ( ~n4407 & n4614 ) ;
  assign n4624 = ( n4621 & ~n4622 ) | ( n4621 & n4623 ) | ( ~n4622 & n4623 ) ;
  assign n4625 = ( n4208 & ~x65 ) | ( n4208 & n4209 ) | ( ~x65 & n4209 ) ;
  assign n4626 = ( n4210 & ~n4209 ) | ( n4210 & n4625 ) | ( ~n4209 & n4625 ) ;
  assign n4627 = ~n4407 & n4626 ;
  assign n4628 = n4208 &  n4406 ;
  assign n4629 = n4405 &  n4628 ;
  assign n4630 = n4627 | n4629 ;
  assign n4631 = ( x64 & ~n4407 ) | ( x64 & 1'b0 ) | ( ~n4407 & 1'b0 ) ;
  assign n4632 = ( x34 & ~n4631 ) | ( x34 & 1'b0 ) | ( ~n4631 & 1'b0 ) ;
  assign n4633 = ( n4209 & ~n4407 ) | ( n4209 & 1'b0 ) | ( ~n4407 & 1'b0 ) ;
  assign n4634 = n4632 | n4633 ;
  assign n4635 = ~x33 & x64 ;
  assign n4636 = ( x65 & ~n4634 ) | ( x65 & n4635 ) | ( ~n4634 & n4635 ) ;
  assign n4637 = ( x66 & ~n4630 ) | ( x66 & n4636 ) | ( ~n4630 & n4636 ) ;
  assign n4638 = ( x67 & ~n4624 ) | ( x67 & n4637 ) | ( ~n4624 & n4637 ) ;
  assign n4639 = ( x68 & ~n4619 ) | ( x68 & n4638 ) | ( ~n4619 & n4638 ) ;
  assign n4640 = ( x69 & ~n4611 ) | ( x69 & n4639 ) | ( ~n4611 & n4639 ) ;
  assign n4641 = ( x70 & ~n4603 ) | ( x70 & n4640 ) | ( ~n4603 & n4640 ) ;
  assign n4642 = ( x71 & ~n4595 ) | ( x71 & n4641 ) | ( ~n4595 & n4641 ) ;
  assign n4643 = ( x72 & ~n4587 ) | ( x72 & n4642 ) | ( ~n4587 & n4642 ) ;
  assign n4644 = ( x73 & ~n4579 ) | ( x73 & n4643 ) | ( ~n4579 & n4643 ) ;
  assign n4645 = ( x74 & ~n4571 ) | ( x74 & n4644 ) | ( ~n4571 & n4644 ) ;
  assign n4646 = ( x75 & ~n4412 ) | ( x75 & n4645 ) | ( ~n4412 & n4645 ) ;
  assign n4647 = ( x76 & ~n4563 ) | ( x76 & n4646 ) | ( ~n4563 & n4646 ) ;
  assign n4648 = ( x77 & ~n4558 ) | ( x77 & n4647 ) | ( ~n4558 & n4647 ) ;
  assign n4649 = ( x78 & ~n4550 ) | ( x78 & n4648 ) | ( ~n4550 & n4648 ) ;
  assign n4650 = ( x79 & ~n4542 ) | ( x79 & n4649 ) | ( ~n4542 & n4649 ) ;
  assign n4651 = ( x80 & ~n4534 ) | ( x80 & n4650 ) | ( ~n4534 & n4650 ) ;
  assign n4652 = ( x81 & ~n4526 ) | ( x81 & n4651 ) | ( ~n4526 & n4651 ) ;
  assign n4653 = ( x82 & ~n4518 ) | ( x82 & n4652 ) | ( ~n4518 & n4652 ) ;
  assign n4654 = ( x83 & ~n4510 ) | ( x83 & n4653 ) | ( ~n4510 & n4653 ) ;
  assign n4655 = ( x84 & ~n4502 ) | ( x84 & n4654 ) | ( ~n4502 & n4654 ) ;
  assign n4656 = ( x85 & ~n4494 ) | ( x85 & n4655 ) | ( ~n4494 & n4655 ) ;
  assign n4657 = ( x86 & ~n4486 ) | ( x86 & n4656 ) | ( ~n4486 & n4656 ) ;
  assign n4658 = ( x87 & ~n4478 ) | ( x87 & n4657 ) | ( ~n4478 & n4657 ) ;
  assign n4659 = ( x88 & ~n4470 ) | ( x88 & n4658 ) | ( ~n4470 & n4658 ) ;
  assign n4660 = ( x89 & ~n4462 ) | ( x89 & n4659 ) | ( ~n4462 & n4659 ) ;
  assign n4661 = ( x90 & ~n4454 ) | ( x90 & n4660 ) | ( ~n4454 & n4660 ) ;
  assign n4662 = ( x91 & ~n4446 ) | ( x91 & n4661 ) | ( ~n4446 & n4661 ) ;
  assign n4663 = ( x92 & ~n4438 ) | ( x92 & n4662 ) | ( ~n4438 & n4662 ) ;
  assign n4664 = ( x93 & ~n4430 ) | ( x93 & n4663 ) | ( ~n4430 & n4663 ) ;
  assign n4665 = ( x94 & ~n4422 ) | ( x94 & n4664 ) | ( ~n4422 & n4664 ) ;
  assign n4666 = n204 | n246 ;
  assign n4667 = ( n428 & ~n425 ) | ( n428 & n4666 ) | ( ~n425 & n4666 ) ;
  assign n4668 = n425 | n4667 ;
  assign n4669 = n4665 | n4668 ;
  assign n4687 = n4430 &  n4669 ;
  assign n4681 = x93 | n4430 ;
  assign n4682 = x93 &  n4430 ;
  assign n4683 = ( n4681 & ~n4682 ) | ( n4681 & 1'b0 ) | ( ~n4682 & 1'b0 ) ;
  assign n4691 = ( n4663 & n4665 ) | ( n4663 & n4683 ) | ( n4665 & n4683 ) ;
  assign n4692 = ( n4663 & ~n4668 ) | ( n4663 & n4683 ) | ( ~n4668 & n4683 ) ;
  assign n4693 = ~n4691 & n4692 ;
  assign n4694 = n4687 | n4693 ;
  assign n4684 = x94 | n4664 ;
  assign n4685 = ( x94 & n4664 ) | ( x94 & n4668 ) | ( n4664 & n4668 ) ;
  assign n4686 = ( n4422 & ~n4684 ) | ( n4422 & n4685 ) | ( ~n4684 & n4685 ) ;
  assign n4695 = n4438 &  n4669 ;
  assign n4688 = x92 | n4438 ;
  assign n4689 = x92 &  n4438 ;
  assign n4690 = ( n4688 & ~n4689 ) | ( n4688 & 1'b0 ) | ( ~n4689 & 1'b0 ) ;
  assign n4699 = ( n4662 & n4665 ) | ( n4662 & n4690 ) | ( n4665 & n4690 ) ;
  assign n4700 = ( n4662 & ~n4668 ) | ( n4662 & n4690 ) | ( ~n4668 & n4690 ) ;
  assign n4701 = ~n4699 & n4700 ;
  assign n4702 = n4695 | n4701 ;
  assign n4703 = n4446 &  n4669 ;
  assign n4696 = x91 | n4446 ;
  assign n4697 = x91 &  n4446 ;
  assign n4698 = ( n4696 & ~n4697 ) | ( n4696 & 1'b0 ) | ( ~n4697 & 1'b0 ) ;
  assign n4707 = ( n4661 & n4665 ) | ( n4661 & n4698 ) | ( n4665 & n4698 ) ;
  assign n4708 = ( n4661 & ~n4668 ) | ( n4661 & n4698 ) | ( ~n4668 & n4698 ) ;
  assign n4709 = ~n4707 & n4708 ;
  assign n4710 = n4703 | n4709 ;
  assign n4711 = n4454 &  n4669 ;
  assign n4704 = x90 | n4454 ;
  assign n4705 = x90 &  n4454 ;
  assign n4706 = ( n4704 & ~n4705 ) | ( n4704 & 1'b0 ) | ( ~n4705 & 1'b0 ) ;
  assign n4715 = ( n4660 & n4665 ) | ( n4660 & n4706 ) | ( n4665 & n4706 ) ;
  assign n4716 = ( n4660 & ~n4668 ) | ( n4660 & n4706 ) | ( ~n4668 & n4706 ) ;
  assign n4717 = ~n4715 & n4716 ;
  assign n4718 = n4711 | n4717 ;
  assign n4719 = n4462 &  n4669 ;
  assign n4712 = x89 | n4462 ;
  assign n4713 = x89 &  n4462 ;
  assign n4714 = ( n4712 & ~n4713 ) | ( n4712 & 1'b0 ) | ( ~n4713 & 1'b0 ) ;
  assign n4723 = ( n4659 & n4665 ) | ( n4659 & n4714 ) | ( n4665 & n4714 ) ;
  assign n4724 = ( n4659 & ~n4668 ) | ( n4659 & n4714 ) | ( ~n4668 & n4714 ) ;
  assign n4725 = ~n4723 & n4724 ;
  assign n4726 = n4719 | n4725 ;
  assign n4727 = n4470 &  n4669 ;
  assign n4720 = x88 | n4470 ;
  assign n4721 = x88 &  n4470 ;
  assign n4722 = ( n4720 & ~n4721 ) | ( n4720 & 1'b0 ) | ( ~n4721 & 1'b0 ) ;
  assign n4731 = ( n4658 & n4665 ) | ( n4658 & n4722 ) | ( n4665 & n4722 ) ;
  assign n4732 = ( n4658 & ~n4668 ) | ( n4658 & n4722 ) | ( ~n4668 & n4722 ) ;
  assign n4733 = ~n4731 & n4732 ;
  assign n4734 = n4727 | n4733 ;
  assign n4735 = n4478 &  n4669 ;
  assign n4728 = x87 | n4478 ;
  assign n4729 = x87 &  n4478 ;
  assign n4730 = ( n4728 & ~n4729 ) | ( n4728 & 1'b0 ) | ( ~n4729 & 1'b0 ) ;
  assign n4739 = ( n4657 & n4665 ) | ( n4657 & n4730 ) | ( n4665 & n4730 ) ;
  assign n4740 = ( n4657 & ~n4668 ) | ( n4657 & n4730 ) | ( ~n4668 & n4730 ) ;
  assign n4741 = ~n4739 & n4740 ;
  assign n4742 = n4735 | n4741 ;
  assign n4743 = n4486 &  n4669 ;
  assign n4736 = x86 | n4486 ;
  assign n4737 = x86 &  n4486 ;
  assign n4738 = ( n4736 & ~n4737 ) | ( n4736 & 1'b0 ) | ( ~n4737 & 1'b0 ) ;
  assign n4747 = ( n4656 & n4665 ) | ( n4656 & n4738 ) | ( n4665 & n4738 ) ;
  assign n4748 = ( n4656 & ~n4668 ) | ( n4656 & n4738 ) | ( ~n4668 & n4738 ) ;
  assign n4749 = ~n4747 & n4748 ;
  assign n4750 = n4743 | n4749 ;
  assign n4751 = n4494 &  n4669 ;
  assign n4744 = x85 | n4494 ;
  assign n4745 = x85 &  n4494 ;
  assign n4746 = ( n4744 & ~n4745 ) | ( n4744 & 1'b0 ) | ( ~n4745 & 1'b0 ) ;
  assign n4755 = ( n4655 & n4665 ) | ( n4655 & n4746 ) | ( n4665 & n4746 ) ;
  assign n4756 = ( n4655 & ~n4668 ) | ( n4655 & n4746 ) | ( ~n4668 & n4746 ) ;
  assign n4757 = ~n4755 & n4756 ;
  assign n4758 = n4751 | n4757 ;
  assign n4759 = n4502 &  n4669 ;
  assign n4752 = x84 | n4502 ;
  assign n4753 = x84 &  n4502 ;
  assign n4754 = ( n4752 & ~n4753 ) | ( n4752 & 1'b0 ) | ( ~n4753 & 1'b0 ) ;
  assign n4763 = ( n4654 & n4665 ) | ( n4654 & n4754 ) | ( n4665 & n4754 ) ;
  assign n4764 = ( n4654 & ~n4668 ) | ( n4654 & n4754 ) | ( ~n4668 & n4754 ) ;
  assign n4765 = ~n4763 & n4764 ;
  assign n4766 = n4759 | n4765 ;
  assign n4767 = n4510 &  n4669 ;
  assign n4760 = x83 | n4510 ;
  assign n4761 = x83 &  n4510 ;
  assign n4762 = ( n4760 & ~n4761 ) | ( n4760 & 1'b0 ) | ( ~n4761 & 1'b0 ) ;
  assign n4771 = ( n4653 & n4665 ) | ( n4653 & n4762 ) | ( n4665 & n4762 ) ;
  assign n4772 = ( n4653 & ~n4668 ) | ( n4653 & n4762 ) | ( ~n4668 & n4762 ) ;
  assign n4773 = ~n4771 & n4772 ;
  assign n4774 = n4767 | n4773 ;
  assign n4775 = n4518 &  n4669 ;
  assign n4768 = x82 | n4518 ;
  assign n4769 = x82 &  n4518 ;
  assign n4770 = ( n4768 & ~n4769 ) | ( n4768 & 1'b0 ) | ( ~n4769 & 1'b0 ) ;
  assign n4779 = ( n4652 & n4665 ) | ( n4652 & n4770 ) | ( n4665 & n4770 ) ;
  assign n4780 = ( n4652 & ~n4668 ) | ( n4652 & n4770 ) | ( ~n4668 & n4770 ) ;
  assign n4781 = ~n4779 & n4780 ;
  assign n4782 = n4775 | n4781 ;
  assign n4783 = n4526 &  n4669 ;
  assign n4776 = x81 | n4526 ;
  assign n4777 = x81 &  n4526 ;
  assign n4778 = ( n4776 & ~n4777 ) | ( n4776 & 1'b0 ) | ( ~n4777 & 1'b0 ) ;
  assign n4787 = ( n4651 & n4665 ) | ( n4651 & n4778 ) | ( n4665 & n4778 ) ;
  assign n4788 = ( n4651 & ~n4668 ) | ( n4651 & n4778 ) | ( ~n4668 & n4778 ) ;
  assign n4789 = ~n4787 & n4788 ;
  assign n4790 = n4783 | n4789 ;
  assign n4791 = n4534 &  n4669 ;
  assign n4784 = x80 | n4534 ;
  assign n4785 = x80 &  n4534 ;
  assign n4786 = ( n4784 & ~n4785 ) | ( n4784 & 1'b0 ) | ( ~n4785 & 1'b0 ) ;
  assign n4795 = ( n4650 & n4665 ) | ( n4650 & n4786 ) | ( n4665 & n4786 ) ;
  assign n4796 = ( n4650 & ~n4668 ) | ( n4650 & n4786 ) | ( ~n4668 & n4786 ) ;
  assign n4797 = ~n4795 & n4796 ;
  assign n4798 = n4791 | n4797 ;
  assign n4799 = n4542 &  n4669 ;
  assign n4792 = x79 | n4542 ;
  assign n4793 = x79 &  n4542 ;
  assign n4794 = ( n4792 & ~n4793 ) | ( n4792 & 1'b0 ) | ( ~n4793 & 1'b0 ) ;
  assign n4803 = ( n4649 & n4665 ) | ( n4649 & n4794 ) | ( n4665 & n4794 ) ;
  assign n4804 = ( n4649 & ~n4668 ) | ( n4649 & n4794 ) | ( ~n4668 & n4794 ) ;
  assign n4805 = ~n4803 & n4804 ;
  assign n4806 = n4799 | n4805 ;
  assign n4807 = n4550 &  n4669 ;
  assign n4800 = x78 | n4550 ;
  assign n4801 = x78 &  n4550 ;
  assign n4802 = ( n4800 & ~n4801 ) | ( n4800 & 1'b0 ) | ( ~n4801 & 1'b0 ) ;
  assign n4811 = ( n4648 & n4665 ) | ( n4648 & n4802 ) | ( n4665 & n4802 ) ;
  assign n4812 = ( n4648 & ~n4668 ) | ( n4648 & n4802 ) | ( ~n4668 & n4802 ) ;
  assign n4813 = ~n4811 & n4812 ;
  assign n4814 = n4807 | n4813 ;
  assign n4815 = n4558 &  n4669 ;
  assign n4808 = x77 | n4558 ;
  assign n4809 = x77 &  n4558 ;
  assign n4810 = ( n4808 & ~n4809 ) | ( n4808 & 1'b0 ) | ( ~n4809 & 1'b0 ) ;
  assign n4819 = ( n4647 & n4665 ) | ( n4647 & n4810 ) | ( n4665 & n4810 ) ;
  assign n4820 = ( n4647 & ~n4668 ) | ( n4647 & n4810 ) | ( ~n4668 & n4810 ) ;
  assign n4821 = ~n4819 & n4820 ;
  assign n4822 = n4815 | n4821 ;
  assign n4823 = n4563 &  n4669 ;
  assign n4816 = x76 | n4563 ;
  assign n4817 = x76 &  n4563 ;
  assign n4818 = ( n4816 & ~n4817 ) | ( n4816 & 1'b0 ) | ( ~n4817 & 1'b0 ) ;
  assign n4824 = ( n4646 & n4665 ) | ( n4646 & n4818 ) | ( n4665 & n4818 ) ;
  assign n4825 = ( n4646 & ~n4668 ) | ( n4646 & n4818 ) | ( ~n4668 & n4818 ) ;
  assign n4826 = ~n4824 & n4825 ;
  assign n4827 = n4823 | n4826 ;
  assign n4670 = n4412 &  n4669 ;
  assign n4674 = x75 | n4412 ;
  assign n4675 = x75 &  n4412 ;
  assign n4676 = ( n4674 & ~n4675 ) | ( n4674 & 1'b0 ) | ( ~n4675 & 1'b0 ) ;
  assign n4677 = ( n4645 & n4665 ) | ( n4645 & n4676 ) | ( n4665 & n4676 ) ;
  assign n4678 = ( n4645 & ~n4668 ) | ( n4645 & n4676 ) | ( ~n4668 & n4676 ) ;
  assign n4679 = ~n4677 & n4678 ;
  assign n4680 = n4670 | n4679 ;
  assign n4828 = n4571 &  n4669 ;
  assign n4671 = x74 | n4571 ;
  assign n4672 = x74 &  n4571 ;
  assign n4673 = ( n4671 & ~n4672 ) | ( n4671 & 1'b0 ) | ( ~n4672 & 1'b0 ) ;
  assign n4832 = ( n4644 & n4665 ) | ( n4644 & n4673 ) | ( n4665 & n4673 ) ;
  assign n4833 = ( n4644 & ~n4668 ) | ( n4644 & n4673 ) | ( ~n4668 & n4673 ) ;
  assign n4834 = ~n4832 & n4833 ;
  assign n4835 = n4828 | n4834 ;
  assign n4836 = n4579 &  n4669 ;
  assign n4829 = x73 | n4579 ;
  assign n4830 = x73 &  n4579 ;
  assign n4831 = ( n4829 & ~n4830 ) | ( n4829 & 1'b0 ) | ( ~n4830 & 1'b0 ) ;
  assign n4840 = ( n4643 & n4665 ) | ( n4643 & n4831 ) | ( n4665 & n4831 ) ;
  assign n4841 = ( n4643 & ~n4668 ) | ( n4643 & n4831 ) | ( ~n4668 & n4831 ) ;
  assign n4842 = ~n4840 & n4841 ;
  assign n4843 = n4836 | n4842 ;
  assign n4844 = n4587 &  n4669 ;
  assign n4837 = x72 | n4587 ;
  assign n4838 = x72 &  n4587 ;
  assign n4839 = ( n4837 & ~n4838 ) | ( n4837 & 1'b0 ) | ( ~n4838 & 1'b0 ) ;
  assign n4848 = ( n4642 & n4665 ) | ( n4642 & n4839 ) | ( n4665 & n4839 ) ;
  assign n4849 = ( n4642 & ~n4668 ) | ( n4642 & n4839 ) | ( ~n4668 & n4839 ) ;
  assign n4850 = ~n4848 & n4849 ;
  assign n4851 = n4844 | n4850 ;
  assign n4852 = n4595 &  n4669 ;
  assign n4845 = x71 | n4595 ;
  assign n4846 = x71 &  n4595 ;
  assign n4847 = ( n4845 & ~n4846 ) | ( n4845 & 1'b0 ) | ( ~n4846 & 1'b0 ) ;
  assign n4856 = ( n4641 & n4665 ) | ( n4641 & n4847 ) | ( n4665 & n4847 ) ;
  assign n4857 = ( n4641 & ~n4668 ) | ( n4641 & n4847 ) | ( ~n4668 & n4847 ) ;
  assign n4858 = ~n4856 & n4857 ;
  assign n4859 = n4852 | n4858 ;
  assign n4860 = n4603 &  n4669 ;
  assign n4853 = x70 | n4603 ;
  assign n4854 = x70 &  n4603 ;
  assign n4855 = ( n4853 & ~n4854 ) | ( n4853 & 1'b0 ) | ( ~n4854 & 1'b0 ) ;
  assign n4864 = ( n4640 & n4665 ) | ( n4640 & n4855 ) | ( n4665 & n4855 ) ;
  assign n4865 = ( n4640 & ~n4668 ) | ( n4640 & n4855 ) | ( ~n4668 & n4855 ) ;
  assign n4866 = ~n4864 & n4865 ;
  assign n4867 = n4860 | n4866 ;
  assign n4868 = n4611 &  n4669 ;
  assign n4861 = x69 | n4611 ;
  assign n4862 = x69 &  n4611 ;
  assign n4863 = ( n4861 & ~n4862 ) | ( n4861 & 1'b0 ) | ( ~n4862 & 1'b0 ) ;
  assign n4872 = ( n4639 & n4665 ) | ( n4639 & n4863 ) | ( n4665 & n4863 ) ;
  assign n4873 = ( n4639 & ~n4668 ) | ( n4639 & n4863 ) | ( ~n4668 & n4863 ) ;
  assign n4874 = ~n4872 & n4873 ;
  assign n4875 = n4868 | n4874 ;
  assign n4876 = n4619 &  n4669 ;
  assign n4869 = x68 | n4619 ;
  assign n4870 = x68 &  n4619 ;
  assign n4871 = ( n4869 & ~n4870 ) | ( n4869 & 1'b0 ) | ( ~n4870 & 1'b0 ) ;
  assign n4880 = ( n4638 & n4665 ) | ( n4638 & n4871 ) | ( n4665 & n4871 ) ;
  assign n4881 = ( n4638 & ~n4668 ) | ( n4638 & n4871 ) | ( ~n4668 & n4871 ) ;
  assign n4882 = ~n4880 & n4881 ;
  assign n4883 = n4876 | n4882 ;
  assign n4884 = n4624 &  n4669 ;
  assign n4877 = x67 | n4624 ;
  assign n4878 = x67 &  n4624 ;
  assign n4879 = ( n4877 & ~n4878 ) | ( n4877 & 1'b0 ) | ( ~n4878 & 1'b0 ) ;
  assign n4888 = ( n4637 & n4665 ) | ( n4637 & n4879 ) | ( n4665 & n4879 ) ;
  assign n4889 = ( n4637 & ~n4668 ) | ( n4637 & n4879 ) | ( ~n4668 & n4879 ) ;
  assign n4890 = ~n4888 & n4889 ;
  assign n4891 = n4884 | n4890 ;
  assign n4892 = n4630 &  n4669 ;
  assign n4885 = x66 | n4630 ;
  assign n4886 = x66 &  n4630 ;
  assign n4887 = ( n4885 & ~n4886 ) | ( n4885 & 1'b0 ) | ( ~n4886 & 1'b0 ) ;
  assign n4897 = ( n4636 & ~n4665 ) | ( n4636 & n4887 ) | ( ~n4665 & n4887 ) ;
  assign n4898 = ( n4636 & n4668 ) | ( n4636 & n4887 ) | ( n4668 & n4887 ) ;
  assign n4899 = ( n4897 & ~n4898 ) | ( n4897 & 1'b0 ) | ( ~n4898 & 1'b0 ) ;
  assign n4900 = n4892 | n4899 ;
  assign n4901 = n4634 &  n4669 ;
  assign n4893 = x65 &  n4634 ;
  assign n4894 = ( n4632 & ~x65 ) | ( n4632 & n4633 ) | ( ~x65 & n4633 ) ;
  assign n4895 = x65 | n4894 ;
  assign n4896 = ( n4635 & ~n4893 ) | ( n4635 & n4895 ) | ( ~n4893 & n4895 ) ;
  assign n4902 = ( x65 & n4634 ) | ( x65 & n4635 ) | ( n4634 & n4635 ) ;
  assign n4903 = ( n4668 & ~n4893 ) | ( n4668 & n4902 ) | ( ~n4893 & n4902 ) ;
  assign n4904 = ( n4665 & n4896 ) | ( n4665 & n4903 ) | ( n4896 & n4903 ) ;
  assign n4905 = ( n4896 & ~n4904 ) | ( n4896 & 1'b0 ) | ( ~n4904 & 1'b0 ) ;
  assign n4906 = n4901 | n4905 ;
  assign n4907 = ( x64 & ~x95 ) | ( x64 & 1'b0 ) | ( ~x95 & 1'b0 ) ;
  assign n4908 = ( n175 & ~n185 ) | ( n175 & n4907 ) | ( ~n185 & n4907 ) ;
  assign n4909 = ~n175 & n4908 ;
  assign n4910 = ~n160 & n4909 ;
  assign n4911 = n4665 &  n4910 ;
  assign n4912 = ( x33 & ~n4910 ) | ( x33 & n4911 ) | ( ~n4910 & n4911 ) ;
  assign n4913 = ~n204 & n4635 ;
  assign n4914 = ( n246 & ~n428 ) | ( n246 & n4913 ) | ( ~n428 & n4913 ) ;
  assign n4915 = ~n246 & n4914 ;
  assign n4916 = ~n425 & n4915 ;
  assign n4917 = ~n4665 & n4916 ;
  assign n4918 = n4912 | n4917 ;
  assign n4919 = ~x32 & x64 ;
  assign n4920 = ( x65 & ~n4918 ) | ( x65 & n4919 ) | ( ~n4918 & n4919 ) ;
  assign n4921 = ( x66 & ~n4906 ) | ( x66 & n4920 ) | ( ~n4906 & n4920 ) ;
  assign n4922 = ( x67 & ~n4900 ) | ( x67 & n4921 ) | ( ~n4900 & n4921 ) ;
  assign n4923 = ( x68 & ~n4891 ) | ( x68 & n4922 ) | ( ~n4891 & n4922 ) ;
  assign n4924 = ( x69 & ~n4883 ) | ( x69 & n4923 ) | ( ~n4883 & n4923 ) ;
  assign n4925 = ( x70 & ~n4875 ) | ( x70 & n4924 ) | ( ~n4875 & n4924 ) ;
  assign n4926 = ( x71 & ~n4867 ) | ( x71 & n4925 ) | ( ~n4867 & n4925 ) ;
  assign n4927 = ( x72 & ~n4859 ) | ( x72 & n4926 ) | ( ~n4859 & n4926 ) ;
  assign n4928 = ( x73 & ~n4851 ) | ( x73 & n4927 ) | ( ~n4851 & n4927 ) ;
  assign n4929 = ( x74 & ~n4843 ) | ( x74 & n4928 ) | ( ~n4843 & n4928 ) ;
  assign n4930 = ( x75 & ~n4835 ) | ( x75 & n4929 ) | ( ~n4835 & n4929 ) ;
  assign n4931 = ( x76 & ~n4680 ) | ( x76 & n4930 ) | ( ~n4680 & n4930 ) ;
  assign n4932 = ( x77 & ~n4827 ) | ( x77 & n4931 ) | ( ~n4827 & n4931 ) ;
  assign n4933 = ( x78 & ~n4822 ) | ( x78 & n4932 ) | ( ~n4822 & n4932 ) ;
  assign n4934 = ( x79 & ~n4814 ) | ( x79 & n4933 ) | ( ~n4814 & n4933 ) ;
  assign n4935 = ( x80 & ~n4806 ) | ( x80 & n4934 ) | ( ~n4806 & n4934 ) ;
  assign n4936 = ( x81 & ~n4798 ) | ( x81 & n4935 ) | ( ~n4798 & n4935 ) ;
  assign n4937 = ( x82 & ~n4790 ) | ( x82 & n4936 ) | ( ~n4790 & n4936 ) ;
  assign n4938 = ( x83 & ~n4782 ) | ( x83 & n4937 ) | ( ~n4782 & n4937 ) ;
  assign n4939 = ( x84 & ~n4774 ) | ( x84 & n4938 ) | ( ~n4774 & n4938 ) ;
  assign n4940 = ( x85 & ~n4766 ) | ( x85 & n4939 ) | ( ~n4766 & n4939 ) ;
  assign n4941 = ( x86 & ~n4758 ) | ( x86 & n4940 ) | ( ~n4758 & n4940 ) ;
  assign n4942 = ( x87 & ~n4750 ) | ( x87 & n4941 ) | ( ~n4750 & n4941 ) ;
  assign n4943 = ( x88 & ~n4742 ) | ( x88 & n4942 ) | ( ~n4742 & n4942 ) ;
  assign n4944 = ( x89 & ~n4734 ) | ( x89 & n4943 ) | ( ~n4734 & n4943 ) ;
  assign n4945 = ( x90 & ~n4726 ) | ( x90 & n4944 ) | ( ~n4726 & n4944 ) ;
  assign n4946 = ( x91 & ~n4718 ) | ( x91 & n4945 ) | ( ~n4718 & n4945 ) ;
  assign n4947 = ( x92 & ~n4710 ) | ( x92 & n4946 ) | ( ~n4710 & n4946 ) ;
  assign n4948 = ( x93 & ~n4702 ) | ( x93 & n4947 ) | ( ~n4702 & n4947 ) ;
  assign n4949 = ( x94 & ~n4694 ) | ( x94 & n4948 ) | ( ~n4694 & n4948 ) ;
  assign n4950 = ( x95 & ~n4686 ) | ( x95 & n4949 ) | ( ~n4686 & n4949 ) ;
  assign n4951 = n274 | n4950 ;
  assign n5088 = n4694 &  n4951 ;
  assign n5092 = x94 | n4694 ;
  assign n5093 = x94 &  n4694 ;
  assign n5094 = ( n5092 & ~n5093 ) | ( n5092 & 1'b0 ) | ( ~n5093 & 1'b0 ) ;
  assign n5095 = ( n274 & n4948 ) | ( n274 & n5094 ) | ( n4948 & n5094 ) ;
  assign n5096 = ( n4948 & ~n4950 ) | ( n4948 & n5094 ) | ( ~n4950 & n5094 ) ;
  assign n5097 = ~n5095 & n5096 ;
  assign n5098 = n5088 | n5097 ;
  assign n5099 = n4702 &  n4951 ;
  assign n5089 = x93 | n4702 ;
  assign n5090 = x93 &  n4702 ;
  assign n5091 = ( n5089 & ~n5090 ) | ( n5089 & 1'b0 ) | ( ~n5090 & 1'b0 ) ;
  assign n5103 = ( n274 & n4947 ) | ( n274 & n5091 ) | ( n4947 & n5091 ) ;
  assign n5104 = ( n4947 & ~n4950 ) | ( n4947 & n5091 ) | ( ~n4950 & n5091 ) ;
  assign n5105 = ~n5103 & n5104 ;
  assign n5106 = n5099 | n5105 ;
  assign n5107 = n4710 &  n4951 ;
  assign n5100 = x92 | n4710 ;
  assign n5101 = x92 &  n4710 ;
  assign n5102 = ( n5100 & ~n5101 ) | ( n5100 & 1'b0 ) | ( ~n5101 & 1'b0 ) ;
  assign n5111 = ( n274 & n4946 ) | ( n274 & n5102 ) | ( n4946 & n5102 ) ;
  assign n5112 = ( n4946 & ~n4950 ) | ( n4946 & n5102 ) | ( ~n4950 & n5102 ) ;
  assign n5113 = ~n5111 & n5112 ;
  assign n5114 = n5107 | n5113 ;
  assign n5115 = n4718 &  n4951 ;
  assign n5108 = x91 | n4718 ;
  assign n5109 = x91 &  n4718 ;
  assign n5110 = ( n5108 & ~n5109 ) | ( n5108 & 1'b0 ) | ( ~n5109 & 1'b0 ) ;
  assign n5119 = ( n274 & n4945 ) | ( n274 & n5110 ) | ( n4945 & n5110 ) ;
  assign n5120 = ( n4945 & ~n4950 ) | ( n4945 & n5110 ) | ( ~n4950 & n5110 ) ;
  assign n5121 = ~n5119 & n5120 ;
  assign n5122 = n5115 | n5121 ;
  assign n5123 = n4726 &  n4951 ;
  assign n5116 = x90 | n4726 ;
  assign n5117 = x90 &  n4726 ;
  assign n5118 = ( n5116 & ~n5117 ) | ( n5116 & 1'b0 ) | ( ~n5117 & 1'b0 ) ;
  assign n5127 = ( n274 & n4944 ) | ( n274 & n5118 ) | ( n4944 & n5118 ) ;
  assign n5128 = ( n4944 & ~n4950 ) | ( n4944 & n5118 ) | ( ~n4950 & n5118 ) ;
  assign n5129 = ~n5127 & n5128 ;
  assign n5130 = n5123 | n5129 ;
  assign n5131 = n4734 &  n4951 ;
  assign n5124 = x89 | n4734 ;
  assign n5125 = x89 &  n4734 ;
  assign n5126 = ( n5124 & ~n5125 ) | ( n5124 & 1'b0 ) | ( ~n5125 & 1'b0 ) ;
  assign n5135 = ( n274 & n4943 ) | ( n274 & n5126 ) | ( n4943 & n5126 ) ;
  assign n5136 = ( n4943 & ~n4950 ) | ( n4943 & n5126 ) | ( ~n4950 & n5126 ) ;
  assign n5137 = ~n5135 & n5136 ;
  assign n5138 = n5131 | n5137 ;
  assign n5139 = n4742 &  n4951 ;
  assign n5132 = x88 | n4742 ;
  assign n5133 = x88 &  n4742 ;
  assign n5134 = ( n5132 & ~n5133 ) | ( n5132 & 1'b0 ) | ( ~n5133 & 1'b0 ) ;
  assign n5143 = ( n274 & n4942 ) | ( n274 & n5134 ) | ( n4942 & n5134 ) ;
  assign n5144 = ( n4942 & ~n4950 ) | ( n4942 & n5134 ) | ( ~n4950 & n5134 ) ;
  assign n5145 = ~n5143 & n5144 ;
  assign n5146 = n5139 | n5145 ;
  assign n5147 = n4750 &  n4951 ;
  assign n5140 = x87 | n4750 ;
  assign n5141 = x87 &  n4750 ;
  assign n5142 = ( n5140 & ~n5141 ) | ( n5140 & 1'b0 ) | ( ~n5141 & 1'b0 ) ;
  assign n5151 = ( n274 & n4941 ) | ( n274 & n5142 ) | ( n4941 & n5142 ) ;
  assign n5152 = ( n4941 & ~n4950 ) | ( n4941 & n5142 ) | ( ~n4950 & n5142 ) ;
  assign n5153 = ~n5151 & n5152 ;
  assign n5154 = n5147 | n5153 ;
  assign n5155 = n4758 &  n4951 ;
  assign n5148 = x86 | n4758 ;
  assign n5149 = x86 &  n4758 ;
  assign n5150 = ( n5148 & ~n5149 ) | ( n5148 & 1'b0 ) | ( ~n5149 & 1'b0 ) ;
  assign n5159 = ( n274 & n4940 ) | ( n274 & n5150 ) | ( n4940 & n5150 ) ;
  assign n5160 = ( n4940 & ~n4950 ) | ( n4940 & n5150 ) | ( ~n4950 & n5150 ) ;
  assign n5161 = ~n5159 & n5160 ;
  assign n5162 = n5155 | n5161 ;
  assign n5163 = n4766 &  n4951 ;
  assign n5156 = x85 | n4766 ;
  assign n5157 = x85 &  n4766 ;
  assign n5158 = ( n5156 & ~n5157 ) | ( n5156 & 1'b0 ) | ( ~n5157 & 1'b0 ) ;
  assign n5167 = ( n274 & n4939 ) | ( n274 & n5158 ) | ( n4939 & n5158 ) ;
  assign n5168 = ( n4939 & ~n4950 ) | ( n4939 & n5158 ) | ( ~n4950 & n5158 ) ;
  assign n5169 = ~n5167 & n5168 ;
  assign n5170 = n5163 | n5169 ;
  assign n5171 = n4774 &  n4951 ;
  assign n5164 = x84 | n4774 ;
  assign n5165 = x84 &  n4774 ;
  assign n5166 = ( n5164 & ~n5165 ) | ( n5164 & 1'b0 ) | ( ~n5165 & 1'b0 ) ;
  assign n5175 = ( n274 & n4938 ) | ( n274 & n5166 ) | ( n4938 & n5166 ) ;
  assign n5176 = ( n4938 & ~n4950 ) | ( n4938 & n5166 ) | ( ~n4950 & n5166 ) ;
  assign n5177 = ~n5175 & n5176 ;
  assign n5178 = n5171 | n5177 ;
  assign n5179 = n4782 &  n4951 ;
  assign n5172 = x83 | n4782 ;
  assign n5173 = x83 &  n4782 ;
  assign n5174 = ( n5172 & ~n5173 ) | ( n5172 & 1'b0 ) | ( ~n5173 & 1'b0 ) ;
  assign n5183 = ( n274 & n4937 ) | ( n274 & n5174 ) | ( n4937 & n5174 ) ;
  assign n5184 = ( n4937 & ~n4950 ) | ( n4937 & n5174 ) | ( ~n4950 & n5174 ) ;
  assign n5185 = ~n5183 & n5184 ;
  assign n5186 = n5179 | n5185 ;
  assign n5187 = n4790 &  n4951 ;
  assign n5180 = x82 | n4790 ;
  assign n5181 = x82 &  n4790 ;
  assign n5182 = ( n5180 & ~n5181 ) | ( n5180 & 1'b0 ) | ( ~n5181 & 1'b0 ) ;
  assign n5191 = ( n274 & n4936 ) | ( n274 & n5182 ) | ( n4936 & n5182 ) ;
  assign n5192 = ( n4936 & ~n4950 ) | ( n4936 & n5182 ) | ( ~n4950 & n5182 ) ;
  assign n5193 = ~n5191 & n5192 ;
  assign n5194 = n5187 | n5193 ;
  assign n5195 = n4798 &  n4951 ;
  assign n5188 = x81 | n4798 ;
  assign n5189 = x81 &  n4798 ;
  assign n5190 = ( n5188 & ~n5189 ) | ( n5188 & 1'b0 ) | ( ~n5189 & 1'b0 ) ;
  assign n5199 = ( n274 & n4935 ) | ( n274 & n5190 ) | ( n4935 & n5190 ) ;
  assign n5200 = ( n4935 & ~n4950 ) | ( n4935 & n5190 ) | ( ~n4950 & n5190 ) ;
  assign n5201 = ~n5199 & n5200 ;
  assign n5202 = n5195 | n5201 ;
  assign n5203 = n4806 &  n4951 ;
  assign n5196 = x80 | n4806 ;
  assign n5197 = x80 &  n4806 ;
  assign n5198 = ( n5196 & ~n5197 ) | ( n5196 & 1'b0 ) | ( ~n5197 & 1'b0 ) ;
  assign n5207 = ( n274 & n4934 ) | ( n274 & n5198 ) | ( n4934 & n5198 ) ;
  assign n5208 = ( n4934 & ~n4950 ) | ( n4934 & n5198 ) | ( ~n4950 & n5198 ) ;
  assign n5209 = ~n5207 & n5208 ;
  assign n5210 = n5203 | n5209 ;
  assign n5211 = n4814 &  n4951 ;
  assign n5204 = x79 | n4814 ;
  assign n5205 = x79 &  n4814 ;
  assign n5206 = ( n5204 & ~n5205 ) | ( n5204 & 1'b0 ) | ( ~n5205 & 1'b0 ) ;
  assign n5215 = ( n274 & n4933 ) | ( n274 & n5206 ) | ( n4933 & n5206 ) ;
  assign n5216 = ( n4933 & ~n4950 ) | ( n4933 & n5206 ) | ( ~n4950 & n5206 ) ;
  assign n5217 = ~n5215 & n5216 ;
  assign n5218 = n5211 | n5217 ;
  assign n5219 = n4822 &  n4951 ;
  assign n5212 = x78 | n4822 ;
  assign n5213 = x78 &  n4822 ;
  assign n5214 = ( n5212 & ~n5213 ) | ( n5212 & 1'b0 ) | ( ~n5213 & 1'b0 ) ;
  assign n5220 = ( n274 & n4932 ) | ( n274 & n5214 ) | ( n4932 & n5214 ) ;
  assign n5221 = ( n4932 & ~n4950 ) | ( n4932 & n5214 ) | ( ~n4950 & n5214 ) ;
  assign n5222 = ~n5220 & n5221 ;
  assign n5223 = n5219 | n5222 ;
  assign n5077 = n4827 &  n4951 ;
  assign n5078 = x77 | n4827 ;
  assign n5079 = x77 &  n4827 ;
  assign n5080 = ( n5078 & ~n5079 ) | ( n5078 & 1'b0 ) | ( ~n5079 & 1'b0 ) ;
  assign n5081 = ( n274 & n4931 ) | ( n274 & n5080 ) | ( n4931 & n5080 ) ;
  assign n5082 = ( n4931 & ~n4950 ) | ( n4931 & n5080 ) | ( ~n4950 & n5080 ) ;
  assign n5083 = ~n5081 & n5082 ;
  assign n5084 = n5077 | n5083 ;
  assign n4952 = n4680 &  n4951 ;
  assign n4956 = x76 | n4680 ;
  assign n4957 = x76 &  n4680 ;
  assign n4958 = ( n4956 & ~n4957 ) | ( n4956 & 1'b0 ) | ( ~n4957 & 1'b0 ) ;
  assign n4959 = ( n274 & n4930 ) | ( n274 & n4958 ) | ( n4930 & n4958 ) ;
  assign n4960 = ( n4930 & ~n4950 ) | ( n4930 & n4958 ) | ( ~n4950 & n4958 ) ;
  assign n4961 = ~n4959 & n4960 ;
  assign n4962 = n4952 | n4961 ;
  assign n4963 = n4835 &  n4951 ;
  assign n4953 = x75 | n4835 ;
  assign n4954 = x75 &  n4835 ;
  assign n4955 = ( n4953 & ~n4954 ) | ( n4953 & 1'b0 ) | ( ~n4954 & 1'b0 ) ;
  assign n4967 = ( n274 & n4929 ) | ( n274 & n4955 ) | ( n4929 & n4955 ) ;
  assign n4968 = ( n4929 & ~n4950 ) | ( n4929 & n4955 ) | ( ~n4950 & n4955 ) ;
  assign n4969 = ~n4967 & n4968 ;
  assign n4970 = n4963 | n4969 ;
  assign n4971 = n4843 &  n4951 ;
  assign n4964 = x74 | n4843 ;
  assign n4965 = x74 &  n4843 ;
  assign n4966 = ( n4964 & ~n4965 ) | ( n4964 & 1'b0 ) | ( ~n4965 & 1'b0 ) ;
  assign n4975 = ( n274 & n4928 ) | ( n274 & n4966 ) | ( n4928 & n4966 ) ;
  assign n4976 = ( n4928 & ~n4950 ) | ( n4928 & n4966 ) | ( ~n4950 & n4966 ) ;
  assign n4977 = ~n4975 & n4976 ;
  assign n4978 = n4971 | n4977 ;
  assign n4979 = n4851 &  n4951 ;
  assign n4972 = x73 | n4851 ;
  assign n4973 = x73 &  n4851 ;
  assign n4974 = ( n4972 & ~n4973 ) | ( n4972 & 1'b0 ) | ( ~n4973 & 1'b0 ) ;
  assign n4983 = ( n274 & n4927 ) | ( n274 & n4974 ) | ( n4927 & n4974 ) ;
  assign n4984 = ( n4927 & ~n4950 ) | ( n4927 & n4974 ) | ( ~n4950 & n4974 ) ;
  assign n4985 = ~n4983 & n4984 ;
  assign n4986 = n4979 | n4985 ;
  assign n4987 = n4859 &  n4951 ;
  assign n4980 = x72 | n4859 ;
  assign n4981 = x72 &  n4859 ;
  assign n4982 = ( n4980 & ~n4981 ) | ( n4980 & 1'b0 ) | ( ~n4981 & 1'b0 ) ;
  assign n4991 = ( n274 & n4926 ) | ( n274 & n4982 ) | ( n4926 & n4982 ) ;
  assign n4992 = ( n4926 & ~n4950 ) | ( n4926 & n4982 ) | ( ~n4950 & n4982 ) ;
  assign n4993 = ~n4991 & n4992 ;
  assign n4994 = n4987 | n4993 ;
  assign n4995 = n4867 &  n4951 ;
  assign n4988 = x71 | n4867 ;
  assign n4989 = x71 &  n4867 ;
  assign n4990 = ( n4988 & ~n4989 ) | ( n4988 & 1'b0 ) | ( ~n4989 & 1'b0 ) ;
  assign n4999 = ( n274 & n4925 ) | ( n274 & n4990 ) | ( n4925 & n4990 ) ;
  assign n5000 = ( n4925 & ~n4950 ) | ( n4925 & n4990 ) | ( ~n4950 & n4990 ) ;
  assign n5001 = ~n4999 & n5000 ;
  assign n5002 = n4995 | n5001 ;
  assign n5003 = n4875 &  n4951 ;
  assign n4996 = x70 | n4875 ;
  assign n4997 = x70 &  n4875 ;
  assign n4998 = ( n4996 & ~n4997 ) | ( n4996 & 1'b0 ) | ( ~n4997 & 1'b0 ) ;
  assign n5007 = ( n274 & n4924 ) | ( n274 & n4998 ) | ( n4924 & n4998 ) ;
  assign n5008 = ( n4924 & ~n4950 ) | ( n4924 & n4998 ) | ( ~n4950 & n4998 ) ;
  assign n5009 = ~n5007 & n5008 ;
  assign n5010 = n5003 | n5009 ;
  assign n5011 = n4883 &  n4951 ;
  assign n5004 = x69 | n4883 ;
  assign n5005 = x69 &  n4883 ;
  assign n5006 = ( n5004 & ~n5005 ) | ( n5004 & 1'b0 ) | ( ~n5005 & 1'b0 ) ;
  assign n5015 = ( n274 & n4923 ) | ( n274 & n5006 ) | ( n4923 & n5006 ) ;
  assign n5016 = ( n4923 & ~n4950 ) | ( n4923 & n5006 ) | ( ~n4950 & n5006 ) ;
  assign n5017 = ~n5015 & n5016 ;
  assign n5018 = n5011 | n5017 ;
  assign n5019 = n4891 &  n4951 ;
  assign n5012 = x68 | n4891 ;
  assign n5013 = x68 &  n4891 ;
  assign n5014 = ( n5012 & ~n5013 ) | ( n5012 & 1'b0 ) | ( ~n5013 & 1'b0 ) ;
  assign n5023 = ( n274 & n4922 ) | ( n274 & n5014 ) | ( n4922 & n5014 ) ;
  assign n5024 = ( n4922 & ~n4950 ) | ( n4922 & n5014 ) | ( ~n4950 & n5014 ) ;
  assign n5025 = ~n5023 & n5024 ;
  assign n5026 = n5019 | n5025 ;
  assign n5027 = n4900 &  n4951 ;
  assign n5020 = x67 | n4900 ;
  assign n5021 = x67 &  n4900 ;
  assign n5022 = ( n5020 & ~n5021 ) | ( n5020 & 1'b0 ) | ( ~n5021 & 1'b0 ) ;
  assign n5031 = ( n274 & n4921 ) | ( n274 & n5022 ) | ( n4921 & n5022 ) ;
  assign n5032 = ( n4921 & ~n4950 ) | ( n4921 & n5022 ) | ( ~n4950 & n5022 ) ;
  assign n5033 = ~n5031 & n5032 ;
  assign n5034 = n5027 | n5033 ;
  assign n5035 = n4906 &  n4951 ;
  assign n5028 = x66 | n4906 ;
  assign n5029 = x66 &  n4906 ;
  assign n5030 = ( n5028 & ~n5029 ) | ( n5028 & 1'b0 ) | ( ~n5029 & 1'b0 ) ;
  assign n5039 = ( n4920 & ~n274 ) | ( n4920 & n5030 ) | ( ~n274 & n5030 ) ;
  assign n5040 = ( n4920 & n4950 ) | ( n4920 & n5030 ) | ( n4950 & n5030 ) ;
  assign n5041 = ( n5039 & ~n5040 ) | ( n5039 & 1'b0 ) | ( ~n5040 & 1'b0 ) ;
  assign n5042 = n5035 | n5041 ;
  assign n5043 = n4918 &  n4951 ;
  assign n5036 = x65 &  n4918 ;
  assign n5037 = x65 | n4917 ;
  assign n5038 = n4912 | n5037 ;
  assign n5044 = ~n5036 & n5038 ;
  assign n5045 = ( n4919 & ~n4950 ) | ( n4919 & n5044 ) | ( ~n4950 & n5044 ) ;
  assign n5046 = ( n274 & n4919 ) | ( n274 & n5044 ) | ( n4919 & n5044 ) ;
  assign n5047 = ( n5045 & ~n5046 ) | ( n5045 & 1'b0 ) | ( ~n5046 & 1'b0 ) ;
  assign n5048 = n5043 | n5047 ;
  assign n5049 = ( x64 & ~x96 ) | ( x64 & 1'b0 ) | ( ~x96 & 1'b0 ) ;
  assign n5050 = ( n246 & ~n428 ) | ( n246 & n5049 ) | ( ~n428 & n5049 ) ;
  assign n5051 = ~n246 & n5050 ;
  assign n5052 = ~n425 & n5051 ;
  assign n5053 = n4950 &  n5052 ;
  assign n5054 = ( x32 & ~n5052 ) | ( x32 & n5053 ) | ( ~n5052 & n5053 ) ;
  assign n5055 = ~n185 & n4919 ;
  assign n5056 = ( n160 & ~n175 ) | ( n160 & n5055 ) | ( ~n175 & n5055 ) ;
  assign n5057 = ~n160 & n5056 ;
  assign n5058 = ~n4950 & n5057 ;
  assign n5059 = n5054 | n5058 ;
  assign n5060 = ~x31 & x64 ;
  assign n5061 = ( x65 & ~n5059 ) | ( x65 & n5060 ) | ( ~n5059 & n5060 ) ;
  assign n5062 = ( x66 & ~n5048 ) | ( x66 & n5061 ) | ( ~n5048 & n5061 ) ;
  assign n5063 = ( x67 & ~n5042 ) | ( x67 & n5062 ) | ( ~n5042 & n5062 ) ;
  assign n5064 = ( x68 & ~n5034 ) | ( x68 & n5063 ) | ( ~n5034 & n5063 ) ;
  assign n5065 = ( x69 & ~n5026 ) | ( x69 & n5064 ) | ( ~n5026 & n5064 ) ;
  assign n5066 = ( x70 & ~n5018 ) | ( x70 & n5065 ) | ( ~n5018 & n5065 ) ;
  assign n5067 = ( x71 & ~n5010 ) | ( x71 & n5066 ) | ( ~n5010 & n5066 ) ;
  assign n5068 = ( x72 & ~n5002 ) | ( x72 & n5067 ) | ( ~n5002 & n5067 ) ;
  assign n5069 = ( x73 & ~n4994 ) | ( x73 & n5068 ) | ( ~n4994 & n5068 ) ;
  assign n5070 = ( x74 & ~n4986 ) | ( x74 & n5069 ) | ( ~n4986 & n5069 ) ;
  assign n5071 = ( x75 & ~n4978 ) | ( x75 & n5070 ) | ( ~n4978 & n5070 ) ;
  assign n5072 = ( x76 & ~n4970 ) | ( x76 & n5071 ) | ( ~n4970 & n5071 ) ;
  assign n5076 = ( x77 & ~n4962 ) | ( x77 & n5072 ) | ( ~n4962 & n5072 ) ;
  assign n5224 = ( x78 & ~n5084 ) | ( x78 & n5076 ) | ( ~n5084 & n5076 ) ;
  assign n5225 = ( x79 & ~n5223 ) | ( x79 & n5224 ) | ( ~n5223 & n5224 ) ;
  assign n5226 = ( x80 & ~n5218 ) | ( x80 & n5225 ) | ( ~n5218 & n5225 ) ;
  assign n5227 = ( x81 & ~n5210 ) | ( x81 & n5226 ) | ( ~n5210 & n5226 ) ;
  assign n5228 = ( x82 & ~n5202 ) | ( x82 & n5227 ) | ( ~n5202 & n5227 ) ;
  assign n5229 = ( x83 & ~n5194 ) | ( x83 & n5228 ) | ( ~n5194 & n5228 ) ;
  assign n5230 = ( x84 & ~n5186 ) | ( x84 & n5229 ) | ( ~n5186 & n5229 ) ;
  assign n5231 = ( x85 & ~n5178 ) | ( x85 & n5230 ) | ( ~n5178 & n5230 ) ;
  assign n5232 = ( x86 & ~n5170 ) | ( x86 & n5231 ) | ( ~n5170 & n5231 ) ;
  assign n5233 = ( x87 & ~n5162 ) | ( x87 & n5232 ) | ( ~n5162 & n5232 ) ;
  assign n5234 = ( x88 & ~n5154 ) | ( x88 & n5233 ) | ( ~n5154 & n5233 ) ;
  assign n5235 = ( x89 & ~n5146 ) | ( x89 & n5234 ) | ( ~n5146 & n5234 ) ;
  assign n5236 = ( x90 & ~n5138 ) | ( x90 & n5235 ) | ( ~n5138 & n5235 ) ;
  assign n5237 = ( x91 & ~n5130 ) | ( x91 & n5236 ) | ( ~n5130 & n5236 ) ;
  assign n5238 = ( x92 & ~n5122 ) | ( x92 & n5237 ) | ( ~n5122 & n5237 ) ;
  assign n5239 = ( x93 & ~n5114 ) | ( x93 & n5238 ) | ( ~n5114 & n5238 ) ;
  assign n5240 = ( x94 & ~n5106 ) | ( x94 & n5239 ) | ( ~n5106 & n5239 ) ;
  assign n5241 = ( x95 & ~n5098 ) | ( x95 & n5240 ) | ( ~n5098 & n5240 ) ;
  assign n5242 = n4686 &  n4951 ;
  assign n5243 = ( n274 & n4686 ) | ( n274 & n4949 ) | ( n4686 & n4949 ) ;
  assign n5244 = ( x95 & ~n5243 ) | ( x95 & n4686 ) | ( ~n5243 & n4686 ) ;
  assign n5245 = ~x95 & n5244 ;
  assign n5246 = n5242 | n5245 ;
  assign n5247 = ~x96 & n5246 ;
  assign n5248 = ( x96 & ~n5242 ) | ( x96 & 1'b0 ) | ( ~n5242 & 1'b0 ) ;
  assign n5249 = ~n5245 & n5248 ;
  assign n5250 = n256 | n5249 ;
  assign n5251 = n5247 | n5250 ;
  assign n5252 = n5241 | n5251 ;
  assign n5253 = ~n5246 |  n274 ;
  assign n5272 = n5098 &  n5253 ;
  assign n5273 = n5252 &  n5272 ;
  assign n5260 = x95 | n5098 ;
  assign n5261 = x95 &  n5098 ;
  assign n5262 = ( n5260 & ~n5261 ) | ( n5260 & 1'b0 ) | ( ~n5261 & 1'b0 ) ;
  assign n5274 = n5240 &  n5262 ;
  assign n5254 = n5252 &  n5253 ;
  assign n5275 = ( n5240 & ~n5254 ) | ( n5240 & n5262 ) | ( ~n5254 & n5262 ) ;
  assign n5276 = ( n5273 & ~n5274 ) | ( n5273 & n5275 ) | ( ~n5274 & n5275 ) ;
  assign n5264 = n274 &  n4686 ;
  assign n5265 = n5252 &  n5264 ;
  assign n5263 = n5247 | n5249 ;
  assign n5267 = ( n5241 & n5254 ) | ( n5241 & n5263 ) | ( n5254 & n5263 ) ;
  assign n5266 = n5241 | n5263 ;
  assign n5268 = ( n5265 & ~n5267 ) | ( n5265 & n5266 ) | ( ~n5267 & n5266 ) ;
  assign n5280 = n5106 &  n5253 ;
  assign n5281 = n5252 &  n5280 ;
  assign n5269 = x94 | n5106 ;
  assign n5270 = x94 &  n5106 ;
  assign n5271 = ( n5269 & ~n5270 ) | ( n5269 & 1'b0 ) | ( ~n5270 & 1'b0 ) ;
  assign n5282 = n5239 &  n5271 ;
  assign n5283 = ( n5239 & ~n5254 ) | ( n5239 & n5271 ) | ( ~n5254 & n5271 ) ;
  assign n5284 = ( n5281 & ~n5282 ) | ( n5281 & n5283 ) | ( ~n5282 & n5283 ) ;
  assign n5288 = n5114 &  n5253 ;
  assign n5289 = n5252 &  n5288 ;
  assign n5277 = x93 | n5114 ;
  assign n5278 = x93 &  n5114 ;
  assign n5279 = ( n5277 & ~n5278 ) | ( n5277 & 1'b0 ) | ( ~n5278 & 1'b0 ) ;
  assign n5290 = n5238 &  n5279 ;
  assign n5291 = ( n5238 & ~n5254 ) | ( n5238 & n5279 ) | ( ~n5254 & n5279 ) ;
  assign n5292 = ( n5289 & ~n5290 ) | ( n5289 & n5291 ) | ( ~n5290 & n5291 ) ;
  assign n5296 = n5122 &  n5253 ;
  assign n5297 = n5252 &  n5296 ;
  assign n5285 = x92 | n5122 ;
  assign n5286 = x92 &  n5122 ;
  assign n5287 = ( n5285 & ~n5286 ) | ( n5285 & 1'b0 ) | ( ~n5286 & 1'b0 ) ;
  assign n5298 = n5237 &  n5287 ;
  assign n5299 = ( n5237 & ~n5254 ) | ( n5237 & n5287 ) | ( ~n5254 & n5287 ) ;
  assign n5300 = ( n5297 & ~n5298 ) | ( n5297 & n5299 ) | ( ~n5298 & n5299 ) ;
  assign n5304 = n5130 &  n5253 ;
  assign n5305 = n5252 &  n5304 ;
  assign n5293 = x91 | n5130 ;
  assign n5294 = x91 &  n5130 ;
  assign n5295 = ( n5293 & ~n5294 ) | ( n5293 & 1'b0 ) | ( ~n5294 & 1'b0 ) ;
  assign n5306 = n5236 &  n5295 ;
  assign n5307 = ( n5236 & ~n5254 ) | ( n5236 & n5295 ) | ( ~n5254 & n5295 ) ;
  assign n5308 = ( n5305 & ~n5306 ) | ( n5305 & n5307 ) | ( ~n5306 & n5307 ) ;
  assign n5312 = n5138 &  n5253 ;
  assign n5313 = n5252 &  n5312 ;
  assign n5301 = x90 | n5138 ;
  assign n5302 = x90 &  n5138 ;
  assign n5303 = ( n5301 & ~n5302 ) | ( n5301 & 1'b0 ) | ( ~n5302 & 1'b0 ) ;
  assign n5315 = ( n5235 & n5254 ) | ( n5235 & n5303 ) | ( n5254 & n5303 ) ;
  assign n5314 = n5235 | n5303 ;
  assign n5316 = ( n5313 & ~n5315 ) | ( n5313 & n5314 ) | ( ~n5315 & n5314 ) ;
  assign n5320 = n5146 &  n5253 ;
  assign n5321 = n5252 &  n5320 ;
  assign n5309 = x89 | n5146 ;
  assign n5310 = x89 &  n5146 ;
  assign n5311 = ( n5309 & ~n5310 ) | ( n5309 & 1'b0 ) | ( ~n5310 & 1'b0 ) ;
  assign n5323 = ( n5234 & n5254 ) | ( n5234 & n5311 ) | ( n5254 & n5311 ) ;
  assign n5322 = n5234 | n5311 ;
  assign n5324 = ( n5321 & ~n5323 ) | ( n5321 & n5322 ) | ( ~n5323 & n5322 ) ;
  assign n5328 = n5154 &  n5253 ;
  assign n5329 = n5252 &  n5328 ;
  assign n5317 = x88 | n5154 ;
  assign n5318 = x88 &  n5154 ;
  assign n5319 = ( n5317 & ~n5318 ) | ( n5317 & 1'b0 ) | ( ~n5318 & 1'b0 ) ;
  assign n5331 = ( n5233 & n5254 ) | ( n5233 & n5319 ) | ( n5254 & n5319 ) ;
  assign n5330 = n5233 | n5319 ;
  assign n5332 = ( n5329 & ~n5331 ) | ( n5329 & n5330 ) | ( ~n5331 & n5330 ) ;
  assign n5336 = n5162 &  n5253 ;
  assign n5337 = n5252 &  n5336 ;
  assign n5325 = x87 | n5162 ;
  assign n5326 = x87 &  n5162 ;
  assign n5327 = ( n5325 & ~n5326 ) | ( n5325 & 1'b0 ) | ( ~n5326 & 1'b0 ) ;
  assign n5339 = ( n5232 & n5254 ) | ( n5232 & n5327 ) | ( n5254 & n5327 ) ;
  assign n5338 = n5232 | n5327 ;
  assign n5340 = ( n5337 & ~n5339 ) | ( n5337 & n5338 ) | ( ~n5339 & n5338 ) ;
  assign n5344 = n5170 &  n5253 ;
  assign n5345 = n5252 &  n5344 ;
  assign n5333 = x86 | n5170 ;
  assign n5334 = x86 &  n5170 ;
  assign n5335 = ( n5333 & ~n5334 ) | ( n5333 & 1'b0 ) | ( ~n5334 & 1'b0 ) ;
  assign n5347 = ( n5231 & n5254 ) | ( n5231 & n5335 ) | ( n5254 & n5335 ) ;
  assign n5346 = n5231 | n5335 ;
  assign n5348 = ( n5345 & ~n5347 ) | ( n5345 & n5346 ) | ( ~n5347 & n5346 ) ;
  assign n5352 = n5178 &  n5253 ;
  assign n5353 = n5252 &  n5352 ;
  assign n5341 = x85 | n5178 ;
  assign n5342 = x85 &  n5178 ;
  assign n5343 = ( n5341 & ~n5342 ) | ( n5341 & 1'b0 ) | ( ~n5342 & 1'b0 ) ;
  assign n5355 = ( n5230 & n5254 ) | ( n5230 & n5343 ) | ( n5254 & n5343 ) ;
  assign n5354 = n5230 | n5343 ;
  assign n5356 = ( n5353 & ~n5355 ) | ( n5353 & n5354 ) | ( ~n5355 & n5354 ) ;
  assign n5360 = n5186 &  n5253 ;
  assign n5361 = n5252 &  n5360 ;
  assign n5349 = x84 | n5186 ;
  assign n5350 = x84 &  n5186 ;
  assign n5351 = ( n5349 & ~n5350 ) | ( n5349 & 1'b0 ) | ( ~n5350 & 1'b0 ) ;
  assign n5363 = ( n5229 & n5254 ) | ( n5229 & n5351 ) | ( n5254 & n5351 ) ;
  assign n5362 = n5229 | n5351 ;
  assign n5364 = ( n5361 & ~n5363 ) | ( n5361 & n5362 ) | ( ~n5363 & n5362 ) ;
  assign n5368 = n5194 &  n5253 ;
  assign n5369 = n5252 &  n5368 ;
  assign n5357 = x83 | n5194 ;
  assign n5358 = x83 &  n5194 ;
  assign n5359 = ( n5357 & ~n5358 ) | ( n5357 & 1'b0 ) | ( ~n5358 & 1'b0 ) ;
  assign n5371 = ( n5228 & n5254 ) | ( n5228 & n5359 ) | ( n5254 & n5359 ) ;
  assign n5370 = n5228 | n5359 ;
  assign n5372 = ( n5369 & ~n5371 ) | ( n5369 & n5370 ) | ( ~n5371 & n5370 ) ;
  assign n5376 = n5202 &  n5253 ;
  assign n5377 = n5252 &  n5376 ;
  assign n5365 = x82 | n5202 ;
  assign n5366 = x82 &  n5202 ;
  assign n5367 = ( n5365 & ~n5366 ) | ( n5365 & 1'b0 ) | ( ~n5366 & 1'b0 ) ;
  assign n5379 = ( n5227 & n5254 ) | ( n5227 & n5367 ) | ( n5254 & n5367 ) ;
  assign n5378 = n5227 | n5367 ;
  assign n5380 = ( n5377 & ~n5379 ) | ( n5377 & n5378 ) | ( ~n5379 & n5378 ) ;
  assign n5384 = n5210 &  n5253 ;
  assign n5385 = n5252 &  n5384 ;
  assign n5373 = x81 | n5210 ;
  assign n5374 = x81 &  n5210 ;
  assign n5375 = ( n5373 & ~n5374 ) | ( n5373 & 1'b0 ) | ( ~n5374 & 1'b0 ) ;
  assign n5387 = ( n5226 & n5254 ) | ( n5226 & n5375 ) | ( n5254 & n5375 ) ;
  assign n5386 = n5226 | n5375 ;
  assign n5388 = ( n5385 & ~n5387 ) | ( n5385 & n5386 ) | ( ~n5387 & n5386 ) ;
  assign n5392 = n5218 &  n5253 ;
  assign n5393 = n5252 &  n5392 ;
  assign n5381 = x80 | n5218 ;
  assign n5382 = x80 &  n5218 ;
  assign n5383 = ( n5381 & ~n5382 ) | ( n5381 & 1'b0 ) | ( ~n5382 & 1'b0 ) ;
  assign n5395 = ( n5225 & n5254 ) | ( n5225 & n5383 ) | ( n5254 & n5383 ) ;
  assign n5394 = n5225 | n5383 ;
  assign n5396 = ( n5393 & ~n5395 ) | ( n5393 & n5394 ) | ( ~n5395 & n5394 ) ;
  assign n5397 = n5223 &  n5253 ;
  assign n5398 = n5252 &  n5397 ;
  assign n5389 = x79 | n5223 ;
  assign n5390 = x79 &  n5223 ;
  assign n5391 = ( n5389 & ~n5390 ) | ( n5389 & 1'b0 ) | ( ~n5390 & 1'b0 ) ;
  assign n5400 = ( n5224 & n5254 ) | ( n5224 & n5391 ) | ( n5254 & n5391 ) ;
  assign n5399 = n5224 | n5391 ;
  assign n5401 = ( n5398 & ~n5400 ) | ( n5398 & n5399 ) | ( ~n5400 & n5399 ) ;
  assign n5255 = n5084 &  n5253 ;
  assign n5256 = n5252 &  n5255 ;
  assign n5085 = x78 | n5084 ;
  assign n5086 = x78 &  n5084 ;
  assign n5087 = ( n5085 & ~n5086 ) | ( n5085 & 1'b0 ) | ( ~n5086 & 1'b0 ) ;
  assign n5258 = ( n5076 & n5087 ) | ( n5076 & n5254 ) | ( n5087 & n5254 ) ;
  assign n5257 = n5076 | n5087 ;
  assign n5259 = ( n5256 & ~n5258 ) | ( n5256 & n5257 ) | ( ~n5258 & n5257 ) ;
  assign n5405 = n4962 &  n5253 ;
  assign n5406 = n5252 &  n5405 ;
  assign n5073 = x77 | n4962 ;
  assign n5074 = x77 &  n4962 ;
  assign n5075 = ( n5073 & ~n5074 ) | ( n5073 & 1'b0 ) | ( ~n5074 & 1'b0 ) ;
  assign n5407 = n5072 &  n5075 ;
  assign n5408 = ( n5072 & ~n5254 ) | ( n5072 & n5075 ) | ( ~n5254 & n5075 ) ;
  assign n5409 = ( n5406 & ~n5407 ) | ( n5406 & n5408 ) | ( ~n5407 & n5408 ) ;
  assign n5413 = n4970 &  n5253 ;
  assign n5414 = n5252 &  n5413 ;
  assign n5402 = x76 | n4970 ;
  assign n5403 = x76 &  n4970 ;
  assign n5404 = ( n5402 & ~n5403 ) | ( n5402 & 1'b0 ) | ( ~n5403 & 1'b0 ) ;
  assign n5416 = ( n5071 & n5254 ) | ( n5071 & n5404 ) | ( n5254 & n5404 ) ;
  assign n5415 = n5071 | n5404 ;
  assign n5417 = ( n5414 & ~n5416 ) | ( n5414 & n5415 ) | ( ~n5416 & n5415 ) ;
  assign n5421 = n4978 &  n5253 ;
  assign n5422 = n5252 &  n5421 ;
  assign n5410 = x75 | n4978 ;
  assign n5411 = x75 &  n4978 ;
  assign n5412 = ( n5410 & ~n5411 ) | ( n5410 & 1'b0 ) | ( ~n5411 & 1'b0 ) ;
  assign n5424 = ( n5070 & n5254 ) | ( n5070 & n5412 ) | ( n5254 & n5412 ) ;
  assign n5423 = n5070 | n5412 ;
  assign n5425 = ( n5422 & ~n5424 ) | ( n5422 & n5423 ) | ( ~n5424 & n5423 ) ;
  assign n5429 = n4986 &  n5253 ;
  assign n5430 = n5252 &  n5429 ;
  assign n5418 = x74 | n4986 ;
  assign n5419 = x74 &  n4986 ;
  assign n5420 = ( n5418 & ~n5419 ) | ( n5418 & 1'b0 ) | ( ~n5419 & 1'b0 ) ;
  assign n5432 = ( n5069 & n5254 ) | ( n5069 & n5420 ) | ( n5254 & n5420 ) ;
  assign n5431 = n5069 | n5420 ;
  assign n5433 = ( n5430 & ~n5432 ) | ( n5430 & n5431 ) | ( ~n5432 & n5431 ) ;
  assign n5437 = n4994 &  n5253 ;
  assign n5438 = n5252 &  n5437 ;
  assign n5426 = x73 | n4994 ;
  assign n5427 = x73 &  n4994 ;
  assign n5428 = ( n5426 & ~n5427 ) | ( n5426 & 1'b0 ) | ( ~n5427 & 1'b0 ) ;
  assign n5440 = ( n5068 & n5254 ) | ( n5068 & n5428 ) | ( n5254 & n5428 ) ;
  assign n5439 = n5068 | n5428 ;
  assign n5441 = ( n5438 & ~n5440 ) | ( n5438 & n5439 ) | ( ~n5440 & n5439 ) ;
  assign n5445 = n5002 &  n5253 ;
  assign n5446 = n5252 &  n5445 ;
  assign n5434 = x72 | n5002 ;
  assign n5435 = x72 &  n5002 ;
  assign n5436 = ( n5434 & ~n5435 ) | ( n5434 & 1'b0 ) | ( ~n5435 & 1'b0 ) ;
  assign n5448 = ( n5067 & n5254 ) | ( n5067 & n5436 ) | ( n5254 & n5436 ) ;
  assign n5447 = n5067 | n5436 ;
  assign n5449 = ( n5446 & ~n5448 ) | ( n5446 & n5447 ) | ( ~n5448 & n5447 ) ;
  assign n5453 = n5010 &  n5253 ;
  assign n5454 = n5252 &  n5453 ;
  assign n5442 = x71 | n5010 ;
  assign n5443 = x71 &  n5010 ;
  assign n5444 = ( n5442 & ~n5443 ) | ( n5442 & 1'b0 ) | ( ~n5443 & 1'b0 ) ;
  assign n5456 = ( n5066 & n5254 ) | ( n5066 & n5444 ) | ( n5254 & n5444 ) ;
  assign n5455 = n5066 | n5444 ;
  assign n5457 = ( n5454 & ~n5456 ) | ( n5454 & n5455 ) | ( ~n5456 & n5455 ) ;
  assign n5461 = n5018 &  n5253 ;
  assign n5462 = n5252 &  n5461 ;
  assign n5450 = x70 | n5018 ;
  assign n5451 = x70 &  n5018 ;
  assign n5452 = ( n5450 & ~n5451 ) | ( n5450 & 1'b0 ) | ( ~n5451 & 1'b0 ) ;
  assign n5464 = ( n5065 & n5254 ) | ( n5065 & n5452 ) | ( n5254 & n5452 ) ;
  assign n5463 = n5065 | n5452 ;
  assign n5465 = ( n5462 & ~n5464 ) | ( n5462 & n5463 ) | ( ~n5464 & n5463 ) ;
  assign n5469 = n5026 &  n5253 ;
  assign n5470 = n5252 &  n5469 ;
  assign n5458 = x69 | n5026 ;
  assign n5459 = x69 &  n5026 ;
  assign n5460 = ( n5458 & ~n5459 ) | ( n5458 & 1'b0 ) | ( ~n5459 & 1'b0 ) ;
  assign n5472 = ( n5064 & n5254 ) | ( n5064 & n5460 ) | ( n5254 & n5460 ) ;
  assign n5471 = n5064 | n5460 ;
  assign n5473 = ( n5470 & ~n5472 ) | ( n5470 & n5471 ) | ( ~n5472 & n5471 ) ;
  assign n5477 = n5034 &  n5253 ;
  assign n5478 = n5252 &  n5477 ;
  assign n5466 = x68 | n5034 ;
  assign n5467 = x68 &  n5034 ;
  assign n5468 = ( n5466 & ~n5467 ) | ( n5466 & 1'b0 ) | ( ~n5467 & 1'b0 ) ;
  assign n5480 = ( n5063 & n5254 ) | ( n5063 & n5468 ) | ( n5254 & n5468 ) ;
  assign n5479 = n5063 | n5468 ;
  assign n5481 = ( n5478 & ~n5480 ) | ( n5478 & n5479 ) | ( ~n5480 & n5479 ) ;
  assign n5485 = n5042 &  n5253 ;
  assign n5486 = n5252 &  n5485 ;
  assign n5474 = x67 | n5042 ;
  assign n5475 = x67 &  n5042 ;
  assign n5476 = ( n5474 & ~n5475 ) | ( n5474 & 1'b0 ) | ( ~n5475 & 1'b0 ) ;
  assign n5488 = ( n5062 & n5254 ) | ( n5062 & n5476 ) | ( n5254 & n5476 ) ;
  assign n5487 = n5062 | n5476 ;
  assign n5489 = ( n5486 & ~n5488 ) | ( n5486 & n5487 ) | ( ~n5488 & n5487 ) ;
  assign n5490 = n5048 &  n5253 ;
  assign n5491 = n5252 &  n5490 ;
  assign n5482 = x66 | n5048 ;
  assign n5483 = x66 &  n5048 ;
  assign n5484 = ( n5482 & ~n5483 ) | ( n5482 & 1'b0 ) | ( ~n5483 & 1'b0 ) ;
  assign n5492 = n5061 &  n5484 ;
  assign n5493 = ( n5061 & ~n5254 ) | ( n5061 & n5484 ) | ( ~n5254 & n5484 ) ;
  assign n5494 = ( n5491 & ~n5492 ) | ( n5491 & n5493 ) | ( ~n5492 & n5493 ) ;
  assign n5495 = ( n5059 & ~x65 ) | ( n5059 & n5060 ) | ( ~x65 & n5060 ) ;
  assign n5496 = ( n5061 & ~n5060 ) | ( n5061 & n5495 ) | ( ~n5060 & n5495 ) ;
  assign n5497 = ~n5254 & n5496 ;
  assign n5498 = n5059 &  n5253 ;
  assign n5499 = n5252 &  n5498 ;
  assign n5500 = n5497 | n5499 ;
  assign n5501 = ( x64 & ~n5254 ) | ( x64 & 1'b0 ) | ( ~n5254 & 1'b0 ) ;
  assign n5502 = ( x31 & ~n5501 ) | ( x31 & 1'b0 ) | ( ~n5501 & 1'b0 ) ;
  assign n5503 = ( n5060 & ~n5254 ) | ( n5060 & 1'b0 ) | ( ~n5254 & 1'b0 ) ;
  assign n5504 = n5502 | n5503 ;
  assign n5505 = ~x30 & x64 ;
  assign n5506 = ( x65 & ~n5504 ) | ( x65 & n5505 ) | ( ~n5504 & n5505 ) ;
  assign n5507 = ( x66 & ~n5500 ) | ( x66 & n5506 ) | ( ~n5500 & n5506 ) ;
  assign n5508 = ( x67 & ~n5494 ) | ( x67 & n5507 ) | ( ~n5494 & n5507 ) ;
  assign n5509 = ( x68 & ~n5489 ) | ( x68 & n5508 ) | ( ~n5489 & n5508 ) ;
  assign n5510 = ( x69 & ~n5481 ) | ( x69 & n5509 ) | ( ~n5481 & n5509 ) ;
  assign n5511 = ( x70 & ~n5473 ) | ( x70 & n5510 ) | ( ~n5473 & n5510 ) ;
  assign n5512 = ( x71 & ~n5465 ) | ( x71 & n5511 ) | ( ~n5465 & n5511 ) ;
  assign n5513 = ( x72 & ~n5457 ) | ( x72 & n5512 ) | ( ~n5457 & n5512 ) ;
  assign n5514 = ( x73 & ~n5449 ) | ( x73 & n5513 ) | ( ~n5449 & n5513 ) ;
  assign n5515 = ( x74 & ~n5441 ) | ( x74 & n5514 ) | ( ~n5441 & n5514 ) ;
  assign n5516 = ( x75 & ~n5433 ) | ( x75 & n5515 ) | ( ~n5433 & n5515 ) ;
  assign n5517 = ( x76 & ~n5425 ) | ( x76 & n5516 ) | ( ~n5425 & n5516 ) ;
  assign n5518 = ( x77 & ~n5417 ) | ( x77 & n5517 ) | ( ~n5417 & n5517 ) ;
  assign n5519 = ( x78 & ~n5409 ) | ( x78 & n5518 ) | ( ~n5409 & n5518 ) ;
  assign n5520 = ( x79 & ~n5259 ) | ( x79 & n5519 ) | ( ~n5259 & n5519 ) ;
  assign n5521 = ( x80 & ~n5401 ) | ( x80 & n5520 ) | ( ~n5401 & n5520 ) ;
  assign n5522 = ( x81 & ~n5396 ) | ( x81 & n5521 ) | ( ~n5396 & n5521 ) ;
  assign n5523 = ( x82 & ~n5388 ) | ( x82 & n5522 ) | ( ~n5388 & n5522 ) ;
  assign n5524 = ( x83 & ~n5380 ) | ( x83 & n5523 ) | ( ~n5380 & n5523 ) ;
  assign n5525 = ( x84 & ~n5372 ) | ( x84 & n5524 ) | ( ~n5372 & n5524 ) ;
  assign n5526 = ( x85 & ~n5364 ) | ( x85 & n5525 ) | ( ~n5364 & n5525 ) ;
  assign n5527 = ( x86 & ~n5356 ) | ( x86 & n5526 ) | ( ~n5356 & n5526 ) ;
  assign n5528 = ( x87 & ~n5348 ) | ( x87 & n5527 ) | ( ~n5348 & n5527 ) ;
  assign n5529 = ( x88 & ~n5340 ) | ( x88 & n5528 ) | ( ~n5340 & n5528 ) ;
  assign n5530 = ( x89 & ~n5332 ) | ( x89 & n5529 ) | ( ~n5332 & n5529 ) ;
  assign n5531 = ( x90 & ~n5324 ) | ( x90 & n5530 ) | ( ~n5324 & n5530 ) ;
  assign n5532 = ( x91 & ~n5316 ) | ( x91 & n5531 ) | ( ~n5316 & n5531 ) ;
  assign n5533 = ( x92 & ~n5308 ) | ( x92 & n5532 ) | ( ~n5308 & n5532 ) ;
  assign n5534 = ( x93 & ~n5300 ) | ( x93 & n5533 ) | ( ~n5300 & n5533 ) ;
  assign n5535 = ( x94 & ~n5292 ) | ( x94 & n5534 ) | ( ~n5292 & n5534 ) ;
  assign n5536 = ( x95 & ~n5284 ) | ( x95 & n5535 ) | ( ~n5284 & n5535 ) ;
  assign n5537 = ( x96 & ~n5276 ) | ( x96 & n5536 ) | ( ~n5276 & n5536 ) ;
  assign n5538 = ( x97 & ~n5268 ) | ( x97 & n5537 ) | ( ~n5268 & n5537 ) ;
  assign n5539 = n166 | n184 ;
  assign n5540 = ( n272 & ~n270 ) | ( n272 & n5539 ) | ( ~n270 & n5539 ) ;
  assign n5541 = n270 | n5540 ;
  assign n5542 = n5538 | n5541 ;
  assign n5560 = n5276 &  n5542 ;
  assign n5554 = x96 | n5276 ;
  assign n5555 = x96 &  n5276 ;
  assign n5556 = ( n5554 & ~n5555 ) | ( n5554 & 1'b0 ) | ( ~n5555 & 1'b0 ) ;
  assign n5564 = ( n5536 & n5538 ) | ( n5536 & n5556 ) | ( n5538 & n5556 ) ;
  assign n5565 = ( n5536 & ~n5541 ) | ( n5536 & n5556 ) | ( ~n5541 & n5556 ) ;
  assign n5566 = ~n5564 & n5565 ;
  assign n5567 = n5560 | n5566 ;
  assign n5557 = x97 | n5537 ;
  assign n5558 = ( x97 & n5537 ) | ( x97 & n5541 ) | ( n5537 & n5541 ) ;
  assign n5559 = ( n5268 & ~n5557 ) | ( n5268 & n5558 ) | ( ~n5557 & n5558 ) ;
  assign n5568 = n5284 &  n5542 ;
  assign n5561 = x95 | n5284 ;
  assign n5562 = x95 &  n5284 ;
  assign n5563 = ( n5561 & ~n5562 ) | ( n5561 & 1'b0 ) | ( ~n5562 & 1'b0 ) ;
  assign n5572 = ( n5535 & n5538 ) | ( n5535 & n5563 ) | ( n5538 & n5563 ) ;
  assign n5573 = ( n5535 & ~n5541 ) | ( n5535 & n5563 ) | ( ~n5541 & n5563 ) ;
  assign n5574 = ~n5572 & n5573 ;
  assign n5575 = n5568 | n5574 ;
  assign n5576 = n5292 &  n5542 ;
  assign n5569 = x94 | n5292 ;
  assign n5570 = x94 &  n5292 ;
  assign n5571 = ( n5569 & ~n5570 ) | ( n5569 & 1'b0 ) | ( ~n5570 & 1'b0 ) ;
  assign n5580 = ( n5534 & n5538 ) | ( n5534 & n5571 ) | ( n5538 & n5571 ) ;
  assign n5581 = ( n5534 & ~n5541 ) | ( n5534 & n5571 ) | ( ~n5541 & n5571 ) ;
  assign n5582 = ~n5580 & n5581 ;
  assign n5583 = n5576 | n5582 ;
  assign n5584 = n5300 &  n5542 ;
  assign n5577 = x93 | n5300 ;
  assign n5578 = x93 &  n5300 ;
  assign n5579 = ( n5577 & ~n5578 ) | ( n5577 & 1'b0 ) | ( ~n5578 & 1'b0 ) ;
  assign n5588 = ( n5533 & n5538 ) | ( n5533 & n5579 ) | ( n5538 & n5579 ) ;
  assign n5589 = ( n5533 & ~n5541 ) | ( n5533 & n5579 ) | ( ~n5541 & n5579 ) ;
  assign n5590 = ~n5588 & n5589 ;
  assign n5591 = n5584 | n5590 ;
  assign n5592 = n5308 &  n5542 ;
  assign n5585 = x92 | n5308 ;
  assign n5586 = x92 &  n5308 ;
  assign n5587 = ( n5585 & ~n5586 ) | ( n5585 & 1'b0 ) | ( ~n5586 & 1'b0 ) ;
  assign n5596 = ( n5532 & n5538 ) | ( n5532 & n5587 ) | ( n5538 & n5587 ) ;
  assign n5597 = ( n5532 & ~n5541 ) | ( n5532 & n5587 ) | ( ~n5541 & n5587 ) ;
  assign n5598 = ~n5596 & n5597 ;
  assign n5599 = n5592 | n5598 ;
  assign n5600 = n5316 &  n5542 ;
  assign n5593 = x91 | n5316 ;
  assign n5594 = x91 &  n5316 ;
  assign n5595 = ( n5593 & ~n5594 ) | ( n5593 & 1'b0 ) | ( ~n5594 & 1'b0 ) ;
  assign n5604 = ( n5531 & n5538 ) | ( n5531 & n5595 ) | ( n5538 & n5595 ) ;
  assign n5605 = ( n5531 & ~n5541 ) | ( n5531 & n5595 ) | ( ~n5541 & n5595 ) ;
  assign n5606 = ~n5604 & n5605 ;
  assign n5607 = n5600 | n5606 ;
  assign n5608 = n5324 &  n5542 ;
  assign n5601 = x90 | n5324 ;
  assign n5602 = x90 &  n5324 ;
  assign n5603 = ( n5601 & ~n5602 ) | ( n5601 & 1'b0 ) | ( ~n5602 & 1'b0 ) ;
  assign n5612 = ( n5530 & n5538 ) | ( n5530 & n5603 ) | ( n5538 & n5603 ) ;
  assign n5613 = ( n5530 & ~n5541 ) | ( n5530 & n5603 ) | ( ~n5541 & n5603 ) ;
  assign n5614 = ~n5612 & n5613 ;
  assign n5615 = n5608 | n5614 ;
  assign n5616 = n5332 &  n5542 ;
  assign n5609 = x89 | n5332 ;
  assign n5610 = x89 &  n5332 ;
  assign n5611 = ( n5609 & ~n5610 ) | ( n5609 & 1'b0 ) | ( ~n5610 & 1'b0 ) ;
  assign n5620 = ( n5529 & n5538 ) | ( n5529 & n5611 ) | ( n5538 & n5611 ) ;
  assign n5621 = ( n5529 & ~n5541 ) | ( n5529 & n5611 ) | ( ~n5541 & n5611 ) ;
  assign n5622 = ~n5620 & n5621 ;
  assign n5623 = n5616 | n5622 ;
  assign n5624 = n5340 &  n5542 ;
  assign n5617 = x88 | n5340 ;
  assign n5618 = x88 &  n5340 ;
  assign n5619 = ( n5617 & ~n5618 ) | ( n5617 & 1'b0 ) | ( ~n5618 & 1'b0 ) ;
  assign n5628 = ( n5528 & n5538 ) | ( n5528 & n5619 ) | ( n5538 & n5619 ) ;
  assign n5629 = ( n5528 & ~n5541 ) | ( n5528 & n5619 ) | ( ~n5541 & n5619 ) ;
  assign n5630 = ~n5628 & n5629 ;
  assign n5631 = n5624 | n5630 ;
  assign n5632 = n5348 &  n5542 ;
  assign n5625 = x87 | n5348 ;
  assign n5626 = x87 &  n5348 ;
  assign n5627 = ( n5625 & ~n5626 ) | ( n5625 & 1'b0 ) | ( ~n5626 & 1'b0 ) ;
  assign n5636 = ( n5527 & n5538 ) | ( n5527 & n5627 ) | ( n5538 & n5627 ) ;
  assign n5637 = ( n5527 & ~n5541 ) | ( n5527 & n5627 ) | ( ~n5541 & n5627 ) ;
  assign n5638 = ~n5636 & n5637 ;
  assign n5639 = n5632 | n5638 ;
  assign n5640 = n5356 &  n5542 ;
  assign n5633 = x86 | n5356 ;
  assign n5634 = x86 &  n5356 ;
  assign n5635 = ( n5633 & ~n5634 ) | ( n5633 & 1'b0 ) | ( ~n5634 & 1'b0 ) ;
  assign n5644 = ( n5526 & n5538 ) | ( n5526 & n5635 ) | ( n5538 & n5635 ) ;
  assign n5645 = ( n5526 & ~n5541 ) | ( n5526 & n5635 ) | ( ~n5541 & n5635 ) ;
  assign n5646 = ~n5644 & n5645 ;
  assign n5647 = n5640 | n5646 ;
  assign n5648 = n5364 &  n5542 ;
  assign n5641 = x85 | n5364 ;
  assign n5642 = x85 &  n5364 ;
  assign n5643 = ( n5641 & ~n5642 ) | ( n5641 & 1'b0 ) | ( ~n5642 & 1'b0 ) ;
  assign n5652 = ( n5525 & n5538 ) | ( n5525 & n5643 ) | ( n5538 & n5643 ) ;
  assign n5653 = ( n5525 & ~n5541 ) | ( n5525 & n5643 ) | ( ~n5541 & n5643 ) ;
  assign n5654 = ~n5652 & n5653 ;
  assign n5655 = n5648 | n5654 ;
  assign n5656 = n5372 &  n5542 ;
  assign n5649 = x84 | n5372 ;
  assign n5650 = x84 &  n5372 ;
  assign n5651 = ( n5649 & ~n5650 ) | ( n5649 & 1'b0 ) | ( ~n5650 & 1'b0 ) ;
  assign n5660 = ( n5524 & n5538 ) | ( n5524 & n5651 ) | ( n5538 & n5651 ) ;
  assign n5661 = ( n5524 & ~n5541 ) | ( n5524 & n5651 ) | ( ~n5541 & n5651 ) ;
  assign n5662 = ~n5660 & n5661 ;
  assign n5663 = n5656 | n5662 ;
  assign n5664 = n5380 &  n5542 ;
  assign n5657 = x83 | n5380 ;
  assign n5658 = x83 &  n5380 ;
  assign n5659 = ( n5657 & ~n5658 ) | ( n5657 & 1'b0 ) | ( ~n5658 & 1'b0 ) ;
  assign n5668 = ( n5523 & n5538 ) | ( n5523 & n5659 ) | ( n5538 & n5659 ) ;
  assign n5669 = ( n5523 & ~n5541 ) | ( n5523 & n5659 ) | ( ~n5541 & n5659 ) ;
  assign n5670 = ~n5668 & n5669 ;
  assign n5671 = n5664 | n5670 ;
  assign n5672 = n5388 &  n5542 ;
  assign n5665 = x82 | n5388 ;
  assign n5666 = x82 &  n5388 ;
  assign n5667 = ( n5665 & ~n5666 ) | ( n5665 & 1'b0 ) | ( ~n5666 & 1'b0 ) ;
  assign n5676 = ( n5522 & n5538 ) | ( n5522 & n5667 ) | ( n5538 & n5667 ) ;
  assign n5677 = ( n5522 & ~n5541 ) | ( n5522 & n5667 ) | ( ~n5541 & n5667 ) ;
  assign n5678 = ~n5676 & n5677 ;
  assign n5679 = n5672 | n5678 ;
  assign n5680 = n5396 &  n5542 ;
  assign n5673 = x81 | n5396 ;
  assign n5674 = x81 &  n5396 ;
  assign n5675 = ( n5673 & ~n5674 ) | ( n5673 & 1'b0 ) | ( ~n5674 & 1'b0 ) ;
  assign n5684 = ( n5521 & n5538 ) | ( n5521 & n5675 ) | ( n5538 & n5675 ) ;
  assign n5685 = ( n5521 & ~n5541 ) | ( n5521 & n5675 ) | ( ~n5541 & n5675 ) ;
  assign n5686 = ~n5684 & n5685 ;
  assign n5687 = n5680 | n5686 ;
  assign n5688 = n5401 &  n5542 ;
  assign n5681 = x80 | n5401 ;
  assign n5682 = x80 &  n5401 ;
  assign n5683 = ( n5681 & ~n5682 ) | ( n5681 & 1'b0 ) | ( ~n5682 & 1'b0 ) ;
  assign n5689 = ( n5520 & n5538 ) | ( n5520 & n5683 ) | ( n5538 & n5683 ) ;
  assign n5690 = ( n5520 & ~n5541 ) | ( n5520 & n5683 ) | ( ~n5541 & n5683 ) ;
  assign n5691 = ~n5689 & n5690 ;
  assign n5692 = n5688 | n5691 ;
  assign n5543 = n5259 &  n5542 ;
  assign n5547 = x79 | n5259 ;
  assign n5548 = x79 &  n5259 ;
  assign n5549 = ( n5547 & ~n5548 ) | ( n5547 & 1'b0 ) | ( ~n5548 & 1'b0 ) ;
  assign n5550 = ( n5519 & n5538 ) | ( n5519 & n5549 ) | ( n5538 & n5549 ) ;
  assign n5551 = ( n5519 & ~n5541 ) | ( n5519 & n5549 ) | ( ~n5541 & n5549 ) ;
  assign n5552 = ~n5550 & n5551 ;
  assign n5553 = n5543 | n5552 ;
  assign n5693 = n5409 &  n5542 ;
  assign n5544 = x78 | n5409 ;
  assign n5545 = x78 &  n5409 ;
  assign n5546 = ( n5544 & ~n5545 ) | ( n5544 & 1'b0 ) | ( ~n5545 & 1'b0 ) ;
  assign n5697 = ( n5518 & n5538 ) | ( n5518 & n5546 ) | ( n5538 & n5546 ) ;
  assign n5698 = ( n5518 & ~n5541 ) | ( n5518 & n5546 ) | ( ~n5541 & n5546 ) ;
  assign n5699 = ~n5697 & n5698 ;
  assign n5700 = n5693 | n5699 ;
  assign n5701 = n5417 &  n5542 ;
  assign n5694 = x77 | n5417 ;
  assign n5695 = x77 &  n5417 ;
  assign n5696 = ( n5694 & ~n5695 ) | ( n5694 & 1'b0 ) | ( ~n5695 & 1'b0 ) ;
  assign n5705 = ( n5517 & n5538 ) | ( n5517 & n5696 ) | ( n5538 & n5696 ) ;
  assign n5706 = ( n5517 & ~n5541 ) | ( n5517 & n5696 ) | ( ~n5541 & n5696 ) ;
  assign n5707 = ~n5705 & n5706 ;
  assign n5708 = n5701 | n5707 ;
  assign n5709 = n5425 &  n5542 ;
  assign n5702 = x76 | n5425 ;
  assign n5703 = x76 &  n5425 ;
  assign n5704 = ( n5702 & ~n5703 ) | ( n5702 & 1'b0 ) | ( ~n5703 & 1'b0 ) ;
  assign n5713 = ( n5516 & n5538 ) | ( n5516 & n5704 ) | ( n5538 & n5704 ) ;
  assign n5714 = ( n5516 & ~n5541 ) | ( n5516 & n5704 ) | ( ~n5541 & n5704 ) ;
  assign n5715 = ~n5713 & n5714 ;
  assign n5716 = n5709 | n5715 ;
  assign n5717 = n5433 &  n5542 ;
  assign n5710 = x75 | n5433 ;
  assign n5711 = x75 &  n5433 ;
  assign n5712 = ( n5710 & ~n5711 ) | ( n5710 & 1'b0 ) | ( ~n5711 & 1'b0 ) ;
  assign n5721 = ( n5515 & n5538 ) | ( n5515 & n5712 ) | ( n5538 & n5712 ) ;
  assign n5722 = ( n5515 & ~n5541 ) | ( n5515 & n5712 ) | ( ~n5541 & n5712 ) ;
  assign n5723 = ~n5721 & n5722 ;
  assign n5724 = n5717 | n5723 ;
  assign n5725 = n5441 &  n5542 ;
  assign n5718 = x74 | n5441 ;
  assign n5719 = x74 &  n5441 ;
  assign n5720 = ( n5718 & ~n5719 ) | ( n5718 & 1'b0 ) | ( ~n5719 & 1'b0 ) ;
  assign n5729 = ( n5514 & n5538 ) | ( n5514 & n5720 ) | ( n5538 & n5720 ) ;
  assign n5730 = ( n5514 & ~n5541 ) | ( n5514 & n5720 ) | ( ~n5541 & n5720 ) ;
  assign n5731 = ~n5729 & n5730 ;
  assign n5732 = n5725 | n5731 ;
  assign n5733 = n5449 &  n5542 ;
  assign n5726 = x73 | n5449 ;
  assign n5727 = x73 &  n5449 ;
  assign n5728 = ( n5726 & ~n5727 ) | ( n5726 & 1'b0 ) | ( ~n5727 & 1'b0 ) ;
  assign n5737 = ( n5513 & n5538 ) | ( n5513 & n5728 ) | ( n5538 & n5728 ) ;
  assign n5738 = ( n5513 & ~n5541 ) | ( n5513 & n5728 ) | ( ~n5541 & n5728 ) ;
  assign n5739 = ~n5737 & n5738 ;
  assign n5740 = n5733 | n5739 ;
  assign n5741 = n5457 &  n5542 ;
  assign n5734 = x72 | n5457 ;
  assign n5735 = x72 &  n5457 ;
  assign n5736 = ( n5734 & ~n5735 ) | ( n5734 & 1'b0 ) | ( ~n5735 & 1'b0 ) ;
  assign n5745 = ( n5512 & n5538 ) | ( n5512 & n5736 ) | ( n5538 & n5736 ) ;
  assign n5746 = ( n5512 & ~n5541 ) | ( n5512 & n5736 ) | ( ~n5541 & n5736 ) ;
  assign n5747 = ~n5745 & n5746 ;
  assign n5748 = n5741 | n5747 ;
  assign n5749 = n5465 &  n5542 ;
  assign n5742 = x71 | n5465 ;
  assign n5743 = x71 &  n5465 ;
  assign n5744 = ( n5742 & ~n5743 ) | ( n5742 & 1'b0 ) | ( ~n5743 & 1'b0 ) ;
  assign n5753 = ( n5511 & n5538 ) | ( n5511 & n5744 ) | ( n5538 & n5744 ) ;
  assign n5754 = ( n5511 & ~n5541 ) | ( n5511 & n5744 ) | ( ~n5541 & n5744 ) ;
  assign n5755 = ~n5753 & n5754 ;
  assign n5756 = n5749 | n5755 ;
  assign n5757 = n5473 &  n5542 ;
  assign n5750 = x70 | n5473 ;
  assign n5751 = x70 &  n5473 ;
  assign n5752 = ( n5750 & ~n5751 ) | ( n5750 & 1'b0 ) | ( ~n5751 & 1'b0 ) ;
  assign n5761 = ( n5510 & n5538 ) | ( n5510 & n5752 ) | ( n5538 & n5752 ) ;
  assign n5762 = ( n5510 & ~n5541 ) | ( n5510 & n5752 ) | ( ~n5541 & n5752 ) ;
  assign n5763 = ~n5761 & n5762 ;
  assign n5764 = n5757 | n5763 ;
  assign n5765 = n5481 &  n5542 ;
  assign n5758 = x69 | n5481 ;
  assign n5759 = x69 &  n5481 ;
  assign n5760 = ( n5758 & ~n5759 ) | ( n5758 & 1'b0 ) | ( ~n5759 & 1'b0 ) ;
  assign n5769 = ( n5509 & n5538 ) | ( n5509 & n5760 ) | ( n5538 & n5760 ) ;
  assign n5770 = ( n5509 & ~n5541 ) | ( n5509 & n5760 ) | ( ~n5541 & n5760 ) ;
  assign n5771 = ~n5769 & n5770 ;
  assign n5772 = n5765 | n5771 ;
  assign n5773 = n5489 &  n5542 ;
  assign n5766 = x68 | n5489 ;
  assign n5767 = x68 &  n5489 ;
  assign n5768 = ( n5766 & ~n5767 ) | ( n5766 & 1'b0 ) | ( ~n5767 & 1'b0 ) ;
  assign n5777 = ( n5508 & n5538 ) | ( n5508 & n5768 ) | ( n5538 & n5768 ) ;
  assign n5778 = ( n5508 & ~n5541 ) | ( n5508 & n5768 ) | ( ~n5541 & n5768 ) ;
  assign n5779 = ~n5777 & n5778 ;
  assign n5780 = n5773 | n5779 ;
  assign n5781 = n5494 &  n5542 ;
  assign n5774 = x67 | n5494 ;
  assign n5775 = x67 &  n5494 ;
  assign n5776 = ( n5774 & ~n5775 ) | ( n5774 & 1'b0 ) | ( ~n5775 & 1'b0 ) ;
  assign n5785 = ( n5507 & n5538 ) | ( n5507 & n5776 ) | ( n5538 & n5776 ) ;
  assign n5786 = ( n5507 & ~n5541 ) | ( n5507 & n5776 ) | ( ~n5541 & n5776 ) ;
  assign n5787 = ~n5785 & n5786 ;
  assign n5788 = n5781 | n5787 ;
  assign n5789 = n5500 &  n5542 ;
  assign n5782 = x66 | n5500 ;
  assign n5783 = x66 &  n5500 ;
  assign n5784 = ( n5782 & ~n5783 ) | ( n5782 & 1'b0 ) | ( ~n5783 & 1'b0 ) ;
  assign n5794 = ( n5506 & ~n5538 ) | ( n5506 & n5784 ) | ( ~n5538 & n5784 ) ;
  assign n5795 = ( n5506 & n5541 ) | ( n5506 & n5784 ) | ( n5541 & n5784 ) ;
  assign n5796 = ( n5794 & ~n5795 ) | ( n5794 & 1'b0 ) | ( ~n5795 & 1'b0 ) ;
  assign n5797 = n5789 | n5796 ;
  assign n5798 = n5504 &  n5542 ;
  assign n5790 = x65 &  n5504 ;
  assign n5791 = ( n5502 & ~x65 ) | ( n5502 & n5503 ) | ( ~x65 & n5503 ) ;
  assign n5792 = x65 | n5791 ;
  assign n5793 = ( n5505 & ~n5790 ) | ( n5505 & n5792 ) | ( ~n5790 & n5792 ) ;
  assign n5799 = ( x65 & n5504 ) | ( x65 & n5505 ) | ( n5504 & n5505 ) ;
  assign n5800 = ( n5541 & ~n5790 ) | ( n5541 & n5799 ) | ( ~n5790 & n5799 ) ;
  assign n5801 = ( n5538 & n5793 ) | ( n5538 & n5800 ) | ( n5793 & n5800 ) ;
  assign n5802 = ( n5793 & ~n5801 ) | ( n5793 & 1'b0 ) | ( ~n5801 & 1'b0 ) ;
  assign n5803 = n5798 | n5802 ;
  assign n5804 = ( x64 & ~x98 ) | ( x64 & 1'b0 ) | ( ~x98 & 1'b0 ) ;
  assign n5805 = ( n243 & ~n245 ) | ( n243 & n5804 ) | ( ~n245 & n5804 ) ;
  assign n5806 = ~n243 & n5805 ;
  assign n5807 = ( n240 & ~n254 ) | ( n240 & n5806 ) | ( ~n254 & n5806 ) ;
  assign n5808 = ~n240 & n5807 ;
  assign n5809 = n5538 &  n5808 ;
  assign n5810 = ( x30 & ~n5808 ) | ( x30 & n5809 ) | ( ~n5808 & n5809 ) ;
  assign n5811 = ~n184 & n5505 ;
  assign n5812 = ( n166 & ~n272 ) | ( n166 & n5811 ) | ( ~n272 & n5811 ) ;
  assign n5813 = ~n166 & n5812 ;
  assign n5814 = ~n270 & n5813 ;
  assign n5815 = ~n5538 & n5814 ;
  assign n5816 = n5810 | n5815 ;
  assign n5817 = ~x29 & x64 ;
  assign n5818 = ( x65 & ~n5816 ) | ( x65 & n5817 ) | ( ~n5816 & n5817 ) ;
  assign n5819 = ( x66 & ~n5803 ) | ( x66 & n5818 ) | ( ~n5803 & n5818 ) ;
  assign n5820 = ( x67 & ~n5797 ) | ( x67 & n5819 ) | ( ~n5797 & n5819 ) ;
  assign n5821 = ( x68 & ~n5788 ) | ( x68 & n5820 ) | ( ~n5788 & n5820 ) ;
  assign n5822 = ( x69 & ~n5780 ) | ( x69 & n5821 ) | ( ~n5780 & n5821 ) ;
  assign n5823 = ( x70 & ~n5772 ) | ( x70 & n5822 ) | ( ~n5772 & n5822 ) ;
  assign n5824 = ( x71 & ~n5764 ) | ( x71 & n5823 ) | ( ~n5764 & n5823 ) ;
  assign n5825 = ( x72 & ~n5756 ) | ( x72 & n5824 ) | ( ~n5756 & n5824 ) ;
  assign n5826 = ( x73 & ~n5748 ) | ( x73 & n5825 ) | ( ~n5748 & n5825 ) ;
  assign n5827 = ( x74 & ~n5740 ) | ( x74 & n5826 ) | ( ~n5740 & n5826 ) ;
  assign n5828 = ( x75 & ~n5732 ) | ( x75 & n5827 ) | ( ~n5732 & n5827 ) ;
  assign n5829 = ( x76 & ~n5724 ) | ( x76 & n5828 ) | ( ~n5724 & n5828 ) ;
  assign n5830 = ( x77 & ~n5716 ) | ( x77 & n5829 ) | ( ~n5716 & n5829 ) ;
  assign n5831 = ( x78 & ~n5708 ) | ( x78 & n5830 ) | ( ~n5708 & n5830 ) ;
  assign n5832 = ( x79 & ~n5700 ) | ( x79 & n5831 ) | ( ~n5700 & n5831 ) ;
  assign n5833 = ( x80 & ~n5553 ) | ( x80 & n5832 ) | ( ~n5553 & n5832 ) ;
  assign n5834 = ( x81 & ~n5692 ) | ( x81 & n5833 ) | ( ~n5692 & n5833 ) ;
  assign n5835 = ( x82 & ~n5687 ) | ( x82 & n5834 ) | ( ~n5687 & n5834 ) ;
  assign n5836 = ( x83 & ~n5679 ) | ( x83 & n5835 ) | ( ~n5679 & n5835 ) ;
  assign n5837 = ( x84 & ~n5671 ) | ( x84 & n5836 ) | ( ~n5671 & n5836 ) ;
  assign n5838 = ( x85 & ~n5663 ) | ( x85 & n5837 ) | ( ~n5663 & n5837 ) ;
  assign n5839 = ( x86 & ~n5655 ) | ( x86 & n5838 ) | ( ~n5655 & n5838 ) ;
  assign n5840 = ( x87 & ~n5647 ) | ( x87 & n5839 ) | ( ~n5647 & n5839 ) ;
  assign n5841 = ( x88 & ~n5639 ) | ( x88 & n5840 ) | ( ~n5639 & n5840 ) ;
  assign n5842 = ( x89 & ~n5631 ) | ( x89 & n5841 ) | ( ~n5631 & n5841 ) ;
  assign n5843 = ( x90 & ~n5623 ) | ( x90 & n5842 ) | ( ~n5623 & n5842 ) ;
  assign n5844 = ( x91 & ~n5615 ) | ( x91 & n5843 ) | ( ~n5615 & n5843 ) ;
  assign n5845 = ( x92 & ~n5607 ) | ( x92 & n5844 ) | ( ~n5607 & n5844 ) ;
  assign n5846 = ( x93 & ~n5599 ) | ( x93 & n5845 ) | ( ~n5599 & n5845 ) ;
  assign n5847 = ( x94 & ~n5591 ) | ( x94 & n5846 ) | ( ~n5591 & n5846 ) ;
  assign n5848 = ( x95 & ~n5583 ) | ( x95 & n5847 ) | ( ~n5583 & n5847 ) ;
  assign n5849 = ( x96 & ~n5575 ) | ( x96 & n5848 ) | ( ~n5575 & n5848 ) ;
  assign n5850 = ( x97 & ~n5567 ) | ( x97 & n5849 ) | ( ~n5567 & n5849 ) ;
  assign n5851 = ( x98 & ~n5559 ) | ( x98 & n5850 ) | ( ~n5559 & n5850 ) ;
  assign n5852 = n243 | n245 ;
  assign n5853 = ( n254 & ~n240 ) | ( n254 & n5852 ) | ( ~n240 & n5852 ) ;
  assign n5854 = n240 | n5853 ;
  assign n5855 = n5851 | n5854 ;
  assign n6030 = n5567 &  n5855 ;
  assign n6034 = x97 | n5567 ;
  assign n6035 = x97 &  n5567 ;
  assign n6036 = ( n6034 & ~n6035 ) | ( n6034 & 1'b0 ) | ( ~n6035 & 1'b0 ) ;
  assign n6037 = ( n5849 & n5851 ) | ( n5849 & n6036 ) | ( n5851 & n6036 ) ;
  assign n6038 = ( n5849 & ~n5854 ) | ( n5849 & n6036 ) | ( ~n5854 & n6036 ) ;
  assign n6039 = ~n6037 & n6038 ;
  assign n6040 = n6030 | n6039 ;
  assign n6041 = n5575 &  n5855 ;
  assign n6031 = x96 | n5575 ;
  assign n6032 = x96 &  n5575 ;
  assign n6033 = ( n6031 & ~n6032 ) | ( n6031 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n6045 = ( n5848 & n5851 ) | ( n5848 & n6033 ) | ( n5851 & n6033 ) ;
  assign n6046 = ( n5848 & ~n5854 ) | ( n5848 & n6033 ) | ( ~n5854 & n6033 ) ;
  assign n6047 = ~n6045 & n6046 ;
  assign n6048 = n6041 | n6047 ;
  assign n6049 = n5583 &  n5855 ;
  assign n6042 = x95 | n5583 ;
  assign n6043 = x95 &  n5583 ;
  assign n6044 = ( n6042 & ~n6043 ) | ( n6042 & 1'b0 ) | ( ~n6043 & 1'b0 ) ;
  assign n6053 = ( n5847 & n5851 ) | ( n5847 & n6044 ) | ( n5851 & n6044 ) ;
  assign n6054 = ( n5847 & ~n5854 ) | ( n5847 & n6044 ) | ( ~n5854 & n6044 ) ;
  assign n6055 = ~n6053 & n6054 ;
  assign n6056 = n6049 | n6055 ;
  assign n6057 = n5591 &  n5855 ;
  assign n6050 = x94 | n5591 ;
  assign n6051 = x94 &  n5591 ;
  assign n6052 = ( n6050 & ~n6051 ) | ( n6050 & 1'b0 ) | ( ~n6051 & 1'b0 ) ;
  assign n6061 = ( n5846 & n5851 ) | ( n5846 & n6052 ) | ( n5851 & n6052 ) ;
  assign n6062 = ( n5846 & ~n5854 ) | ( n5846 & n6052 ) | ( ~n5854 & n6052 ) ;
  assign n6063 = ~n6061 & n6062 ;
  assign n6064 = n6057 | n6063 ;
  assign n6065 = n5599 &  n5855 ;
  assign n6058 = x93 | n5599 ;
  assign n6059 = x93 &  n5599 ;
  assign n6060 = ( n6058 & ~n6059 ) | ( n6058 & 1'b0 ) | ( ~n6059 & 1'b0 ) ;
  assign n6069 = ( n5845 & n5851 ) | ( n5845 & n6060 ) | ( n5851 & n6060 ) ;
  assign n6070 = ( n5845 & ~n5854 ) | ( n5845 & n6060 ) | ( ~n5854 & n6060 ) ;
  assign n6071 = ~n6069 & n6070 ;
  assign n6072 = n6065 | n6071 ;
  assign n6073 = n5607 &  n5855 ;
  assign n6066 = x92 | n5607 ;
  assign n6067 = x92 &  n5607 ;
  assign n6068 = ( n6066 & ~n6067 ) | ( n6066 & 1'b0 ) | ( ~n6067 & 1'b0 ) ;
  assign n6077 = ( n5844 & n5851 ) | ( n5844 & n6068 ) | ( n5851 & n6068 ) ;
  assign n6078 = ( n5844 & ~n5854 ) | ( n5844 & n6068 ) | ( ~n5854 & n6068 ) ;
  assign n6079 = ~n6077 & n6078 ;
  assign n6080 = n6073 | n6079 ;
  assign n6081 = n5615 &  n5855 ;
  assign n6074 = x91 | n5615 ;
  assign n6075 = x91 &  n5615 ;
  assign n6076 = ( n6074 & ~n6075 ) | ( n6074 & 1'b0 ) | ( ~n6075 & 1'b0 ) ;
  assign n6085 = ( n5843 & n5851 ) | ( n5843 & n6076 ) | ( n5851 & n6076 ) ;
  assign n6086 = ( n5843 & ~n5854 ) | ( n5843 & n6076 ) | ( ~n5854 & n6076 ) ;
  assign n6087 = ~n6085 & n6086 ;
  assign n6088 = n6081 | n6087 ;
  assign n6089 = n5623 &  n5855 ;
  assign n6082 = x90 | n5623 ;
  assign n6083 = x90 &  n5623 ;
  assign n6084 = ( n6082 & ~n6083 ) | ( n6082 & 1'b0 ) | ( ~n6083 & 1'b0 ) ;
  assign n6093 = ( n5842 & n5851 ) | ( n5842 & n6084 ) | ( n5851 & n6084 ) ;
  assign n6094 = ( n5842 & ~n5854 ) | ( n5842 & n6084 ) | ( ~n5854 & n6084 ) ;
  assign n6095 = ~n6093 & n6094 ;
  assign n6096 = n6089 | n6095 ;
  assign n6097 = n5631 &  n5855 ;
  assign n6090 = x89 | n5631 ;
  assign n6091 = x89 &  n5631 ;
  assign n6092 = ( n6090 & ~n6091 ) | ( n6090 & 1'b0 ) | ( ~n6091 & 1'b0 ) ;
  assign n6101 = ( n5841 & n5851 ) | ( n5841 & n6092 ) | ( n5851 & n6092 ) ;
  assign n6102 = ( n5841 & ~n5854 ) | ( n5841 & n6092 ) | ( ~n5854 & n6092 ) ;
  assign n6103 = ~n6101 & n6102 ;
  assign n6104 = n6097 | n6103 ;
  assign n6105 = n5639 &  n5855 ;
  assign n6098 = x88 | n5639 ;
  assign n6099 = x88 &  n5639 ;
  assign n6100 = ( n6098 & ~n6099 ) | ( n6098 & 1'b0 ) | ( ~n6099 & 1'b0 ) ;
  assign n6109 = ( n5840 & n5851 ) | ( n5840 & n6100 ) | ( n5851 & n6100 ) ;
  assign n6110 = ( n5840 & ~n5854 ) | ( n5840 & n6100 ) | ( ~n5854 & n6100 ) ;
  assign n6111 = ~n6109 & n6110 ;
  assign n6112 = n6105 | n6111 ;
  assign n6113 = n5647 &  n5855 ;
  assign n6106 = x87 | n5647 ;
  assign n6107 = x87 &  n5647 ;
  assign n6108 = ( n6106 & ~n6107 ) | ( n6106 & 1'b0 ) | ( ~n6107 & 1'b0 ) ;
  assign n6117 = ( n5839 & n5851 ) | ( n5839 & n6108 ) | ( n5851 & n6108 ) ;
  assign n6118 = ( n5839 & ~n5854 ) | ( n5839 & n6108 ) | ( ~n5854 & n6108 ) ;
  assign n6119 = ~n6117 & n6118 ;
  assign n6120 = n6113 | n6119 ;
  assign n6121 = n5655 &  n5855 ;
  assign n6114 = x86 | n5655 ;
  assign n6115 = x86 &  n5655 ;
  assign n6116 = ( n6114 & ~n6115 ) | ( n6114 & 1'b0 ) | ( ~n6115 & 1'b0 ) ;
  assign n6125 = ( n5838 & n5851 ) | ( n5838 & n6116 ) | ( n5851 & n6116 ) ;
  assign n6126 = ( n5838 & ~n5854 ) | ( n5838 & n6116 ) | ( ~n5854 & n6116 ) ;
  assign n6127 = ~n6125 & n6126 ;
  assign n6128 = n6121 | n6127 ;
  assign n6129 = n5663 &  n5855 ;
  assign n6122 = x85 | n5663 ;
  assign n6123 = x85 &  n5663 ;
  assign n6124 = ( n6122 & ~n6123 ) | ( n6122 & 1'b0 ) | ( ~n6123 & 1'b0 ) ;
  assign n6133 = ( n5837 & n5851 ) | ( n5837 & n6124 ) | ( n5851 & n6124 ) ;
  assign n6134 = ( n5837 & ~n5854 ) | ( n5837 & n6124 ) | ( ~n5854 & n6124 ) ;
  assign n6135 = ~n6133 & n6134 ;
  assign n6136 = n6129 | n6135 ;
  assign n6137 = n5671 &  n5855 ;
  assign n6130 = x84 | n5671 ;
  assign n6131 = x84 &  n5671 ;
  assign n6132 = ( n6130 & ~n6131 ) | ( n6130 & 1'b0 ) | ( ~n6131 & 1'b0 ) ;
  assign n6141 = ( n5836 & n5851 ) | ( n5836 & n6132 ) | ( n5851 & n6132 ) ;
  assign n6142 = ( n5836 & ~n5854 ) | ( n5836 & n6132 ) | ( ~n5854 & n6132 ) ;
  assign n6143 = ~n6141 & n6142 ;
  assign n6144 = n6137 | n6143 ;
  assign n6145 = n5679 &  n5855 ;
  assign n6138 = x83 | n5679 ;
  assign n6139 = x83 &  n5679 ;
  assign n6140 = ( n6138 & ~n6139 ) | ( n6138 & 1'b0 ) | ( ~n6139 & 1'b0 ) ;
  assign n6149 = ( n5835 & n5851 ) | ( n5835 & n6140 ) | ( n5851 & n6140 ) ;
  assign n6150 = ( n5835 & ~n5854 ) | ( n5835 & n6140 ) | ( ~n5854 & n6140 ) ;
  assign n6151 = ~n6149 & n6150 ;
  assign n6152 = n6145 | n6151 ;
  assign n6153 = n5687 &  n5855 ;
  assign n6146 = x82 | n5687 ;
  assign n6147 = x82 &  n5687 ;
  assign n6148 = ( n6146 & ~n6147 ) | ( n6146 & 1'b0 ) | ( ~n6147 & 1'b0 ) ;
  assign n6154 = ( n5834 & n5851 ) | ( n5834 & n6148 ) | ( n5851 & n6148 ) ;
  assign n6155 = ( n5834 & ~n5854 ) | ( n5834 & n6148 ) | ( ~n5854 & n6148 ) ;
  assign n6156 = ~n6154 & n6155 ;
  assign n6157 = n6153 | n6156 ;
  assign n6019 = n5692 &  n5855 ;
  assign n6020 = x81 | n5692 ;
  assign n6021 = x81 &  n5692 ;
  assign n6022 = ( n6020 & ~n6021 ) | ( n6020 & 1'b0 ) | ( ~n6021 & 1'b0 ) ;
  assign n6023 = ( n5833 & n5851 ) | ( n5833 & n6022 ) | ( n5851 & n6022 ) ;
  assign n6024 = ( n5833 & ~n5854 ) | ( n5833 & n6022 ) | ( ~n5854 & n6022 ) ;
  assign n6025 = ~n6023 & n6024 ;
  assign n6026 = n6019 | n6025 ;
  assign n5856 = n5553 &  n5855 ;
  assign n5860 = x80 | n5553 ;
  assign n5861 = x80 &  n5553 ;
  assign n5862 = ( n5860 & ~n5861 ) | ( n5860 & 1'b0 ) | ( ~n5861 & 1'b0 ) ;
  assign n5863 = ( n5832 & n5851 ) | ( n5832 & n5862 ) | ( n5851 & n5862 ) ;
  assign n5864 = ( n5832 & ~n5854 ) | ( n5832 & n5862 ) | ( ~n5854 & n5862 ) ;
  assign n5865 = ~n5863 & n5864 ;
  assign n5866 = n5856 | n5865 ;
  assign n5867 = n5700 &  n5855 ;
  assign n5857 = x79 | n5700 ;
  assign n5858 = x79 &  n5700 ;
  assign n5859 = ( n5857 & ~n5858 ) | ( n5857 & 1'b0 ) | ( ~n5858 & 1'b0 ) ;
  assign n5871 = ( n5831 & n5851 ) | ( n5831 & n5859 ) | ( n5851 & n5859 ) ;
  assign n5872 = ( n5831 & ~n5854 ) | ( n5831 & n5859 ) | ( ~n5854 & n5859 ) ;
  assign n5873 = ~n5871 & n5872 ;
  assign n5874 = n5867 | n5873 ;
  assign n5875 = n5708 &  n5855 ;
  assign n5868 = x78 | n5708 ;
  assign n5869 = x78 &  n5708 ;
  assign n5870 = ( n5868 & ~n5869 ) | ( n5868 & 1'b0 ) | ( ~n5869 & 1'b0 ) ;
  assign n5879 = ( n5830 & n5851 ) | ( n5830 & n5870 ) | ( n5851 & n5870 ) ;
  assign n5880 = ( n5830 & ~n5854 ) | ( n5830 & n5870 ) | ( ~n5854 & n5870 ) ;
  assign n5881 = ~n5879 & n5880 ;
  assign n5882 = n5875 | n5881 ;
  assign n5883 = n5716 &  n5855 ;
  assign n5876 = x77 | n5716 ;
  assign n5877 = x77 &  n5716 ;
  assign n5878 = ( n5876 & ~n5877 ) | ( n5876 & 1'b0 ) | ( ~n5877 & 1'b0 ) ;
  assign n5887 = ( n5829 & n5851 ) | ( n5829 & n5878 ) | ( n5851 & n5878 ) ;
  assign n5888 = ( n5829 & ~n5854 ) | ( n5829 & n5878 ) | ( ~n5854 & n5878 ) ;
  assign n5889 = ~n5887 & n5888 ;
  assign n5890 = n5883 | n5889 ;
  assign n5891 = n5724 &  n5855 ;
  assign n5884 = x76 | n5724 ;
  assign n5885 = x76 &  n5724 ;
  assign n5886 = ( n5884 & ~n5885 ) | ( n5884 & 1'b0 ) | ( ~n5885 & 1'b0 ) ;
  assign n5895 = ( n5828 & n5851 ) | ( n5828 & n5886 ) | ( n5851 & n5886 ) ;
  assign n5896 = ( n5828 & ~n5854 ) | ( n5828 & n5886 ) | ( ~n5854 & n5886 ) ;
  assign n5897 = ~n5895 & n5896 ;
  assign n5898 = n5891 | n5897 ;
  assign n5899 = n5732 &  n5855 ;
  assign n5892 = x75 | n5732 ;
  assign n5893 = x75 &  n5732 ;
  assign n5894 = ( n5892 & ~n5893 ) | ( n5892 & 1'b0 ) | ( ~n5893 & 1'b0 ) ;
  assign n5903 = ( n5827 & n5851 ) | ( n5827 & n5894 ) | ( n5851 & n5894 ) ;
  assign n5904 = ( n5827 & ~n5854 ) | ( n5827 & n5894 ) | ( ~n5854 & n5894 ) ;
  assign n5905 = ~n5903 & n5904 ;
  assign n5906 = n5899 | n5905 ;
  assign n5907 = n5740 &  n5855 ;
  assign n5900 = x74 | n5740 ;
  assign n5901 = x74 &  n5740 ;
  assign n5902 = ( n5900 & ~n5901 ) | ( n5900 & 1'b0 ) | ( ~n5901 & 1'b0 ) ;
  assign n5911 = ( n5826 & n5851 ) | ( n5826 & n5902 ) | ( n5851 & n5902 ) ;
  assign n5912 = ( n5826 & ~n5854 ) | ( n5826 & n5902 ) | ( ~n5854 & n5902 ) ;
  assign n5913 = ~n5911 & n5912 ;
  assign n5914 = n5907 | n5913 ;
  assign n5915 = n5748 &  n5855 ;
  assign n5908 = x73 | n5748 ;
  assign n5909 = x73 &  n5748 ;
  assign n5910 = ( n5908 & ~n5909 ) | ( n5908 & 1'b0 ) | ( ~n5909 & 1'b0 ) ;
  assign n5919 = ( n5825 & n5851 ) | ( n5825 & n5910 ) | ( n5851 & n5910 ) ;
  assign n5920 = ( n5825 & ~n5854 ) | ( n5825 & n5910 ) | ( ~n5854 & n5910 ) ;
  assign n5921 = ~n5919 & n5920 ;
  assign n5922 = n5915 | n5921 ;
  assign n5923 = n5756 &  n5855 ;
  assign n5916 = x72 | n5756 ;
  assign n5917 = x72 &  n5756 ;
  assign n5918 = ( n5916 & ~n5917 ) | ( n5916 & 1'b0 ) | ( ~n5917 & 1'b0 ) ;
  assign n5927 = ( n5824 & n5851 ) | ( n5824 & n5918 ) | ( n5851 & n5918 ) ;
  assign n5928 = ( n5824 & ~n5854 ) | ( n5824 & n5918 ) | ( ~n5854 & n5918 ) ;
  assign n5929 = ~n5927 & n5928 ;
  assign n5930 = n5923 | n5929 ;
  assign n5931 = n5764 &  n5855 ;
  assign n5924 = x71 | n5764 ;
  assign n5925 = x71 &  n5764 ;
  assign n5926 = ( n5924 & ~n5925 ) | ( n5924 & 1'b0 ) | ( ~n5925 & 1'b0 ) ;
  assign n5935 = ( n5823 & n5851 ) | ( n5823 & n5926 ) | ( n5851 & n5926 ) ;
  assign n5936 = ( n5823 & ~n5854 ) | ( n5823 & n5926 ) | ( ~n5854 & n5926 ) ;
  assign n5937 = ~n5935 & n5936 ;
  assign n5938 = n5931 | n5937 ;
  assign n5939 = n5772 &  n5855 ;
  assign n5932 = x70 | n5772 ;
  assign n5933 = x70 &  n5772 ;
  assign n5934 = ( n5932 & ~n5933 ) | ( n5932 & 1'b0 ) | ( ~n5933 & 1'b0 ) ;
  assign n5943 = ( n5822 & n5851 ) | ( n5822 & n5934 ) | ( n5851 & n5934 ) ;
  assign n5944 = ( n5822 & ~n5854 ) | ( n5822 & n5934 ) | ( ~n5854 & n5934 ) ;
  assign n5945 = ~n5943 & n5944 ;
  assign n5946 = n5939 | n5945 ;
  assign n5947 = n5780 &  n5855 ;
  assign n5940 = x69 | n5780 ;
  assign n5941 = x69 &  n5780 ;
  assign n5942 = ( n5940 & ~n5941 ) | ( n5940 & 1'b0 ) | ( ~n5941 & 1'b0 ) ;
  assign n5951 = ( n5821 & n5851 ) | ( n5821 & n5942 ) | ( n5851 & n5942 ) ;
  assign n5952 = ( n5821 & ~n5854 ) | ( n5821 & n5942 ) | ( ~n5854 & n5942 ) ;
  assign n5953 = ~n5951 & n5952 ;
  assign n5954 = n5947 | n5953 ;
  assign n5955 = n5788 &  n5855 ;
  assign n5948 = x68 | n5788 ;
  assign n5949 = x68 &  n5788 ;
  assign n5950 = ( n5948 & ~n5949 ) | ( n5948 & 1'b0 ) | ( ~n5949 & 1'b0 ) ;
  assign n5959 = ( n5820 & n5851 ) | ( n5820 & n5950 ) | ( n5851 & n5950 ) ;
  assign n5960 = ( n5820 & ~n5854 ) | ( n5820 & n5950 ) | ( ~n5854 & n5950 ) ;
  assign n5961 = ~n5959 & n5960 ;
  assign n5962 = n5955 | n5961 ;
  assign n5963 = n5797 &  n5855 ;
  assign n5956 = x67 | n5797 ;
  assign n5957 = x67 &  n5797 ;
  assign n5958 = ( n5956 & ~n5957 ) | ( n5956 & 1'b0 ) | ( ~n5957 & 1'b0 ) ;
  assign n5967 = ( n5819 & n5851 ) | ( n5819 & n5958 ) | ( n5851 & n5958 ) ;
  assign n5968 = ( n5819 & ~n5854 ) | ( n5819 & n5958 ) | ( ~n5854 & n5958 ) ;
  assign n5969 = ~n5967 & n5968 ;
  assign n5970 = n5963 | n5969 ;
  assign n5971 = n5803 &  n5855 ;
  assign n5964 = x66 | n5803 ;
  assign n5965 = x66 &  n5803 ;
  assign n5966 = ( n5964 & ~n5965 ) | ( n5964 & 1'b0 ) | ( ~n5965 & 1'b0 ) ;
  assign n5976 = ( n5818 & ~n5851 ) | ( n5818 & n5966 ) | ( ~n5851 & n5966 ) ;
  assign n5977 = ( n5818 & n5854 ) | ( n5818 & n5966 ) | ( n5854 & n5966 ) ;
  assign n5978 = ( n5976 & ~n5977 ) | ( n5976 & 1'b0 ) | ( ~n5977 & 1'b0 ) ;
  assign n5979 = n5971 | n5978 ;
  assign n5980 = n5816 &  n5855 ;
  assign n5972 = x65 &  n5816 ;
  assign n5973 = x65 | n5815 ;
  assign n5974 = n5810 | n5973 ;
  assign n5975 = ( n5817 & ~n5972 ) | ( n5817 & n5974 ) | ( ~n5972 & n5974 ) ;
  assign n5981 = ( x65 & n5816 ) | ( x65 & n5817 ) | ( n5816 & n5817 ) ;
  assign n5982 = ( n5854 & ~n5972 ) | ( n5854 & n5981 ) | ( ~n5972 & n5981 ) ;
  assign n5983 = ( n5851 & n5975 ) | ( n5851 & n5982 ) | ( n5975 & n5982 ) ;
  assign n5984 = ( n5975 & ~n5983 ) | ( n5975 & 1'b0 ) | ( ~n5983 & 1'b0 ) ;
  assign n5985 = n5980 | n5984 ;
  assign n5986 = ( x64 & ~x99 ) | ( x64 & 1'b0 ) | ( ~x99 & 1'b0 ) ;
  assign n5987 = ( n166 & ~n272 ) | ( n166 & n5986 ) | ( ~n272 & n5986 ) ;
  assign n5988 = ~n166 & n5987 ;
  assign n5989 = ~n270 & n5988 ;
  assign n5990 = n5851 &  n5989 ;
  assign n5991 = ( x29 & ~n5989 ) | ( x29 & n5990 ) | ( ~n5989 & n5990 ) ;
  assign n5992 = ~n245 & n5817 ;
  assign n5993 = ( n243 & ~n254 ) | ( n243 & n5992 ) | ( ~n254 & n5992 ) ;
  assign n5994 = ~n243 & n5993 ;
  assign n5995 = ~n240 & n5994 ;
  assign n5996 = ~n5851 & n5995 ;
  assign n5997 = n5991 | n5996 ;
  assign n5998 = ~x28 & x64 ;
  assign n5999 = ( x65 & ~n5997 ) | ( x65 & n5998 ) | ( ~n5997 & n5998 ) ;
  assign n6000 = ( x66 & ~n5985 ) | ( x66 & n5999 ) | ( ~n5985 & n5999 ) ;
  assign n6001 = ( x67 & ~n5979 ) | ( x67 & n6000 ) | ( ~n5979 & n6000 ) ;
  assign n6002 = ( x68 & ~n5970 ) | ( x68 & n6001 ) | ( ~n5970 & n6001 ) ;
  assign n6003 = ( x69 & ~n5962 ) | ( x69 & n6002 ) | ( ~n5962 & n6002 ) ;
  assign n6004 = ( x70 & ~n5954 ) | ( x70 & n6003 ) | ( ~n5954 & n6003 ) ;
  assign n6005 = ( x71 & ~n5946 ) | ( x71 & n6004 ) | ( ~n5946 & n6004 ) ;
  assign n6006 = ( x72 & ~n5938 ) | ( x72 & n6005 ) | ( ~n5938 & n6005 ) ;
  assign n6007 = ( x73 & ~n5930 ) | ( x73 & n6006 ) | ( ~n5930 & n6006 ) ;
  assign n6008 = ( x74 & ~n5922 ) | ( x74 & n6007 ) | ( ~n5922 & n6007 ) ;
  assign n6009 = ( x75 & ~n5914 ) | ( x75 & n6008 ) | ( ~n5914 & n6008 ) ;
  assign n6010 = ( x76 & ~n5906 ) | ( x76 & n6009 ) | ( ~n5906 & n6009 ) ;
  assign n6011 = ( x77 & ~n5898 ) | ( x77 & n6010 ) | ( ~n5898 & n6010 ) ;
  assign n6012 = ( x78 & ~n5890 ) | ( x78 & n6011 ) | ( ~n5890 & n6011 ) ;
  assign n6013 = ( x79 & ~n5882 ) | ( x79 & n6012 ) | ( ~n5882 & n6012 ) ;
  assign n6014 = ( x80 & ~n5874 ) | ( x80 & n6013 ) | ( ~n5874 & n6013 ) ;
  assign n6018 = ( x81 & ~n5866 ) | ( x81 & n6014 ) | ( ~n5866 & n6014 ) ;
  assign n6158 = ( x82 & ~n6026 ) | ( x82 & n6018 ) | ( ~n6026 & n6018 ) ;
  assign n6159 = ( x83 & ~n6157 ) | ( x83 & n6158 ) | ( ~n6157 & n6158 ) ;
  assign n6160 = ( x84 & ~n6152 ) | ( x84 & n6159 ) | ( ~n6152 & n6159 ) ;
  assign n6161 = ( x85 & ~n6144 ) | ( x85 & n6160 ) | ( ~n6144 & n6160 ) ;
  assign n6162 = ( x86 & ~n6136 ) | ( x86 & n6161 ) | ( ~n6136 & n6161 ) ;
  assign n6163 = ( x87 & ~n6128 ) | ( x87 & n6162 ) | ( ~n6128 & n6162 ) ;
  assign n6164 = ( x88 & ~n6120 ) | ( x88 & n6163 ) | ( ~n6120 & n6163 ) ;
  assign n6165 = ( x89 & ~n6112 ) | ( x89 & n6164 ) | ( ~n6112 & n6164 ) ;
  assign n6166 = ( x90 & ~n6104 ) | ( x90 & n6165 ) | ( ~n6104 & n6165 ) ;
  assign n6167 = ( x91 & ~n6096 ) | ( x91 & n6166 ) | ( ~n6096 & n6166 ) ;
  assign n6168 = ( x92 & ~n6088 ) | ( x92 & n6167 ) | ( ~n6088 & n6167 ) ;
  assign n6169 = ( x93 & ~n6080 ) | ( x93 & n6168 ) | ( ~n6080 & n6168 ) ;
  assign n6170 = ( x94 & ~n6072 ) | ( x94 & n6169 ) | ( ~n6072 & n6169 ) ;
  assign n6171 = ( x95 & ~n6064 ) | ( x95 & n6170 ) | ( ~n6064 & n6170 ) ;
  assign n6172 = ( x96 & ~n6056 ) | ( x96 & n6171 ) | ( ~n6056 & n6171 ) ;
  assign n6173 = ( x97 & ~n6048 ) | ( x97 & n6172 ) | ( ~n6048 & n6172 ) ;
  assign n6174 = ( x98 & ~n6040 ) | ( x98 & n6173 ) | ( ~n6040 & n6173 ) ;
  assign n6175 = n5559 &  n5855 ;
  assign n6176 = ( n5559 & ~n5854 ) | ( n5559 & n5850 ) | ( ~n5854 & n5850 ) ;
  assign n6177 = ( x98 & ~n5850 ) | ( x98 & n6176 ) | ( ~n5850 & n6176 ) ;
  assign n6178 = ~x98 & n6177 ;
  assign n6179 = n6175 | n6178 ;
  assign n6180 = ~x99 & n6179 ;
  assign n6181 = ( x99 & ~n6175 ) | ( x99 & 1'b0 ) | ( ~n6175 & 1'b0 ) ;
  assign n6182 = ~n6178 & n6181 ;
  assign n6183 = n356 | n6182 ;
  assign n6184 = n6180 | n6183 ;
  assign n6185 = n6174 | n6184 ;
  assign n6186 = ~n6179 |  n5854 ;
  assign n6205 = n6040 &  n6186 ;
  assign n6206 = n6185 &  n6205 ;
  assign n6193 = x98 | n6040 ;
  assign n6194 = x98 &  n6040 ;
  assign n6195 = ( n6193 & ~n6194 ) | ( n6193 & 1'b0 ) | ( ~n6194 & 1'b0 ) ;
  assign n6207 = n6173 &  n6195 ;
  assign n6187 = n6185 &  n6186 ;
  assign n6208 = ( n6173 & ~n6187 ) | ( n6173 & n6195 ) | ( ~n6187 & n6195 ) ;
  assign n6209 = ( n6206 & ~n6207 ) | ( n6206 & n6208 ) | ( ~n6207 & n6208 ) ;
  assign n6197 = n5559 &  n5854 ;
  assign n6198 = n6185 &  n6197 ;
  assign n6196 = n6180 | n6182 ;
  assign n6200 = ( n6174 & n6187 ) | ( n6174 & n6196 ) | ( n6187 & n6196 ) ;
  assign n6199 = n6174 | n6196 ;
  assign n6201 = ( n6198 & ~n6200 ) | ( n6198 & n6199 ) | ( ~n6200 & n6199 ) ;
  assign n6213 = n6048 &  n6186 ;
  assign n6214 = n6185 &  n6213 ;
  assign n6202 = x97 | n6048 ;
  assign n6203 = x97 &  n6048 ;
  assign n6204 = ( n6202 & ~n6203 ) | ( n6202 & 1'b0 ) | ( ~n6203 & 1'b0 ) ;
  assign n6215 = n6172 &  n6204 ;
  assign n6216 = ( n6172 & ~n6187 ) | ( n6172 & n6204 ) | ( ~n6187 & n6204 ) ;
  assign n6217 = ( n6214 & ~n6215 ) | ( n6214 & n6216 ) | ( ~n6215 & n6216 ) ;
  assign n6221 = n6056 &  n6186 ;
  assign n6222 = n6185 &  n6221 ;
  assign n6210 = x96 | n6056 ;
  assign n6211 = x96 &  n6056 ;
  assign n6212 = ( n6210 & ~n6211 ) | ( n6210 & 1'b0 ) | ( ~n6211 & 1'b0 ) ;
  assign n6223 = n6171 &  n6212 ;
  assign n6224 = ( n6171 & ~n6187 ) | ( n6171 & n6212 ) | ( ~n6187 & n6212 ) ;
  assign n6225 = ( n6222 & ~n6223 ) | ( n6222 & n6224 ) | ( ~n6223 & n6224 ) ;
  assign n6229 = n6064 &  n6186 ;
  assign n6230 = n6185 &  n6229 ;
  assign n6218 = x95 | n6064 ;
  assign n6219 = x95 &  n6064 ;
  assign n6220 = ( n6218 & ~n6219 ) | ( n6218 & 1'b0 ) | ( ~n6219 & 1'b0 ) ;
  assign n6231 = n6170 &  n6220 ;
  assign n6232 = ( n6170 & ~n6187 ) | ( n6170 & n6220 ) | ( ~n6187 & n6220 ) ;
  assign n6233 = ( n6230 & ~n6231 ) | ( n6230 & n6232 ) | ( ~n6231 & n6232 ) ;
  assign n6237 = n6072 &  n6186 ;
  assign n6238 = n6185 &  n6237 ;
  assign n6226 = x94 | n6072 ;
  assign n6227 = x94 &  n6072 ;
  assign n6228 = ( n6226 & ~n6227 ) | ( n6226 & 1'b0 ) | ( ~n6227 & 1'b0 ) ;
  assign n6239 = n6169 &  n6228 ;
  assign n6240 = ( n6169 & ~n6187 ) | ( n6169 & n6228 ) | ( ~n6187 & n6228 ) ;
  assign n6241 = ( n6238 & ~n6239 ) | ( n6238 & n6240 ) | ( ~n6239 & n6240 ) ;
  assign n6245 = n6080 &  n6186 ;
  assign n6246 = n6185 &  n6245 ;
  assign n6234 = x93 | n6080 ;
  assign n6235 = x93 &  n6080 ;
  assign n6236 = ( n6234 & ~n6235 ) | ( n6234 & 1'b0 ) | ( ~n6235 & 1'b0 ) ;
  assign n6248 = ( n6168 & n6187 ) | ( n6168 & n6236 ) | ( n6187 & n6236 ) ;
  assign n6247 = n6168 | n6236 ;
  assign n6249 = ( n6246 & ~n6248 ) | ( n6246 & n6247 ) | ( ~n6248 & n6247 ) ;
  assign n6253 = n6088 &  n6186 ;
  assign n6254 = n6185 &  n6253 ;
  assign n6242 = x92 | n6088 ;
  assign n6243 = x92 &  n6088 ;
  assign n6244 = ( n6242 & ~n6243 ) | ( n6242 & 1'b0 ) | ( ~n6243 & 1'b0 ) ;
  assign n6256 = ( n6167 & n6187 ) | ( n6167 & n6244 ) | ( n6187 & n6244 ) ;
  assign n6255 = n6167 | n6244 ;
  assign n6257 = ( n6254 & ~n6256 ) | ( n6254 & n6255 ) | ( ~n6256 & n6255 ) ;
  assign n6261 = n6096 &  n6186 ;
  assign n6262 = n6185 &  n6261 ;
  assign n6250 = x91 | n6096 ;
  assign n6251 = x91 &  n6096 ;
  assign n6252 = ( n6250 & ~n6251 ) | ( n6250 & 1'b0 ) | ( ~n6251 & 1'b0 ) ;
  assign n6264 = ( n6166 & n6187 ) | ( n6166 & n6252 ) | ( n6187 & n6252 ) ;
  assign n6263 = n6166 | n6252 ;
  assign n6265 = ( n6262 & ~n6264 ) | ( n6262 & n6263 ) | ( ~n6264 & n6263 ) ;
  assign n6269 = n6104 &  n6186 ;
  assign n6270 = n6185 &  n6269 ;
  assign n6258 = x90 | n6104 ;
  assign n6259 = x90 &  n6104 ;
  assign n6260 = ( n6258 & ~n6259 ) | ( n6258 & 1'b0 ) | ( ~n6259 & 1'b0 ) ;
  assign n6272 = ( n6165 & n6187 ) | ( n6165 & n6260 ) | ( n6187 & n6260 ) ;
  assign n6271 = n6165 | n6260 ;
  assign n6273 = ( n6270 & ~n6272 ) | ( n6270 & n6271 ) | ( ~n6272 & n6271 ) ;
  assign n6277 = n6112 &  n6186 ;
  assign n6278 = n6185 &  n6277 ;
  assign n6266 = x89 | n6112 ;
  assign n6267 = x89 &  n6112 ;
  assign n6268 = ( n6266 & ~n6267 ) | ( n6266 & 1'b0 ) | ( ~n6267 & 1'b0 ) ;
  assign n6280 = ( n6164 & n6187 ) | ( n6164 & n6268 ) | ( n6187 & n6268 ) ;
  assign n6279 = n6164 | n6268 ;
  assign n6281 = ( n6278 & ~n6280 ) | ( n6278 & n6279 ) | ( ~n6280 & n6279 ) ;
  assign n6285 = n6120 &  n6186 ;
  assign n6286 = n6185 &  n6285 ;
  assign n6274 = x88 | n6120 ;
  assign n6275 = x88 &  n6120 ;
  assign n6276 = ( n6274 & ~n6275 ) | ( n6274 & 1'b0 ) | ( ~n6275 & 1'b0 ) ;
  assign n6288 = ( n6163 & n6187 ) | ( n6163 & n6276 ) | ( n6187 & n6276 ) ;
  assign n6287 = n6163 | n6276 ;
  assign n6289 = ( n6286 & ~n6288 ) | ( n6286 & n6287 ) | ( ~n6288 & n6287 ) ;
  assign n6293 = n6128 &  n6186 ;
  assign n6294 = n6185 &  n6293 ;
  assign n6282 = x87 | n6128 ;
  assign n6283 = x87 &  n6128 ;
  assign n6284 = ( n6282 & ~n6283 ) | ( n6282 & 1'b0 ) | ( ~n6283 & 1'b0 ) ;
  assign n6296 = ( n6162 & n6187 ) | ( n6162 & n6284 ) | ( n6187 & n6284 ) ;
  assign n6295 = n6162 | n6284 ;
  assign n6297 = ( n6294 & ~n6296 ) | ( n6294 & n6295 ) | ( ~n6296 & n6295 ) ;
  assign n6301 = n6136 &  n6186 ;
  assign n6302 = n6185 &  n6301 ;
  assign n6290 = x86 | n6136 ;
  assign n6291 = x86 &  n6136 ;
  assign n6292 = ( n6290 & ~n6291 ) | ( n6290 & 1'b0 ) | ( ~n6291 & 1'b0 ) ;
  assign n6304 = ( n6161 & n6187 ) | ( n6161 & n6292 ) | ( n6187 & n6292 ) ;
  assign n6303 = n6161 | n6292 ;
  assign n6305 = ( n6302 & ~n6304 ) | ( n6302 & n6303 ) | ( ~n6304 & n6303 ) ;
  assign n6309 = n6144 &  n6186 ;
  assign n6310 = n6185 &  n6309 ;
  assign n6298 = x85 | n6144 ;
  assign n6299 = x85 &  n6144 ;
  assign n6300 = ( n6298 & ~n6299 ) | ( n6298 & 1'b0 ) | ( ~n6299 & 1'b0 ) ;
  assign n6312 = ( n6160 & n6187 ) | ( n6160 & n6300 ) | ( n6187 & n6300 ) ;
  assign n6311 = n6160 | n6300 ;
  assign n6313 = ( n6310 & ~n6312 ) | ( n6310 & n6311 ) | ( ~n6312 & n6311 ) ;
  assign n6317 = n6152 &  n6186 ;
  assign n6318 = n6185 &  n6317 ;
  assign n6306 = x84 | n6152 ;
  assign n6307 = x84 &  n6152 ;
  assign n6308 = ( n6306 & ~n6307 ) | ( n6306 & 1'b0 ) | ( ~n6307 & 1'b0 ) ;
  assign n6320 = ( n6159 & n6187 ) | ( n6159 & n6308 ) | ( n6187 & n6308 ) ;
  assign n6319 = n6159 | n6308 ;
  assign n6321 = ( n6318 & ~n6320 ) | ( n6318 & n6319 ) | ( ~n6320 & n6319 ) ;
  assign n6322 = n6157 &  n6186 ;
  assign n6323 = n6185 &  n6322 ;
  assign n6314 = x83 | n6157 ;
  assign n6315 = x83 &  n6157 ;
  assign n6316 = ( n6314 & ~n6315 ) | ( n6314 & 1'b0 ) | ( ~n6315 & 1'b0 ) ;
  assign n6325 = ( n6158 & n6187 ) | ( n6158 & n6316 ) | ( n6187 & n6316 ) ;
  assign n6324 = n6158 | n6316 ;
  assign n6326 = ( n6323 & ~n6325 ) | ( n6323 & n6324 ) | ( ~n6325 & n6324 ) ;
  assign n6188 = n6026 &  n6186 ;
  assign n6189 = n6185 &  n6188 ;
  assign n6027 = x82 | n6026 ;
  assign n6028 = x82 &  n6026 ;
  assign n6029 = ( n6027 & ~n6028 ) | ( n6027 & 1'b0 ) | ( ~n6028 & 1'b0 ) ;
  assign n6191 = ( n6018 & n6029 ) | ( n6018 & n6187 ) | ( n6029 & n6187 ) ;
  assign n6190 = n6018 | n6029 ;
  assign n6192 = ( n6189 & ~n6191 ) | ( n6189 & n6190 ) | ( ~n6191 & n6190 ) ;
  assign n6330 = n5866 &  n6186 ;
  assign n6331 = n6185 &  n6330 ;
  assign n6015 = x81 | n5866 ;
  assign n6016 = x81 &  n5866 ;
  assign n6017 = ( n6015 & ~n6016 ) | ( n6015 & 1'b0 ) | ( ~n6016 & 1'b0 ) ;
  assign n6332 = n6014 &  n6017 ;
  assign n6333 = ( n6014 & ~n6187 ) | ( n6014 & n6017 ) | ( ~n6187 & n6017 ) ;
  assign n6334 = ( n6331 & ~n6332 ) | ( n6331 & n6333 ) | ( ~n6332 & n6333 ) ;
  assign n6338 = n5874 &  n6186 ;
  assign n6339 = n6185 &  n6338 ;
  assign n6327 = x80 | n5874 ;
  assign n6328 = x80 &  n5874 ;
  assign n6329 = ( n6327 & ~n6328 ) | ( n6327 & 1'b0 ) | ( ~n6328 & 1'b0 ) ;
  assign n6341 = ( n6013 & n6187 ) | ( n6013 & n6329 ) | ( n6187 & n6329 ) ;
  assign n6340 = n6013 | n6329 ;
  assign n6342 = ( n6339 & ~n6341 ) | ( n6339 & n6340 ) | ( ~n6341 & n6340 ) ;
  assign n6346 = n5882 &  n6186 ;
  assign n6347 = n6185 &  n6346 ;
  assign n6335 = x79 | n5882 ;
  assign n6336 = x79 &  n5882 ;
  assign n6337 = ( n6335 & ~n6336 ) | ( n6335 & 1'b0 ) | ( ~n6336 & 1'b0 ) ;
  assign n6349 = ( n6012 & n6187 ) | ( n6012 & n6337 ) | ( n6187 & n6337 ) ;
  assign n6348 = n6012 | n6337 ;
  assign n6350 = ( n6347 & ~n6349 ) | ( n6347 & n6348 ) | ( ~n6349 & n6348 ) ;
  assign n6354 = n5890 &  n6186 ;
  assign n6355 = n6185 &  n6354 ;
  assign n6343 = x78 | n5890 ;
  assign n6344 = x78 &  n5890 ;
  assign n6345 = ( n6343 & ~n6344 ) | ( n6343 & 1'b0 ) | ( ~n6344 & 1'b0 ) ;
  assign n6357 = ( n6011 & n6187 ) | ( n6011 & n6345 ) | ( n6187 & n6345 ) ;
  assign n6356 = n6011 | n6345 ;
  assign n6358 = ( n6355 & ~n6357 ) | ( n6355 & n6356 ) | ( ~n6357 & n6356 ) ;
  assign n6362 = n5898 &  n6186 ;
  assign n6363 = n6185 &  n6362 ;
  assign n6351 = x77 | n5898 ;
  assign n6352 = x77 &  n5898 ;
  assign n6353 = ( n6351 & ~n6352 ) | ( n6351 & 1'b0 ) | ( ~n6352 & 1'b0 ) ;
  assign n6365 = ( n6010 & n6187 ) | ( n6010 & n6353 ) | ( n6187 & n6353 ) ;
  assign n6364 = n6010 | n6353 ;
  assign n6366 = ( n6363 & ~n6365 ) | ( n6363 & n6364 ) | ( ~n6365 & n6364 ) ;
  assign n6370 = n5906 &  n6186 ;
  assign n6371 = n6185 &  n6370 ;
  assign n6359 = x76 | n5906 ;
  assign n6360 = x76 &  n5906 ;
  assign n6361 = ( n6359 & ~n6360 ) | ( n6359 & 1'b0 ) | ( ~n6360 & 1'b0 ) ;
  assign n6373 = ( n6009 & n6187 ) | ( n6009 & n6361 ) | ( n6187 & n6361 ) ;
  assign n6372 = n6009 | n6361 ;
  assign n6374 = ( n6371 & ~n6373 ) | ( n6371 & n6372 ) | ( ~n6373 & n6372 ) ;
  assign n6378 = n5914 &  n6186 ;
  assign n6379 = n6185 &  n6378 ;
  assign n6367 = x75 | n5914 ;
  assign n6368 = x75 &  n5914 ;
  assign n6369 = ( n6367 & ~n6368 ) | ( n6367 & 1'b0 ) | ( ~n6368 & 1'b0 ) ;
  assign n6381 = ( n6008 & n6187 ) | ( n6008 & n6369 ) | ( n6187 & n6369 ) ;
  assign n6380 = n6008 | n6369 ;
  assign n6382 = ( n6379 & ~n6381 ) | ( n6379 & n6380 ) | ( ~n6381 & n6380 ) ;
  assign n6386 = n5922 &  n6186 ;
  assign n6387 = n6185 &  n6386 ;
  assign n6375 = x74 | n5922 ;
  assign n6376 = x74 &  n5922 ;
  assign n6377 = ( n6375 & ~n6376 ) | ( n6375 & 1'b0 ) | ( ~n6376 & 1'b0 ) ;
  assign n6389 = ( n6007 & n6187 ) | ( n6007 & n6377 ) | ( n6187 & n6377 ) ;
  assign n6388 = n6007 | n6377 ;
  assign n6390 = ( n6387 & ~n6389 ) | ( n6387 & n6388 ) | ( ~n6389 & n6388 ) ;
  assign n6394 = n5930 &  n6186 ;
  assign n6395 = n6185 &  n6394 ;
  assign n6383 = x73 | n5930 ;
  assign n6384 = x73 &  n5930 ;
  assign n6385 = ( n6383 & ~n6384 ) | ( n6383 & 1'b0 ) | ( ~n6384 & 1'b0 ) ;
  assign n6397 = ( n6006 & n6187 ) | ( n6006 & n6385 ) | ( n6187 & n6385 ) ;
  assign n6396 = n6006 | n6385 ;
  assign n6398 = ( n6395 & ~n6397 ) | ( n6395 & n6396 ) | ( ~n6397 & n6396 ) ;
  assign n6402 = n5938 &  n6186 ;
  assign n6403 = n6185 &  n6402 ;
  assign n6391 = x72 | n5938 ;
  assign n6392 = x72 &  n5938 ;
  assign n6393 = ( n6391 & ~n6392 ) | ( n6391 & 1'b0 ) | ( ~n6392 & 1'b0 ) ;
  assign n6405 = ( n6005 & n6187 ) | ( n6005 & n6393 ) | ( n6187 & n6393 ) ;
  assign n6404 = n6005 | n6393 ;
  assign n6406 = ( n6403 & ~n6405 ) | ( n6403 & n6404 ) | ( ~n6405 & n6404 ) ;
  assign n6410 = n5946 &  n6186 ;
  assign n6411 = n6185 &  n6410 ;
  assign n6399 = x71 | n5946 ;
  assign n6400 = x71 &  n5946 ;
  assign n6401 = ( n6399 & ~n6400 ) | ( n6399 & 1'b0 ) | ( ~n6400 & 1'b0 ) ;
  assign n6413 = ( n6004 & n6187 ) | ( n6004 & n6401 ) | ( n6187 & n6401 ) ;
  assign n6412 = n6004 | n6401 ;
  assign n6414 = ( n6411 & ~n6413 ) | ( n6411 & n6412 ) | ( ~n6413 & n6412 ) ;
  assign n6418 = n5954 &  n6186 ;
  assign n6419 = n6185 &  n6418 ;
  assign n6407 = x70 | n5954 ;
  assign n6408 = x70 &  n5954 ;
  assign n6409 = ( n6407 & ~n6408 ) | ( n6407 & 1'b0 ) | ( ~n6408 & 1'b0 ) ;
  assign n6421 = ( n6003 & n6187 ) | ( n6003 & n6409 ) | ( n6187 & n6409 ) ;
  assign n6420 = n6003 | n6409 ;
  assign n6422 = ( n6419 & ~n6421 ) | ( n6419 & n6420 ) | ( ~n6421 & n6420 ) ;
  assign n6426 = n5962 &  n6186 ;
  assign n6427 = n6185 &  n6426 ;
  assign n6415 = x69 | n5962 ;
  assign n6416 = x69 &  n5962 ;
  assign n6417 = ( n6415 & ~n6416 ) | ( n6415 & 1'b0 ) | ( ~n6416 & 1'b0 ) ;
  assign n6429 = ( n6002 & n6187 ) | ( n6002 & n6417 ) | ( n6187 & n6417 ) ;
  assign n6428 = n6002 | n6417 ;
  assign n6430 = ( n6427 & ~n6429 ) | ( n6427 & n6428 ) | ( ~n6429 & n6428 ) ;
  assign n6434 = n5970 &  n6186 ;
  assign n6435 = n6185 &  n6434 ;
  assign n6423 = x68 | n5970 ;
  assign n6424 = x68 &  n5970 ;
  assign n6425 = ( n6423 & ~n6424 ) | ( n6423 & 1'b0 ) | ( ~n6424 & 1'b0 ) ;
  assign n6437 = ( n6001 & n6187 ) | ( n6001 & n6425 ) | ( n6187 & n6425 ) ;
  assign n6436 = n6001 | n6425 ;
  assign n6438 = ( n6435 & ~n6437 ) | ( n6435 & n6436 ) | ( ~n6437 & n6436 ) ;
  assign n6442 = n5979 &  n6186 ;
  assign n6443 = n6185 &  n6442 ;
  assign n6431 = x67 | n5979 ;
  assign n6432 = x67 &  n5979 ;
  assign n6433 = ( n6431 & ~n6432 ) | ( n6431 & 1'b0 ) | ( ~n6432 & 1'b0 ) ;
  assign n6445 = ( n6000 & n6187 ) | ( n6000 & n6433 ) | ( n6187 & n6433 ) ;
  assign n6444 = n6000 | n6433 ;
  assign n6446 = ( n6443 & ~n6445 ) | ( n6443 & n6444 ) | ( ~n6445 & n6444 ) ;
  assign n6447 = n5985 &  n6186 ;
  assign n6448 = n6185 &  n6447 ;
  assign n6439 = x66 | n5985 ;
  assign n6440 = x66 &  n5985 ;
  assign n6441 = ( n6439 & ~n6440 ) | ( n6439 & 1'b0 ) | ( ~n6440 & 1'b0 ) ;
  assign n6449 = n5999 &  n6441 ;
  assign n6450 = ( n5999 & ~n6187 ) | ( n5999 & n6441 ) | ( ~n6187 & n6441 ) ;
  assign n6451 = ( n6448 & ~n6449 ) | ( n6448 & n6450 ) | ( ~n6449 & n6450 ) ;
  assign n6452 = ( n5997 & ~x65 ) | ( n5997 & n5998 ) | ( ~x65 & n5998 ) ;
  assign n6453 = ( n5999 & ~n5998 ) | ( n5999 & n6452 ) | ( ~n5998 & n6452 ) ;
  assign n6454 = ~n6187 & n6453 ;
  assign n6455 = n5997 &  n6186 ;
  assign n6456 = n6185 &  n6455 ;
  assign n6457 = n6454 | n6456 ;
  assign n6458 = ( x64 & ~n6187 ) | ( x64 & 1'b0 ) | ( ~n6187 & 1'b0 ) ;
  assign n6459 = ( x28 & ~n6458 ) | ( x28 & 1'b0 ) | ( ~n6458 & 1'b0 ) ;
  assign n6460 = ( n5998 & ~n6187 ) | ( n5998 & 1'b0 ) | ( ~n6187 & 1'b0 ) ;
  assign n6461 = n6459 | n6460 ;
  assign n6462 = ~x27 & x64 ;
  assign n6463 = ( x65 & ~n6461 ) | ( x65 & n6462 ) | ( ~n6461 & n6462 ) ;
  assign n6464 = ( x66 & ~n6457 ) | ( x66 & n6463 ) | ( ~n6457 & n6463 ) ;
  assign n6465 = ( x67 & ~n6451 ) | ( x67 & n6464 ) | ( ~n6451 & n6464 ) ;
  assign n6466 = ( x68 & ~n6446 ) | ( x68 & n6465 ) | ( ~n6446 & n6465 ) ;
  assign n6467 = ( x69 & ~n6438 ) | ( x69 & n6466 ) | ( ~n6438 & n6466 ) ;
  assign n6468 = ( x70 & ~n6430 ) | ( x70 & n6467 ) | ( ~n6430 & n6467 ) ;
  assign n6469 = ( x71 & ~n6422 ) | ( x71 & n6468 ) | ( ~n6422 & n6468 ) ;
  assign n6470 = ( x72 & ~n6414 ) | ( x72 & n6469 ) | ( ~n6414 & n6469 ) ;
  assign n6471 = ( x73 & ~n6406 ) | ( x73 & n6470 ) | ( ~n6406 & n6470 ) ;
  assign n6472 = ( x74 & ~n6398 ) | ( x74 & n6471 ) | ( ~n6398 & n6471 ) ;
  assign n6473 = ( x75 & ~n6390 ) | ( x75 & n6472 ) | ( ~n6390 & n6472 ) ;
  assign n6474 = ( x76 & ~n6382 ) | ( x76 & n6473 ) | ( ~n6382 & n6473 ) ;
  assign n6475 = ( x77 & ~n6374 ) | ( x77 & n6474 ) | ( ~n6374 & n6474 ) ;
  assign n6476 = ( x78 & ~n6366 ) | ( x78 & n6475 ) | ( ~n6366 & n6475 ) ;
  assign n6477 = ( x79 & ~n6358 ) | ( x79 & n6476 ) | ( ~n6358 & n6476 ) ;
  assign n6478 = ( x80 & ~n6350 ) | ( x80 & n6477 ) | ( ~n6350 & n6477 ) ;
  assign n6479 = ( x81 & ~n6342 ) | ( x81 & n6478 ) | ( ~n6342 & n6478 ) ;
  assign n6480 = ( x82 & ~n6334 ) | ( x82 & n6479 ) | ( ~n6334 & n6479 ) ;
  assign n6481 = ( x83 & ~n6192 ) | ( x83 & n6480 ) | ( ~n6192 & n6480 ) ;
  assign n6482 = ( x84 & ~n6326 ) | ( x84 & n6481 ) | ( ~n6326 & n6481 ) ;
  assign n6483 = ( x85 & ~n6321 ) | ( x85 & n6482 ) | ( ~n6321 & n6482 ) ;
  assign n6484 = ( x86 & ~n6313 ) | ( x86 & n6483 ) | ( ~n6313 & n6483 ) ;
  assign n6485 = ( x87 & ~n6305 ) | ( x87 & n6484 ) | ( ~n6305 & n6484 ) ;
  assign n6486 = ( x88 & ~n6297 ) | ( x88 & n6485 ) | ( ~n6297 & n6485 ) ;
  assign n6487 = ( x89 & ~n6289 ) | ( x89 & n6486 ) | ( ~n6289 & n6486 ) ;
  assign n6488 = ( x90 & ~n6281 ) | ( x90 & n6487 ) | ( ~n6281 & n6487 ) ;
  assign n6489 = ( x91 & ~n6273 ) | ( x91 & n6488 ) | ( ~n6273 & n6488 ) ;
  assign n6490 = ( x92 & ~n6265 ) | ( x92 & n6489 ) | ( ~n6265 & n6489 ) ;
  assign n6491 = ( x93 & ~n6257 ) | ( x93 & n6490 ) | ( ~n6257 & n6490 ) ;
  assign n6492 = ( x94 & ~n6249 ) | ( x94 & n6491 ) | ( ~n6249 & n6491 ) ;
  assign n6493 = ( x95 & ~n6241 ) | ( x95 & n6492 ) | ( ~n6241 & n6492 ) ;
  assign n6494 = ( x96 & ~n6233 ) | ( x96 & n6493 ) | ( ~n6233 & n6493 ) ;
  assign n6495 = ( x97 & ~n6225 ) | ( x97 & n6494 ) | ( ~n6225 & n6494 ) ;
  assign n6496 = ( x98 & ~n6217 ) | ( x98 & n6495 ) | ( ~n6217 & n6495 ) ;
  assign n6497 = ( x99 & ~n6209 ) | ( x99 & n6496 ) | ( ~n6209 & n6496 ) ;
  assign n6498 = ( x100 & ~n6201 ) | ( x100 & n6497 ) | ( ~n6201 & n6497 ) ;
  assign n6499 = n429 | n6498 ;
  assign n6517 = n6209 &  n6499 ;
  assign n6511 = x99 | n6209 ;
  assign n6512 = x99 &  n6209 ;
  assign n6513 = ( n6511 & ~n6512 ) | ( n6511 & 1'b0 ) | ( ~n6512 & 1'b0 ) ;
  assign n6521 = ( n429 & n6496 ) | ( n429 & n6513 ) | ( n6496 & n6513 ) ;
  assign n6522 = ( n6496 & ~n6498 ) | ( n6496 & n6513 ) | ( ~n6498 & n6513 ) ;
  assign n6523 = ~n6521 & n6522 ;
  assign n6524 = n6517 | n6523 ;
  assign n6515 = ( x100 & ~n429 ) | ( x100 & n6497 ) | ( ~n429 & n6497 ) ;
  assign n6514 = x100 &  n6497 ;
  assign n6516 = ( n6201 & ~n6515 ) | ( n6201 & n6514 ) | ( ~n6515 & n6514 ) ;
  assign n6525 = n6217 &  n6499 ;
  assign n6518 = x98 | n6217 ;
  assign n6519 = x98 &  n6217 ;
  assign n6520 = ( n6518 & ~n6519 ) | ( n6518 & 1'b0 ) | ( ~n6519 & 1'b0 ) ;
  assign n6529 = ( n429 & n6495 ) | ( n429 & n6520 ) | ( n6495 & n6520 ) ;
  assign n6530 = ( n6495 & ~n6498 ) | ( n6495 & n6520 ) | ( ~n6498 & n6520 ) ;
  assign n6531 = ~n6529 & n6530 ;
  assign n6532 = n6525 | n6531 ;
  assign n6533 = n6225 &  n6499 ;
  assign n6526 = x97 | n6225 ;
  assign n6527 = x97 &  n6225 ;
  assign n6528 = ( n6526 & ~n6527 ) | ( n6526 & 1'b0 ) | ( ~n6527 & 1'b0 ) ;
  assign n6537 = ( n429 & n6494 ) | ( n429 & n6528 ) | ( n6494 & n6528 ) ;
  assign n6538 = ( n6494 & ~n6498 ) | ( n6494 & n6528 ) | ( ~n6498 & n6528 ) ;
  assign n6539 = ~n6537 & n6538 ;
  assign n6540 = n6533 | n6539 ;
  assign n6541 = n6233 &  n6499 ;
  assign n6534 = x96 | n6233 ;
  assign n6535 = x96 &  n6233 ;
  assign n6536 = ( n6534 & ~n6535 ) | ( n6534 & 1'b0 ) | ( ~n6535 & 1'b0 ) ;
  assign n6545 = ( n429 & n6493 ) | ( n429 & n6536 ) | ( n6493 & n6536 ) ;
  assign n6546 = ( n6493 & ~n6498 ) | ( n6493 & n6536 ) | ( ~n6498 & n6536 ) ;
  assign n6547 = ~n6545 & n6546 ;
  assign n6548 = n6541 | n6547 ;
  assign n6549 = n6241 &  n6499 ;
  assign n6542 = x95 | n6241 ;
  assign n6543 = x95 &  n6241 ;
  assign n6544 = ( n6542 & ~n6543 ) | ( n6542 & 1'b0 ) | ( ~n6543 & 1'b0 ) ;
  assign n6553 = ( n429 & n6492 ) | ( n429 & n6544 ) | ( n6492 & n6544 ) ;
  assign n6554 = ( n6492 & ~n6498 ) | ( n6492 & n6544 ) | ( ~n6498 & n6544 ) ;
  assign n6555 = ~n6553 & n6554 ;
  assign n6556 = n6549 | n6555 ;
  assign n6557 = n6249 &  n6499 ;
  assign n6550 = x94 | n6249 ;
  assign n6551 = x94 &  n6249 ;
  assign n6552 = ( n6550 & ~n6551 ) | ( n6550 & 1'b0 ) | ( ~n6551 & 1'b0 ) ;
  assign n6561 = ( n429 & n6491 ) | ( n429 & n6552 ) | ( n6491 & n6552 ) ;
  assign n6562 = ( n6491 & ~n6498 ) | ( n6491 & n6552 ) | ( ~n6498 & n6552 ) ;
  assign n6563 = ~n6561 & n6562 ;
  assign n6564 = n6557 | n6563 ;
  assign n6565 = n6257 &  n6499 ;
  assign n6558 = x93 | n6257 ;
  assign n6559 = x93 &  n6257 ;
  assign n6560 = ( n6558 & ~n6559 ) | ( n6558 & 1'b0 ) | ( ~n6559 & 1'b0 ) ;
  assign n6569 = ( n429 & n6490 ) | ( n429 & n6560 ) | ( n6490 & n6560 ) ;
  assign n6570 = ( n6490 & ~n6498 ) | ( n6490 & n6560 ) | ( ~n6498 & n6560 ) ;
  assign n6571 = ~n6569 & n6570 ;
  assign n6572 = n6565 | n6571 ;
  assign n6573 = n6265 &  n6499 ;
  assign n6566 = x92 | n6265 ;
  assign n6567 = x92 &  n6265 ;
  assign n6568 = ( n6566 & ~n6567 ) | ( n6566 & 1'b0 ) | ( ~n6567 & 1'b0 ) ;
  assign n6577 = ( n429 & n6489 ) | ( n429 & n6568 ) | ( n6489 & n6568 ) ;
  assign n6578 = ( n6489 & ~n6498 ) | ( n6489 & n6568 ) | ( ~n6498 & n6568 ) ;
  assign n6579 = ~n6577 & n6578 ;
  assign n6580 = n6573 | n6579 ;
  assign n6581 = n6273 &  n6499 ;
  assign n6574 = x91 | n6273 ;
  assign n6575 = x91 &  n6273 ;
  assign n6576 = ( n6574 & ~n6575 ) | ( n6574 & 1'b0 ) | ( ~n6575 & 1'b0 ) ;
  assign n6585 = ( n429 & n6488 ) | ( n429 & n6576 ) | ( n6488 & n6576 ) ;
  assign n6586 = ( n6488 & ~n6498 ) | ( n6488 & n6576 ) | ( ~n6498 & n6576 ) ;
  assign n6587 = ~n6585 & n6586 ;
  assign n6588 = n6581 | n6587 ;
  assign n6589 = n6281 &  n6499 ;
  assign n6582 = x90 | n6281 ;
  assign n6583 = x90 &  n6281 ;
  assign n6584 = ( n6582 & ~n6583 ) | ( n6582 & 1'b0 ) | ( ~n6583 & 1'b0 ) ;
  assign n6593 = ( n429 & n6487 ) | ( n429 & n6584 ) | ( n6487 & n6584 ) ;
  assign n6594 = ( n6487 & ~n6498 ) | ( n6487 & n6584 ) | ( ~n6498 & n6584 ) ;
  assign n6595 = ~n6593 & n6594 ;
  assign n6596 = n6589 | n6595 ;
  assign n6597 = n6289 &  n6499 ;
  assign n6590 = x89 | n6289 ;
  assign n6591 = x89 &  n6289 ;
  assign n6592 = ( n6590 & ~n6591 ) | ( n6590 & 1'b0 ) | ( ~n6591 & 1'b0 ) ;
  assign n6601 = ( n429 & n6486 ) | ( n429 & n6592 ) | ( n6486 & n6592 ) ;
  assign n6602 = ( n6486 & ~n6498 ) | ( n6486 & n6592 ) | ( ~n6498 & n6592 ) ;
  assign n6603 = ~n6601 & n6602 ;
  assign n6604 = n6597 | n6603 ;
  assign n6605 = n6297 &  n6499 ;
  assign n6598 = x88 | n6297 ;
  assign n6599 = x88 &  n6297 ;
  assign n6600 = ( n6598 & ~n6599 ) | ( n6598 & 1'b0 ) | ( ~n6599 & 1'b0 ) ;
  assign n6609 = ( n429 & n6485 ) | ( n429 & n6600 ) | ( n6485 & n6600 ) ;
  assign n6610 = ( n6485 & ~n6498 ) | ( n6485 & n6600 ) | ( ~n6498 & n6600 ) ;
  assign n6611 = ~n6609 & n6610 ;
  assign n6612 = n6605 | n6611 ;
  assign n6613 = n6305 &  n6499 ;
  assign n6606 = x87 | n6305 ;
  assign n6607 = x87 &  n6305 ;
  assign n6608 = ( n6606 & ~n6607 ) | ( n6606 & 1'b0 ) | ( ~n6607 & 1'b0 ) ;
  assign n6617 = ( n429 & n6484 ) | ( n429 & n6608 ) | ( n6484 & n6608 ) ;
  assign n6618 = ( n6484 & ~n6498 ) | ( n6484 & n6608 ) | ( ~n6498 & n6608 ) ;
  assign n6619 = ~n6617 & n6618 ;
  assign n6620 = n6613 | n6619 ;
  assign n6621 = n6313 &  n6499 ;
  assign n6614 = x86 | n6313 ;
  assign n6615 = x86 &  n6313 ;
  assign n6616 = ( n6614 & ~n6615 ) | ( n6614 & 1'b0 ) | ( ~n6615 & 1'b0 ) ;
  assign n6625 = ( n429 & n6483 ) | ( n429 & n6616 ) | ( n6483 & n6616 ) ;
  assign n6626 = ( n6483 & ~n6498 ) | ( n6483 & n6616 ) | ( ~n6498 & n6616 ) ;
  assign n6627 = ~n6625 & n6626 ;
  assign n6628 = n6621 | n6627 ;
  assign n6629 = n6321 &  n6499 ;
  assign n6622 = x85 | n6321 ;
  assign n6623 = x85 &  n6321 ;
  assign n6624 = ( n6622 & ~n6623 ) | ( n6622 & 1'b0 ) | ( ~n6623 & 1'b0 ) ;
  assign n6633 = ( n429 & n6482 ) | ( n429 & n6624 ) | ( n6482 & n6624 ) ;
  assign n6634 = ( n6482 & ~n6498 ) | ( n6482 & n6624 ) | ( ~n6498 & n6624 ) ;
  assign n6635 = ~n6633 & n6634 ;
  assign n6636 = n6629 | n6635 ;
  assign n6637 = n6326 &  n6499 ;
  assign n6630 = x84 | n6326 ;
  assign n6631 = x84 &  n6326 ;
  assign n6632 = ( n6630 & ~n6631 ) | ( n6630 & 1'b0 ) | ( ~n6631 & 1'b0 ) ;
  assign n6638 = ( n429 & n6481 ) | ( n429 & n6632 ) | ( n6481 & n6632 ) ;
  assign n6639 = ( n6481 & ~n6498 ) | ( n6481 & n6632 ) | ( ~n6498 & n6632 ) ;
  assign n6640 = ~n6638 & n6639 ;
  assign n6641 = n6637 | n6640 ;
  assign n6500 = n6192 &  n6499 ;
  assign n6504 = x83 | n6192 ;
  assign n6505 = x83 &  n6192 ;
  assign n6506 = ( n6504 & ~n6505 ) | ( n6504 & 1'b0 ) | ( ~n6505 & 1'b0 ) ;
  assign n6507 = ( n429 & n6480 ) | ( n429 & n6506 ) | ( n6480 & n6506 ) ;
  assign n6508 = ( n6480 & ~n6498 ) | ( n6480 & n6506 ) | ( ~n6498 & n6506 ) ;
  assign n6509 = ~n6507 & n6508 ;
  assign n6510 = n6500 | n6509 ;
  assign n6642 = n6334 &  n6499 ;
  assign n6501 = x82 | n6334 ;
  assign n6502 = x82 &  n6334 ;
  assign n6503 = ( n6501 & ~n6502 ) | ( n6501 & 1'b0 ) | ( ~n6502 & 1'b0 ) ;
  assign n6646 = ( n429 & n6479 ) | ( n429 & n6503 ) | ( n6479 & n6503 ) ;
  assign n6647 = ( n6479 & ~n6498 ) | ( n6479 & n6503 ) | ( ~n6498 & n6503 ) ;
  assign n6648 = ~n6646 & n6647 ;
  assign n6649 = n6642 | n6648 ;
  assign n6650 = n6342 &  n6499 ;
  assign n6643 = x81 | n6342 ;
  assign n6644 = x81 &  n6342 ;
  assign n6645 = ( n6643 & ~n6644 ) | ( n6643 & 1'b0 ) | ( ~n6644 & 1'b0 ) ;
  assign n6654 = ( n429 & n6478 ) | ( n429 & n6645 ) | ( n6478 & n6645 ) ;
  assign n6655 = ( n6478 & ~n6498 ) | ( n6478 & n6645 ) | ( ~n6498 & n6645 ) ;
  assign n6656 = ~n6654 & n6655 ;
  assign n6657 = n6650 | n6656 ;
  assign n6658 = n6350 &  n6499 ;
  assign n6651 = x80 | n6350 ;
  assign n6652 = x80 &  n6350 ;
  assign n6653 = ( n6651 & ~n6652 ) | ( n6651 & 1'b0 ) | ( ~n6652 & 1'b0 ) ;
  assign n6662 = ( n429 & n6477 ) | ( n429 & n6653 ) | ( n6477 & n6653 ) ;
  assign n6663 = ( n6477 & ~n6498 ) | ( n6477 & n6653 ) | ( ~n6498 & n6653 ) ;
  assign n6664 = ~n6662 & n6663 ;
  assign n6665 = n6658 | n6664 ;
  assign n6666 = n6358 &  n6499 ;
  assign n6659 = x79 | n6358 ;
  assign n6660 = x79 &  n6358 ;
  assign n6661 = ( n6659 & ~n6660 ) | ( n6659 & 1'b0 ) | ( ~n6660 & 1'b0 ) ;
  assign n6670 = ( n429 & n6476 ) | ( n429 & n6661 ) | ( n6476 & n6661 ) ;
  assign n6671 = ( n6476 & ~n6498 ) | ( n6476 & n6661 ) | ( ~n6498 & n6661 ) ;
  assign n6672 = ~n6670 & n6671 ;
  assign n6673 = n6666 | n6672 ;
  assign n6674 = n6366 &  n6499 ;
  assign n6667 = x78 | n6366 ;
  assign n6668 = x78 &  n6366 ;
  assign n6669 = ( n6667 & ~n6668 ) | ( n6667 & 1'b0 ) | ( ~n6668 & 1'b0 ) ;
  assign n6678 = ( n429 & n6475 ) | ( n429 & n6669 ) | ( n6475 & n6669 ) ;
  assign n6679 = ( n6475 & ~n6498 ) | ( n6475 & n6669 ) | ( ~n6498 & n6669 ) ;
  assign n6680 = ~n6678 & n6679 ;
  assign n6681 = n6674 | n6680 ;
  assign n6682 = n6374 &  n6499 ;
  assign n6675 = x77 | n6374 ;
  assign n6676 = x77 &  n6374 ;
  assign n6677 = ( n6675 & ~n6676 ) | ( n6675 & 1'b0 ) | ( ~n6676 & 1'b0 ) ;
  assign n6686 = ( n429 & n6474 ) | ( n429 & n6677 ) | ( n6474 & n6677 ) ;
  assign n6687 = ( n6474 & ~n6498 ) | ( n6474 & n6677 ) | ( ~n6498 & n6677 ) ;
  assign n6688 = ~n6686 & n6687 ;
  assign n6689 = n6682 | n6688 ;
  assign n6690 = n6382 &  n6499 ;
  assign n6683 = x76 | n6382 ;
  assign n6684 = x76 &  n6382 ;
  assign n6685 = ( n6683 & ~n6684 ) | ( n6683 & 1'b0 ) | ( ~n6684 & 1'b0 ) ;
  assign n6694 = ( n429 & n6473 ) | ( n429 & n6685 ) | ( n6473 & n6685 ) ;
  assign n6695 = ( n6473 & ~n6498 ) | ( n6473 & n6685 ) | ( ~n6498 & n6685 ) ;
  assign n6696 = ~n6694 & n6695 ;
  assign n6697 = n6690 | n6696 ;
  assign n6698 = n6390 &  n6499 ;
  assign n6691 = x75 | n6390 ;
  assign n6692 = x75 &  n6390 ;
  assign n6693 = ( n6691 & ~n6692 ) | ( n6691 & 1'b0 ) | ( ~n6692 & 1'b0 ) ;
  assign n6702 = ( n429 & n6472 ) | ( n429 & n6693 ) | ( n6472 & n6693 ) ;
  assign n6703 = ( n6472 & ~n6498 ) | ( n6472 & n6693 ) | ( ~n6498 & n6693 ) ;
  assign n6704 = ~n6702 & n6703 ;
  assign n6705 = n6698 | n6704 ;
  assign n6706 = n6398 &  n6499 ;
  assign n6699 = x74 | n6398 ;
  assign n6700 = x74 &  n6398 ;
  assign n6701 = ( n6699 & ~n6700 ) | ( n6699 & 1'b0 ) | ( ~n6700 & 1'b0 ) ;
  assign n6710 = ( n429 & n6471 ) | ( n429 & n6701 ) | ( n6471 & n6701 ) ;
  assign n6711 = ( n6471 & ~n6498 ) | ( n6471 & n6701 ) | ( ~n6498 & n6701 ) ;
  assign n6712 = ~n6710 & n6711 ;
  assign n6713 = n6706 | n6712 ;
  assign n6714 = n6406 &  n6499 ;
  assign n6707 = x73 | n6406 ;
  assign n6708 = x73 &  n6406 ;
  assign n6709 = ( n6707 & ~n6708 ) | ( n6707 & 1'b0 ) | ( ~n6708 & 1'b0 ) ;
  assign n6718 = ( n429 & n6470 ) | ( n429 & n6709 ) | ( n6470 & n6709 ) ;
  assign n6719 = ( n6470 & ~n6498 ) | ( n6470 & n6709 ) | ( ~n6498 & n6709 ) ;
  assign n6720 = ~n6718 & n6719 ;
  assign n6721 = n6714 | n6720 ;
  assign n6722 = n6414 &  n6499 ;
  assign n6715 = x72 | n6414 ;
  assign n6716 = x72 &  n6414 ;
  assign n6717 = ( n6715 & ~n6716 ) | ( n6715 & 1'b0 ) | ( ~n6716 & 1'b0 ) ;
  assign n6726 = ( n429 & n6469 ) | ( n429 & n6717 ) | ( n6469 & n6717 ) ;
  assign n6727 = ( n6469 & ~n6498 ) | ( n6469 & n6717 ) | ( ~n6498 & n6717 ) ;
  assign n6728 = ~n6726 & n6727 ;
  assign n6729 = n6722 | n6728 ;
  assign n6730 = n6422 &  n6499 ;
  assign n6723 = x71 | n6422 ;
  assign n6724 = x71 &  n6422 ;
  assign n6725 = ( n6723 & ~n6724 ) | ( n6723 & 1'b0 ) | ( ~n6724 & 1'b0 ) ;
  assign n6734 = ( n429 & n6468 ) | ( n429 & n6725 ) | ( n6468 & n6725 ) ;
  assign n6735 = ( n6468 & ~n6498 ) | ( n6468 & n6725 ) | ( ~n6498 & n6725 ) ;
  assign n6736 = ~n6734 & n6735 ;
  assign n6737 = n6730 | n6736 ;
  assign n6738 = n6430 &  n6499 ;
  assign n6731 = x70 | n6430 ;
  assign n6732 = x70 &  n6430 ;
  assign n6733 = ( n6731 & ~n6732 ) | ( n6731 & 1'b0 ) | ( ~n6732 & 1'b0 ) ;
  assign n6742 = ( n429 & n6467 ) | ( n429 & n6733 ) | ( n6467 & n6733 ) ;
  assign n6743 = ( n6467 & ~n6498 ) | ( n6467 & n6733 ) | ( ~n6498 & n6733 ) ;
  assign n6744 = ~n6742 & n6743 ;
  assign n6745 = n6738 | n6744 ;
  assign n6746 = n6438 &  n6499 ;
  assign n6739 = x69 | n6438 ;
  assign n6740 = x69 &  n6438 ;
  assign n6741 = ( n6739 & ~n6740 ) | ( n6739 & 1'b0 ) | ( ~n6740 & 1'b0 ) ;
  assign n6750 = ( n429 & n6466 ) | ( n429 & n6741 ) | ( n6466 & n6741 ) ;
  assign n6751 = ( n6466 & ~n6498 ) | ( n6466 & n6741 ) | ( ~n6498 & n6741 ) ;
  assign n6752 = ~n6750 & n6751 ;
  assign n6753 = n6746 | n6752 ;
  assign n6754 = n6446 &  n6499 ;
  assign n6747 = x68 | n6446 ;
  assign n6748 = x68 &  n6446 ;
  assign n6749 = ( n6747 & ~n6748 ) | ( n6747 & 1'b0 ) | ( ~n6748 & 1'b0 ) ;
  assign n6758 = ( n429 & n6465 ) | ( n429 & n6749 ) | ( n6465 & n6749 ) ;
  assign n6759 = ( n6465 & ~n6498 ) | ( n6465 & n6749 ) | ( ~n6498 & n6749 ) ;
  assign n6760 = ~n6758 & n6759 ;
  assign n6761 = n6754 | n6760 ;
  assign n6762 = n6451 &  n6499 ;
  assign n6755 = x67 | n6451 ;
  assign n6756 = x67 &  n6451 ;
  assign n6757 = ( n6755 & ~n6756 ) | ( n6755 & 1'b0 ) | ( ~n6756 & 1'b0 ) ;
  assign n6766 = ( n429 & n6464 ) | ( n429 & n6757 ) | ( n6464 & n6757 ) ;
  assign n6767 = ( n6464 & ~n6498 ) | ( n6464 & n6757 ) | ( ~n6498 & n6757 ) ;
  assign n6768 = ~n6766 & n6767 ;
  assign n6769 = n6762 | n6768 ;
  assign n6770 = n6457 &  n6499 ;
  assign n6763 = x66 | n6457 ;
  assign n6764 = x66 &  n6457 ;
  assign n6765 = ( n6763 & ~n6764 ) | ( n6763 & 1'b0 ) | ( ~n6764 & 1'b0 ) ;
  assign n6771 = ( n6463 & ~n429 ) | ( n6463 & n6765 ) | ( ~n429 & n6765 ) ;
  assign n6772 = ( n6463 & n6498 ) | ( n6463 & n6765 ) | ( n6498 & n6765 ) ;
  assign n6773 = ( n6771 & ~n6772 ) | ( n6771 & 1'b0 ) | ( ~n6772 & 1'b0 ) ;
  assign n6774 = n6770 | n6773 ;
  assign n6775 = n6461 &  n6499 ;
  assign n6776 = ( x65 & ~x28 ) | ( x65 & n6458 ) | ( ~x28 & n6458 ) ;
  assign n6777 = ( x28 & ~n6458 ) | ( x28 & x65 ) | ( ~n6458 & x65 ) ;
  assign n6778 = ( n6776 & ~x65 ) | ( n6776 & n6777 ) | ( ~x65 & n6777 ) ;
  assign n6779 = ( n6462 & ~n6498 ) | ( n6462 & n6778 ) | ( ~n6498 & n6778 ) ;
  assign n6780 = ( n429 & n6462 ) | ( n429 & n6778 ) | ( n6462 & n6778 ) ;
  assign n6781 = ( n6779 & ~n6780 ) | ( n6779 & 1'b0 ) | ( ~n6780 & 1'b0 ) ;
  assign n6782 = n6775 | n6781 ;
  assign n6783 = ( x64 & ~x101 ) | ( x64 & 1'b0 ) | ( ~x101 & 1'b0 ) ;
  assign n6784 = ( n163 & ~n165 ) | ( n163 & n6783 ) | ( ~n165 & n6783 ) ;
  assign n6785 = ~n163 & n6784 ;
  assign n6786 = ( n160 & ~n174 ) | ( n160 & n6785 ) | ( ~n174 & n6785 ) ;
  assign n6787 = ~n160 & n6786 ;
  assign n6788 = n6498 &  n6787 ;
  assign n6789 = ( x27 & ~n6787 ) | ( x27 & n6788 ) | ( ~n6787 & n6788 ) ;
  assign n6790 = ~n243 & n6462 ;
  assign n6791 = ( n240 & ~n254 ) | ( n240 & n6790 ) | ( ~n254 & n6790 ) ;
  assign n6792 = ~n240 & n6791 ;
  assign n6793 = ~n6498 & n6792 ;
  assign n6794 = n6789 | n6793 ;
  assign n6795 = ~x26 & x64 ;
  assign n6796 = ( x65 & ~n6794 ) | ( x65 & n6795 ) | ( ~n6794 & n6795 ) ;
  assign n6797 = ( x66 & ~n6782 ) | ( x66 & n6796 ) | ( ~n6782 & n6796 ) ;
  assign n6798 = ( x67 & ~n6774 ) | ( x67 & n6797 ) | ( ~n6774 & n6797 ) ;
  assign n6799 = ( x68 & ~n6769 ) | ( x68 & n6798 ) | ( ~n6769 & n6798 ) ;
  assign n6800 = ( x69 & ~n6761 ) | ( x69 & n6799 ) | ( ~n6761 & n6799 ) ;
  assign n6801 = ( x70 & ~n6753 ) | ( x70 & n6800 ) | ( ~n6753 & n6800 ) ;
  assign n6802 = ( x71 & ~n6745 ) | ( x71 & n6801 ) | ( ~n6745 & n6801 ) ;
  assign n6803 = ( x72 & ~n6737 ) | ( x72 & n6802 ) | ( ~n6737 & n6802 ) ;
  assign n6804 = ( x73 & ~n6729 ) | ( x73 & n6803 ) | ( ~n6729 & n6803 ) ;
  assign n6805 = ( x74 & ~n6721 ) | ( x74 & n6804 ) | ( ~n6721 & n6804 ) ;
  assign n6806 = ( x75 & ~n6713 ) | ( x75 & n6805 ) | ( ~n6713 & n6805 ) ;
  assign n6807 = ( x76 & ~n6705 ) | ( x76 & n6806 ) | ( ~n6705 & n6806 ) ;
  assign n6808 = ( x77 & ~n6697 ) | ( x77 & n6807 ) | ( ~n6697 & n6807 ) ;
  assign n6809 = ( x78 & ~n6689 ) | ( x78 & n6808 ) | ( ~n6689 & n6808 ) ;
  assign n6810 = ( x79 & ~n6681 ) | ( x79 & n6809 ) | ( ~n6681 & n6809 ) ;
  assign n6811 = ( x80 & ~n6673 ) | ( x80 & n6810 ) | ( ~n6673 & n6810 ) ;
  assign n6812 = ( x81 & ~n6665 ) | ( x81 & n6811 ) | ( ~n6665 & n6811 ) ;
  assign n6813 = ( x82 & ~n6657 ) | ( x82 & n6812 ) | ( ~n6657 & n6812 ) ;
  assign n6814 = ( x83 & ~n6649 ) | ( x83 & n6813 ) | ( ~n6649 & n6813 ) ;
  assign n6815 = ( x84 & ~n6510 ) | ( x84 & n6814 ) | ( ~n6510 & n6814 ) ;
  assign n6816 = ( x85 & ~n6641 ) | ( x85 & n6815 ) | ( ~n6641 & n6815 ) ;
  assign n6817 = ( x86 & ~n6636 ) | ( x86 & n6816 ) | ( ~n6636 & n6816 ) ;
  assign n6818 = ( x87 & ~n6628 ) | ( x87 & n6817 ) | ( ~n6628 & n6817 ) ;
  assign n6819 = ( x88 & ~n6620 ) | ( x88 & n6818 ) | ( ~n6620 & n6818 ) ;
  assign n6820 = ( x89 & ~n6612 ) | ( x89 & n6819 ) | ( ~n6612 & n6819 ) ;
  assign n6821 = ( x90 & ~n6604 ) | ( x90 & n6820 ) | ( ~n6604 & n6820 ) ;
  assign n6822 = ( x91 & ~n6596 ) | ( x91 & n6821 ) | ( ~n6596 & n6821 ) ;
  assign n6823 = ( x92 & ~n6588 ) | ( x92 & n6822 ) | ( ~n6588 & n6822 ) ;
  assign n6824 = ( x93 & ~n6580 ) | ( x93 & n6823 ) | ( ~n6580 & n6823 ) ;
  assign n6825 = ( x94 & ~n6572 ) | ( x94 & n6824 ) | ( ~n6572 & n6824 ) ;
  assign n6826 = ( x95 & ~n6564 ) | ( x95 & n6825 ) | ( ~n6564 & n6825 ) ;
  assign n6827 = ( x96 & ~n6556 ) | ( x96 & n6826 ) | ( ~n6556 & n6826 ) ;
  assign n6828 = ( x97 & ~n6548 ) | ( x97 & n6827 ) | ( ~n6548 & n6827 ) ;
  assign n6829 = ( x98 & ~n6540 ) | ( x98 & n6828 ) | ( ~n6540 & n6828 ) ;
  assign n6830 = ( x99 & ~n6532 ) | ( x99 & n6829 ) | ( ~n6532 & n6829 ) ;
  assign n6831 = ( x100 & ~n6524 ) | ( x100 & n6830 ) | ( ~n6524 & n6830 ) ;
  assign n6832 = ( x101 & ~n6516 ) | ( x101 & n6831 ) | ( ~n6516 & n6831 ) ;
  assign n6833 = n163 | n165 ;
  assign n6834 = ( n174 & ~n160 ) | ( n174 & n6833 ) | ( ~n160 & n6833 ) ;
  assign n6835 = n160 | n6834 ;
  assign n6836 = n6832 | n6835 ;
  assign n7048 = n6524 &  n6836 ;
  assign n7052 = x100 | n6524 ;
  assign n7053 = x100 &  n6524 ;
  assign n7054 = ( n7052 & ~n7053 ) | ( n7052 & 1'b0 ) | ( ~n7053 & 1'b0 ) ;
  assign n7055 = ( n6830 & n6832 ) | ( n6830 & n7054 ) | ( n6832 & n7054 ) ;
  assign n7056 = ( n6830 & ~n6835 ) | ( n6830 & n7054 ) | ( ~n6835 & n7054 ) ;
  assign n7057 = ~n7055 & n7056 ;
  assign n7058 = n7048 | n7057 ;
  assign n7059 = n6532 &  n6836 ;
  assign n7049 = x99 | n6532 ;
  assign n7050 = x99 &  n6532 ;
  assign n7051 = ( n7049 & ~n7050 ) | ( n7049 & 1'b0 ) | ( ~n7050 & 1'b0 ) ;
  assign n7063 = ( n6829 & n6832 ) | ( n6829 & n7051 ) | ( n6832 & n7051 ) ;
  assign n7064 = ( n6829 & ~n6835 ) | ( n6829 & n7051 ) | ( ~n6835 & n7051 ) ;
  assign n7065 = ~n7063 & n7064 ;
  assign n7066 = n7059 | n7065 ;
  assign n7067 = n6540 &  n6836 ;
  assign n7060 = x98 | n6540 ;
  assign n7061 = x98 &  n6540 ;
  assign n7062 = ( n7060 & ~n7061 ) | ( n7060 & 1'b0 ) | ( ~n7061 & 1'b0 ) ;
  assign n7071 = ( n6828 & n6832 ) | ( n6828 & n7062 ) | ( n6832 & n7062 ) ;
  assign n7072 = ( n6828 & ~n6835 ) | ( n6828 & n7062 ) | ( ~n6835 & n7062 ) ;
  assign n7073 = ~n7071 & n7072 ;
  assign n7074 = n7067 | n7073 ;
  assign n7075 = n6548 &  n6836 ;
  assign n7068 = x97 | n6548 ;
  assign n7069 = x97 &  n6548 ;
  assign n7070 = ( n7068 & ~n7069 ) | ( n7068 & 1'b0 ) | ( ~n7069 & 1'b0 ) ;
  assign n7079 = ( n6827 & n6832 ) | ( n6827 & n7070 ) | ( n6832 & n7070 ) ;
  assign n7080 = ( n6827 & ~n6835 ) | ( n6827 & n7070 ) | ( ~n6835 & n7070 ) ;
  assign n7081 = ~n7079 & n7080 ;
  assign n7082 = n7075 | n7081 ;
  assign n7083 = n6556 &  n6836 ;
  assign n7076 = x96 | n6556 ;
  assign n7077 = x96 &  n6556 ;
  assign n7078 = ( n7076 & ~n7077 ) | ( n7076 & 1'b0 ) | ( ~n7077 & 1'b0 ) ;
  assign n7087 = ( n6826 & n6832 ) | ( n6826 & n7078 ) | ( n6832 & n7078 ) ;
  assign n7088 = ( n6826 & ~n6835 ) | ( n6826 & n7078 ) | ( ~n6835 & n7078 ) ;
  assign n7089 = ~n7087 & n7088 ;
  assign n7090 = n7083 | n7089 ;
  assign n7091 = n6564 &  n6836 ;
  assign n7084 = x95 | n6564 ;
  assign n7085 = x95 &  n6564 ;
  assign n7086 = ( n7084 & ~n7085 ) | ( n7084 & 1'b0 ) | ( ~n7085 & 1'b0 ) ;
  assign n7095 = ( n6825 & n6832 ) | ( n6825 & n7086 ) | ( n6832 & n7086 ) ;
  assign n7096 = ( n6825 & ~n6835 ) | ( n6825 & n7086 ) | ( ~n6835 & n7086 ) ;
  assign n7097 = ~n7095 & n7096 ;
  assign n7098 = n7091 | n7097 ;
  assign n7099 = n6572 &  n6836 ;
  assign n7092 = x94 | n6572 ;
  assign n7093 = x94 &  n6572 ;
  assign n7094 = ( n7092 & ~n7093 ) | ( n7092 & 1'b0 ) | ( ~n7093 & 1'b0 ) ;
  assign n7103 = ( n6824 & n6832 ) | ( n6824 & n7094 ) | ( n6832 & n7094 ) ;
  assign n7104 = ( n6824 & ~n6835 ) | ( n6824 & n7094 ) | ( ~n6835 & n7094 ) ;
  assign n7105 = ~n7103 & n7104 ;
  assign n7106 = n7099 | n7105 ;
  assign n7107 = n6580 &  n6836 ;
  assign n7100 = x93 | n6580 ;
  assign n7101 = x93 &  n6580 ;
  assign n7102 = ( n7100 & ~n7101 ) | ( n7100 & 1'b0 ) | ( ~n7101 & 1'b0 ) ;
  assign n7111 = ( n6823 & n6832 ) | ( n6823 & n7102 ) | ( n6832 & n7102 ) ;
  assign n7112 = ( n6823 & ~n6835 ) | ( n6823 & n7102 ) | ( ~n6835 & n7102 ) ;
  assign n7113 = ~n7111 & n7112 ;
  assign n7114 = n7107 | n7113 ;
  assign n7115 = n6588 &  n6836 ;
  assign n7108 = x92 | n6588 ;
  assign n7109 = x92 &  n6588 ;
  assign n7110 = ( n7108 & ~n7109 ) | ( n7108 & 1'b0 ) | ( ~n7109 & 1'b0 ) ;
  assign n7119 = ( n6822 & n6832 ) | ( n6822 & n7110 ) | ( n6832 & n7110 ) ;
  assign n7120 = ( n6822 & ~n6835 ) | ( n6822 & n7110 ) | ( ~n6835 & n7110 ) ;
  assign n7121 = ~n7119 & n7120 ;
  assign n7122 = n7115 | n7121 ;
  assign n7123 = n6596 &  n6836 ;
  assign n7116 = x91 | n6596 ;
  assign n7117 = x91 &  n6596 ;
  assign n7118 = ( n7116 & ~n7117 ) | ( n7116 & 1'b0 ) | ( ~n7117 & 1'b0 ) ;
  assign n7127 = ( n6821 & n6832 ) | ( n6821 & n7118 ) | ( n6832 & n7118 ) ;
  assign n7128 = ( n6821 & ~n6835 ) | ( n6821 & n7118 ) | ( ~n6835 & n7118 ) ;
  assign n7129 = ~n7127 & n7128 ;
  assign n7130 = n7123 | n7129 ;
  assign n7131 = n6604 &  n6836 ;
  assign n7124 = x90 | n6604 ;
  assign n7125 = x90 &  n6604 ;
  assign n7126 = ( n7124 & ~n7125 ) | ( n7124 & 1'b0 ) | ( ~n7125 & 1'b0 ) ;
  assign n7135 = ( n6820 & n6832 ) | ( n6820 & n7126 ) | ( n6832 & n7126 ) ;
  assign n7136 = ( n6820 & ~n6835 ) | ( n6820 & n7126 ) | ( ~n6835 & n7126 ) ;
  assign n7137 = ~n7135 & n7136 ;
  assign n7138 = n7131 | n7137 ;
  assign n7139 = n6612 &  n6836 ;
  assign n7132 = x89 | n6612 ;
  assign n7133 = x89 &  n6612 ;
  assign n7134 = ( n7132 & ~n7133 ) | ( n7132 & 1'b0 ) | ( ~n7133 & 1'b0 ) ;
  assign n7143 = ( n6819 & n6832 ) | ( n6819 & n7134 ) | ( n6832 & n7134 ) ;
  assign n7144 = ( n6819 & ~n6835 ) | ( n6819 & n7134 ) | ( ~n6835 & n7134 ) ;
  assign n7145 = ~n7143 & n7144 ;
  assign n7146 = n7139 | n7145 ;
  assign n7147 = n6620 &  n6836 ;
  assign n7140 = x88 | n6620 ;
  assign n7141 = x88 &  n6620 ;
  assign n7142 = ( n7140 & ~n7141 ) | ( n7140 & 1'b0 ) | ( ~n7141 & 1'b0 ) ;
  assign n7151 = ( n6818 & n6832 ) | ( n6818 & n7142 ) | ( n6832 & n7142 ) ;
  assign n7152 = ( n6818 & ~n6835 ) | ( n6818 & n7142 ) | ( ~n6835 & n7142 ) ;
  assign n7153 = ~n7151 & n7152 ;
  assign n7154 = n7147 | n7153 ;
  assign n7155 = n6628 &  n6836 ;
  assign n7148 = x87 | n6628 ;
  assign n7149 = x87 &  n6628 ;
  assign n7150 = ( n7148 & ~n7149 ) | ( n7148 & 1'b0 ) | ( ~n7149 & 1'b0 ) ;
  assign n7159 = ( n6817 & n6832 ) | ( n6817 & n7150 ) | ( n6832 & n7150 ) ;
  assign n7160 = ( n6817 & ~n6835 ) | ( n6817 & n7150 ) | ( ~n6835 & n7150 ) ;
  assign n7161 = ~n7159 & n7160 ;
  assign n7162 = n7155 | n7161 ;
  assign n7163 = n6636 &  n6836 ;
  assign n7156 = x86 | n6636 ;
  assign n7157 = x86 &  n6636 ;
  assign n7158 = ( n7156 & ~n7157 ) | ( n7156 & 1'b0 ) | ( ~n7157 & 1'b0 ) ;
  assign n7164 = ( n6816 & n6832 ) | ( n6816 & n7158 ) | ( n6832 & n7158 ) ;
  assign n7165 = ( n6816 & ~n6835 ) | ( n6816 & n7158 ) | ( ~n6835 & n7158 ) ;
  assign n7166 = ~n7164 & n7165 ;
  assign n7167 = n7163 | n7166 ;
  assign n7037 = n6641 &  n6836 ;
  assign n7038 = x85 | n6641 ;
  assign n7039 = x85 &  n6641 ;
  assign n7040 = ( n7038 & ~n7039 ) | ( n7038 & 1'b0 ) | ( ~n7039 & 1'b0 ) ;
  assign n7041 = ( n6815 & n6832 ) | ( n6815 & n7040 ) | ( n6832 & n7040 ) ;
  assign n7042 = ( n6815 & ~n6835 ) | ( n6815 & n7040 ) | ( ~n6835 & n7040 ) ;
  assign n7043 = ~n7041 & n7042 ;
  assign n7044 = n7037 | n7043 ;
  assign n6837 = n6510 &  n6836 ;
  assign n6841 = x84 | n6510 ;
  assign n6842 = x84 &  n6510 ;
  assign n6843 = ( n6841 & ~n6842 ) | ( n6841 & 1'b0 ) | ( ~n6842 & 1'b0 ) ;
  assign n6844 = ( n6814 & n6832 ) | ( n6814 & n6843 ) | ( n6832 & n6843 ) ;
  assign n6845 = ( n6814 & ~n6835 ) | ( n6814 & n6843 ) | ( ~n6835 & n6843 ) ;
  assign n6846 = ~n6844 & n6845 ;
  assign n6847 = n6837 | n6846 ;
  assign n6848 = n6649 &  n6836 ;
  assign n6838 = x83 | n6649 ;
  assign n6839 = x83 &  n6649 ;
  assign n6840 = ( n6838 & ~n6839 ) | ( n6838 & 1'b0 ) | ( ~n6839 & 1'b0 ) ;
  assign n6852 = ( n6813 & n6832 ) | ( n6813 & n6840 ) | ( n6832 & n6840 ) ;
  assign n6853 = ( n6813 & ~n6835 ) | ( n6813 & n6840 ) | ( ~n6835 & n6840 ) ;
  assign n6854 = ~n6852 & n6853 ;
  assign n6855 = n6848 | n6854 ;
  assign n6856 = n6657 &  n6836 ;
  assign n6849 = x82 | n6657 ;
  assign n6850 = x82 &  n6657 ;
  assign n6851 = ( n6849 & ~n6850 ) | ( n6849 & 1'b0 ) | ( ~n6850 & 1'b0 ) ;
  assign n6860 = ( n6812 & n6832 ) | ( n6812 & n6851 ) | ( n6832 & n6851 ) ;
  assign n6861 = ( n6812 & ~n6835 ) | ( n6812 & n6851 ) | ( ~n6835 & n6851 ) ;
  assign n6862 = ~n6860 & n6861 ;
  assign n6863 = n6856 | n6862 ;
  assign n6864 = n6665 &  n6836 ;
  assign n6857 = x81 | n6665 ;
  assign n6858 = x81 &  n6665 ;
  assign n6859 = ( n6857 & ~n6858 ) | ( n6857 & 1'b0 ) | ( ~n6858 & 1'b0 ) ;
  assign n6868 = ( n6811 & n6832 ) | ( n6811 & n6859 ) | ( n6832 & n6859 ) ;
  assign n6869 = ( n6811 & ~n6835 ) | ( n6811 & n6859 ) | ( ~n6835 & n6859 ) ;
  assign n6870 = ~n6868 & n6869 ;
  assign n6871 = n6864 | n6870 ;
  assign n6872 = n6673 &  n6836 ;
  assign n6865 = x80 | n6673 ;
  assign n6866 = x80 &  n6673 ;
  assign n6867 = ( n6865 & ~n6866 ) | ( n6865 & 1'b0 ) | ( ~n6866 & 1'b0 ) ;
  assign n6876 = ( n6810 & n6832 ) | ( n6810 & n6867 ) | ( n6832 & n6867 ) ;
  assign n6877 = ( n6810 & ~n6835 ) | ( n6810 & n6867 ) | ( ~n6835 & n6867 ) ;
  assign n6878 = ~n6876 & n6877 ;
  assign n6879 = n6872 | n6878 ;
  assign n6880 = n6681 &  n6836 ;
  assign n6873 = x79 | n6681 ;
  assign n6874 = x79 &  n6681 ;
  assign n6875 = ( n6873 & ~n6874 ) | ( n6873 & 1'b0 ) | ( ~n6874 & 1'b0 ) ;
  assign n6884 = ( n6809 & n6832 ) | ( n6809 & n6875 ) | ( n6832 & n6875 ) ;
  assign n6885 = ( n6809 & ~n6835 ) | ( n6809 & n6875 ) | ( ~n6835 & n6875 ) ;
  assign n6886 = ~n6884 & n6885 ;
  assign n6887 = n6880 | n6886 ;
  assign n6888 = n6689 &  n6836 ;
  assign n6881 = x78 | n6689 ;
  assign n6882 = x78 &  n6689 ;
  assign n6883 = ( n6881 & ~n6882 ) | ( n6881 & 1'b0 ) | ( ~n6882 & 1'b0 ) ;
  assign n6892 = ( n6808 & n6832 ) | ( n6808 & n6883 ) | ( n6832 & n6883 ) ;
  assign n6893 = ( n6808 & ~n6835 ) | ( n6808 & n6883 ) | ( ~n6835 & n6883 ) ;
  assign n6894 = ~n6892 & n6893 ;
  assign n6895 = n6888 | n6894 ;
  assign n6896 = n6697 &  n6836 ;
  assign n6889 = x77 | n6697 ;
  assign n6890 = x77 &  n6697 ;
  assign n6891 = ( n6889 & ~n6890 ) | ( n6889 & 1'b0 ) | ( ~n6890 & 1'b0 ) ;
  assign n6900 = ( n6807 & n6832 ) | ( n6807 & n6891 ) | ( n6832 & n6891 ) ;
  assign n6901 = ( n6807 & ~n6835 ) | ( n6807 & n6891 ) | ( ~n6835 & n6891 ) ;
  assign n6902 = ~n6900 & n6901 ;
  assign n6903 = n6896 | n6902 ;
  assign n6904 = n6705 &  n6836 ;
  assign n6897 = x76 | n6705 ;
  assign n6898 = x76 &  n6705 ;
  assign n6899 = ( n6897 & ~n6898 ) | ( n6897 & 1'b0 ) | ( ~n6898 & 1'b0 ) ;
  assign n6908 = ( n6806 & n6832 ) | ( n6806 & n6899 ) | ( n6832 & n6899 ) ;
  assign n6909 = ( n6806 & ~n6835 ) | ( n6806 & n6899 ) | ( ~n6835 & n6899 ) ;
  assign n6910 = ~n6908 & n6909 ;
  assign n6911 = n6904 | n6910 ;
  assign n6912 = n6713 &  n6836 ;
  assign n6905 = x75 | n6713 ;
  assign n6906 = x75 &  n6713 ;
  assign n6907 = ( n6905 & ~n6906 ) | ( n6905 & 1'b0 ) | ( ~n6906 & 1'b0 ) ;
  assign n6916 = ( n6805 & n6832 ) | ( n6805 & n6907 ) | ( n6832 & n6907 ) ;
  assign n6917 = ( n6805 & ~n6835 ) | ( n6805 & n6907 ) | ( ~n6835 & n6907 ) ;
  assign n6918 = ~n6916 & n6917 ;
  assign n6919 = n6912 | n6918 ;
  assign n6920 = n6721 &  n6836 ;
  assign n6913 = x74 | n6721 ;
  assign n6914 = x74 &  n6721 ;
  assign n6915 = ( n6913 & ~n6914 ) | ( n6913 & 1'b0 ) | ( ~n6914 & 1'b0 ) ;
  assign n6924 = ( n6804 & n6832 ) | ( n6804 & n6915 ) | ( n6832 & n6915 ) ;
  assign n6925 = ( n6804 & ~n6835 ) | ( n6804 & n6915 ) | ( ~n6835 & n6915 ) ;
  assign n6926 = ~n6924 & n6925 ;
  assign n6927 = n6920 | n6926 ;
  assign n6928 = n6729 &  n6836 ;
  assign n6921 = x73 | n6729 ;
  assign n6922 = x73 &  n6729 ;
  assign n6923 = ( n6921 & ~n6922 ) | ( n6921 & 1'b0 ) | ( ~n6922 & 1'b0 ) ;
  assign n6932 = ( n6803 & n6832 ) | ( n6803 & n6923 ) | ( n6832 & n6923 ) ;
  assign n6933 = ( n6803 & ~n6835 ) | ( n6803 & n6923 ) | ( ~n6835 & n6923 ) ;
  assign n6934 = ~n6932 & n6933 ;
  assign n6935 = n6928 | n6934 ;
  assign n6936 = n6737 &  n6836 ;
  assign n6929 = x72 | n6737 ;
  assign n6930 = x72 &  n6737 ;
  assign n6931 = ( n6929 & ~n6930 ) | ( n6929 & 1'b0 ) | ( ~n6930 & 1'b0 ) ;
  assign n6940 = ( n6802 & n6832 ) | ( n6802 & n6931 ) | ( n6832 & n6931 ) ;
  assign n6941 = ( n6802 & ~n6835 ) | ( n6802 & n6931 ) | ( ~n6835 & n6931 ) ;
  assign n6942 = ~n6940 & n6941 ;
  assign n6943 = n6936 | n6942 ;
  assign n6944 = n6745 &  n6836 ;
  assign n6937 = x71 | n6745 ;
  assign n6938 = x71 &  n6745 ;
  assign n6939 = ( n6937 & ~n6938 ) | ( n6937 & 1'b0 ) | ( ~n6938 & 1'b0 ) ;
  assign n6948 = ( n6801 & n6832 ) | ( n6801 & n6939 ) | ( n6832 & n6939 ) ;
  assign n6949 = ( n6801 & ~n6835 ) | ( n6801 & n6939 ) | ( ~n6835 & n6939 ) ;
  assign n6950 = ~n6948 & n6949 ;
  assign n6951 = n6944 | n6950 ;
  assign n6952 = n6753 &  n6836 ;
  assign n6945 = x70 | n6753 ;
  assign n6946 = x70 &  n6753 ;
  assign n6947 = ( n6945 & ~n6946 ) | ( n6945 & 1'b0 ) | ( ~n6946 & 1'b0 ) ;
  assign n6956 = ( n6800 & n6832 ) | ( n6800 & n6947 ) | ( n6832 & n6947 ) ;
  assign n6957 = ( n6800 & ~n6835 ) | ( n6800 & n6947 ) | ( ~n6835 & n6947 ) ;
  assign n6958 = ~n6956 & n6957 ;
  assign n6959 = n6952 | n6958 ;
  assign n6960 = n6761 &  n6836 ;
  assign n6953 = x69 | n6761 ;
  assign n6954 = x69 &  n6761 ;
  assign n6955 = ( n6953 & ~n6954 ) | ( n6953 & 1'b0 ) | ( ~n6954 & 1'b0 ) ;
  assign n6964 = ( n6799 & n6832 ) | ( n6799 & n6955 ) | ( n6832 & n6955 ) ;
  assign n6965 = ( n6799 & ~n6835 ) | ( n6799 & n6955 ) | ( ~n6835 & n6955 ) ;
  assign n6966 = ~n6964 & n6965 ;
  assign n6967 = n6960 | n6966 ;
  assign n6968 = n6769 &  n6836 ;
  assign n6961 = x68 | n6769 ;
  assign n6962 = x68 &  n6769 ;
  assign n6963 = ( n6961 & ~n6962 ) | ( n6961 & 1'b0 ) | ( ~n6962 & 1'b0 ) ;
  assign n6972 = ( n6798 & n6832 ) | ( n6798 & n6963 ) | ( n6832 & n6963 ) ;
  assign n6973 = ( n6798 & ~n6835 ) | ( n6798 & n6963 ) | ( ~n6835 & n6963 ) ;
  assign n6974 = ~n6972 & n6973 ;
  assign n6975 = n6968 | n6974 ;
  assign n6976 = n6774 &  n6836 ;
  assign n6969 = x67 | n6774 ;
  assign n6970 = x67 &  n6774 ;
  assign n6971 = ( n6969 & ~n6970 ) | ( n6969 & 1'b0 ) | ( ~n6970 & 1'b0 ) ;
  assign n6980 = ( n6797 & n6832 ) | ( n6797 & n6971 ) | ( n6832 & n6971 ) ;
  assign n6981 = ( n6797 & ~n6835 ) | ( n6797 & n6971 ) | ( ~n6835 & n6971 ) ;
  assign n6982 = ~n6980 & n6981 ;
  assign n6983 = n6976 | n6982 ;
  assign n6984 = n6782 &  n6836 ;
  assign n6977 = x66 | n6782 ;
  assign n6978 = x66 &  n6782 ;
  assign n6979 = ( n6977 & ~n6978 ) | ( n6977 & 1'b0 ) | ( ~n6978 & 1'b0 ) ;
  assign n6989 = ( n6796 & ~n6832 ) | ( n6796 & n6979 ) | ( ~n6832 & n6979 ) ;
  assign n6990 = ( n6796 & n6835 ) | ( n6796 & n6979 ) | ( n6835 & n6979 ) ;
  assign n6991 = ( n6989 & ~n6990 ) | ( n6989 & 1'b0 ) | ( ~n6990 & 1'b0 ) ;
  assign n6992 = n6984 | n6991 ;
  assign n6993 = n6794 &  n6836 ;
  assign n6985 = x65 &  n6794 ;
  assign n6986 = x65 | n6793 ;
  assign n6987 = n6789 | n6986 ;
  assign n6988 = ( n6795 & ~n6985 ) | ( n6795 & n6987 ) | ( ~n6985 & n6987 ) ;
  assign n6994 = ( x65 & n6794 ) | ( x65 & n6795 ) | ( n6794 & n6795 ) ;
  assign n6995 = ( n6835 & ~n6985 ) | ( n6835 & n6994 ) | ( ~n6985 & n6994 ) ;
  assign n6996 = ( n6832 & n6988 ) | ( n6832 & n6995 ) | ( n6988 & n6995 ) ;
  assign n6997 = ( n6988 & ~n6996 ) | ( n6988 & 1'b0 ) | ( ~n6996 & 1'b0 ) ;
  assign n6998 = n6993 | n6997 ;
  assign n6999 = ( x64 & ~x102 ) | ( x64 & 1'b0 ) | ( ~x102 & 1'b0 ) ;
  assign n7000 = ( n242 & ~n253 ) | ( n242 & n6999 ) | ( ~n253 & n6999 ) ;
  assign n7001 = ~n242 & n7000 ;
  assign n7002 = ( n425 & ~n427 ) | ( n425 & n7001 ) | ( ~n427 & n7001 ) ;
  assign n7003 = ~n425 & n7002 ;
  assign n7004 = n6832 &  n7003 ;
  assign n7005 = ( x26 & ~n7003 ) | ( x26 & n7004 ) | ( ~n7003 & n7004 ) ;
  assign n7006 = ~n165 & n6795 ;
  assign n7007 = ( n163 & ~n174 ) | ( n163 & n7006 ) | ( ~n174 & n7006 ) ;
  assign n7008 = ~n163 & n7007 ;
  assign n7009 = ~n160 & n7008 ;
  assign n7010 = ~n6832 & n7009 ;
  assign n7011 = n7005 | n7010 ;
  assign n7012 = ~x25 & x64 ;
  assign n7013 = ( x65 & ~n7011 ) | ( x65 & n7012 ) | ( ~n7011 & n7012 ) ;
  assign n7014 = ( x66 & ~n6998 ) | ( x66 & n7013 ) | ( ~n6998 & n7013 ) ;
  assign n7015 = ( x67 & ~n6992 ) | ( x67 & n7014 ) | ( ~n6992 & n7014 ) ;
  assign n7016 = ( x68 & ~n6983 ) | ( x68 & n7015 ) | ( ~n6983 & n7015 ) ;
  assign n7017 = ( x69 & ~n6975 ) | ( x69 & n7016 ) | ( ~n6975 & n7016 ) ;
  assign n7018 = ( x70 & ~n6967 ) | ( x70 & n7017 ) | ( ~n6967 & n7017 ) ;
  assign n7019 = ( x71 & ~n6959 ) | ( x71 & n7018 ) | ( ~n6959 & n7018 ) ;
  assign n7020 = ( x72 & ~n6951 ) | ( x72 & n7019 ) | ( ~n6951 & n7019 ) ;
  assign n7021 = ( x73 & ~n6943 ) | ( x73 & n7020 ) | ( ~n6943 & n7020 ) ;
  assign n7022 = ( x74 & ~n6935 ) | ( x74 & n7021 ) | ( ~n6935 & n7021 ) ;
  assign n7023 = ( x75 & ~n6927 ) | ( x75 & n7022 ) | ( ~n6927 & n7022 ) ;
  assign n7024 = ( x76 & ~n6919 ) | ( x76 & n7023 ) | ( ~n6919 & n7023 ) ;
  assign n7025 = ( x77 & ~n6911 ) | ( x77 & n7024 ) | ( ~n6911 & n7024 ) ;
  assign n7026 = ( x78 & ~n6903 ) | ( x78 & n7025 ) | ( ~n6903 & n7025 ) ;
  assign n7027 = ( x79 & ~n6895 ) | ( x79 & n7026 ) | ( ~n6895 & n7026 ) ;
  assign n7028 = ( x80 & ~n6887 ) | ( x80 & n7027 ) | ( ~n6887 & n7027 ) ;
  assign n7029 = ( x81 & ~n6879 ) | ( x81 & n7028 ) | ( ~n6879 & n7028 ) ;
  assign n7030 = ( x82 & ~n6871 ) | ( x82 & n7029 ) | ( ~n6871 & n7029 ) ;
  assign n7031 = ( x83 & ~n6863 ) | ( x83 & n7030 ) | ( ~n6863 & n7030 ) ;
  assign n7032 = ( x84 & ~n6855 ) | ( x84 & n7031 ) | ( ~n6855 & n7031 ) ;
  assign n7036 = ( x85 & ~n6847 ) | ( x85 & n7032 ) | ( ~n6847 & n7032 ) ;
  assign n7168 = ( x86 & ~n7044 ) | ( x86 & n7036 ) | ( ~n7044 & n7036 ) ;
  assign n7169 = ( x87 & ~n7167 ) | ( x87 & n7168 ) | ( ~n7167 & n7168 ) ;
  assign n7170 = ( x88 & ~n7162 ) | ( x88 & n7169 ) | ( ~n7162 & n7169 ) ;
  assign n7171 = ( x89 & ~n7154 ) | ( x89 & n7170 ) | ( ~n7154 & n7170 ) ;
  assign n7172 = ( x90 & ~n7146 ) | ( x90 & n7171 ) | ( ~n7146 & n7171 ) ;
  assign n7173 = ( x91 & ~n7138 ) | ( x91 & n7172 ) | ( ~n7138 & n7172 ) ;
  assign n7174 = ( x92 & ~n7130 ) | ( x92 & n7173 ) | ( ~n7130 & n7173 ) ;
  assign n7175 = ( x93 & ~n7122 ) | ( x93 & n7174 ) | ( ~n7122 & n7174 ) ;
  assign n7176 = ( x94 & ~n7114 ) | ( x94 & n7175 ) | ( ~n7114 & n7175 ) ;
  assign n7177 = ( x95 & ~n7106 ) | ( x95 & n7176 ) | ( ~n7106 & n7176 ) ;
  assign n7178 = ( x96 & ~n7098 ) | ( x96 & n7177 ) | ( ~n7098 & n7177 ) ;
  assign n7179 = ( x97 & ~n7090 ) | ( x97 & n7178 ) | ( ~n7090 & n7178 ) ;
  assign n7180 = ( x98 & ~n7082 ) | ( x98 & n7179 ) | ( ~n7082 & n7179 ) ;
  assign n7181 = ( x99 & ~n7074 ) | ( x99 & n7180 ) | ( ~n7074 & n7180 ) ;
  assign n7182 = ( x100 & ~n7066 ) | ( x100 & n7181 ) | ( ~n7066 & n7181 ) ;
  assign n7183 = ( x101 & ~n7058 ) | ( x101 & n7182 ) | ( ~n7058 & n7182 ) ;
  assign n7187 = n242 | n253 ;
  assign n7188 = ( n427 & ~n425 ) | ( n427 & n7187 ) | ( ~n425 & n7187 ) ;
  assign n7189 = n425 | n7188 ;
  assign n7184 = x101 | n6831 ;
  assign n7185 = ( x101 & n6831 ) | ( x101 & n6835 ) | ( n6831 & n6835 ) ;
  assign n7186 = ( n6516 & ~n7184 ) | ( n6516 & n7185 ) | ( ~n7184 & n7185 ) ;
  assign n7191 = x102 &  n7186 ;
  assign n7190 = x102 | n7186 ;
  assign n7192 = ( n7189 & ~n7191 ) | ( n7189 & n7190 ) | ( ~n7191 & n7190 ) ;
  assign n7193 = n7183 | n7192 ;
  assign n7194 = ~n7186 |  n6835 ;
  assign n7214 = n7058 &  n7194 ;
  assign n7215 = n7193 &  n7214 ;
  assign n7201 = x101 | n7058 ;
  assign n7202 = x101 &  n7058 ;
  assign n7203 = ( n7201 & ~n7202 ) | ( n7201 & 1'b0 ) | ( ~n7202 & 1'b0 ) ;
  assign n7216 = n7182 &  n7203 ;
  assign n7195 = n7193 &  n7194 ;
  assign n7217 = ( n7182 & ~n7195 ) | ( n7182 & n7203 ) | ( ~n7195 & n7203 ) ;
  assign n7218 = ( n7215 & ~n7216 ) | ( n7215 & n7217 ) | ( ~n7216 & n7217 ) ;
  assign n7205 = ( x102 & n7183 ) | ( x102 & n7186 ) | ( n7183 & n7186 ) ;
  assign n7204 = ( x102 & ~n7183 ) | ( x102 & n7186 ) | ( ~n7183 & n7186 ) ;
  assign n7206 = ( n7183 & ~n7205 ) | ( n7183 & n7204 ) | ( ~n7205 & n7204 ) ;
  assign n7207 = ~n7195 & n7206 ;
  assign n7208 = n6516 &  n6835 ;
  assign n7209 = n7193 &  n7208 ;
  assign n7210 = n7207 | n7209 ;
  assign n7222 = n7066 &  n7194 ;
  assign n7223 = n7193 &  n7222 ;
  assign n7211 = x100 | n7066 ;
  assign n7212 = x100 &  n7066 ;
  assign n7213 = ( n7211 & ~n7212 ) | ( n7211 & 1'b0 ) | ( ~n7212 & 1'b0 ) ;
  assign n7224 = n7181 &  n7213 ;
  assign n7225 = ( n7181 & ~n7195 ) | ( n7181 & n7213 ) | ( ~n7195 & n7213 ) ;
  assign n7226 = ( n7223 & ~n7224 ) | ( n7223 & n7225 ) | ( ~n7224 & n7225 ) ;
  assign n7230 = n7074 &  n7194 ;
  assign n7231 = n7193 &  n7230 ;
  assign n7219 = x99 | n7074 ;
  assign n7220 = x99 &  n7074 ;
  assign n7221 = ( n7219 & ~n7220 ) | ( n7219 & 1'b0 ) | ( ~n7220 & 1'b0 ) ;
  assign n7232 = n7180 &  n7221 ;
  assign n7233 = ( n7180 & ~n7195 ) | ( n7180 & n7221 ) | ( ~n7195 & n7221 ) ;
  assign n7234 = ( n7231 & ~n7232 ) | ( n7231 & n7233 ) | ( ~n7232 & n7233 ) ;
  assign n7238 = n7082 &  n7194 ;
  assign n7239 = n7193 &  n7238 ;
  assign n7227 = x98 | n7082 ;
  assign n7228 = x98 &  n7082 ;
  assign n7229 = ( n7227 & ~n7228 ) | ( n7227 & 1'b0 ) | ( ~n7228 & 1'b0 ) ;
  assign n7240 = n7179 &  n7229 ;
  assign n7241 = ( n7179 & ~n7195 ) | ( n7179 & n7229 ) | ( ~n7195 & n7229 ) ;
  assign n7242 = ( n7239 & ~n7240 ) | ( n7239 & n7241 ) | ( ~n7240 & n7241 ) ;
  assign n7246 = n7090 &  n7194 ;
  assign n7247 = n7193 &  n7246 ;
  assign n7235 = x97 | n7090 ;
  assign n7236 = x97 &  n7090 ;
  assign n7237 = ( n7235 & ~n7236 ) | ( n7235 & 1'b0 ) | ( ~n7236 & 1'b0 ) ;
  assign n7248 = n7178 &  n7237 ;
  assign n7249 = ( n7178 & ~n7195 ) | ( n7178 & n7237 ) | ( ~n7195 & n7237 ) ;
  assign n7250 = ( n7247 & ~n7248 ) | ( n7247 & n7249 ) | ( ~n7248 & n7249 ) ;
  assign n7254 = n7098 &  n7194 ;
  assign n7255 = n7193 &  n7254 ;
  assign n7243 = x96 | n7098 ;
  assign n7244 = x96 &  n7098 ;
  assign n7245 = ( n7243 & ~n7244 ) | ( n7243 & 1'b0 ) | ( ~n7244 & 1'b0 ) ;
  assign n7257 = ( n7177 & n7195 ) | ( n7177 & n7245 ) | ( n7195 & n7245 ) ;
  assign n7256 = n7177 | n7245 ;
  assign n7258 = ( n7255 & ~n7257 ) | ( n7255 & n7256 ) | ( ~n7257 & n7256 ) ;
  assign n7262 = n7106 &  n7194 ;
  assign n7263 = n7193 &  n7262 ;
  assign n7251 = x95 | n7106 ;
  assign n7252 = x95 &  n7106 ;
  assign n7253 = ( n7251 & ~n7252 ) | ( n7251 & 1'b0 ) | ( ~n7252 & 1'b0 ) ;
  assign n7265 = ( n7176 & n7195 ) | ( n7176 & n7253 ) | ( n7195 & n7253 ) ;
  assign n7264 = n7176 | n7253 ;
  assign n7266 = ( n7263 & ~n7265 ) | ( n7263 & n7264 ) | ( ~n7265 & n7264 ) ;
  assign n7270 = n7114 &  n7194 ;
  assign n7271 = n7193 &  n7270 ;
  assign n7259 = x94 | n7114 ;
  assign n7260 = x94 &  n7114 ;
  assign n7261 = ( n7259 & ~n7260 ) | ( n7259 & 1'b0 ) | ( ~n7260 & 1'b0 ) ;
  assign n7273 = ( n7175 & n7195 ) | ( n7175 & n7261 ) | ( n7195 & n7261 ) ;
  assign n7272 = n7175 | n7261 ;
  assign n7274 = ( n7271 & ~n7273 ) | ( n7271 & n7272 ) | ( ~n7273 & n7272 ) ;
  assign n7278 = n7122 &  n7194 ;
  assign n7279 = n7193 &  n7278 ;
  assign n7267 = x93 | n7122 ;
  assign n7268 = x93 &  n7122 ;
  assign n7269 = ( n7267 & ~n7268 ) | ( n7267 & 1'b0 ) | ( ~n7268 & 1'b0 ) ;
  assign n7281 = ( n7174 & n7195 ) | ( n7174 & n7269 ) | ( n7195 & n7269 ) ;
  assign n7280 = n7174 | n7269 ;
  assign n7282 = ( n7279 & ~n7281 ) | ( n7279 & n7280 ) | ( ~n7281 & n7280 ) ;
  assign n7286 = n7130 &  n7194 ;
  assign n7287 = n7193 &  n7286 ;
  assign n7275 = x92 | n7130 ;
  assign n7276 = x92 &  n7130 ;
  assign n7277 = ( n7275 & ~n7276 ) | ( n7275 & 1'b0 ) | ( ~n7276 & 1'b0 ) ;
  assign n7289 = ( n7173 & n7195 ) | ( n7173 & n7277 ) | ( n7195 & n7277 ) ;
  assign n7288 = n7173 | n7277 ;
  assign n7290 = ( n7287 & ~n7289 ) | ( n7287 & n7288 ) | ( ~n7289 & n7288 ) ;
  assign n7294 = n7138 &  n7194 ;
  assign n7295 = n7193 &  n7294 ;
  assign n7283 = x91 | n7138 ;
  assign n7284 = x91 &  n7138 ;
  assign n7285 = ( n7283 & ~n7284 ) | ( n7283 & 1'b0 ) | ( ~n7284 & 1'b0 ) ;
  assign n7297 = ( n7172 & n7195 ) | ( n7172 & n7285 ) | ( n7195 & n7285 ) ;
  assign n7296 = n7172 | n7285 ;
  assign n7298 = ( n7295 & ~n7297 ) | ( n7295 & n7296 ) | ( ~n7297 & n7296 ) ;
  assign n7302 = n7146 &  n7194 ;
  assign n7303 = n7193 &  n7302 ;
  assign n7291 = x90 | n7146 ;
  assign n7292 = x90 &  n7146 ;
  assign n7293 = ( n7291 & ~n7292 ) | ( n7291 & 1'b0 ) | ( ~n7292 & 1'b0 ) ;
  assign n7305 = ( n7171 & n7195 ) | ( n7171 & n7293 ) | ( n7195 & n7293 ) ;
  assign n7304 = n7171 | n7293 ;
  assign n7306 = ( n7303 & ~n7305 ) | ( n7303 & n7304 ) | ( ~n7305 & n7304 ) ;
  assign n7310 = n7154 &  n7194 ;
  assign n7311 = n7193 &  n7310 ;
  assign n7299 = x89 | n7154 ;
  assign n7300 = x89 &  n7154 ;
  assign n7301 = ( n7299 & ~n7300 ) | ( n7299 & 1'b0 ) | ( ~n7300 & 1'b0 ) ;
  assign n7313 = ( n7170 & n7195 ) | ( n7170 & n7301 ) | ( n7195 & n7301 ) ;
  assign n7312 = n7170 | n7301 ;
  assign n7314 = ( n7311 & ~n7313 ) | ( n7311 & n7312 ) | ( ~n7313 & n7312 ) ;
  assign n7318 = n7162 &  n7194 ;
  assign n7319 = n7193 &  n7318 ;
  assign n7307 = x88 | n7162 ;
  assign n7308 = x88 &  n7162 ;
  assign n7309 = ( n7307 & ~n7308 ) | ( n7307 & 1'b0 ) | ( ~n7308 & 1'b0 ) ;
  assign n7321 = ( n7169 & n7195 ) | ( n7169 & n7309 ) | ( n7195 & n7309 ) ;
  assign n7320 = n7169 | n7309 ;
  assign n7322 = ( n7319 & ~n7321 ) | ( n7319 & n7320 ) | ( ~n7321 & n7320 ) ;
  assign n7323 = n7167 &  n7194 ;
  assign n7324 = n7193 &  n7323 ;
  assign n7315 = x87 | n7167 ;
  assign n7316 = x87 &  n7167 ;
  assign n7317 = ( n7315 & ~n7316 ) | ( n7315 & 1'b0 ) | ( ~n7316 & 1'b0 ) ;
  assign n7326 = ( n7168 & n7195 ) | ( n7168 & n7317 ) | ( n7195 & n7317 ) ;
  assign n7325 = n7168 | n7317 ;
  assign n7327 = ( n7324 & ~n7326 ) | ( n7324 & n7325 ) | ( ~n7326 & n7325 ) ;
  assign n7196 = n7044 &  n7194 ;
  assign n7197 = n7193 &  n7196 ;
  assign n7045 = x86 | n7044 ;
  assign n7046 = x86 &  n7044 ;
  assign n7047 = ( n7045 & ~n7046 ) | ( n7045 & 1'b0 ) | ( ~n7046 & 1'b0 ) ;
  assign n7199 = ( n7036 & n7047 ) | ( n7036 & n7195 ) | ( n7047 & n7195 ) ;
  assign n7198 = n7036 | n7047 ;
  assign n7200 = ( n7197 & ~n7199 ) | ( n7197 & n7198 ) | ( ~n7199 & n7198 ) ;
  assign n7331 = n6847 &  n7194 ;
  assign n7332 = n7193 &  n7331 ;
  assign n7033 = x85 | n6847 ;
  assign n7034 = x85 &  n6847 ;
  assign n7035 = ( n7033 & ~n7034 ) | ( n7033 & 1'b0 ) | ( ~n7034 & 1'b0 ) ;
  assign n7333 = n7032 &  n7035 ;
  assign n7334 = ( n7032 & ~n7195 ) | ( n7032 & n7035 ) | ( ~n7195 & n7035 ) ;
  assign n7335 = ( n7332 & ~n7333 ) | ( n7332 & n7334 ) | ( ~n7333 & n7334 ) ;
  assign n7339 = n6855 &  n7194 ;
  assign n7340 = n7193 &  n7339 ;
  assign n7328 = x84 | n6855 ;
  assign n7329 = x84 &  n6855 ;
  assign n7330 = ( n7328 & ~n7329 ) | ( n7328 & 1'b0 ) | ( ~n7329 & 1'b0 ) ;
  assign n7342 = ( n7031 & n7195 ) | ( n7031 & n7330 ) | ( n7195 & n7330 ) ;
  assign n7341 = n7031 | n7330 ;
  assign n7343 = ( n7340 & ~n7342 ) | ( n7340 & n7341 ) | ( ~n7342 & n7341 ) ;
  assign n7347 = n6863 &  n7194 ;
  assign n7348 = n7193 &  n7347 ;
  assign n7336 = x83 | n6863 ;
  assign n7337 = x83 &  n6863 ;
  assign n7338 = ( n7336 & ~n7337 ) | ( n7336 & 1'b0 ) | ( ~n7337 & 1'b0 ) ;
  assign n7350 = ( n7030 & n7195 ) | ( n7030 & n7338 ) | ( n7195 & n7338 ) ;
  assign n7349 = n7030 | n7338 ;
  assign n7351 = ( n7348 & ~n7350 ) | ( n7348 & n7349 ) | ( ~n7350 & n7349 ) ;
  assign n7355 = n6871 &  n7194 ;
  assign n7356 = n7193 &  n7355 ;
  assign n7344 = x82 | n6871 ;
  assign n7345 = x82 &  n6871 ;
  assign n7346 = ( n7344 & ~n7345 ) | ( n7344 & 1'b0 ) | ( ~n7345 & 1'b0 ) ;
  assign n7358 = ( n7029 & n7195 ) | ( n7029 & n7346 ) | ( n7195 & n7346 ) ;
  assign n7357 = n7029 | n7346 ;
  assign n7359 = ( n7356 & ~n7358 ) | ( n7356 & n7357 ) | ( ~n7358 & n7357 ) ;
  assign n7363 = n6879 &  n7194 ;
  assign n7364 = n7193 &  n7363 ;
  assign n7352 = x81 | n6879 ;
  assign n7353 = x81 &  n6879 ;
  assign n7354 = ( n7352 & ~n7353 ) | ( n7352 & 1'b0 ) | ( ~n7353 & 1'b0 ) ;
  assign n7366 = ( n7028 & n7195 ) | ( n7028 & n7354 ) | ( n7195 & n7354 ) ;
  assign n7365 = n7028 | n7354 ;
  assign n7367 = ( n7364 & ~n7366 ) | ( n7364 & n7365 ) | ( ~n7366 & n7365 ) ;
  assign n7371 = n6887 &  n7194 ;
  assign n7372 = n7193 &  n7371 ;
  assign n7360 = x80 | n6887 ;
  assign n7361 = x80 &  n6887 ;
  assign n7362 = ( n7360 & ~n7361 ) | ( n7360 & 1'b0 ) | ( ~n7361 & 1'b0 ) ;
  assign n7374 = ( n7027 & n7195 ) | ( n7027 & n7362 ) | ( n7195 & n7362 ) ;
  assign n7373 = n7027 | n7362 ;
  assign n7375 = ( n7372 & ~n7374 ) | ( n7372 & n7373 ) | ( ~n7374 & n7373 ) ;
  assign n7379 = n6895 &  n7194 ;
  assign n7380 = n7193 &  n7379 ;
  assign n7368 = x79 | n6895 ;
  assign n7369 = x79 &  n6895 ;
  assign n7370 = ( n7368 & ~n7369 ) | ( n7368 & 1'b0 ) | ( ~n7369 & 1'b0 ) ;
  assign n7382 = ( n7026 & n7195 ) | ( n7026 & n7370 ) | ( n7195 & n7370 ) ;
  assign n7381 = n7026 | n7370 ;
  assign n7383 = ( n7380 & ~n7382 ) | ( n7380 & n7381 ) | ( ~n7382 & n7381 ) ;
  assign n7387 = n6903 &  n7194 ;
  assign n7388 = n7193 &  n7387 ;
  assign n7376 = x78 | n6903 ;
  assign n7377 = x78 &  n6903 ;
  assign n7378 = ( n7376 & ~n7377 ) | ( n7376 & 1'b0 ) | ( ~n7377 & 1'b0 ) ;
  assign n7390 = ( n7025 & n7195 ) | ( n7025 & n7378 ) | ( n7195 & n7378 ) ;
  assign n7389 = n7025 | n7378 ;
  assign n7391 = ( n7388 & ~n7390 ) | ( n7388 & n7389 ) | ( ~n7390 & n7389 ) ;
  assign n7395 = n6911 &  n7194 ;
  assign n7396 = n7193 &  n7395 ;
  assign n7384 = x77 | n6911 ;
  assign n7385 = x77 &  n6911 ;
  assign n7386 = ( n7384 & ~n7385 ) | ( n7384 & 1'b0 ) | ( ~n7385 & 1'b0 ) ;
  assign n7398 = ( n7024 & n7195 ) | ( n7024 & n7386 ) | ( n7195 & n7386 ) ;
  assign n7397 = n7024 | n7386 ;
  assign n7399 = ( n7396 & ~n7398 ) | ( n7396 & n7397 ) | ( ~n7398 & n7397 ) ;
  assign n7403 = n6919 &  n7194 ;
  assign n7404 = n7193 &  n7403 ;
  assign n7392 = x76 | n6919 ;
  assign n7393 = x76 &  n6919 ;
  assign n7394 = ( n7392 & ~n7393 ) | ( n7392 & 1'b0 ) | ( ~n7393 & 1'b0 ) ;
  assign n7406 = ( n7023 & n7195 ) | ( n7023 & n7394 ) | ( n7195 & n7394 ) ;
  assign n7405 = n7023 | n7394 ;
  assign n7407 = ( n7404 & ~n7406 ) | ( n7404 & n7405 ) | ( ~n7406 & n7405 ) ;
  assign n7411 = n6927 &  n7194 ;
  assign n7412 = n7193 &  n7411 ;
  assign n7400 = x75 | n6927 ;
  assign n7401 = x75 &  n6927 ;
  assign n7402 = ( n7400 & ~n7401 ) | ( n7400 & 1'b0 ) | ( ~n7401 & 1'b0 ) ;
  assign n7414 = ( n7022 & n7195 ) | ( n7022 & n7402 ) | ( n7195 & n7402 ) ;
  assign n7413 = n7022 | n7402 ;
  assign n7415 = ( n7412 & ~n7414 ) | ( n7412 & n7413 ) | ( ~n7414 & n7413 ) ;
  assign n7419 = n6935 &  n7194 ;
  assign n7420 = n7193 &  n7419 ;
  assign n7408 = x74 | n6935 ;
  assign n7409 = x74 &  n6935 ;
  assign n7410 = ( n7408 & ~n7409 ) | ( n7408 & 1'b0 ) | ( ~n7409 & 1'b0 ) ;
  assign n7422 = ( n7021 & n7195 ) | ( n7021 & n7410 ) | ( n7195 & n7410 ) ;
  assign n7421 = n7021 | n7410 ;
  assign n7423 = ( n7420 & ~n7422 ) | ( n7420 & n7421 ) | ( ~n7422 & n7421 ) ;
  assign n7427 = n6943 &  n7194 ;
  assign n7428 = n7193 &  n7427 ;
  assign n7416 = x73 | n6943 ;
  assign n7417 = x73 &  n6943 ;
  assign n7418 = ( n7416 & ~n7417 ) | ( n7416 & 1'b0 ) | ( ~n7417 & 1'b0 ) ;
  assign n7430 = ( n7020 & n7195 ) | ( n7020 & n7418 ) | ( n7195 & n7418 ) ;
  assign n7429 = n7020 | n7418 ;
  assign n7431 = ( n7428 & ~n7430 ) | ( n7428 & n7429 ) | ( ~n7430 & n7429 ) ;
  assign n7435 = n6951 &  n7194 ;
  assign n7436 = n7193 &  n7435 ;
  assign n7424 = x72 | n6951 ;
  assign n7425 = x72 &  n6951 ;
  assign n7426 = ( n7424 & ~n7425 ) | ( n7424 & 1'b0 ) | ( ~n7425 & 1'b0 ) ;
  assign n7438 = ( n7019 & n7195 ) | ( n7019 & n7426 ) | ( n7195 & n7426 ) ;
  assign n7437 = n7019 | n7426 ;
  assign n7439 = ( n7436 & ~n7438 ) | ( n7436 & n7437 ) | ( ~n7438 & n7437 ) ;
  assign n7443 = n6959 &  n7194 ;
  assign n7444 = n7193 &  n7443 ;
  assign n7432 = x71 | n6959 ;
  assign n7433 = x71 &  n6959 ;
  assign n7434 = ( n7432 & ~n7433 ) | ( n7432 & 1'b0 ) | ( ~n7433 & 1'b0 ) ;
  assign n7446 = ( n7018 & n7195 ) | ( n7018 & n7434 ) | ( n7195 & n7434 ) ;
  assign n7445 = n7018 | n7434 ;
  assign n7447 = ( n7444 & ~n7446 ) | ( n7444 & n7445 ) | ( ~n7446 & n7445 ) ;
  assign n7451 = n6967 &  n7194 ;
  assign n7452 = n7193 &  n7451 ;
  assign n7440 = x70 | n6967 ;
  assign n7441 = x70 &  n6967 ;
  assign n7442 = ( n7440 & ~n7441 ) | ( n7440 & 1'b0 ) | ( ~n7441 & 1'b0 ) ;
  assign n7454 = ( n7017 & n7195 ) | ( n7017 & n7442 ) | ( n7195 & n7442 ) ;
  assign n7453 = n7017 | n7442 ;
  assign n7455 = ( n7452 & ~n7454 ) | ( n7452 & n7453 ) | ( ~n7454 & n7453 ) ;
  assign n7459 = n6975 &  n7194 ;
  assign n7460 = n7193 &  n7459 ;
  assign n7448 = x69 | n6975 ;
  assign n7449 = x69 &  n6975 ;
  assign n7450 = ( n7448 & ~n7449 ) | ( n7448 & 1'b0 ) | ( ~n7449 & 1'b0 ) ;
  assign n7462 = ( n7016 & n7195 ) | ( n7016 & n7450 ) | ( n7195 & n7450 ) ;
  assign n7461 = n7016 | n7450 ;
  assign n7463 = ( n7460 & ~n7462 ) | ( n7460 & n7461 ) | ( ~n7462 & n7461 ) ;
  assign n7467 = n6983 &  n7194 ;
  assign n7468 = n7193 &  n7467 ;
  assign n7456 = x68 | n6983 ;
  assign n7457 = x68 &  n6983 ;
  assign n7458 = ( n7456 & ~n7457 ) | ( n7456 & 1'b0 ) | ( ~n7457 & 1'b0 ) ;
  assign n7470 = ( n7015 & n7195 ) | ( n7015 & n7458 ) | ( n7195 & n7458 ) ;
  assign n7469 = n7015 | n7458 ;
  assign n7471 = ( n7468 & ~n7470 ) | ( n7468 & n7469 ) | ( ~n7470 & n7469 ) ;
  assign n7475 = n6992 &  n7194 ;
  assign n7476 = n7193 &  n7475 ;
  assign n7464 = x67 | n6992 ;
  assign n7465 = x67 &  n6992 ;
  assign n7466 = ( n7464 & ~n7465 ) | ( n7464 & 1'b0 ) | ( ~n7465 & 1'b0 ) ;
  assign n7478 = ( n7014 & n7195 ) | ( n7014 & n7466 ) | ( n7195 & n7466 ) ;
  assign n7477 = n7014 | n7466 ;
  assign n7479 = ( n7476 & ~n7478 ) | ( n7476 & n7477 ) | ( ~n7478 & n7477 ) ;
  assign n7480 = n6998 &  n7194 ;
  assign n7481 = n7193 &  n7480 ;
  assign n7472 = x66 | n6998 ;
  assign n7473 = x66 &  n6998 ;
  assign n7474 = ( n7472 & ~n7473 ) | ( n7472 & 1'b0 ) | ( ~n7473 & 1'b0 ) ;
  assign n7482 = n7013 &  n7474 ;
  assign n7483 = ( n7013 & ~n7195 ) | ( n7013 & n7474 ) | ( ~n7195 & n7474 ) ;
  assign n7484 = ( n7481 & ~n7482 ) | ( n7481 & n7483 ) | ( ~n7482 & n7483 ) ;
  assign n7485 = ( n7011 & ~x65 ) | ( n7011 & n7012 ) | ( ~x65 & n7012 ) ;
  assign n7486 = ( n7013 & ~n7012 ) | ( n7013 & n7485 ) | ( ~n7012 & n7485 ) ;
  assign n7487 = ~n7195 & n7486 ;
  assign n7488 = n7011 &  n7194 ;
  assign n7489 = n7193 &  n7488 ;
  assign n7490 = n7487 | n7489 ;
  assign n7491 = ( x64 & ~n7195 ) | ( x64 & 1'b0 ) | ( ~n7195 & 1'b0 ) ;
  assign n7492 = ( x25 & ~n7491 ) | ( x25 & 1'b0 ) | ( ~n7491 & 1'b0 ) ;
  assign n7493 = ( n7012 & ~n7195 ) | ( n7012 & 1'b0 ) | ( ~n7195 & 1'b0 ) ;
  assign n7494 = n7492 | n7493 ;
  assign n7495 = ~x24 & x64 ;
  assign n7496 = ( x65 & ~n7494 ) | ( x65 & n7495 ) | ( ~n7494 & n7495 ) ;
  assign n7497 = ( x66 & ~n7490 ) | ( x66 & n7496 ) | ( ~n7490 & n7496 ) ;
  assign n7498 = ( x67 & ~n7484 ) | ( x67 & n7497 ) | ( ~n7484 & n7497 ) ;
  assign n7499 = ( x68 & ~n7479 ) | ( x68 & n7498 ) | ( ~n7479 & n7498 ) ;
  assign n7500 = ( x69 & ~n7471 ) | ( x69 & n7499 ) | ( ~n7471 & n7499 ) ;
  assign n7501 = ( x70 & ~n7463 ) | ( x70 & n7500 ) | ( ~n7463 & n7500 ) ;
  assign n7502 = ( x71 & ~n7455 ) | ( x71 & n7501 ) | ( ~n7455 & n7501 ) ;
  assign n7503 = ( x72 & ~n7447 ) | ( x72 & n7502 ) | ( ~n7447 & n7502 ) ;
  assign n7504 = ( x73 & ~n7439 ) | ( x73 & n7503 ) | ( ~n7439 & n7503 ) ;
  assign n7505 = ( x74 & ~n7431 ) | ( x74 & n7504 ) | ( ~n7431 & n7504 ) ;
  assign n7506 = ( x75 & ~n7423 ) | ( x75 & n7505 ) | ( ~n7423 & n7505 ) ;
  assign n7507 = ( x76 & ~n7415 ) | ( x76 & n7506 ) | ( ~n7415 & n7506 ) ;
  assign n7508 = ( x77 & ~n7407 ) | ( x77 & n7507 ) | ( ~n7407 & n7507 ) ;
  assign n7509 = ( x78 & ~n7399 ) | ( x78 & n7508 ) | ( ~n7399 & n7508 ) ;
  assign n7510 = ( x79 & ~n7391 ) | ( x79 & n7509 ) | ( ~n7391 & n7509 ) ;
  assign n7511 = ( x80 & ~n7383 ) | ( x80 & n7510 ) | ( ~n7383 & n7510 ) ;
  assign n7512 = ( x81 & ~n7375 ) | ( x81 & n7511 ) | ( ~n7375 & n7511 ) ;
  assign n7513 = ( x82 & ~n7367 ) | ( x82 & n7512 ) | ( ~n7367 & n7512 ) ;
  assign n7514 = ( x83 & ~n7359 ) | ( x83 & n7513 ) | ( ~n7359 & n7513 ) ;
  assign n7515 = ( x84 & ~n7351 ) | ( x84 & n7514 ) | ( ~n7351 & n7514 ) ;
  assign n7516 = ( x85 & ~n7343 ) | ( x85 & n7515 ) | ( ~n7343 & n7515 ) ;
  assign n7517 = ( x86 & ~n7335 ) | ( x86 & n7516 ) | ( ~n7335 & n7516 ) ;
  assign n7518 = ( x87 & ~n7200 ) | ( x87 & n7517 ) | ( ~n7200 & n7517 ) ;
  assign n7519 = ( x88 & ~n7327 ) | ( x88 & n7518 ) | ( ~n7327 & n7518 ) ;
  assign n7520 = ( x89 & ~n7322 ) | ( x89 & n7519 ) | ( ~n7322 & n7519 ) ;
  assign n7521 = ( x90 & ~n7314 ) | ( x90 & n7520 ) | ( ~n7314 & n7520 ) ;
  assign n7522 = ( x91 & ~n7306 ) | ( x91 & n7521 ) | ( ~n7306 & n7521 ) ;
  assign n7523 = ( x92 & ~n7298 ) | ( x92 & n7522 ) | ( ~n7298 & n7522 ) ;
  assign n7524 = ( x93 & ~n7290 ) | ( x93 & n7523 ) | ( ~n7290 & n7523 ) ;
  assign n7525 = ( x94 & ~n7282 ) | ( x94 & n7524 ) | ( ~n7282 & n7524 ) ;
  assign n7526 = ( x95 & ~n7274 ) | ( x95 & n7525 ) | ( ~n7274 & n7525 ) ;
  assign n7527 = ( x96 & ~n7266 ) | ( x96 & n7526 ) | ( ~n7266 & n7526 ) ;
  assign n7528 = ( x97 & ~n7258 ) | ( x97 & n7527 ) | ( ~n7258 & n7527 ) ;
  assign n7529 = ( x98 & ~n7250 ) | ( x98 & n7528 ) | ( ~n7250 & n7528 ) ;
  assign n7530 = ( x99 & ~n7242 ) | ( x99 & n7529 ) | ( ~n7242 & n7529 ) ;
  assign n7531 = ( x100 & ~n7234 ) | ( x100 & n7530 ) | ( ~n7234 & n7530 ) ;
  assign n7532 = ( x101 & ~n7226 ) | ( x101 & n7531 ) | ( ~n7226 & n7531 ) ;
  assign n7533 = ( x102 & ~n7218 ) | ( x102 & n7532 ) | ( ~n7218 & n7532 ) ;
  assign n7534 = ( x103 & ~n7210 ) | ( x103 & n7533 ) | ( ~n7210 & n7533 ) ;
  assign n7535 = n270 | n272 ;
  assign n7536 = n7534 | n7535 ;
  assign n7554 = n7218 &  n7536 ;
  assign n7548 = x102 | n7218 ;
  assign n7549 = x102 &  n7218 ;
  assign n7550 = ( n7548 & ~n7549 ) | ( n7548 & 1'b0 ) | ( ~n7549 & 1'b0 ) ;
  assign n7558 = ( n7532 & n7534 ) | ( n7532 & n7550 ) | ( n7534 & n7550 ) ;
  assign n7559 = ( n7532 & ~n7535 ) | ( n7532 & n7550 ) | ( ~n7535 & n7550 ) ;
  assign n7560 = ~n7558 & n7559 ;
  assign n7561 = n7554 | n7560 ;
  assign n7551 = x103 | n7533 ;
  assign n7552 = ( x103 & n7533 ) | ( x103 & n7535 ) | ( n7533 & n7535 ) ;
  assign n7553 = ( n7210 & ~n7551 ) | ( n7210 & n7552 ) | ( ~n7551 & n7552 ) ;
  assign n7562 = n7226 &  n7536 ;
  assign n7555 = x101 | n7226 ;
  assign n7556 = x101 &  n7226 ;
  assign n7557 = ( n7555 & ~n7556 ) | ( n7555 & 1'b0 ) | ( ~n7556 & 1'b0 ) ;
  assign n7566 = ( n7531 & n7534 ) | ( n7531 & n7557 ) | ( n7534 & n7557 ) ;
  assign n7567 = ( n7531 & ~n7535 ) | ( n7531 & n7557 ) | ( ~n7535 & n7557 ) ;
  assign n7568 = ~n7566 & n7567 ;
  assign n7569 = n7562 | n7568 ;
  assign n7570 = n7234 &  n7536 ;
  assign n7563 = x100 | n7234 ;
  assign n7564 = x100 &  n7234 ;
  assign n7565 = ( n7563 & ~n7564 ) | ( n7563 & 1'b0 ) | ( ~n7564 & 1'b0 ) ;
  assign n7574 = ( n7530 & n7534 ) | ( n7530 & n7565 ) | ( n7534 & n7565 ) ;
  assign n7575 = ( n7530 & ~n7535 ) | ( n7530 & n7565 ) | ( ~n7535 & n7565 ) ;
  assign n7576 = ~n7574 & n7575 ;
  assign n7577 = n7570 | n7576 ;
  assign n7578 = n7242 &  n7536 ;
  assign n7571 = x99 | n7242 ;
  assign n7572 = x99 &  n7242 ;
  assign n7573 = ( n7571 & ~n7572 ) | ( n7571 & 1'b0 ) | ( ~n7572 & 1'b0 ) ;
  assign n7582 = ( n7529 & n7534 ) | ( n7529 & n7573 ) | ( n7534 & n7573 ) ;
  assign n7583 = ( n7529 & ~n7535 ) | ( n7529 & n7573 ) | ( ~n7535 & n7573 ) ;
  assign n7584 = ~n7582 & n7583 ;
  assign n7585 = n7578 | n7584 ;
  assign n7586 = n7250 &  n7536 ;
  assign n7579 = x98 | n7250 ;
  assign n7580 = x98 &  n7250 ;
  assign n7581 = ( n7579 & ~n7580 ) | ( n7579 & 1'b0 ) | ( ~n7580 & 1'b0 ) ;
  assign n7590 = ( n7528 & n7534 ) | ( n7528 & n7581 ) | ( n7534 & n7581 ) ;
  assign n7591 = ( n7528 & ~n7535 ) | ( n7528 & n7581 ) | ( ~n7535 & n7581 ) ;
  assign n7592 = ~n7590 & n7591 ;
  assign n7593 = n7586 | n7592 ;
  assign n7594 = n7258 &  n7536 ;
  assign n7587 = x97 | n7258 ;
  assign n7588 = x97 &  n7258 ;
  assign n7589 = ( n7587 & ~n7588 ) | ( n7587 & 1'b0 ) | ( ~n7588 & 1'b0 ) ;
  assign n7598 = ( n7527 & n7534 ) | ( n7527 & n7589 ) | ( n7534 & n7589 ) ;
  assign n7599 = ( n7527 & ~n7535 ) | ( n7527 & n7589 ) | ( ~n7535 & n7589 ) ;
  assign n7600 = ~n7598 & n7599 ;
  assign n7601 = n7594 | n7600 ;
  assign n7602 = n7266 &  n7536 ;
  assign n7595 = x96 | n7266 ;
  assign n7596 = x96 &  n7266 ;
  assign n7597 = ( n7595 & ~n7596 ) | ( n7595 & 1'b0 ) | ( ~n7596 & 1'b0 ) ;
  assign n7606 = ( n7526 & n7534 ) | ( n7526 & n7597 ) | ( n7534 & n7597 ) ;
  assign n7607 = ( n7526 & ~n7535 ) | ( n7526 & n7597 ) | ( ~n7535 & n7597 ) ;
  assign n7608 = ~n7606 & n7607 ;
  assign n7609 = n7602 | n7608 ;
  assign n7610 = n7274 &  n7536 ;
  assign n7603 = x95 | n7274 ;
  assign n7604 = x95 &  n7274 ;
  assign n7605 = ( n7603 & ~n7604 ) | ( n7603 & 1'b0 ) | ( ~n7604 & 1'b0 ) ;
  assign n7614 = ( n7525 & n7534 ) | ( n7525 & n7605 ) | ( n7534 & n7605 ) ;
  assign n7615 = ( n7525 & ~n7535 ) | ( n7525 & n7605 ) | ( ~n7535 & n7605 ) ;
  assign n7616 = ~n7614 & n7615 ;
  assign n7617 = n7610 | n7616 ;
  assign n7618 = n7282 &  n7536 ;
  assign n7611 = x94 | n7282 ;
  assign n7612 = x94 &  n7282 ;
  assign n7613 = ( n7611 & ~n7612 ) | ( n7611 & 1'b0 ) | ( ~n7612 & 1'b0 ) ;
  assign n7622 = ( n7524 & n7534 ) | ( n7524 & n7613 ) | ( n7534 & n7613 ) ;
  assign n7623 = ( n7524 & ~n7535 ) | ( n7524 & n7613 ) | ( ~n7535 & n7613 ) ;
  assign n7624 = ~n7622 & n7623 ;
  assign n7625 = n7618 | n7624 ;
  assign n7626 = n7290 &  n7536 ;
  assign n7619 = x93 | n7290 ;
  assign n7620 = x93 &  n7290 ;
  assign n7621 = ( n7619 & ~n7620 ) | ( n7619 & 1'b0 ) | ( ~n7620 & 1'b0 ) ;
  assign n7630 = ( n7523 & n7534 ) | ( n7523 & n7621 ) | ( n7534 & n7621 ) ;
  assign n7631 = ( n7523 & ~n7535 ) | ( n7523 & n7621 ) | ( ~n7535 & n7621 ) ;
  assign n7632 = ~n7630 & n7631 ;
  assign n7633 = n7626 | n7632 ;
  assign n7634 = n7298 &  n7536 ;
  assign n7627 = x92 | n7298 ;
  assign n7628 = x92 &  n7298 ;
  assign n7629 = ( n7627 & ~n7628 ) | ( n7627 & 1'b0 ) | ( ~n7628 & 1'b0 ) ;
  assign n7638 = ( n7522 & n7534 ) | ( n7522 & n7629 ) | ( n7534 & n7629 ) ;
  assign n7639 = ( n7522 & ~n7535 ) | ( n7522 & n7629 ) | ( ~n7535 & n7629 ) ;
  assign n7640 = ~n7638 & n7639 ;
  assign n7641 = n7634 | n7640 ;
  assign n7642 = n7306 &  n7536 ;
  assign n7635 = x91 | n7306 ;
  assign n7636 = x91 &  n7306 ;
  assign n7637 = ( n7635 & ~n7636 ) | ( n7635 & 1'b0 ) | ( ~n7636 & 1'b0 ) ;
  assign n7646 = ( n7521 & n7534 ) | ( n7521 & n7637 ) | ( n7534 & n7637 ) ;
  assign n7647 = ( n7521 & ~n7535 ) | ( n7521 & n7637 ) | ( ~n7535 & n7637 ) ;
  assign n7648 = ~n7646 & n7647 ;
  assign n7649 = n7642 | n7648 ;
  assign n7650 = n7314 &  n7536 ;
  assign n7643 = x90 | n7314 ;
  assign n7644 = x90 &  n7314 ;
  assign n7645 = ( n7643 & ~n7644 ) | ( n7643 & 1'b0 ) | ( ~n7644 & 1'b0 ) ;
  assign n7654 = ( n7520 & n7534 ) | ( n7520 & n7645 ) | ( n7534 & n7645 ) ;
  assign n7655 = ( n7520 & ~n7535 ) | ( n7520 & n7645 ) | ( ~n7535 & n7645 ) ;
  assign n7656 = ~n7654 & n7655 ;
  assign n7657 = n7650 | n7656 ;
  assign n7658 = n7322 &  n7536 ;
  assign n7651 = x89 | n7322 ;
  assign n7652 = x89 &  n7322 ;
  assign n7653 = ( n7651 & ~n7652 ) | ( n7651 & 1'b0 ) | ( ~n7652 & 1'b0 ) ;
  assign n7662 = ( n7519 & n7534 ) | ( n7519 & n7653 ) | ( n7534 & n7653 ) ;
  assign n7663 = ( n7519 & ~n7535 ) | ( n7519 & n7653 ) | ( ~n7535 & n7653 ) ;
  assign n7664 = ~n7662 & n7663 ;
  assign n7665 = n7658 | n7664 ;
  assign n7666 = n7327 &  n7536 ;
  assign n7659 = x88 | n7327 ;
  assign n7660 = x88 &  n7327 ;
  assign n7661 = ( n7659 & ~n7660 ) | ( n7659 & 1'b0 ) | ( ~n7660 & 1'b0 ) ;
  assign n7667 = ( n7518 & n7534 ) | ( n7518 & n7661 ) | ( n7534 & n7661 ) ;
  assign n7668 = ( n7518 & ~n7535 ) | ( n7518 & n7661 ) | ( ~n7535 & n7661 ) ;
  assign n7669 = ~n7667 & n7668 ;
  assign n7670 = n7666 | n7669 ;
  assign n7537 = n7200 &  n7536 ;
  assign n7541 = x87 | n7200 ;
  assign n7542 = x87 &  n7200 ;
  assign n7543 = ( n7541 & ~n7542 ) | ( n7541 & 1'b0 ) | ( ~n7542 & 1'b0 ) ;
  assign n7544 = ( n7517 & n7534 ) | ( n7517 & n7543 ) | ( n7534 & n7543 ) ;
  assign n7545 = ( n7517 & ~n7535 ) | ( n7517 & n7543 ) | ( ~n7535 & n7543 ) ;
  assign n7546 = ~n7544 & n7545 ;
  assign n7547 = n7537 | n7546 ;
  assign n7671 = n7335 &  n7536 ;
  assign n7538 = x86 | n7335 ;
  assign n7539 = x86 &  n7335 ;
  assign n7540 = ( n7538 & ~n7539 ) | ( n7538 & 1'b0 ) | ( ~n7539 & 1'b0 ) ;
  assign n7675 = ( n7516 & n7534 ) | ( n7516 & n7540 ) | ( n7534 & n7540 ) ;
  assign n7676 = ( n7516 & ~n7535 ) | ( n7516 & n7540 ) | ( ~n7535 & n7540 ) ;
  assign n7677 = ~n7675 & n7676 ;
  assign n7678 = n7671 | n7677 ;
  assign n7679 = n7343 &  n7536 ;
  assign n7672 = x85 | n7343 ;
  assign n7673 = x85 &  n7343 ;
  assign n7674 = ( n7672 & ~n7673 ) | ( n7672 & 1'b0 ) | ( ~n7673 & 1'b0 ) ;
  assign n7683 = ( n7515 & n7534 ) | ( n7515 & n7674 ) | ( n7534 & n7674 ) ;
  assign n7684 = ( n7515 & ~n7535 ) | ( n7515 & n7674 ) | ( ~n7535 & n7674 ) ;
  assign n7685 = ~n7683 & n7684 ;
  assign n7686 = n7679 | n7685 ;
  assign n7687 = n7351 &  n7536 ;
  assign n7680 = x84 | n7351 ;
  assign n7681 = x84 &  n7351 ;
  assign n7682 = ( n7680 & ~n7681 ) | ( n7680 & 1'b0 ) | ( ~n7681 & 1'b0 ) ;
  assign n7691 = ( n7514 & n7534 ) | ( n7514 & n7682 ) | ( n7534 & n7682 ) ;
  assign n7692 = ( n7514 & ~n7535 ) | ( n7514 & n7682 ) | ( ~n7535 & n7682 ) ;
  assign n7693 = ~n7691 & n7692 ;
  assign n7694 = n7687 | n7693 ;
  assign n7695 = n7359 &  n7536 ;
  assign n7688 = x83 | n7359 ;
  assign n7689 = x83 &  n7359 ;
  assign n7690 = ( n7688 & ~n7689 ) | ( n7688 & 1'b0 ) | ( ~n7689 & 1'b0 ) ;
  assign n7699 = ( n7513 & n7534 ) | ( n7513 & n7690 ) | ( n7534 & n7690 ) ;
  assign n7700 = ( n7513 & ~n7535 ) | ( n7513 & n7690 ) | ( ~n7535 & n7690 ) ;
  assign n7701 = ~n7699 & n7700 ;
  assign n7702 = n7695 | n7701 ;
  assign n7703 = n7367 &  n7536 ;
  assign n7696 = x82 | n7367 ;
  assign n7697 = x82 &  n7367 ;
  assign n7698 = ( n7696 & ~n7697 ) | ( n7696 & 1'b0 ) | ( ~n7697 & 1'b0 ) ;
  assign n7707 = ( n7512 & n7534 ) | ( n7512 & n7698 ) | ( n7534 & n7698 ) ;
  assign n7708 = ( n7512 & ~n7535 ) | ( n7512 & n7698 ) | ( ~n7535 & n7698 ) ;
  assign n7709 = ~n7707 & n7708 ;
  assign n7710 = n7703 | n7709 ;
  assign n7711 = n7375 &  n7536 ;
  assign n7704 = x81 | n7375 ;
  assign n7705 = x81 &  n7375 ;
  assign n7706 = ( n7704 & ~n7705 ) | ( n7704 & 1'b0 ) | ( ~n7705 & 1'b0 ) ;
  assign n7715 = ( n7511 & n7534 ) | ( n7511 & n7706 ) | ( n7534 & n7706 ) ;
  assign n7716 = ( n7511 & ~n7535 ) | ( n7511 & n7706 ) | ( ~n7535 & n7706 ) ;
  assign n7717 = ~n7715 & n7716 ;
  assign n7718 = n7711 | n7717 ;
  assign n7719 = n7383 &  n7536 ;
  assign n7712 = x80 | n7383 ;
  assign n7713 = x80 &  n7383 ;
  assign n7714 = ( n7712 & ~n7713 ) | ( n7712 & 1'b0 ) | ( ~n7713 & 1'b0 ) ;
  assign n7723 = ( n7510 & n7534 ) | ( n7510 & n7714 ) | ( n7534 & n7714 ) ;
  assign n7724 = ( n7510 & ~n7535 ) | ( n7510 & n7714 ) | ( ~n7535 & n7714 ) ;
  assign n7725 = ~n7723 & n7724 ;
  assign n7726 = n7719 | n7725 ;
  assign n7727 = n7391 &  n7536 ;
  assign n7720 = x79 | n7391 ;
  assign n7721 = x79 &  n7391 ;
  assign n7722 = ( n7720 & ~n7721 ) | ( n7720 & 1'b0 ) | ( ~n7721 & 1'b0 ) ;
  assign n7731 = ( n7509 & n7534 ) | ( n7509 & n7722 ) | ( n7534 & n7722 ) ;
  assign n7732 = ( n7509 & ~n7535 ) | ( n7509 & n7722 ) | ( ~n7535 & n7722 ) ;
  assign n7733 = ~n7731 & n7732 ;
  assign n7734 = n7727 | n7733 ;
  assign n7735 = n7399 &  n7536 ;
  assign n7728 = x78 | n7399 ;
  assign n7729 = x78 &  n7399 ;
  assign n7730 = ( n7728 & ~n7729 ) | ( n7728 & 1'b0 ) | ( ~n7729 & 1'b0 ) ;
  assign n7739 = ( n7508 & n7534 ) | ( n7508 & n7730 ) | ( n7534 & n7730 ) ;
  assign n7740 = ( n7508 & ~n7535 ) | ( n7508 & n7730 ) | ( ~n7535 & n7730 ) ;
  assign n7741 = ~n7739 & n7740 ;
  assign n7742 = n7735 | n7741 ;
  assign n7743 = n7407 &  n7536 ;
  assign n7736 = x77 | n7407 ;
  assign n7737 = x77 &  n7407 ;
  assign n7738 = ( n7736 & ~n7737 ) | ( n7736 & 1'b0 ) | ( ~n7737 & 1'b0 ) ;
  assign n7747 = ( n7507 & n7534 ) | ( n7507 & n7738 ) | ( n7534 & n7738 ) ;
  assign n7748 = ( n7507 & ~n7535 ) | ( n7507 & n7738 ) | ( ~n7535 & n7738 ) ;
  assign n7749 = ~n7747 & n7748 ;
  assign n7750 = n7743 | n7749 ;
  assign n7751 = n7415 &  n7536 ;
  assign n7744 = x76 | n7415 ;
  assign n7745 = x76 &  n7415 ;
  assign n7746 = ( n7744 & ~n7745 ) | ( n7744 & 1'b0 ) | ( ~n7745 & 1'b0 ) ;
  assign n7755 = ( n7506 & n7534 ) | ( n7506 & n7746 ) | ( n7534 & n7746 ) ;
  assign n7756 = ( n7506 & ~n7535 ) | ( n7506 & n7746 ) | ( ~n7535 & n7746 ) ;
  assign n7757 = ~n7755 & n7756 ;
  assign n7758 = n7751 | n7757 ;
  assign n7759 = n7423 &  n7536 ;
  assign n7752 = x75 | n7423 ;
  assign n7753 = x75 &  n7423 ;
  assign n7754 = ( n7752 & ~n7753 ) | ( n7752 & 1'b0 ) | ( ~n7753 & 1'b0 ) ;
  assign n7763 = ( n7505 & n7534 ) | ( n7505 & n7754 ) | ( n7534 & n7754 ) ;
  assign n7764 = ( n7505 & ~n7535 ) | ( n7505 & n7754 ) | ( ~n7535 & n7754 ) ;
  assign n7765 = ~n7763 & n7764 ;
  assign n7766 = n7759 | n7765 ;
  assign n7767 = n7431 &  n7536 ;
  assign n7760 = x74 | n7431 ;
  assign n7761 = x74 &  n7431 ;
  assign n7762 = ( n7760 & ~n7761 ) | ( n7760 & 1'b0 ) | ( ~n7761 & 1'b0 ) ;
  assign n7771 = ( n7504 & n7534 ) | ( n7504 & n7762 ) | ( n7534 & n7762 ) ;
  assign n7772 = ( n7504 & ~n7535 ) | ( n7504 & n7762 ) | ( ~n7535 & n7762 ) ;
  assign n7773 = ~n7771 & n7772 ;
  assign n7774 = n7767 | n7773 ;
  assign n7775 = n7439 &  n7536 ;
  assign n7768 = x73 | n7439 ;
  assign n7769 = x73 &  n7439 ;
  assign n7770 = ( n7768 & ~n7769 ) | ( n7768 & 1'b0 ) | ( ~n7769 & 1'b0 ) ;
  assign n7779 = ( n7503 & n7534 ) | ( n7503 & n7770 ) | ( n7534 & n7770 ) ;
  assign n7780 = ( n7503 & ~n7535 ) | ( n7503 & n7770 ) | ( ~n7535 & n7770 ) ;
  assign n7781 = ~n7779 & n7780 ;
  assign n7782 = n7775 | n7781 ;
  assign n7783 = n7447 &  n7536 ;
  assign n7776 = x72 | n7447 ;
  assign n7777 = x72 &  n7447 ;
  assign n7778 = ( n7776 & ~n7777 ) | ( n7776 & 1'b0 ) | ( ~n7777 & 1'b0 ) ;
  assign n7787 = ( n7502 & n7534 ) | ( n7502 & n7778 ) | ( n7534 & n7778 ) ;
  assign n7788 = ( n7502 & ~n7535 ) | ( n7502 & n7778 ) | ( ~n7535 & n7778 ) ;
  assign n7789 = ~n7787 & n7788 ;
  assign n7790 = n7783 | n7789 ;
  assign n7791 = n7455 &  n7536 ;
  assign n7784 = x71 | n7455 ;
  assign n7785 = x71 &  n7455 ;
  assign n7786 = ( n7784 & ~n7785 ) | ( n7784 & 1'b0 ) | ( ~n7785 & 1'b0 ) ;
  assign n7795 = ( n7501 & n7534 ) | ( n7501 & n7786 ) | ( n7534 & n7786 ) ;
  assign n7796 = ( n7501 & ~n7535 ) | ( n7501 & n7786 ) | ( ~n7535 & n7786 ) ;
  assign n7797 = ~n7795 & n7796 ;
  assign n7798 = n7791 | n7797 ;
  assign n7799 = n7463 &  n7536 ;
  assign n7792 = x70 | n7463 ;
  assign n7793 = x70 &  n7463 ;
  assign n7794 = ( n7792 & ~n7793 ) | ( n7792 & 1'b0 ) | ( ~n7793 & 1'b0 ) ;
  assign n7803 = ( n7500 & n7534 ) | ( n7500 & n7794 ) | ( n7534 & n7794 ) ;
  assign n7804 = ( n7500 & ~n7535 ) | ( n7500 & n7794 ) | ( ~n7535 & n7794 ) ;
  assign n7805 = ~n7803 & n7804 ;
  assign n7806 = n7799 | n7805 ;
  assign n7807 = n7471 &  n7536 ;
  assign n7800 = x69 | n7471 ;
  assign n7801 = x69 &  n7471 ;
  assign n7802 = ( n7800 & ~n7801 ) | ( n7800 & 1'b0 ) | ( ~n7801 & 1'b0 ) ;
  assign n7811 = ( n7499 & n7534 ) | ( n7499 & n7802 ) | ( n7534 & n7802 ) ;
  assign n7812 = ( n7499 & ~n7535 ) | ( n7499 & n7802 ) | ( ~n7535 & n7802 ) ;
  assign n7813 = ~n7811 & n7812 ;
  assign n7814 = n7807 | n7813 ;
  assign n7815 = n7479 &  n7536 ;
  assign n7808 = x68 | n7479 ;
  assign n7809 = x68 &  n7479 ;
  assign n7810 = ( n7808 & ~n7809 ) | ( n7808 & 1'b0 ) | ( ~n7809 & 1'b0 ) ;
  assign n7819 = ( n7498 & n7534 ) | ( n7498 & n7810 ) | ( n7534 & n7810 ) ;
  assign n7820 = ( n7498 & ~n7535 ) | ( n7498 & n7810 ) | ( ~n7535 & n7810 ) ;
  assign n7821 = ~n7819 & n7820 ;
  assign n7822 = n7815 | n7821 ;
  assign n7823 = n7484 &  n7536 ;
  assign n7816 = x67 | n7484 ;
  assign n7817 = x67 &  n7484 ;
  assign n7818 = ( n7816 & ~n7817 ) | ( n7816 & 1'b0 ) | ( ~n7817 & 1'b0 ) ;
  assign n7827 = ( n7497 & n7534 ) | ( n7497 & n7818 ) | ( n7534 & n7818 ) ;
  assign n7828 = ( n7497 & ~n7535 ) | ( n7497 & n7818 ) | ( ~n7535 & n7818 ) ;
  assign n7829 = ~n7827 & n7828 ;
  assign n7830 = n7823 | n7829 ;
  assign n7831 = n7490 &  n7536 ;
  assign n7824 = x66 | n7490 ;
  assign n7825 = x66 &  n7490 ;
  assign n7826 = ( n7824 & ~n7825 ) | ( n7824 & 1'b0 ) | ( ~n7825 & 1'b0 ) ;
  assign n7836 = ( n7496 & ~n7534 ) | ( n7496 & n7826 ) | ( ~n7534 & n7826 ) ;
  assign n7837 = ( n7496 & n7535 ) | ( n7496 & n7826 ) | ( n7535 & n7826 ) ;
  assign n7838 = ( n7836 & ~n7837 ) | ( n7836 & 1'b0 ) | ( ~n7837 & 1'b0 ) ;
  assign n7839 = n7831 | n7838 ;
  assign n7840 = n7494 &  n7536 ;
  assign n7832 = x65 &  n7494 ;
  assign n7833 = ( n7492 & ~x65 ) | ( n7492 & n7493 ) | ( ~x65 & n7493 ) ;
  assign n7834 = x65 | n7833 ;
  assign n7835 = ( n7495 & ~n7832 ) | ( n7495 & n7834 ) | ( ~n7832 & n7834 ) ;
  assign n7841 = ( x65 & n7494 ) | ( x65 & n7495 ) | ( n7494 & n7495 ) ;
  assign n7842 = ( n7535 & ~n7832 ) | ( n7535 & n7841 ) | ( ~n7832 & n7841 ) ;
  assign n7843 = ( n7534 & n7835 ) | ( n7534 & n7842 ) | ( n7835 & n7842 ) ;
  assign n7844 = ( n7835 & ~n7843 ) | ( n7835 & 1'b0 ) | ( ~n7843 & 1'b0 ) ;
  assign n7845 = n7840 | n7844 ;
  assign n7846 = ( x64 & ~x104 ) | ( x64 & 1'b0 ) | ( ~x104 & 1'b0 ) ;
  assign n7847 = ( n253 & ~n427 ) | ( n253 & n7846 ) | ( ~n427 & n7846 ) ;
  assign n7848 = ~n253 & n7847 ;
  assign n7849 = ~n425 & n7848 ;
  assign n7850 = n7534 &  n7849 ;
  assign n7851 = ( x24 & ~n7849 ) | ( x24 & n7850 ) | ( ~n7849 & n7850 ) ;
  assign n7852 = ~n163 & n7495 ;
  assign n7853 = ( n160 & ~n174 ) | ( n160 & n7852 ) | ( ~n174 & n7852 ) ;
  assign n7854 = ~n160 & n7853 ;
  assign n7855 = ~n7534 & n7854 ;
  assign n7856 = n7851 | n7855 ;
  assign n7857 = ~x23 & x64 ;
  assign n7858 = ( x65 & ~n7856 ) | ( x65 & n7857 ) | ( ~n7856 & n7857 ) ;
  assign n7859 = ( x66 & ~n7845 ) | ( x66 & n7858 ) | ( ~n7845 & n7858 ) ;
  assign n7860 = ( x67 & ~n7839 ) | ( x67 & n7859 ) | ( ~n7839 & n7859 ) ;
  assign n7861 = ( x68 & ~n7830 ) | ( x68 & n7860 ) | ( ~n7830 & n7860 ) ;
  assign n7862 = ( x69 & ~n7822 ) | ( x69 & n7861 ) | ( ~n7822 & n7861 ) ;
  assign n7863 = ( x70 & ~n7814 ) | ( x70 & n7862 ) | ( ~n7814 & n7862 ) ;
  assign n7864 = ( x71 & ~n7806 ) | ( x71 & n7863 ) | ( ~n7806 & n7863 ) ;
  assign n7865 = ( x72 & ~n7798 ) | ( x72 & n7864 ) | ( ~n7798 & n7864 ) ;
  assign n7866 = ( x73 & ~n7790 ) | ( x73 & n7865 ) | ( ~n7790 & n7865 ) ;
  assign n7867 = ( x74 & ~n7782 ) | ( x74 & n7866 ) | ( ~n7782 & n7866 ) ;
  assign n7868 = ( x75 & ~n7774 ) | ( x75 & n7867 ) | ( ~n7774 & n7867 ) ;
  assign n7869 = ( x76 & ~n7766 ) | ( x76 & n7868 ) | ( ~n7766 & n7868 ) ;
  assign n7870 = ( x77 & ~n7758 ) | ( x77 & n7869 ) | ( ~n7758 & n7869 ) ;
  assign n7871 = ( x78 & ~n7750 ) | ( x78 & n7870 ) | ( ~n7750 & n7870 ) ;
  assign n7872 = ( x79 & ~n7742 ) | ( x79 & n7871 ) | ( ~n7742 & n7871 ) ;
  assign n7873 = ( x80 & ~n7734 ) | ( x80 & n7872 ) | ( ~n7734 & n7872 ) ;
  assign n7874 = ( x81 & ~n7726 ) | ( x81 & n7873 ) | ( ~n7726 & n7873 ) ;
  assign n7875 = ( x82 & ~n7718 ) | ( x82 & n7874 ) | ( ~n7718 & n7874 ) ;
  assign n7876 = ( x83 & ~n7710 ) | ( x83 & n7875 ) | ( ~n7710 & n7875 ) ;
  assign n7877 = ( x84 & ~n7702 ) | ( x84 & n7876 ) | ( ~n7702 & n7876 ) ;
  assign n7878 = ( x85 & ~n7694 ) | ( x85 & n7877 ) | ( ~n7694 & n7877 ) ;
  assign n7879 = ( x86 & ~n7686 ) | ( x86 & n7878 ) | ( ~n7686 & n7878 ) ;
  assign n7880 = ( x87 & ~n7678 ) | ( x87 & n7879 ) | ( ~n7678 & n7879 ) ;
  assign n7881 = ( x88 & ~n7547 ) | ( x88 & n7880 ) | ( ~n7547 & n7880 ) ;
  assign n7882 = ( x89 & ~n7670 ) | ( x89 & n7881 ) | ( ~n7670 & n7881 ) ;
  assign n7883 = ( x90 & ~n7665 ) | ( x90 & n7882 ) | ( ~n7665 & n7882 ) ;
  assign n7884 = ( x91 & ~n7657 ) | ( x91 & n7883 ) | ( ~n7657 & n7883 ) ;
  assign n7885 = ( x92 & ~n7649 ) | ( x92 & n7884 ) | ( ~n7649 & n7884 ) ;
  assign n7886 = ( x93 & ~n7641 ) | ( x93 & n7885 ) | ( ~n7641 & n7885 ) ;
  assign n7887 = ( x94 & ~n7633 ) | ( x94 & n7886 ) | ( ~n7633 & n7886 ) ;
  assign n7888 = ( x95 & ~n7625 ) | ( x95 & n7887 ) | ( ~n7625 & n7887 ) ;
  assign n7889 = ( x96 & ~n7617 ) | ( x96 & n7888 ) | ( ~n7617 & n7888 ) ;
  assign n7890 = ( x97 & ~n7609 ) | ( x97 & n7889 ) | ( ~n7609 & n7889 ) ;
  assign n7891 = ( x98 & ~n7601 ) | ( x98 & n7890 ) | ( ~n7601 & n7890 ) ;
  assign n7892 = ( x99 & ~n7593 ) | ( x99 & n7891 ) | ( ~n7593 & n7891 ) ;
  assign n7893 = ( x100 & ~n7585 ) | ( x100 & n7892 ) | ( ~n7585 & n7892 ) ;
  assign n7894 = ( x101 & ~n7577 ) | ( x101 & n7893 ) | ( ~n7577 & n7893 ) ;
  assign n7895 = ( x102 & ~n7569 ) | ( x102 & n7894 ) | ( ~n7569 & n7894 ) ;
  assign n7896 = ( x103 & ~n7561 ) | ( x103 & n7895 ) | ( ~n7561 & n7895 ) ;
  assign n7897 = ( x104 & ~n7553 ) | ( x104 & n7896 ) | ( ~n7553 & n7896 ) ;
  assign n7898 = n240 | n254 ;
  assign n7899 = n7897 | n7898 ;
  assign n8145 = n7561 &  n7899 ;
  assign n8149 = x103 | n7561 ;
  assign n8150 = x103 &  n7561 ;
  assign n8151 = ( n8149 & ~n8150 ) | ( n8149 & 1'b0 ) | ( ~n8150 & 1'b0 ) ;
  assign n8152 = ( n7895 & n7897 ) | ( n7895 & n8151 ) | ( n7897 & n8151 ) ;
  assign n8153 = ( n7895 & ~n7898 ) | ( n7895 & n8151 ) | ( ~n7898 & n8151 ) ;
  assign n8154 = ~n8152 & n8153 ;
  assign n8155 = n8145 | n8154 ;
  assign n8156 = n7569 &  n7899 ;
  assign n8146 = x102 | n7569 ;
  assign n8147 = x102 &  n7569 ;
  assign n8148 = ( n8146 & ~n8147 ) | ( n8146 & 1'b0 ) | ( ~n8147 & 1'b0 ) ;
  assign n8160 = ( n7894 & n7897 ) | ( n7894 & n8148 ) | ( n7897 & n8148 ) ;
  assign n8161 = ( n7894 & ~n7898 ) | ( n7894 & n8148 ) | ( ~n7898 & n8148 ) ;
  assign n8162 = ~n8160 & n8161 ;
  assign n8163 = n8156 | n8162 ;
  assign n8164 = n7577 &  n7899 ;
  assign n8157 = x101 | n7577 ;
  assign n8158 = x101 &  n7577 ;
  assign n8159 = ( n8157 & ~n8158 ) | ( n8157 & 1'b0 ) | ( ~n8158 & 1'b0 ) ;
  assign n8168 = ( n7893 & n7897 ) | ( n7893 & n8159 ) | ( n7897 & n8159 ) ;
  assign n8169 = ( n7893 & ~n7898 ) | ( n7893 & n8159 ) | ( ~n7898 & n8159 ) ;
  assign n8170 = ~n8168 & n8169 ;
  assign n8171 = n8164 | n8170 ;
  assign n8172 = n7585 &  n7899 ;
  assign n8165 = x100 | n7585 ;
  assign n8166 = x100 &  n7585 ;
  assign n8167 = ( n8165 & ~n8166 ) | ( n8165 & 1'b0 ) | ( ~n8166 & 1'b0 ) ;
  assign n8176 = ( n7892 & n7897 ) | ( n7892 & n8167 ) | ( n7897 & n8167 ) ;
  assign n8177 = ( n7892 & ~n7898 ) | ( n7892 & n8167 ) | ( ~n7898 & n8167 ) ;
  assign n8178 = ~n8176 & n8177 ;
  assign n8179 = n8172 | n8178 ;
  assign n8180 = n7593 &  n7899 ;
  assign n8173 = x99 | n7593 ;
  assign n8174 = x99 &  n7593 ;
  assign n8175 = ( n8173 & ~n8174 ) | ( n8173 & 1'b0 ) | ( ~n8174 & 1'b0 ) ;
  assign n8184 = ( n7891 & n7897 ) | ( n7891 & n8175 ) | ( n7897 & n8175 ) ;
  assign n8185 = ( n7891 & ~n7898 ) | ( n7891 & n8175 ) | ( ~n7898 & n8175 ) ;
  assign n8186 = ~n8184 & n8185 ;
  assign n8187 = n8180 | n8186 ;
  assign n8188 = n7601 &  n7899 ;
  assign n8181 = x98 | n7601 ;
  assign n8182 = x98 &  n7601 ;
  assign n8183 = ( n8181 & ~n8182 ) | ( n8181 & 1'b0 ) | ( ~n8182 & 1'b0 ) ;
  assign n8192 = ( n7890 & n7897 ) | ( n7890 & n8183 ) | ( n7897 & n8183 ) ;
  assign n8193 = ( n7890 & ~n7898 ) | ( n7890 & n8183 ) | ( ~n7898 & n8183 ) ;
  assign n8194 = ~n8192 & n8193 ;
  assign n8195 = n8188 | n8194 ;
  assign n8196 = n7609 &  n7899 ;
  assign n8189 = x97 | n7609 ;
  assign n8190 = x97 &  n7609 ;
  assign n8191 = ( n8189 & ~n8190 ) | ( n8189 & 1'b0 ) | ( ~n8190 & 1'b0 ) ;
  assign n8200 = ( n7889 & n7897 ) | ( n7889 & n8191 ) | ( n7897 & n8191 ) ;
  assign n8201 = ( n7889 & ~n7898 ) | ( n7889 & n8191 ) | ( ~n7898 & n8191 ) ;
  assign n8202 = ~n8200 & n8201 ;
  assign n8203 = n8196 | n8202 ;
  assign n8204 = n7617 &  n7899 ;
  assign n8197 = x96 | n7617 ;
  assign n8198 = x96 &  n7617 ;
  assign n8199 = ( n8197 & ~n8198 ) | ( n8197 & 1'b0 ) | ( ~n8198 & 1'b0 ) ;
  assign n8208 = ( n7888 & n7897 ) | ( n7888 & n8199 ) | ( n7897 & n8199 ) ;
  assign n8209 = ( n7888 & ~n7898 ) | ( n7888 & n8199 ) | ( ~n7898 & n8199 ) ;
  assign n8210 = ~n8208 & n8209 ;
  assign n8211 = n8204 | n8210 ;
  assign n8212 = n7625 &  n7899 ;
  assign n8205 = x95 | n7625 ;
  assign n8206 = x95 &  n7625 ;
  assign n8207 = ( n8205 & ~n8206 ) | ( n8205 & 1'b0 ) | ( ~n8206 & 1'b0 ) ;
  assign n8216 = ( n7887 & n7897 ) | ( n7887 & n8207 ) | ( n7897 & n8207 ) ;
  assign n8217 = ( n7887 & ~n7898 ) | ( n7887 & n8207 ) | ( ~n7898 & n8207 ) ;
  assign n8218 = ~n8216 & n8217 ;
  assign n8219 = n8212 | n8218 ;
  assign n8220 = n7633 &  n7899 ;
  assign n8213 = x94 | n7633 ;
  assign n8214 = x94 &  n7633 ;
  assign n8215 = ( n8213 & ~n8214 ) | ( n8213 & 1'b0 ) | ( ~n8214 & 1'b0 ) ;
  assign n8224 = ( n7886 & n7897 ) | ( n7886 & n8215 ) | ( n7897 & n8215 ) ;
  assign n8225 = ( n7886 & ~n7898 ) | ( n7886 & n8215 ) | ( ~n7898 & n8215 ) ;
  assign n8226 = ~n8224 & n8225 ;
  assign n8227 = n8220 | n8226 ;
  assign n8228 = n7641 &  n7899 ;
  assign n8221 = x93 | n7641 ;
  assign n8222 = x93 &  n7641 ;
  assign n8223 = ( n8221 & ~n8222 ) | ( n8221 & 1'b0 ) | ( ~n8222 & 1'b0 ) ;
  assign n8232 = ( n7885 & n7897 ) | ( n7885 & n8223 ) | ( n7897 & n8223 ) ;
  assign n8233 = ( n7885 & ~n7898 ) | ( n7885 & n8223 ) | ( ~n7898 & n8223 ) ;
  assign n8234 = ~n8232 & n8233 ;
  assign n8235 = n8228 | n8234 ;
  assign n8236 = n7649 &  n7899 ;
  assign n8229 = x92 | n7649 ;
  assign n8230 = x92 &  n7649 ;
  assign n8231 = ( n8229 & ~n8230 ) | ( n8229 & 1'b0 ) | ( ~n8230 & 1'b0 ) ;
  assign n8240 = ( n7884 & n7897 ) | ( n7884 & n8231 ) | ( n7897 & n8231 ) ;
  assign n8241 = ( n7884 & ~n7898 ) | ( n7884 & n8231 ) | ( ~n7898 & n8231 ) ;
  assign n8242 = ~n8240 & n8241 ;
  assign n8243 = n8236 | n8242 ;
  assign n8244 = n7657 &  n7899 ;
  assign n8237 = x91 | n7657 ;
  assign n8238 = x91 &  n7657 ;
  assign n8239 = ( n8237 & ~n8238 ) | ( n8237 & 1'b0 ) | ( ~n8238 & 1'b0 ) ;
  assign n8248 = ( n7883 & n7897 ) | ( n7883 & n8239 ) | ( n7897 & n8239 ) ;
  assign n8249 = ( n7883 & ~n7898 ) | ( n7883 & n8239 ) | ( ~n7898 & n8239 ) ;
  assign n8250 = ~n8248 & n8249 ;
  assign n8251 = n8244 | n8250 ;
  assign n8252 = n7665 &  n7899 ;
  assign n8245 = x90 | n7665 ;
  assign n8246 = x90 &  n7665 ;
  assign n8247 = ( n8245 & ~n8246 ) | ( n8245 & 1'b0 ) | ( ~n8246 & 1'b0 ) ;
  assign n8253 = ( n7882 & n7897 ) | ( n7882 & n8247 ) | ( n7897 & n8247 ) ;
  assign n8254 = ( n7882 & ~n7898 ) | ( n7882 & n8247 ) | ( ~n7898 & n8247 ) ;
  assign n8255 = ~n8253 & n8254 ;
  assign n8256 = n8252 | n8255 ;
  assign n8134 = n7670 &  n7899 ;
  assign n8135 = x89 | n7670 ;
  assign n8136 = x89 &  n7670 ;
  assign n8137 = ( n8135 & ~n8136 ) | ( n8135 & 1'b0 ) | ( ~n8136 & 1'b0 ) ;
  assign n8138 = ( n7881 & n7897 ) | ( n7881 & n8137 ) | ( n7897 & n8137 ) ;
  assign n8139 = ( n7881 & ~n7898 ) | ( n7881 & n8137 ) | ( ~n7898 & n8137 ) ;
  assign n8140 = ~n8138 & n8139 ;
  assign n8141 = n8134 | n8140 ;
  assign n7900 = n7547 &  n7899 ;
  assign n7904 = x88 | n7547 ;
  assign n7905 = x88 &  n7547 ;
  assign n7906 = ( n7904 & ~n7905 ) | ( n7904 & 1'b0 ) | ( ~n7905 & 1'b0 ) ;
  assign n7907 = ( n7880 & n7897 ) | ( n7880 & n7906 ) | ( n7897 & n7906 ) ;
  assign n7908 = ( n7880 & ~n7898 ) | ( n7880 & n7906 ) | ( ~n7898 & n7906 ) ;
  assign n7909 = ~n7907 & n7908 ;
  assign n7910 = n7900 | n7909 ;
  assign n7911 = n7678 &  n7899 ;
  assign n7901 = x87 | n7678 ;
  assign n7902 = x87 &  n7678 ;
  assign n7903 = ( n7901 & ~n7902 ) | ( n7901 & 1'b0 ) | ( ~n7902 & 1'b0 ) ;
  assign n7915 = ( n7879 & n7897 ) | ( n7879 & n7903 ) | ( n7897 & n7903 ) ;
  assign n7916 = ( n7879 & ~n7898 ) | ( n7879 & n7903 ) | ( ~n7898 & n7903 ) ;
  assign n7917 = ~n7915 & n7916 ;
  assign n7918 = n7911 | n7917 ;
  assign n7919 = n7686 &  n7899 ;
  assign n7912 = x86 | n7686 ;
  assign n7913 = x86 &  n7686 ;
  assign n7914 = ( n7912 & ~n7913 ) | ( n7912 & 1'b0 ) | ( ~n7913 & 1'b0 ) ;
  assign n7923 = ( n7878 & n7897 ) | ( n7878 & n7914 ) | ( n7897 & n7914 ) ;
  assign n7924 = ( n7878 & ~n7898 ) | ( n7878 & n7914 ) | ( ~n7898 & n7914 ) ;
  assign n7925 = ~n7923 & n7924 ;
  assign n7926 = n7919 | n7925 ;
  assign n7927 = n7694 &  n7899 ;
  assign n7920 = x85 | n7694 ;
  assign n7921 = x85 &  n7694 ;
  assign n7922 = ( n7920 & ~n7921 ) | ( n7920 & 1'b0 ) | ( ~n7921 & 1'b0 ) ;
  assign n7931 = ( n7877 & n7897 ) | ( n7877 & n7922 ) | ( n7897 & n7922 ) ;
  assign n7932 = ( n7877 & ~n7898 ) | ( n7877 & n7922 ) | ( ~n7898 & n7922 ) ;
  assign n7933 = ~n7931 & n7932 ;
  assign n7934 = n7927 | n7933 ;
  assign n7935 = n7702 &  n7899 ;
  assign n7928 = x84 | n7702 ;
  assign n7929 = x84 &  n7702 ;
  assign n7930 = ( n7928 & ~n7929 ) | ( n7928 & 1'b0 ) | ( ~n7929 & 1'b0 ) ;
  assign n7939 = ( n7876 & n7897 ) | ( n7876 & n7930 ) | ( n7897 & n7930 ) ;
  assign n7940 = ( n7876 & ~n7898 ) | ( n7876 & n7930 ) | ( ~n7898 & n7930 ) ;
  assign n7941 = ~n7939 & n7940 ;
  assign n7942 = n7935 | n7941 ;
  assign n7943 = n7710 &  n7899 ;
  assign n7936 = x83 | n7710 ;
  assign n7937 = x83 &  n7710 ;
  assign n7938 = ( n7936 & ~n7937 ) | ( n7936 & 1'b0 ) | ( ~n7937 & 1'b0 ) ;
  assign n7947 = ( n7875 & n7897 ) | ( n7875 & n7938 ) | ( n7897 & n7938 ) ;
  assign n7948 = ( n7875 & ~n7898 ) | ( n7875 & n7938 ) | ( ~n7898 & n7938 ) ;
  assign n7949 = ~n7947 & n7948 ;
  assign n7950 = n7943 | n7949 ;
  assign n7951 = n7718 &  n7899 ;
  assign n7944 = x82 | n7718 ;
  assign n7945 = x82 &  n7718 ;
  assign n7946 = ( n7944 & ~n7945 ) | ( n7944 & 1'b0 ) | ( ~n7945 & 1'b0 ) ;
  assign n7955 = ( n7874 & n7897 ) | ( n7874 & n7946 ) | ( n7897 & n7946 ) ;
  assign n7956 = ( n7874 & ~n7898 ) | ( n7874 & n7946 ) | ( ~n7898 & n7946 ) ;
  assign n7957 = ~n7955 & n7956 ;
  assign n7958 = n7951 | n7957 ;
  assign n7959 = n7726 &  n7899 ;
  assign n7952 = x81 | n7726 ;
  assign n7953 = x81 &  n7726 ;
  assign n7954 = ( n7952 & ~n7953 ) | ( n7952 & 1'b0 ) | ( ~n7953 & 1'b0 ) ;
  assign n7963 = ( n7873 & n7897 ) | ( n7873 & n7954 ) | ( n7897 & n7954 ) ;
  assign n7964 = ( n7873 & ~n7898 ) | ( n7873 & n7954 ) | ( ~n7898 & n7954 ) ;
  assign n7965 = ~n7963 & n7964 ;
  assign n7966 = n7959 | n7965 ;
  assign n7967 = n7734 &  n7899 ;
  assign n7960 = x80 | n7734 ;
  assign n7961 = x80 &  n7734 ;
  assign n7962 = ( n7960 & ~n7961 ) | ( n7960 & 1'b0 ) | ( ~n7961 & 1'b0 ) ;
  assign n7971 = ( n7872 & n7897 ) | ( n7872 & n7962 ) | ( n7897 & n7962 ) ;
  assign n7972 = ( n7872 & ~n7898 ) | ( n7872 & n7962 ) | ( ~n7898 & n7962 ) ;
  assign n7973 = ~n7971 & n7972 ;
  assign n7974 = n7967 | n7973 ;
  assign n7975 = n7742 &  n7899 ;
  assign n7968 = x79 | n7742 ;
  assign n7969 = x79 &  n7742 ;
  assign n7970 = ( n7968 & ~n7969 ) | ( n7968 & 1'b0 ) | ( ~n7969 & 1'b0 ) ;
  assign n7979 = ( n7871 & n7897 ) | ( n7871 & n7970 ) | ( n7897 & n7970 ) ;
  assign n7980 = ( n7871 & ~n7898 ) | ( n7871 & n7970 ) | ( ~n7898 & n7970 ) ;
  assign n7981 = ~n7979 & n7980 ;
  assign n7982 = n7975 | n7981 ;
  assign n7983 = n7750 &  n7899 ;
  assign n7976 = x78 | n7750 ;
  assign n7977 = x78 &  n7750 ;
  assign n7978 = ( n7976 & ~n7977 ) | ( n7976 & 1'b0 ) | ( ~n7977 & 1'b0 ) ;
  assign n7987 = ( n7870 & n7897 ) | ( n7870 & n7978 ) | ( n7897 & n7978 ) ;
  assign n7988 = ( n7870 & ~n7898 ) | ( n7870 & n7978 ) | ( ~n7898 & n7978 ) ;
  assign n7989 = ~n7987 & n7988 ;
  assign n7990 = n7983 | n7989 ;
  assign n7991 = n7758 &  n7899 ;
  assign n7984 = x77 | n7758 ;
  assign n7985 = x77 &  n7758 ;
  assign n7986 = ( n7984 & ~n7985 ) | ( n7984 & 1'b0 ) | ( ~n7985 & 1'b0 ) ;
  assign n7995 = ( n7869 & n7897 ) | ( n7869 & n7986 ) | ( n7897 & n7986 ) ;
  assign n7996 = ( n7869 & ~n7898 ) | ( n7869 & n7986 ) | ( ~n7898 & n7986 ) ;
  assign n7997 = ~n7995 & n7996 ;
  assign n7998 = n7991 | n7997 ;
  assign n7999 = n7766 &  n7899 ;
  assign n7992 = x76 | n7766 ;
  assign n7993 = x76 &  n7766 ;
  assign n7994 = ( n7992 & ~n7993 ) | ( n7992 & 1'b0 ) | ( ~n7993 & 1'b0 ) ;
  assign n8003 = ( n7868 & n7897 ) | ( n7868 & n7994 ) | ( n7897 & n7994 ) ;
  assign n8004 = ( n7868 & ~n7898 ) | ( n7868 & n7994 ) | ( ~n7898 & n7994 ) ;
  assign n8005 = ~n8003 & n8004 ;
  assign n8006 = n7999 | n8005 ;
  assign n8007 = n7774 &  n7899 ;
  assign n8000 = x75 | n7774 ;
  assign n8001 = x75 &  n7774 ;
  assign n8002 = ( n8000 & ~n8001 ) | ( n8000 & 1'b0 ) | ( ~n8001 & 1'b0 ) ;
  assign n8011 = ( n7867 & n7897 ) | ( n7867 & n8002 ) | ( n7897 & n8002 ) ;
  assign n8012 = ( n7867 & ~n7898 ) | ( n7867 & n8002 ) | ( ~n7898 & n8002 ) ;
  assign n8013 = ~n8011 & n8012 ;
  assign n8014 = n8007 | n8013 ;
  assign n8015 = n7782 &  n7899 ;
  assign n8008 = x74 | n7782 ;
  assign n8009 = x74 &  n7782 ;
  assign n8010 = ( n8008 & ~n8009 ) | ( n8008 & 1'b0 ) | ( ~n8009 & 1'b0 ) ;
  assign n8019 = ( n7866 & n7897 ) | ( n7866 & n8010 ) | ( n7897 & n8010 ) ;
  assign n8020 = ( n7866 & ~n7898 ) | ( n7866 & n8010 ) | ( ~n7898 & n8010 ) ;
  assign n8021 = ~n8019 & n8020 ;
  assign n8022 = n8015 | n8021 ;
  assign n8023 = n7790 &  n7899 ;
  assign n8016 = x73 | n7790 ;
  assign n8017 = x73 &  n7790 ;
  assign n8018 = ( n8016 & ~n8017 ) | ( n8016 & 1'b0 ) | ( ~n8017 & 1'b0 ) ;
  assign n8027 = ( n7865 & n7897 ) | ( n7865 & n8018 ) | ( n7897 & n8018 ) ;
  assign n8028 = ( n7865 & ~n7898 ) | ( n7865 & n8018 ) | ( ~n7898 & n8018 ) ;
  assign n8029 = ~n8027 & n8028 ;
  assign n8030 = n8023 | n8029 ;
  assign n8031 = n7798 &  n7899 ;
  assign n8024 = x72 | n7798 ;
  assign n8025 = x72 &  n7798 ;
  assign n8026 = ( n8024 & ~n8025 ) | ( n8024 & 1'b0 ) | ( ~n8025 & 1'b0 ) ;
  assign n8035 = ( n7864 & n7897 ) | ( n7864 & n8026 ) | ( n7897 & n8026 ) ;
  assign n8036 = ( n7864 & ~n7898 ) | ( n7864 & n8026 ) | ( ~n7898 & n8026 ) ;
  assign n8037 = ~n8035 & n8036 ;
  assign n8038 = n8031 | n8037 ;
  assign n8039 = n7806 &  n7899 ;
  assign n8032 = x71 | n7806 ;
  assign n8033 = x71 &  n7806 ;
  assign n8034 = ( n8032 & ~n8033 ) | ( n8032 & 1'b0 ) | ( ~n8033 & 1'b0 ) ;
  assign n8043 = ( n7863 & n7897 ) | ( n7863 & n8034 ) | ( n7897 & n8034 ) ;
  assign n8044 = ( n7863 & ~n7898 ) | ( n7863 & n8034 ) | ( ~n7898 & n8034 ) ;
  assign n8045 = ~n8043 & n8044 ;
  assign n8046 = n8039 | n8045 ;
  assign n8047 = n7814 &  n7899 ;
  assign n8040 = x70 | n7814 ;
  assign n8041 = x70 &  n7814 ;
  assign n8042 = ( n8040 & ~n8041 ) | ( n8040 & 1'b0 ) | ( ~n8041 & 1'b0 ) ;
  assign n8051 = ( n7862 & n7897 ) | ( n7862 & n8042 ) | ( n7897 & n8042 ) ;
  assign n8052 = ( n7862 & ~n7898 ) | ( n7862 & n8042 ) | ( ~n7898 & n8042 ) ;
  assign n8053 = ~n8051 & n8052 ;
  assign n8054 = n8047 | n8053 ;
  assign n8055 = n7822 &  n7899 ;
  assign n8048 = x69 | n7822 ;
  assign n8049 = x69 &  n7822 ;
  assign n8050 = ( n8048 & ~n8049 ) | ( n8048 & 1'b0 ) | ( ~n8049 & 1'b0 ) ;
  assign n8059 = ( n7861 & n7897 ) | ( n7861 & n8050 ) | ( n7897 & n8050 ) ;
  assign n8060 = ( n7861 & ~n7898 ) | ( n7861 & n8050 ) | ( ~n7898 & n8050 ) ;
  assign n8061 = ~n8059 & n8060 ;
  assign n8062 = n8055 | n8061 ;
  assign n8063 = n7830 &  n7899 ;
  assign n8056 = x68 | n7830 ;
  assign n8057 = x68 &  n7830 ;
  assign n8058 = ( n8056 & ~n8057 ) | ( n8056 & 1'b0 ) | ( ~n8057 & 1'b0 ) ;
  assign n8067 = ( n7860 & n7897 ) | ( n7860 & n8058 ) | ( n7897 & n8058 ) ;
  assign n8068 = ( n7860 & ~n7898 ) | ( n7860 & n8058 ) | ( ~n7898 & n8058 ) ;
  assign n8069 = ~n8067 & n8068 ;
  assign n8070 = n8063 | n8069 ;
  assign n8071 = n7839 &  n7899 ;
  assign n8064 = x67 | n7839 ;
  assign n8065 = x67 &  n7839 ;
  assign n8066 = ( n8064 & ~n8065 ) | ( n8064 & 1'b0 ) | ( ~n8065 & 1'b0 ) ;
  assign n8075 = ( n7859 & n7897 ) | ( n7859 & n8066 ) | ( n7897 & n8066 ) ;
  assign n8076 = ( n7859 & ~n7898 ) | ( n7859 & n8066 ) | ( ~n7898 & n8066 ) ;
  assign n8077 = ~n8075 & n8076 ;
  assign n8078 = n8071 | n8077 ;
  assign n8079 = n7845 &  n7899 ;
  assign n8072 = x66 | n7845 ;
  assign n8073 = x66 &  n7845 ;
  assign n8074 = ( n8072 & ~n8073 ) | ( n8072 & 1'b0 ) | ( ~n8073 & 1'b0 ) ;
  assign n8084 = ( n7858 & ~n7897 ) | ( n7858 & n8074 ) | ( ~n7897 & n8074 ) ;
  assign n8085 = ( n7858 & n7898 ) | ( n7858 & n8074 ) | ( n7898 & n8074 ) ;
  assign n8086 = ( n8084 & ~n8085 ) | ( n8084 & 1'b0 ) | ( ~n8085 & 1'b0 ) ;
  assign n8087 = n8079 | n8086 ;
  assign n8088 = n7856 &  n7899 ;
  assign n8080 = x65 &  n7856 ;
  assign n8081 = x65 | n7855 ;
  assign n8082 = n7851 | n8081 ;
  assign n8083 = ( n7857 & ~n8080 ) | ( n7857 & n8082 ) | ( ~n8080 & n8082 ) ;
  assign n8089 = ( x65 & n7856 ) | ( x65 & n7857 ) | ( n7856 & n7857 ) ;
  assign n8090 = ( n7898 & ~n8080 ) | ( n7898 & n8089 ) | ( ~n8080 & n8089 ) ;
  assign n8091 = ( n7897 & n8083 ) | ( n7897 & n8090 ) | ( n8083 & n8090 ) ;
  assign n8092 = ( n8083 & ~n8091 ) | ( n8083 & 1'b0 ) | ( ~n8091 & 1'b0 ) ;
  assign n8093 = n8088 | n8092 ;
  assign n8094 = ( x64 & ~x105 ) | ( x64 & 1'b0 ) | ( ~x105 & 1'b0 ) ;
  assign n8095 = ( n162 & ~n173 ) | ( n162 & n8094 ) | ( ~n173 & n8094 ) ;
  assign n8096 = ~n162 & n8095 ;
  assign n8097 = ~n270 & n8096 ;
  assign n8098 = n7897 &  n8097 ;
  assign n8099 = ( x23 & ~n8097 ) | ( x23 & n8098 ) | ( ~n8097 & n8098 ) ;
  assign n8100 = ~n253 & n7857 ;
  assign n8101 = ( n425 & ~n427 ) | ( n425 & n8100 ) | ( ~n427 & n8100 ) ;
  assign n8102 = ~n425 & n8101 ;
  assign n8103 = ~n7897 & n8102 ;
  assign n8104 = n8099 | n8103 ;
  assign n8105 = ~x22 & x64 ;
  assign n8106 = ( x65 & ~n8104 ) | ( x65 & n8105 ) | ( ~n8104 & n8105 ) ;
  assign n8107 = ( x66 & ~n8093 ) | ( x66 & n8106 ) | ( ~n8093 & n8106 ) ;
  assign n8108 = ( x67 & ~n8087 ) | ( x67 & n8107 ) | ( ~n8087 & n8107 ) ;
  assign n8109 = ( x68 & ~n8078 ) | ( x68 & n8108 ) | ( ~n8078 & n8108 ) ;
  assign n8110 = ( x69 & ~n8070 ) | ( x69 & n8109 ) | ( ~n8070 & n8109 ) ;
  assign n8111 = ( x70 & ~n8062 ) | ( x70 & n8110 ) | ( ~n8062 & n8110 ) ;
  assign n8112 = ( x71 & ~n8054 ) | ( x71 & n8111 ) | ( ~n8054 & n8111 ) ;
  assign n8113 = ( x72 & ~n8046 ) | ( x72 & n8112 ) | ( ~n8046 & n8112 ) ;
  assign n8114 = ( x73 & ~n8038 ) | ( x73 & n8113 ) | ( ~n8038 & n8113 ) ;
  assign n8115 = ( x74 & ~n8030 ) | ( x74 & n8114 ) | ( ~n8030 & n8114 ) ;
  assign n8116 = ( x75 & ~n8022 ) | ( x75 & n8115 ) | ( ~n8022 & n8115 ) ;
  assign n8117 = ( x76 & ~n8014 ) | ( x76 & n8116 ) | ( ~n8014 & n8116 ) ;
  assign n8118 = ( x77 & ~n8006 ) | ( x77 & n8117 ) | ( ~n8006 & n8117 ) ;
  assign n8119 = ( x78 & ~n7998 ) | ( x78 & n8118 ) | ( ~n7998 & n8118 ) ;
  assign n8120 = ( x79 & ~n7990 ) | ( x79 & n8119 ) | ( ~n7990 & n8119 ) ;
  assign n8121 = ( x80 & ~n7982 ) | ( x80 & n8120 ) | ( ~n7982 & n8120 ) ;
  assign n8122 = ( x81 & ~n7974 ) | ( x81 & n8121 ) | ( ~n7974 & n8121 ) ;
  assign n8123 = ( x82 & ~n7966 ) | ( x82 & n8122 ) | ( ~n7966 & n8122 ) ;
  assign n8124 = ( x83 & ~n7958 ) | ( x83 & n8123 ) | ( ~n7958 & n8123 ) ;
  assign n8125 = ( x84 & ~n7950 ) | ( x84 & n8124 ) | ( ~n7950 & n8124 ) ;
  assign n8126 = ( x85 & ~n7942 ) | ( x85 & n8125 ) | ( ~n7942 & n8125 ) ;
  assign n8127 = ( x86 & ~n7934 ) | ( x86 & n8126 ) | ( ~n7934 & n8126 ) ;
  assign n8128 = ( x87 & ~n7926 ) | ( x87 & n8127 ) | ( ~n7926 & n8127 ) ;
  assign n8129 = ( x88 & ~n7918 ) | ( x88 & n8128 ) | ( ~n7918 & n8128 ) ;
  assign n8133 = ( x89 & ~n7910 ) | ( x89 & n8129 ) | ( ~n7910 & n8129 ) ;
  assign n8257 = ( x90 & ~n8141 ) | ( x90 & n8133 ) | ( ~n8141 & n8133 ) ;
  assign n8258 = ( x91 & ~n8256 ) | ( x91 & n8257 ) | ( ~n8256 & n8257 ) ;
  assign n8259 = ( x92 & ~n8251 ) | ( x92 & n8258 ) | ( ~n8251 & n8258 ) ;
  assign n8260 = ( x93 & ~n8243 ) | ( x93 & n8259 ) | ( ~n8243 & n8259 ) ;
  assign n8261 = ( x94 & ~n8235 ) | ( x94 & n8260 ) | ( ~n8235 & n8260 ) ;
  assign n8262 = ( x95 & ~n8227 ) | ( x95 & n8261 ) | ( ~n8227 & n8261 ) ;
  assign n8263 = ( x96 & ~n8219 ) | ( x96 & n8262 ) | ( ~n8219 & n8262 ) ;
  assign n8264 = ( x97 & ~n8211 ) | ( x97 & n8263 ) | ( ~n8211 & n8263 ) ;
  assign n8265 = ( x98 & ~n8203 ) | ( x98 & n8264 ) | ( ~n8203 & n8264 ) ;
  assign n8266 = ( x99 & ~n8195 ) | ( x99 & n8265 ) | ( ~n8195 & n8265 ) ;
  assign n8267 = ( x100 & ~n8187 ) | ( x100 & n8266 ) | ( ~n8187 & n8266 ) ;
  assign n8268 = ( x101 & ~n8179 ) | ( x101 & n8267 ) | ( ~n8179 & n8267 ) ;
  assign n8269 = ( x102 & ~n8171 ) | ( x102 & n8268 ) | ( ~n8171 & n8268 ) ;
  assign n8270 = ( x103 & ~n8163 ) | ( x103 & n8269 ) | ( ~n8163 & n8269 ) ;
  assign n8271 = ( x104 & ~n8155 ) | ( x104 & n8270 ) | ( ~n8155 & n8270 ) ;
  assign n8275 = n162 | n173 ;
  assign n8276 = n270 | n8275 ;
  assign n8272 = x104 | n7896 ;
  assign n8273 = ( x104 & n7896 ) | ( x104 & n7898 ) | ( n7896 & n7898 ) ;
  assign n8274 = ( n7553 & ~n8272 ) | ( n7553 & n8273 ) | ( ~n8272 & n8273 ) ;
  assign n8278 = x105 &  n8274 ;
  assign n8277 = x105 | n8274 ;
  assign n8279 = ( n8276 & ~n8278 ) | ( n8276 & n8277 ) | ( ~n8278 & n8277 ) ;
  assign n8280 = n8271 | n8279 ;
  assign n8281 = ~n8274 |  n7898 ;
  assign n8301 = n8155 &  n8281 ;
  assign n8302 = n8280 &  n8301 ;
  assign n8288 = x104 | n8155 ;
  assign n8289 = x104 &  n8155 ;
  assign n8290 = ( n8288 & ~n8289 ) | ( n8288 & 1'b0 ) | ( ~n8289 & 1'b0 ) ;
  assign n8303 = n8270 &  n8290 ;
  assign n8282 = n8280 &  n8281 ;
  assign n8304 = ( n8270 & ~n8282 ) | ( n8270 & n8290 ) | ( ~n8282 & n8290 ) ;
  assign n8305 = ( n8302 & ~n8303 ) | ( n8302 & n8304 ) | ( ~n8303 & n8304 ) ;
  assign n8292 = ( x105 & n8271 ) | ( x105 & n8274 ) | ( n8271 & n8274 ) ;
  assign n8291 = ( x105 & ~n8271 ) | ( x105 & n8274 ) | ( ~n8271 & n8274 ) ;
  assign n8293 = ( n8271 & ~n8292 ) | ( n8271 & n8291 ) | ( ~n8292 & n8291 ) ;
  assign n8294 = ~n8282 & n8293 ;
  assign n8295 = n7553 &  n7898 ;
  assign n8296 = n8280 &  n8295 ;
  assign n8297 = n8294 | n8296 ;
  assign n8309 = n8163 &  n8281 ;
  assign n8310 = n8280 &  n8309 ;
  assign n8298 = x103 | n8163 ;
  assign n8299 = x103 &  n8163 ;
  assign n8300 = ( n8298 & ~n8299 ) | ( n8298 & 1'b0 ) | ( ~n8299 & 1'b0 ) ;
  assign n8311 = n8269 &  n8300 ;
  assign n8312 = ( n8269 & ~n8282 ) | ( n8269 & n8300 ) | ( ~n8282 & n8300 ) ;
  assign n8313 = ( n8310 & ~n8311 ) | ( n8310 & n8312 ) | ( ~n8311 & n8312 ) ;
  assign n8317 = n8171 &  n8281 ;
  assign n8318 = n8280 &  n8317 ;
  assign n8306 = x102 | n8171 ;
  assign n8307 = x102 &  n8171 ;
  assign n8308 = ( n8306 & ~n8307 ) | ( n8306 & 1'b0 ) | ( ~n8307 & 1'b0 ) ;
  assign n8319 = n8268 &  n8308 ;
  assign n8320 = ( n8268 & ~n8282 ) | ( n8268 & n8308 ) | ( ~n8282 & n8308 ) ;
  assign n8321 = ( n8318 & ~n8319 ) | ( n8318 & n8320 ) | ( ~n8319 & n8320 ) ;
  assign n8325 = n8179 &  n8281 ;
  assign n8326 = n8280 &  n8325 ;
  assign n8314 = x101 | n8179 ;
  assign n8315 = x101 &  n8179 ;
  assign n8316 = ( n8314 & ~n8315 ) | ( n8314 & 1'b0 ) | ( ~n8315 & 1'b0 ) ;
  assign n8327 = n8267 &  n8316 ;
  assign n8328 = ( n8267 & ~n8282 ) | ( n8267 & n8316 ) | ( ~n8282 & n8316 ) ;
  assign n8329 = ( n8326 & ~n8327 ) | ( n8326 & n8328 ) | ( ~n8327 & n8328 ) ;
  assign n8333 = n8187 &  n8281 ;
  assign n8334 = n8280 &  n8333 ;
  assign n8322 = x100 | n8187 ;
  assign n8323 = x100 &  n8187 ;
  assign n8324 = ( n8322 & ~n8323 ) | ( n8322 & 1'b0 ) | ( ~n8323 & 1'b0 ) ;
  assign n8335 = n8266 &  n8324 ;
  assign n8336 = ( n8266 & ~n8282 ) | ( n8266 & n8324 ) | ( ~n8282 & n8324 ) ;
  assign n8337 = ( n8334 & ~n8335 ) | ( n8334 & n8336 ) | ( ~n8335 & n8336 ) ;
  assign n8341 = n8195 &  n8281 ;
  assign n8342 = n8280 &  n8341 ;
  assign n8330 = x99 | n8195 ;
  assign n8331 = x99 &  n8195 ;
  assign n8332 = ( n8330 & ~n8331 ) | ( n8330 & 1'b0 ) | ( ~n8331 & 1'b0 ) ;
  assign n8344 = ( n8265 & n8282 ) | ( n8265 & n8332 ) | ( n8282 & n8332 ) ;
  assign n8343 = n8265 | n8332 ;
  assign n8345 = ( n8342 & ~n8344 ) | ( n8342 & n8343 ) | ( ~n8344 & n8343 ) ;
  assign n8349 = n8203 &  n8281 ;
  assign n8350 = n8280 &  n8349 ;
  assign n8338 = x98 | n8203 ;
  assign n8339 = x98 &  n8203 ;
  assign n8340 = ( n8338 & ~n8339 ) | ( n8338 & 1'b0 ) | ( ~n8339 & 1'b0 ) ;
  assign n8352 = ( n8264 & n8282 ) | ( n8264 & n8340 ) | ( n8282 & n8340 ) ;
  assign n8351 = n8264 | n8340 ;
  assign n8353 = ( n8350 & ~n8352 ) | ( n8350 & n8351 ) | ( ~n8352 & n8351 ) ;
  assign n8357 = n8211 &  n8281 ;
  assign n8358 = n8280 &  n8357 ;
  assign n8346 = x97 | n8211 ;
  assign n8347 = x97 &  n8211 ;
  assign n8348 = ( n8346 & ~n8347 ) | ( n8346 & 1'b0 ) | ( ~n8347 & 1'b0 ) ;
  assign n8360 = ( n8263 & n8282 ) | ( n8263 & n8348 ) | ( n8282 & n8348 ) ;
  assign n8359 = n8263 | n8348 ;
  assign n8361 = ( n8358 & ~n8360 ) | ( n8358 & n8359 ) | ( ~n8360 & n8359 ) ;
  assign n8365 = n8219 &  n8281 ;
  assign n8366 = n8280 &  n8365 ;
  assign n8354 = x96 | n8219 ;
  assign n8355 = x96 &  n8219 ;
  assign n8356 = ( n8354 & ~n8355 ) | ( n8354 & 1'b0 ) | ( ~n8355 & 1'b0 ) ;
  assign n8368 = ( n8262 & n8282 ) | ( n8262 & n8356 ) | ( n8282 & n8356 ) ;
  assign n8367 = n8262 | n8356 ;
  assign n8369 = ( n8366 & ~n8368 ) | ( n8366 & n8367 ) | ( ~n8368 & n8367 ) ;
  assign n8373 = n8227 &  n8281 ;
  assign n8374 = n8280 &  n8373 ;
  assign n8362 = x95 | n8227 ;
  assign n8363 = x95 &  n8227 ;
  assign n8364 = ( n8362 & ~n8363 ) | ( n8362 & 1'b0 ) | ( ~n8363 & 1'b0 ) ;
  assign n8376 = ( n8261 & n8282 ) | ( n8261 & n8364 ) | ( n8282 & n8364 ) ;
  assign n8375 = n8261 | n8364 ;
  assign n8377 = ( n8374 & ~n8376 ) | ( n8374 & n8375 ) | ( ~n8376 & n8375 ) ;
  assign n8381 = n8235 &  n8281 ;
  assign n8382 = n8280 &  n8381 ;
  assign n8370 = x94 | n8235 ;
  assign n8371 = x94 &  n8235 ;
  assign n8372 = ( n8370 & ~n8371 ) | ( n8370 & 1'b0 ) | ( ~n8371 & 1'b0 ) ;
  assign n8384 = ( n8260 & n8282 ) | ( n8260 & n8372 ) | ( n8282 & n8372 ) ;
  assign n8383 = n8260 | n8372 ;
  assign n8385 = ( n8382 & ~n8384 ) | ( n8382 & n8383 ) | ( ~n8384 & n8383 ) ;
  assign n8389 = n8243 &  n8281 ;
  assign n8390 = n8280 &  n8389 ;
  assign n8378 = x93 | n8243 ;
  assign n8379 = x93 &  n8243 ;
  assign n8380 = ( n8378 & ~n8379 ) | ( n8378 & 1'b0 ) | ( ~n8379 & 1'b0 ) ;
  assign n8392 = ( n8259 & n8282 ) | ( n8259 & n8380 ) | ( n8282 & n8380 ) ;
  assign n8391 = n8259 | n8380 ;
  assign n8393 = ( n8390 & ~n8392 ) | ( n8390 & n8391 ) | ( ~n8392 & n8391 ) ;
  assign n8397 = n8251 &  n8281 ;
  assign n8398 = n8280 &  n8397 ;
  assign n8386 = x92 | n8251 ;
  assign n8387 = x92 &  n8251 ;
  assign n8388 = ( n8386 & ~n8387 ) | ( n8386 & 1'b0 ) | ( ~n8387 & 1'b0 ) ;
  assign n8400 = ( n8258 & n8282 ) | ( n8258 & n8388 ) | ( n8282 & n8388 ) ;
  assign n8399 = n8258 | n8388 ;
  assign n8401 = ( n8398 & ~n8400 ) | ( n8398 & n8399 ) | ( ~n8400 & n8399 ) ;
  assign n8402 = n8256 &  n8281 ;
  assign n8403 = n8280 &  n8402 ;
  assign n8394 = x91 | n8256 ;
  assign n8395 = x91 &  n8256 ;
  assign n8396 = ( n8394 & ~n8395 ) | ( n8394 & 1'b0 ) | ( ~n8395 & 1'b0 ) ;
  assign n8405 = ( n8257 & n8282 ) | ( n8257 & n8396 ) | ( n8282 & n8396 ) ;
  assign n8404 = n8257 | n8396 ;
  assign n8406 = ( n8403 & ~n8405 ) | ( n8403 & n8404 ) | ( ~n8405 & n8404 ) ;
  assign n8283 = n8141 &  n8281 ;
  assign n8284 = n8280 &  n8283 ;
  assign n8142 = x90 | n8141 ;
  assign n8143 = x90 &  n8141 ;
  assign n8144 = ( n8142 & ~n8143 ) | ( n8142 & 1'b0 ) | ( ~n8143 & 1'b0 ) ;
  assign n8286 = ( n8133 & n8144 ) | ( n8133 & n8282 ) | ( n8144 & n8282 ) ;
  assign n8285 = n8133 | n8144 ;
  assign n8287 = ( n8284 & ~n8286 ) | ( n8284 & n8285 ) | ( ~n8286 & n8285 ) ;
  assign n8410 = n7910 &  n8281 ;
  assign n8411 = n8280 &  n8410 ;
  assign n8130 = x89 | n7910 ;
  assign n8131 = x89 &  n7910 ;
  assign n8132 = ( n8130 & ~n8131 ) | ( n8130 & 1'b0 ) | ( ~n8131 & 1'b0 ) ;
  assign n8412 = n8129 &  n8132 ;
  assign n8413 = ( n8129 & ~n8282 ) | ( n8129 & n8132 ) | ( ~n8282 & n8132 ) ;
  assign n8414 = ( n8411 & ~n8412 ) | ( n8411 & n8413 ) | ( ~n8412 & n8413 ) ;
  assign n8418 = n7918 &  n8281 ;
  assign n8419 = n8280 &  n8418 ;
  assign n8407 = x88 | n7918 ;
  assign n8408 = x88 &  n7918 ;
  assign n8409 = ( n8407 & ~n8408 ) | ( n8407 & 1'b0 ) | ( ~n8408 & 1'b0 ) ;
  assign n8421 = ( n8128 & n8282 ) | ( n8128 & n8409 ) | ( n8282 & n8409 ) ;
  assign n8420 = n8128 | n8409 ;
  assign n8422 = ( n8419 & ~n8421 ) | ( n8419 & n8420 ) | ( ~n8421 & n8420 ) ;
  assign n8426 = n7926 &  n8281 ;
  assign n8427 = n8280 &  n8426 ;
  assign n8415 = x87 | n7926 ;
  assign n8416 = x87 &  n7926 ;
  assign n8417 = ( n8415 & ~n8416 ) | ( n8415 & 1'b0 ) | ( ~n8416 & 1'b0 ) ;
  assign n8429 = ( n8127 & n8282 ) | ( n8127 & n8417 ) | ( n8282 & n8417 ) ;
  assign n8428 = n8127 | n8417 ;
  assign n8430 = ( n8427 & ~n8429 ) | ( n8427 & n8428 ) | ( ~n8429 & n8428 ) ;
  assign n8434 = n7934 &  n8281 ;
  assign n8435 = n8280 &  n8434 ;
  assign n8423 = x86 | n7934 ;
  assign n8424 = x86 &  n7934 ;
  assign n8425 = ( n8423 & ~n8424 ) | ( n8423 & 1'b0 ) | ( ~n8424 & 1'b0 ) ;
  assign n8437 = ( n8126 & n8282 ) | ( n8126 & n8425 ) | ( n8282 & n8425 ) ;
  assign n8436 = n8126 | n8425 ;
  assign n8438 = ( n8435 & ~n8437 ) | ( n8435 & n8436 ) | ( ~n8437 & n8436 ) ;
  assign n8442 = n7942 &  n8281 ;
  assign n8443 = n8280 &  n8442 ;
  assign n8431 = x85 | n7942 ;
  assign n8432 = x85 &  n7942 ;
  assign n8433 = ( n8431 & ~n8432 ) | ( n8431 & 1'b0 ) | ( ~n8432 & 1'b0 ) ;
  assign n8445 = ( n8125 & n8282 ) | ( n8125 & n8433 ) | ( n8282 & n8433 ) ;
  assign n8444 = n8125 | n8433 ;
  assign n8446 = ( n8443 & ~n8445 ) | ( n8443 & n8444 ) | ( ~n8445 & n8444 ) ;
  assign n8450 = n7950 &  n8281 ;
  assign n8451 = n8280 &  n8450 ;
  assign n8439 = x84 | n7950 ;
  assign n8440 = x84 &  n7950 ;
  assign n8441 = ( n8439 & ~n8440 ) | ( n8439 & 1'b0 ) | ( ~n8440 & 1'b0 ) ;
  assign n8453 = ( n8124 & n8282 ) | ( n8124 & n8441 ) | ( n8282 & n8441 ) ;
  assign n8452 = n8124 | n8441 ;
  assign n8454 = ( n8451 & ~n8453 ) | ( n8451 & n8452 ) | ( ~n8453 & n8452 ) ;
  assign n8458 = n7958 &  n8281 ;
  assign n8459 = n8280 &  n8458 ;
  assign n8447 = x83 | n7958 ;
  assign n8448 = x83 &  n7958 ;
  assign n8449 = ( n8447 & ~n8448 ) | ( n8447 & 1'b0 ) | ( ~n8448 & 1'b0 ) ;
  assign n8461 = ( n8123 & n8282 ) | ( n8123 & n8449 ) | ( n8282 & n8449 ) ;
  assign n8460 = n8123 | n8449 ;
  assign n8462 = ( n8459 & ~n8461 ) | ( n8459 & n8460 ) | ( ~n8461 & n8460 ) ;
  assign n8466 = n7966 &  n8281 ;
  assign n8467 = n8280 &  n8466 ;
  assign n8455 = x82 | n7966 ;
  assign n8456 = x82 &  n7966 ;
  assign n8457 = ( n8455 & ~n8456 ) | ( n8455 & 1'b0 ) | ( ~n8456 & 1'b0 ) ;
  assign n8469 = ( n8122 & n8282 ) | ( n8122 & n8457 ) | ( n8282 & n8457 ) ;
  assign n8468 = n8122 | n8457 ;
  assign n8470 = ( n8467 & ~n8469 ) | ( n8467 & n8468 ) | ( ~n8469 & n8468 ) ;
  assign n8474 = n7974 &  n8281 ;
  assign n8475 = n8280 &  n8474 ;
  assign n8463 = x81 | n7974 ;
  assign n8464 = x81 &  n7974 ;
  assign n8465 = ( n8463 & ~n8464 ) | ( n8463 & 1'b0 ) | ( ~n8464 & 1'b0 ) ;
  assign n8477 = ( n8121 & n8282 ) | ( n8121 & n8465 ) | ( n8282 & n8465 ) ;
  assign n8476 = n8121 | n8465 ;
  assign n8478 = ( n8475 & ~n8477 ) | ( n8475 & n8476 ) | ( ~n8477 & n8476 ) ;
  assign n8482 = n7982 &  n8281 ;
  assign n8483 = n8280 &  n8482 ;
  assign n8471 = x80 | n7982 ;
  assign n8472 = x80 &  n7982 ;
  assign n8473 = ( n8471 & ~n8472 ) | ( n8471 & 1'b0 ) | ( ~n8472 & 1'b0 ) ;
  assign n8485 = ( n8120 & n8282 ) | ( n8120 & n8473 ) | ( n8282 & n8473 ) ;
  assign n8484 = n8120 | n8473 ;
  assign n8486 = ( n8483 & ~n8485 ) | ( n8483 & n8484 ) | ( ~n8485 & n8484 ) ;
  assign n8490 = n7990 &  n8281 ;
  assign n8491 = n8280 &  n8490 ;
  assign n8479 = x79 | n7990 ;
  assign n8480 = x79 &  n7990 ;
  assign n8481 = ( n8479 & ~n8480 ) | ( n8479 & 1'b0 ) | ( ~n8480 & 1'b0 ) ;
  assign n8493 = ( n8119 & n8282 ) | ( n8119 & n8481 ) | ( n8282 & n8481 ) ;
  assign n8492 = n8119 | n8481 ;
  assign n8494 = ( n8491 & ~n8493 ) | ( n8491 & n8492 ) | ( ~n8493 & n8492 ) ;
  assign n8498 = n7998 &  n8281 ;
  assign n8499 = n8280 &  n8498 ;
  assign n8487 = x78 | n7998 ;
  assign n8488 = x78 &  n7998 ;
  assign n8489 = ( n8487 & ~n8488 ) | ( n8487 & 1'b0 ) | ( ~n8488 & 1'b0 ) ;
  assign n8501 = ( n8118 & n8282 ) | ( n8118 & n8489 ) | ( n8282 & n8489 ) ;
  assign n8500 = n8118 | n8489 ;
  assign n8502 = ( n8499 & ~n8501 ) | ( n8499 & n8500 ) | ( ~n8501 & n8500 ) ;
  assign n8506 = n8006 &  n8281 ;
  assign n8507 = n8280 &  n8506 ;
  assign n8495 = x77 | n8006 ;
  assign n8496 = x77 &  n8006 ;
  assign n8497 = ( n8495 & ~n8496 ) | ( n8495 & 1'b0 ) | ( ~n8496 & 1'b0 ) ;
  assign n8509 = ( n8117 & n8282 ) | ( n8117 & n8497 ) | ( n8282 & n8497 ) ;
  assign n8508 = n8117 | n8497 ;
  assign n8510 = ( n8507 & ~n8509 ) | ( n8507 & n8508 ) | ( ~n8509 & n8508 ) ;
  assign n8514 = n8014 &  n8281 ;
  assign n8515 = n8280 &  n8514 ;
  assign n8503 = x76 | n8014 ;
  assign n8504 = x76 &  n8014 ;
  assign n8505 = ( n8503 & ~n8504 ) | ( n8503 & 1'b0 ) | ( ~n8504 & 1'b0 ) ;
  assign n8517 = ( n8116 & n8282 ) | ( n8116 & n8505 ) | ( n8282 & n8505 ) ;
  assign n8516 = n8116 | n8505 ;
  assign n8518 = ( n8515 & ~n8517 ) | ( n8515 & n8516 ) | ( ~n8517 & n8516 ) ;
  assign n8522 = n8022 &  n8281 ;
  assign n8523 = n8280 &  n8522 ;
  assign n8511 = x75 | n8022 ;
  assign n8512 = x75 &  n8022 ;
  assign n8513 = ( n8511 & ~n8512 ) | ( n8511 & 1'b0 ) | ( ~n8512 & 1'b0 ) ;
  assign n8525 = ( n8115 & n8282 ) | ( n8115 & n8513 ) | ( n8282 & n8513 ) ;
  assign n8524 = n8115 | n8513 ;
  assign n8526 = ( n8523 & ~n8525 ) | ( n8523 & n8524 ) | ( ~n8525 & n8524 ) ;
  assign n8530 = n8030 &  n8281 ;
  assign n8531 = n8280 &  n8530 ;
  assign n8519 = x74 | n8030 ;
  assign n8520 = x74 &  n8030 ;
  assign n8521 = ( n8519 & ~n8520 ) | ( n8519 & 1'b0 ) | ( ~n8520 & 1'b0 ) ;
  assign n8533 = ( n8114 & n8282 ) | ( n8114 & n8521 ) | ( n8282 & n8521 ) ;
  assign n8532 = n8114 | n8521 ;
  assign n8534 = ( n8531 & ~n8533 ) | ( n8531 & n8532 ) | ( ~n8533 & n8532 ) ;
  assign n8538 = n8038 &  n8281 ;
  assign n8539 = n8280 &  n8538 ;
  assign n8527 = x73 | n8038 ;
  assign n8528 = x73 &  n8038 ;
  assign n8529 = ( n8527 & ~n8528 ) | ( n8527 & 1'b0 ) | ( ~n8528 & 1'b0 ) ;
  assign n8541 = ( n8113 & n8282 ) | ( n8113 & n8529 ) | ( n8282 & n8529 ) ;
  assign n8540 = n8113 | n8529 ;
  assign n8542 = ( n8539 & ~n8541 ) | ( n8539 & n8540 ) | ( ~n8541 & n8540 ) ;
  assign n8546 = n8046 &  n8281 ;
  assign n8547 = n8280 &  n8546 ;
  assign n8535 = x72 | n8046 ;
  assign n8536 = x72 &  n8046 ;
  assign n8537 = ( n8535 & ~n8536 ) | ( n8535 & 1'b0 ) | ( ~n8536 & 1'b0 ) ;
  assign n8549 = ( n8112 & n8282 ) | ( n8112 & n8537 ) | ( n8282 & n8537 ) ;
  assign n8548 = n8112 | n8537 ;
  assign n8550 = ( n8547 & ~n8549 ) | ( n8547 & n8548 ) | ( ~n8549 & n8548 ) ;
  assign n8554 = n8054 &  n8281 ;
  assign n8555 = n8280 &  n8554 ;
  assign n8543 = x71 | n8054 ;
  assign n8544 = x71 &  n8054 ;
  assign n8545 = ( n8543 & ~n8544 ) | ( n8543 & 1'b0 ) | ( ~n8544 & 1'b0 ) ;
  assign n8557 = ( n8111 & n8282 ) | ( n8111 & n8545 ) | ( n8282 & n8545 ) ;
  assign n8556 = n8111 | n8545 ;
  assign n8558 = ( n8555 & ~n8557 ) | ( n8555 & n8556 ) | ( ~n8557 & n8556 ) ;
  assign n8562 = n8062 &  n8281 ;
  assign n8563 = n8280 &  n8562 ;
  assign n8551 = x70 | n8062 ;
  assign n8552 = x70 &  n8062 ;
  assign n8553 = ( n8551 & ~n8552 ) | ( n8551 & 1'b0 ) | ( ~n8552 & 1'b0 ) ;
  assign n8565 = ( n8110 & n8282 ) | ( n8110 & n8553 ) | ( n8282 & n8553 ) ;
  assign n8564 = n8110 | n8553 ;
  assign n8566 = ( n8563 & ~n8565 ) | ( n8563 & n8564 ) | ( ~n8565 & n8564 ) ;
  assign n8570 = n8070 &  n8281 ;
  assign n8571 = n8280 &  n8570 ;
  assign n8559 = x69 | n8070 ;
  assign n8560 = x69 &  n8070 ;
  assign n8561 = ( n8559 & ~n8560 ) | ( n8559 & 1'b0 ) | ( ~n8560 & 1'b0 ) ;
  assign n8573 = ( n8109 & n8282 ) | ( n8109 & n8561 ) | ( n8282 & n8561 ) ;
  assign n8572 = n8109 | n8561 ;
  assign n8574 = ( n8571 & ~n8573 ) | ( n8571 & n8572 ) | ( ~n8573 & n8572 ) ;
  assign n8578 = n8078 &  n8281 ;
  assign n8579 = n8280 &  n8578 ;
  assign n8567 = x68 | n8078 ;
  assign n8568 = x68 &  n8078 ;
  assign n8569 = ( n8567 & ~n8568 ) | ( n8567 & 1'b0 ) | ( ~n8568 & 1'b0 ) ;
  assign n8581 = ( n8108 & n8282 ) | ( n8108 & n8569 ) | ( n8282 & n8569 ) ;
  assign n8580 = n8108 | n8569 ;
  assign n8582 = ( n8579 & ~n8581 ) | ( n8579 & n8580 ) | ( ~n8581 & n8580 ) ;
  assign n8586 = n8087 &  n8281 ;
  assign n8587 = n8280 &  n8586 ;
  assign n8575 = x67 | n8087 ;
  assign n8576 = x67 &  n8087 ;
  assign n8577 = ( n8575 & ~n8576 ) | ( n8575 & 1'b0 ) | ( ~n8576 & 1'b0 ) ;
  assign n8589 = ( n8107 & n8282 ) | ( n8107 & n8577 ) | ( n8282 & n8577 ) ;
  assign n8588 = n8107 | n8577 ;
  assign n8590 = ( n8587 & ~n8589 ) | ( n8587 & n8588 ) | ( ~n8589 & n8588 ) ;
  assign n8591 = n8093 &  n8281 ;
  assign n8592 = n8280 &  n8591 ;
  assign n8583 = x66 | n8093 ;
  assign n8584 = x66 &  n8093 ;
  assign n8585 = ( n8583 & ~n8584 ) | ( n8583 & 1'b0 ) | ( ~n8584 & 1'b0 ) ;
  assign n8593 = n8106 &  n8585 ;
  assign n8594 = ( n8106 & ~n8282 ) | ( n8106 & n8585 ) | ( ~n8282 & n8585 ) ;
  assign n8595 = ( n8592 & ~n8593 ) | ( n8592 & n8594 ) | ( ~n8593 & n8594 ) ;
  assign n8596 = ( n8104 & ~x65 ) | ( n8104 & n8105 ) | ( ~x65 & n8105 ) ;
  assign n8597 = ( n8106 & ~n8105 ) | ( n8106 & n8596 ) | ( ~n8105 & n8596 ) ;
  assign n8598 = ~n8282 & n8597 ;
  assign n8599 = n8104 &  n8281 ;
  assign n8600 = n8280 &  n8599 ;
  assign n8601 = n8598 | n8600 ;
  assign n8602 = ( x64 & ~n8282 ) | ( x64 & 1'b0 ) | ( ~n8282 & 1'b0 ) ;
  assign n8603 = ( x22 & ~n8602 ) | ( x22 & 1'b0 ) | ( ~n8602 & 1'b0 ) ;
  assign n8604 = ( n8105 & ~n8282 ) | ( n8105 & 1'b0 ) | ( ~n8282 & 1'b0 ) ;
  assign n8605 = n8603 | n8604 ;
  assign n8606 = ~x21 & x64 ;
  assign n8607 = ( x65 & ~n8605 ) | ( x65 & n8606 ) | ( ~n8605 & n8606 ) ;
  assign n8608 = ( x66 & ~n8601 ) | ( x66 & n8607 ) | ( ~n8601 & n8607 ) ;
  assign n8609 = ( x67 & ~n8595 ) | ( x67 & n8608 ) | ( ~n8595 & n8608 ) ;
  assign n8610 = ( x68 & ~n8590 ) | ( x68 & n8609 ) | ( ~n8590 & n8609 ) ;
  assign n8611 = ( x69 & ~n8582 ) | ( x69 & n8610 ) | ( ~n8582 & n8610 ) ;
  assign n8612 = ( x70 & ~n8574 ) | ( x70 & n8611 ) | ( ~n8574 & n8611 ) ;
  assign n8613 = ( x71 & ~n8566 ) | ( x71 & n8612 ) | ( ~n8566 & n8612 ) ;
  assign n8614 = ( x72 & ~n8558 ) | ( x72 & n8613 ) | ( ~n8558 & n8613 ) ;
  assign n8615 = ( x73 & ~n8550 ) | ( x73 & n8614 ) | ( ~n8550 & n8614 ) ;
  assign n8616 = ( x74 & ~n8542 ) | ( x74 & n8615 ) | ( ~n8542 & n8615 ) ;
  assign n8617 = ( x75 & ~n8534 ) | ( x75 & n8616 ) | ( ~n8534 & n8616 ) ;
  assign n8618 = ( x76 & ~n8526 ) | ( x76 & n8617 ) | ( ~n8526 & n8617 ) ;
  assign n8619 = ( x77 & ~n8518 ) | ( x77 & n8618 ) | ( ~n8518 & n8618 ) ;
  assign n8620 = ( x78 & ~n8510 ) | ( x78 & n8619 ) | ( ~n8510 & n8619 ) ;
  assign n8621 = ( x79 & ~n8502 ) | ( x79 & n8620 ) | ( ~n8502 & n8620 ) ;
  assign n8622 = ( x80 & ~n8494 ) | ( x80 & n8621 ) | ( ~n8494 & n8621 ) ;
  assign n8623 = ( x81 & ~n8486 ) | ( x81 & n8622 ) | ( ~n8486 & n8622 ) ;
  assign n8624 = ( x82 & ~n8478 ) | ( x82 & n8623 ) | ( ~n8478 & n8623 ) ;
  assign n8625 = ( x83 & ~n8470 ) | ( x83 & n8624 ) | ( ~n8470 & n8624 ) ;
  assign n8626 = ( x84 & ~n8462 ) | ( x84 & n8625 ) | ( ~n8462 & n8625 ) ;
  assign n8627 = ( x85 & ~n8454 ) | ( x85 & n8626 ) | ( ~n8454 & n8626 ) ;
  assign n8628 = ( x86 & ~n8446 ) | ( x86 & n8627 ) | ( ~n8446 & n8627 ) ;
  assign n8629 = ( x87 & ~n8438 ) | ( x87 & n8628 ) | ( ~n8438 & n8628 ) ;
  assign n8630 = ( x88 & ~n8430 ) | ( x88 & n8629 ) | ( ~n8430 & n8629 ) ;
  assign n8631 = ( x89 & ~n8422 ) | ( x89 & n8630 ) | ( ~n8422 & n8630 ) ;
  assign n8632 = ( x90 & ~n8414 ) | ( x90 & n8631 ) | ( ~n8414 & n8631 ) ;
  assign n8633 = ( x91 & ~n8287 ) | ( x91 & n8632 ) | ( ~n8287 & n8632 ) ;
  assign n8634 = ( x92 & ~n8406 ) | ( x92 & n8633 ) | ( ~n8406 & n8633 ) ;
  assign n8635 = ( x93 & ~n8401 ) | ( x93 & n8634 ) | ( ~n8401 & n8634 ) ;
  assign n8636 = ( x94 & ~n8393 ) | ( x94 & n8635 ) | ( ~n8393 & n8635 ) ;
  assign n8637 = ( x95 & ~n8385 ) | ( x95 & n8636 ) | ( ~n8385 & n8636 ) ;
  assign n8638 = ( x96 & ~n8377 ) | ( x96 & n8637 ) | ( ~n8377 & n8637 ) ;
  assign n8639 = ( x97 & ~n8369 ) | ( x97 & n8638 ) | ( ~n8369 & n8638 ) ;
  assign n8640 = ( x98 & ~n8361 ) | ( x98 & n8639 ) | ( ~n8361 & n8639 ) ;
  assign n8641 = ( x99 & ~n8353 ) | ( x99 & n8640 ) | ( ~n8353 & n8640 ) ;
  assign n8642 = ( x100 & ~n8345 ) | ( x100 & n8641 ) | ( ~n8345 & n8641 ) ;
  assign n8643 = ( x101 & ~n8337 ) | ( x101 & n8642 ) | ( ~n8337 & n8642 ) ;
  assign n8644 = ( x102 & ~n8329 ) | ( x102 & n8643 ) | ( ~n8329 & n8643 ) ;
  assign n8645 = ( x103 & ~n8321 ) | ( x103 & n8644 ) | ( ~n8321 & n8644 ) ;
  assign n8646 = ( x104 & ~n8313 ) | ( x104 & n8645 ) | ( ~n8313 & n8645 ) ;
  assign n8647 = ( x105 & ~n8305 ) | ( x105 & n8646 ) | ( ~n8305 & n8646 ) ;
  assign n8648 = ( x106 & ~n8297 ) | ( x106 & n8647 ) | ( ~n8297 & n8647 ) ;
  assign n8649 = n250 | n252 ;
  assign n8650 = n240 | n8649 ;
  assign n8651 = n8648 | n8650 ;
  assign n8923 = n8305 &  n8651 ;
  assign n8927 = x105 | n8305 ;
  assign n8928 = x105 &  n8305 ;
  assign n8929 = ( n8927 & ~n8928 ) | ( n8927 & 1'b0 ) | ( ~n8928 & 1'b0 ) ;
  assign n8930 = ( n8646 & n8648 ) | ( n8646 & n8929 ) | ( n8648 & n8929 ) ;
  assign n8931 = ( n8646 & ~n8650 ) | ( n8646 & n8929 ) | ( ~n8650 & n8929 ) ;
  assign n8932 = ~n8930 & n8931 ;
  assign n8933 = n8923 | n8932 ;
  assign n8934 = n8313 &  n8651 ;
  assign n8924 = x104 | n8313 ;
  assign n8925 = x104 &  n8313 ;
  assign n8926 = ( n8924 & ~n8925 ) | ( n8924 & 1'b0 ) | ( ~n8925 & 1'b0 ) ;
  assign n8938 = ( n8645 & n8648 ) | ( n8645 & n8926 ) | ( n8648 & n8926 ) ;
  assign n8939 = ( n8645 & ~n8650 ) | ( n8645 & n8926 ) | ( ~n8650 & n8926 ) ;
  assign n8940 = ~n8938 & n8939 ;
  assign n8941 = n8934 | n8940 ;
  assign n8942 = n8321 &  n8651 ;
  assign n8935 = x103 | n8321 ;
  assign n8936 = x103 &  n8321 ;
  assign n8937 = ( n8935 & ~n8936 ) | ( n8935 & 1'b0 ) | ( ~n8936 & 1'b0 ) ;
  assign n8946 = ( n8644 & n8648 ) | ( n8644 & n8937 ) | ( n8648 & n8937 ) ;
  assign n8947 = ( n8644 & ~n8650 ) | ( n8644 & n8937 ) | ( ~n8650 & n8937 ) ;
  assign n8948 = ~n8946 & n8947 ;
  assign n8949 = n8942 | n8948 ;
  assign n8950 = n8329 &  n8651 ;
  assign n8943 = x102 | n8329 ;
  assign n8944 = x102 &  n8329 ;
  assign n8945 = ( n8943 & ~n8944 ) | ( n8943 & 1'b0 ) | ( ~n8944 & 1'b0 ) ;
  assign n8954 = ( n8643 & n8648 ) | ( n8643 & n8945 ) | ( n8648 & n8945 ) ;
  assign n8955 = ( n8643 & ~n8650 ) | ( n8643 & n8945 ) | ( ~n8650 & n8945 ) ;
  assign n8956 = ~n8954 & n8955 ;
  assign n8957 = n8950 | n8956 ;
  assign n8958 = n8337 &  n8651 ;
  assign n8951 = x101 | n8337 ;
  assign n8952 = x101 &  n8337 ;
  assign n8953 = ( n8951 & ~n8952 ) | ( n8951 & 1'b0 ) | ( ~n8952 & 1'b0 ) ;
  assign n8962 = ( n8642 & n8648 ) | ( n8642 & n8953 ) | ( n8648 & n8953 ) ;
  assign n8963 = ( n8642 & ~n8650 ) | ( n8642 & n8953 ) | ( ~n8650 & n8953 ) ;
  assign n8964 = ~n8962 & n8963 ;
  assign n8965 = n8958 | n8964 ;
  assign n8966 = n8345 &  n8651 ;
  assign n8959 = x100 | n8345 ;
  assign n8960 = x100 &  n8345 ;
  assign n8961 = ( n8959 & ~n8960 ) | ( n8959 & 1'b0 ) | ( ~n8960 & 1'b0 ) ;
  assign n8970 = ( n8641 & n8648 ) | ( n8641 & n8961 ) | ( n8648 & n8961 ) ;
  assign n8971 = ( n8641 & ~n8650 ) | ( n8641 & n8961 ) | ( ~n8650 & n8961 ) ;
  assign n8972 = ~n8970 & n8971 ;
  assign n8973 = n8966 | n8972 ;
  assign n8974 = n8353 &  n8651 ;
  assign n8967 = x99 | n8353 ;
  assign n8968 = x99 &  n8353 ;
  assign n8969 = ( n8967 & ~n8968 ) | ( n8967 & 1'b0 ) | ( ~n8968 & 1'b0 ) ;
  assign n8978 = ( n8640 & n8648 ) | ( n8640 & n8969 ) | ( n8648 & n8969 ) ;
  assign n8979 = ( n8640 & ~n8650 ) | ( n8640 & n8969 ) | ( ~n8650 & n8969 ) ;
  assign n8980 = ~n8978 & n8979 ;
  assign n8981 = n8974 | n8980 ;
  assign n8982 = n8361 &  n8651 ;
  assign n8975 = x98 | n8361 ;
  assign n8976 = x98 &  n8361 ;
  assign n8977 = ( n8975 & ~n8976 ) | ( n8975 & 1'b0 ) | ( ~n8976 & 1'b0 ) ;
  assign n8986 = ( n8639 & n8648 ) | ( n8639 & n8977 ) | ( n8648 & n8977 ) ;
  assign n8987 = ( n8639 & ~n8650 ) | ( n8639 & n8977 ) | ( ~n8650 & n8977 ) ;
  assign n8988 = ~n8986 & n8987 ;
  assign n8989 = n8982 | n8988 ;
  assign n8990 = n8369 &  n8651 ;
  assign n8983 = x97 | n8369 ;
  assign n8984 = x97 &  n8369 ;
  assign n8985 = ( n8983 & ~n8984 ) | ( n8983 & 1'b0 ) | ( ~n8984 & 1'b0 ) ;
  assign n8994 = ( n8638 & n8648 ) | ( n8638 & n8985 ) | ( n8648 & n8985 ) ;
  assign n8995 = ( n8638 & ~n8650 ) | ( n8638 & n8985 ) | ( ~n8650 & n8985 ) ;
  assign n8996 = ~n8994 & n8995 ;
  assign n8997 = n8990 | n8996 ;
  assign n8998 = n8377 &  n8651 ;
  assign n8991 = x96 | n8377 ;
  assign n8992 = x96 &  n8377 ;
  assign n8993 = ( n8991 & ~n8992 ) | ( n8991 & 1'b0 ) | ( ~n8992 & 1'b0 ) ;
  assign n9002 = ( n8637 & n8648 ) | ( n8637 & n8993 ) | ( n8648 & n8993 ) ;
  assign n9003 = ( n8637 & ~n8650 ) | ( n8637 & n8993 ) | ( ~n8650 & n8993 ) ;
  assign n9004 = ~n9002 & n9003 ;
  assign n9005 = n8998 | n9004 ;
  assign n9006 = n8385 &  n8651 ;
  assign n8999 = x95 | n8385 ;
  assign n9000 = x95 &  n8385 ;
  assign n9001 = ( n8999 & ~n9000 ) | ( n8999 & 1'b0 ) | ( ~n9000 & 1'b0 ) ;
  assign n9010 = ( n8636 & n8648 ) | ( n8636 & n9001 ) | ( n8648 & n9001 ) ;
  assign n9011 = ( n8636 & ~n8650 ) | ( n8636 & n9001 ) | ( ~n8650 & n9001 ) ;
  assign n9012 = ~n9010 & n9011 ;
  assign n9013 = n9006 | n9012 ;
  assign n9014 = n8393 &  n8651 ;
  assign n9007 = x94 | n8393 ;
  assign n9008 = x94 &  n8393 ;
  assign n9009 = ( n9007 & ~n9008 ) | ( n9007 & 1'b0 ) | ( ~n9008 & 1'b0 ) ;
  assign n9018 = ( n8635 & n8648 ) | ( n8635 & n9009 ) | ( n8648 & n9009 ) ;
  assign n9019 = ( n8635 & ~n8650 ) | ( n8635 & n9009 ) | ( ~n8650 & n9009 ) ;
  assign n9020 = ~n9018 & n9019 ;
  assign n9021 = n9014 | n9020 ;
  assign n9022 = n8401 &  n8651 ;
  assign n9015 = x93 | n8401 ;
  assign n9016 = x93 &  n8401 ;
  assign n9017 = ( n9015 & ~n9016 ) | ( n9015 & 1'b0 ) | ( ~n9016 & 1'b0 ) ;
  assign n9023 = ( n8634 & n8648 ) | ( n8634 & n9017 ) | ( n8648 & n9017 ) ;
  assign n9024 = ( n8634 & ~n8650 ) | ( n8634 & n9017 ) | ( ~n8650 & n9017 ) ;
  assign n9025 = ~n9023 & n9024 ;
  assign n9026 = n9022 | n9025 ;
  assign n8912 = n8406 &  n8651 ;
  assign n8913 = x92 | n8406 ;
  assign n8914 = x92 &  n8406 ;
  assign n8915 = ( n8913 & ~n8914 ) | ( n8913 & 1'b0 ) | ( ~n8914 & 1'b0 ) ;
  assign n8916 = ( n8633 & n8648 ) | ( n8633 & n8915 ) | ( n8648 & n8915 ) ;
  assign n8917 = ( n8633 & ~n8650 ) | ( n8633 & n8915 ) | ( ~n8650 & n8915 ) ;
  assign n8918 = ~n8916 & n8917 ;
  assign n8919 = n8912 | n8918 ;
  assign n8652 = n8287 &  n8651 ;
  assign n8656 = x91 | n8287 ;
  assign n8657 = x91 &  n8287 ;
  assign n8658 = ( n8656 & ~n8657 ) | ( n8656 & 1'b0 ) | ( ~n8657 & 1'b0 ) ;
  assign n8659 = ( n8632 & n8648 ) | ( n8632 & n8658 ) | ( n8648 & n8658 ) ;
  assign n8660 = ( n8632 & ~n8650 ) | ( n8632 & n8658 ) | ( ~n8650 & n8658 ) ;
  assign n8661 = ~n8659 & n8660 ;
  assign n8662 = n8652 | n8661 ;
  assign n8663 = n8414 &  n8651 ;
  assign n8653 = x90 | n8414 ;
  assign n8654 = x90 &  n8414 ;
  assign n8655 = ( n8653 & ~n8654 ) | ( n8653 & 1'b0 ) | ( ~n8654 & 1'b0 ) ;
  assign n8667 = ( n8631 & n8648 ) | ( n8631 & n8655 ) | ( n8648 & n8655 ) ;
  assign n8668 = ( n8631 & ~n8650 ) | ( n8631 & n8655 ) | ( ~n8650 & n8655 ) ;
  assign n8669 = ~n8667 & n8668 ;
  assign n8670 = n8663 | n8669 ;
  assign n8671 = n8422 &  n8651 ;
  assign n8664 = x89 | n8422 ;
  assign n8665 = x89 &  n8422 ;
  assign n8666 = ( n8664 & ~n8665 ) | ( n8664 & 1'b0 ) | ( ~n8665 & 1'b0 ) ;
  assign n8675 = ( n8630 & n8648 ) | ( n8630 & n8666 ) | ( n8648 & n8666 ) ;
  assign n8676 = ( n8630 & ~n8650 ) | ( n8630 & n8666 ) | ( ~n8650 & n8666 ) ;
  assign n8677 = ~n8675 & n8676 ;
  assign n8678 = n8671 | n8677 ;
  assign n8679 = n8430 &  n8651 ;
  assign n8672 = x88 | n8430 ;
  assign n8673 = x88 &  n8430 ;
  assign n8674 = ( n8672 & ~n8673 ) | ( n8672 & 1'b0 ) | ( ~n8673 & 1'b0 ) ;
  assign n8683 = ( n8629 & n8648 ) | ( n8629 & n8674 ) | ( n8648 & n8674 ) ;
  assign n8684 = ( n8629 & ~n8650 ) | ( n8629 & n8674 ) | ( ~n8650 & n8674 ) ;
  assign n8685 = ~n8683 & n8684 ;
  assign n8686 = n8679 | n8685 ;
  assign n8687 = n8438 &  n8651 ;
  assign n8680 = x87 | n8438 ;
  assign n8681 = x87 &  n8438 ;
  assign n8682 = ( n8680 & ~n8681 ) | ( n8680 & 1'b0 ) | ( ~n8681 & 1'b0 ) ;
  assign n8691 = ( n8628 & n8648 ) | ( n8628 & n8682 ) | ( n8648 & n8682 ) ;
  assign n8692 = ( n8628 & ~n8650 ) | ( n8628 & n8682 ) | ( ~n8650 & n8682 ) ;
  assign n8693 = ~n8691 & n8692 ;
  assign n8694 = n8687 | n8693 ;
  assign n8695 = n8446 &  n8651 ;
  assign n8688 = x86 | n8446 ;
  assign n8689 = x86 &  n8446 ;
  assign n8690 = ( n8688 & ~n8689 ) | ( n8688 & 1'b0 ) | ( ~n8689 & 1'b0 ) ;
  assign n8699 = ( n8627 & n8648 ) | ( n8627 & n8690 ) | ( n8648 & n8690 ) ;
  assign n8700 = ( n8627 & ~n8650 ) | ( n8627 & n8690 ) | ( ~n8650 & n8690 ) ;
  assign n8701 = ~n8699 & n8700 ;
  assign n8702 = n8695 | n8701 ;
  assign n8703 = n8454 &  n8651 ;
  assign n8696 = x85 | n8454 ;
  assign n8697 = x85 &  n8454 ;
  assign n8698 = ( n8696 & ~n8697 ) | ( n8696 & 1'b0 ) | ( ~n8697 & 1'b0 ) ;
  assign n8707 = ( n8626 & n8648 ) | ( n8626 & n8698 ) | ( n8648 & n8698 ) ;
  assign n8708 = ( n8626 & ~n8650 ) | ( n8626 & n8698 ) | ( ~n8650 & n8698 ) ;
  assign n8709 = ~n8707 & n8708 ;
  assign n8710 = n8703 | n8709 ;
  assign n8711 = n8462 &  n8651 ;
  assign n8704 = x84 | n8462 ;
  assign n8705 = x84 &  n8462 ;
  assign n8706 = ( n8704 & ~n8705 ) | ( n8704 & 1'b0 ) | ( ~n8705 & 1'b0 ) ;
  assign n8715 = ( n8625 & n8648 ) | ( n8625 & n8706 ) | ( n8648 & n8706 ) ;
  assign n8716 = ( n8625 & ~n8650 ) | ( n8625 & n8706 ) | ( ~n8650 & n8706 ) ;
  assign n8717 = ~n8715 & n8716 ;
  assign n8718 = n8711 | n8717 ;
  assign n8719 = n8470 &  n8651 ;
  assign n8712 = x83 | n8470 ;
  assign n8713 = x83 &  n8470 ;
  assign n8714 = ( n8712 & ~n8713 ) | ( n8712 & 1'b0 ) | ( ~n8713 & 1'b0 ) ;
  assign n8723 = ( n8624 & n8648 ) | ( n8624 & n8714 ) | ( n8648 & n8714 ) ;
  assign n8724 = ( n8624 & ~n8650 ) | ( n8624 & n8714 ) | ( ~n8650 & n8714 ) ;
  assign n8725 = ~n8723 & n8724 ;
  assign n8726 = n8719 | n8725 ;
  assign n8727 = n8478 &  n8651 ;
  assign n8720 = x82 | n8478 ;
  assign n8721 = x82 &  n8478 ;
  assign n8722 = ( n8720 & ~n8721 ) | ( n8720 & 1'b0 ) | ( ~n8721 & 1'b0 ) ;
  assign n8731 = ( n8623 & n8648 ) | ( n8623 & n8722 ) | ( n8648 & n8722 ) ;
  assign n8732 = ( n8623 & ~n8650 ) | ( n8623 & n8722 ) | ( ~n8650 & n8722 ) ;
  assign n8733 = ~n8731 & n8732 ;
  assign n8734 = n8727 | n8733 ;
  assign n8735 = n8486 &  n8651 ;
  assign n8728 = x81 | n8486 ;
  assign n8729 = x81 &  n8486 ;
  assign n8730 = ( n8728 & ~n8729 ) | ( n8728 & 1'b0 ) | ( ~n8729 & 1'b0 ) ;
  assign n8739 = ( n8622 & n8648 ) | ( n8622 & n8730 ) | ( n8648 & n8730 ) ;
  assign n8740 = ( n8622 & ~n8650 ) | ( n8622 & n8730 ) | ( ~n8650 & n8730 ) ;
  assign n8741 = ~n8739 & n8740 ;
  assign n8742 = n8735 | n8741 ;
  assign n8743 = n8494 &  n8651 ;
  assign n8736 = x80 | n8494 ;
  assign n8737 = x80 &  n8494 ;
  assign n8738 = ( n8736 & ~n8737 ) | ( n8736 & 1'b0 ) | ( ~n8737 & 1'b0 ) ;
  assign n8747 = ( n8621 & n8648 ) | ( n8621 & n8738 ) | ( n8648 & n8738 ) ;
  assign n8748 = ( n8621 & ~n8650 ) | ( n8621 & n8738 ) | ( ~n8650 & n8738 ) ;
  assign n8749 = ~n8747 & n8748 ;
  assign n8750 = n8743 | n8749 ;
  assign n8751 = n8502 &  n8651 ;
  assign n8744 = x79 | n8502 ;
  assign n8745 = x79 &  n8502 ;
  assign n8746 = ( n8744 & ~n8745 ) | ( n8744 & 1'b0 ) | ( ~n8745 & 1'b0 ) ;
  assign n8755 = ( n8620 & n8648 ) | ( n8620 & n8746 ) | ( n8648 & n8746 ) ;
  assign n8756 = ( n8620 & ~n8650 ) | ( n8620 & n8746 ) | ( ~n8650 & n8746 ) ;
  assign n8757 = ~n8755 & n8756 ;
  assign n8758 = n8751 | n8757 ;
  assign n8759 = n8510 &  n8651 ;
  assign n8752 = x78 | n8510 ;
  assign n8753 = x78 &  n8510 ;
  assign n8754 = ( n8752 & ~n8753 ) | ( n8752 & 1'b0 ) | ( ~n8753 & 1'b0 ) ;
  assign n8763 = ( n8619 & n8648 ) | ( n8619 & n8754 ) | ( n8648 & n8754 ) ;
  assign n8764 = ( n8619 & ~n8650 ) | ( n8619 & n8754 ) | ( ~n8650 & n8754 ) ;
  assign n8765 = ~n8763 & n8764 ;
  assign n8766 = n8759 | n8765 ;
  assign n8767 = n8518 &  n8651 ;
  assign n8760 = x77 | n8518 ;
  assign n8761 = x77 &  n8518 ;
  assign n8762 = ( n8760 & ~n8761 ) | ( n8760 & 1'b0 ) | ( ~n8761 & 1'b0 ) ;
  assign n8771 = ( n8618 & n8648 ) | ( n8618 & n8762 ) | ( n8648 & n8762 ) ;
  assign n8772 = ( n8618 & ~n8650 ) | ( n8618 & n8762 ) | ( ~n8650 & n8762 ) ;
  assign n8773 = ~n8771 & n8772 ;
  assign n8774 = n8767 | n8773 ;
  assign n8775 = n8526 &  n8651 ;
  assign n8768 = x76 | n8526 ;
  assign n8769 = x76 &  n8526 ;
  assign n8770 = ( n8768 & ~n8769 ) | ( n8768 & 1'b0 ) | ( ~n8769 & 1'b0 ) ;
  assign n8779 = ( n8617 & n8648 ) | ( n8617 & n8770 ) | ( n8648 & n8770 ) ;
  assign n8780 = ( n8617 & ~n8650 ) | ( n8617 & n8770 ) | ( ~n8650 & n8770 ) ;
  assign n8781 = ~n8779 & n8780 ;
  assign n8782 = n8775 | n8781 ;
  assign n8783 = n8534 &  n8651 ;
  assign n8776 = x75 | n8534 ;
  assign n8777 = x75 &  n8534 ;
  assign n8778 = ( n8776 & ~n8777 ) | ( n8776 & 1'b0 ) | ( ~n8777 & 1'b0 ) ;
  assign n8787 = ( n8616 & n8648 ) | ( n8616 & n8778 ) | ( n8648 & n8778 ) ;
  assign n8788 = ( n8616 & ~n8650 ) | ( n8616 & n8778 ) | ( ~n8650 & n8778 ) ;
  assign n8789 = ~n8787 & n8788 ;
  assign n8790 = n8783 | n8789 ;
  assign n8791 = n8542 &  n8651 ;
  assign n8784 = x74 | n8542 ;
  assign n8785 = x74 &  n8542 ;
  assign n8786 = ( n8784 & ~n8785 ) | ( n8784 & 1'b0 ) | ( ~n8785 & 1'b0 ) ;
  assign n8795 = ( n8615 & n8648 ) | ( n8615 & n8786 ) | ( n8648 & n8786 ) ;
  assign n8796 = ( n8615 & ~n8650 ) | ( n8615 & n8786 ) | ( ~n8650 & n8786 ) ;
  assign n8797 = ~n8795 & n8796 ;
  assign n8798 = n8791 | n8797 ;
  assign n8799 = n8550 &  n8651 ;
  assign n8792 = x73 | n8550 ;
  assign n8793 = x73 &  n8550 ;
  assign n8794 = ( n8792 & ~n8793 ) | ( n8792 & 1'b0 ) | ( ~n8793 & 1'b0 ) ;
  assign n8803 = ( n8614 & n8648 ) | ( n8614 & n8794 ) | ( n8648 & n8794 ) ;
  assign n8804 = ( n8614 & ~n8650 ) | ( n8614 & n8794 ) | ( ~n8650 & n8794 ) ;
  assign n8805 = ~n8803 & n8804 ;
  assign n8806 = n8799 | n8805 ;
  assign n8807 = n8558 &  n8651 ;
  assign n8800 = x72 | n8558 ;
  assign n8801 = x72 &  n8558 ;
  assign n8802 = ( n8800 & ~n8801 ) | ( n8800 & 1'b0 ) | ( ~n8801 & 1'b0 ) ;
  assign n8811 = ( n8613 & n8648 ) | ( n8613 & n8802 ) | ( n8648 & n8802 ) ;
  assign n8812 = ( n8613 & ~n8650 ) | ( n8613 & n8802 ) | ( ~n8650 & n8802 ) ;
  assign n8813 = ~n8811 & n8812 ;
  assign n8814 = n8807 | n8813 ;
  assign n8815 = n8566 &  n8651 ;
  assign n8808 = x71 | n8566 ;
  assign n8809 = x71 &  n8566 ;
  assign n8810 = ( n8808 & ~n8809 ) | ( n8808 & 1'b0 ) | ( ~n8809 & 1'b0 ) ;
  assign n8819 = ( n8612 & n8648 ) | ( n8612 & n8810 ) | ( n8648 & n8810 ) ;
  assign n8820 = ( n8612 & ~n8650 ) | ( n8612 & n8810 ) | ( ~n8650 & n8810 ) ;
  assign n8821 = ~n8819 & n8820 ;
  assign n8822 = n8815 | n8821 ;
  assign n8823 = n8574 &  n8651 ;
  assign n8816 = x70 | n8574 ;
  assign n8817 = x70 &  n8574 ;
  assign n8818 = ( n8816 & ~n8817 ) | ( n8816 & 1'b0 ) | ( ~n8817 & 1'b0 ) ;
  assign n8827 = ( n8611 & n8648 ) | ( n8611 & n8818 ) | ( n8648 & n8818 ) ;
  assign n8828 = ( n8611 & ~n8650 ) | ( n8611 & n8818 ) | ( ~n8650 & n8818 ) ;
  assign n8829 = ~n8827 & n8828 ;
  assign n8830 = n8823 | n8829 ;
  assign n8831 = n8582 &  n8651 ;
  assign n8824 = x69 | n8582 ;
  assign n8825 = x69 &  n8582 ;
  assign n8826 = ( n8824 & ~n8825 ) | ( n8824 & 1'b0 ) | ( ~n8825 & 1'b0 ) ;
  assign n8835 = ( n8610 & n8648 ) | ( n8610 & n8826 ) | ( n8648 & n8826 ) ;
  assign n8836 = ( n8610 & ~n8650 ) | ( n8610 & n8826 ) | ( ~n8650 & n8826 ) ;
  assign n8837 = ~n8835 & n8836 ;
  assign n8838 = n8831 | n8837 ;
  assign n8839 = n8590 &  n8651 ;
  assign n8832 = x68 | n8590 ;
  assign n8833 = x68 &  n8590 ;
  assign n8834 = ( n8832 & ~n8833 ) | ( n8832 & 1'b0 ) | ( ~n8833 & 1'b0 ) ;
  assign n8843 = ( n8609 & n8648 ) | ( n8609 & n8834 ) | ( n8648 & n8834 ) ;
  assign n8844 = ( n8609 & ~n8650 ) | ( n8609 & n8834 ) | ( ~n8650 & n8834 ) ;
  assign n8845 = ~n8843 & n8844 ;
  assign n8846 = n8839 | n8845 ;
  assign n8847 = n8595 &  n8651 ;
  assign n8840 = x67 | n8595 ;
  assign n8841 = x67 &  n8595 ;
  assign n8842 = ( n8840 & ~n8841 ) | ( n8840 & 1'b0 ) | ( ~n8841 & 1'b0 ) ;
  assign n8851 = ( n8608 & n8648 ) | ( n8608 & n8842 ) | ( n8648 & n8842 ) ;
  assign n8852 = ( n8608 & ~n8650 ) | ( n8608 & n8842 ) | ( ~n8650 & n8842 ) ;
  assign n8853 = ~n8851 & n8852 ;
  assign n8854 = n8847 | n8853 ;
  assign n8855 = n8601 &  n8651 ;
  assign n8848 = x66 | n8601 ;
  assign n8849 = x66 &  n8601 ;
  assign n8850 = ( n8848 & ~n8849 ) | ( n8848 & 1'b0 ) | ( ~n8849 & 1'b0 ) ;
  assign n8860 = ( n8607 & ~n8648 ) | ( n8607 & n8850 ) | ( ~n8648 & n8850 ) ;
  assign n8861 = ( n8607 & n8650 ) | ( n8607 & n8850 ) | ( n8650 & n8850 ) ;
  assign n8862 = ( n8860 & ~n8861 ) | ( n8860 & 1'b0 ) | ( ~n8861 & 1'b0 ) ;
  assign n8863 = n8855 | n8862 ;
  assign n8864 = n8605 &  n8651 ;
  assign n8856 = x65 &  n8605 ;
  assign n8857 = ( n8603 & ~x65 ) | ( n8603 & n8604 ) | ( ~x65 & n8604 ) ;
  assign n8858 = x65 | n8857 ;
  assign n8859 = ( n8606 & ~n8856 ) | ( n8606 & n8858 ) | ( ~n8856 & n8858 ) ;
  assign n8865 = ( x65 & n8605 ) | ( x65 & n8606 ) | ( n8605 & n8606 ) ;
  assign n8866 = ( n8650 & ~n8856 ) | ( n8650 & n8865 ) | ( ~n8856 & n8865 ) ;
  assign n8867 = ( n8648 & n8859 ) | ( n8648 & n8866 ) | ( n8859 & n8866 ) ;
  assign n8868 = ( n8859 & ~n8867 ) | ( n8859 & 1'b0 ) | ( ~n8867 & 1'b0 ) ;
  assign n8869 = n8864 | n8868 ;
  assign n8870 = ( x64 & ~x107 ) | ( x64 & 1'b0 ) | ( ~x107 & 1'b0 ) ;
  assign n8871 = ( n173 & ~n270 ) | ( n173 & n8870 ) | ( ~n270 & n8870 ) ;
  assign n8872 = ~n173 & n8871 ;
  assign n8873 = n8648 &  n8872 ;
  assign n8874 = ( x21 & ~n8872 ) | ( x21 & n8873 ) | ( ~n8872 & n8873 ) ;
  assign n8875 = ~n252 & n8606 ;
  assign n8876 = ( n240 & ~n250 ) | ( n240 & n8875 ) | ( ~n250 & n8875 ) ;
  assign n8877 = ~n240 & n8876 ;
  assign n8878 = ~n8648 & n8877 ;
  assign n8879 = n8874 | n8878 ;
  assign n8880 = ~x20 & x64 ;
  assign n8881 = ( x65 & ~n8879 ) | ( x65 & n8880 ) | ( ~n8879 & n8880 ) ;
  assign n8882 = ( x66 & ~n8869 ) | ( x66 & n8881 ) | ( ~n8869 & n8881 ) ;
  assign n8883 = ( x67 & ~n8863 ) | ( x67 & n8882 ) | ( ~n8863 & n8882 ) ;
  assign n8884 = ( x68 & ~n8854 ) | ( x68 & n8883 ) | ( ~n8854 & n8883 ) ;
  assign n8885 = ( x69 & ~n8846 ) | ( x69 & n8884 ) | ( ~n8846 & n8884 ) ;
  assign n8886 = ( x70 & ~n8838 ) | ( x70 & n8885 ) | ( ~n8838 & n8885 ) ;
  assign n8887 = ( x71 & ~n8830 ) | ( x71 & n8886 ) | ( ~n8830 & n8886 ) ;
  assign n8888 = ( x72 & ~n8822 ) | ( x72 & n8887 ) | ( ~n8822 & n8887 ) ;
  assign n8889 = ( x73 & ~n8814 ) | ( x73 & n8888 ) | ( ~n8814 & n8888 ) ;
  assign n8890 = ( x74 & ~n8806 ) | ( x74 & n8889 ) | ( ~n8806 & n8889 ) ;
  assign n8891 = ( x75 & ~n8798 ) | ( x75 & n8890 ) | ( ~n8798 & n8890 ) ;
  assign n8892 = ( x76 & ~n8790 ) | ( x76 & n8891 ) | ( ~n8790 & n8891 ) ;
  assign n8893 = ( x77 & ~n8782 ) | ( x77 & n8892 ) | ( ~n8782 & n8892 ) ;
  assign n8894 = ( x78 & ~n8774 ) | ( x78 & n8893 ) | ( ~n8774 & n8893 ) ;
  assign n8895 = ( x79 & ~n8766 ) | ( x79 & n8894 ) | ( ~n8766 & n8894 ) ;
  assign n8896 = ( x80 & ~n8758 ) | ( x80 & n8895 ) | ( ~n8758 & n8895 ) ;
  assign n8897 = ( x81 & ~n8750 ) | ( x81 & n8896 ) | ( ~n8750 & n8896 ) ;
  assign n8898 = ( x82 & ~n8742 ) | ( x82 & n8897 ) | ( ~n8742 & n8897 ) ;
  assign n8899 = ( x83 & ~n8734 ) | ( x83 & n8898 ) | ( ~n8734 & n8898 ) ;
  assign n8900 = ( x84 & ~n8726 ) | ( x84 & n8899 ) | ( ~n8726 & n8899 ) ;
  assign n8901 = ( x85 & ~n8718 ) | ( x85 & n8900 ) | ( ~n8718 & n8900 ) ;
  assign n8902 = ( x86 & ~n8710 ) | ( x86 & n8901 ) | ( ~n8710 & n8901 ) ;
  assign n8903 = ( x87 & ~n8702 ) | ( x87 & n8902 ) | ( ~n8702 & n8902 ) ;
  assign n8904 = ( x88 & ~n8694 ) | ( x88 & n8903 ) | ( ~n8694 & n8903 ) ;
  assign n8905 = ( x89 & ~n8686 ) | ( x89 & n8904 ) | ( ~n8686 & n8904 ) ;
  assign n8906 = ( x90 & ~n8678 ) | ( x90 & n8905 ) | ( ~n8678 & n8905 ) ;
  assign n8907 = ( x91 & ~n8670 ) | ( x91 & n8906 ) | ( ~n8670 & n8906 ) ;
  assign n8911 = ( x92 & ~n8662 ) | ( x92 & n8907 ) | ( ~n8662 & n8907 ) ;
  assign n9027 = ( x93 & ~n8919 ) | ( x93 & n8911 ) | ( ~n8919 & n8911 ) ;
  assign n9028 = ( x94 & ~n9026 ) | ( x94 & n9027 ) | ( ~n9026 & n9027 ) ;
  assign n9029 = ( x95 & ~n9021 ) | ( x95 & n9028 ) | ( ~n9021 & n9028 ) ;
  assign n9030 = ( x96 & ~n9013 ) | ( x96 & n9029 ) | ( ~n9013 & n9029 ) ;
  assign n9031 = ( x97 & ~n9005 ) | ( x97 & n9030 ) | ( ~n9005 & n9030 ) ;
  assign n9032 = ( x98 & ~n8997 ) | ( x98 & n9031 ) | ( ~n8997 & n9031 ) ;
  assign n9033 = ( x99 & ~n8989 ) | ( x99 & n9032 ) | ( ~n8989 & n9032 ) ;
  assign n9034 = ( x100 & ~n8981 ) | ( x100 & n9033 ) | ( ~n8981 & n9033 ) ;
  assign n9035 = ( x101 & ~n8973 ) | ( x101 & n9034 ) | ( ~n8973 & n9034 ) ;
  assign n9036 = ( x102 & ~n8965 ) | ( x102 & n9035 ) | ( ~n8965 & n9035 ) ;
  assign n9037 = ( x103 & ~n8957 ) | ( x103 & n9036 ) | ( ~n8957 & n9036 ) ;
  assign n9038 = ( x104 & ~n8949 ) | ( x104 & n9037 ) | ( ~n8949 & n9037 ) ;
  assign n9039 = ( x105 & ~n8941 ) | ( x105 & n9038 ) | ( ~n8941 & n9038 ) ;
  assign n9040 = ( x106 & ~n8933 ) | ( x106 & n9039 ) | ( ~n8933 & n9039 ) ;
  assign n9044 = n160 | n174 ;
  assign n9041 = x106 | n8647 ;
  assign n9042 = ( x106 & n8647 ) | ( x106 & n8650 ) | ( n8647 & n8650 ) ;
  assign n9043 = ( n8297 & ~n9041 ) | ( n8297 & n9042 ) | ( ~n9041 & n9042 ) ;
  assign n9046 = x107 &  n9043 ;
  assign n9045 = x107 | n9043 ;
  assign n9047 = ( n9044 & ~n9046 ) | ( n9044 & n9045 ) | ( ~n9046 & n9045 ) ;
  assign n9048 = n9040 | n9047 ;
  assign n9049 = ~n9043 |  n8650 ;
  assign n9330 = n8933 &  n9049 ;
  assign n9331 = n9048 &  n9330 ;
  assign n9327 = x106 | n8933 ;
  assign n9328 = x106 &  n8933 ;
  assign n9329 = ( n9327 & ~n9328 ) | ( n9327 & 1'b0 ) | ( ~n9328 & 1'b0 ) ;
  assign n9332 = n9039 &  n9329 ;
  assign n9050 = n9048 &  n9049 ;
  assign n9333 = ( n9039 & ~n9050 ) | ( n9039 & n9329 ) | ( ~n9050 & n9329 ) ;
  assign n9334 = ( n9331 & ~n9332 ) | ( n9331 & n9333 ) | ( ~n9332 & n9333 ) ;
  assign n9338 = n8941 &  n9049 ;
  assign n9339 = n9048 &  n9338 ;
  assign n9324 = x105 | n8941 ;
  assign n9325 = x105 &  n8941 ;
  assign n9326 = ( n9324 & ~n9325 ) | ( n9324 & 1'b0 ) | ( ~n9325 & 1'b0 ) ;
  assign n9340 = n9038 &  n9326 ;
  assign n9341 = ( n9038 & ~n9050 ) | ( n9038 & n9326 ) | ( ~n9050 & n9326 ) ;
  assign n9342 = ( n9339 & ~n9340 ) | ( n9339 & n9341 ) | ( ~n9340 & n9341 ) ;
  assign n9346 = n8949 &  n9049 ;
  assign n9347 = n9048 &  n9346 ;
  assign n9335 = x104 | n8949 ;
  assign n9336 = x104 &  n8949 ;
  assign n9337 = ( n9335 & ~n9336 ) | ( n9335 & 1'b0 ) | ( ~n9336 & 1'b0 ) ;
  assign n9348 = n9037 &  n9337 ;
  assign n9349 = ( n9037 & ~n9050 ) | ( n9037 & n9337 ) | ( ~n9050 & n9337 ) ;
  assign n9350 = ( n9347 & ~n9348 ) | ( n9347 & n9349 ) | ( ~n9348 & n9349 ) ;
  assign n9354 = n8957 &  n9049 ;
  assign n9355 = n9048 &  n9354 ;
  assign n9343 = x103 | n8957 ;
  assign n9344 = x103 &  n8957 ;
  assign n9345 = ( n9343 & ~n9344 ) | ( n9343 & 1'b0 ) | ( ~n9344 & 1'b0 ) ;
  assign n9356 = n9036 &  n9345 ;
  assign n9357 = ( n9036 & ~n9050 ) | ( n9036 & n9345 ) | ( ~n9050 & n9345 ) ;
  assign n9358 = ( n9355 & ~n9356 ) | ( n9355 & n9357 ) | ( ~n9356 & n9357 ) ;
  assign n9362 = n8965 &  n9049 ;
  assign n9363 = n9048 &  n9362 ;
  assign n9351 = x102 | n8965 ;
  assign n9352 = x102 &  n8965 ;
  assign n9353 = ( n9351 & ~n9352 ) | ( n9351 & 1'b0 ) | ( ~n9352 & 1'b0 ) ;
  assign n9364 = n9035 &  n9353 ;
  assign n9365 = ( n9035 & ~n9050 ) | ( n9035 & n9353 ) | ( ~n9050 & n9353 ) ;
  assign n9366 = ( n9363 & ~n9364 ) | ( n9363 & n9365 ) | ( ~n9364 & n9365 ) ;
  assign n9370 = n8973 &  n9049 ;
  assign n9371 = n9048 &  n9370 ;
  assign n9359 = x101 | n8973 ;
  assign n9360 = x101 &  n8973 ;
  assign n9361 = ( n9359 & ~n9360 ) | ( n9359 & 1'b0 ) | ( ~n9360 & 1'b0 ) ;
  assign n9373 = ( n9034 & n9050 ) | ( n9034 & n9361 ) | ( n9050 & n9361 ) ;
  assign n9372 = n9034 | n9361 ;
  assign n9374 = ( n9371 & ~n9373 ) | ( n9371 & n9372 ) | ( ~n9373 & n9372 ) ;
  assign n9378 = n8981 &  n9049 ;
  assign n9379 = n9048 &  n9378 ;
  assign n9367 = x100 | n8981 ;
  assign n9368 = x100 &  n8981 ;
  assign n9369 = ( n9367 & ~n9368 ) | ( n9367 & 1'b0 ) | ( ~n9368 & 1'b0 ) ;
  assign n9381 = ( n9033 & n9050 ) | ( n9033 & n9369 ) | ( n9050 & n9369 ) ;
  assign n9380 = n9033 | n9369 ;
  assign n9382 = ( n9379 & ~n9381 ) | ( n9379 & n9380 ) | ( ~n9381 & n9380 ) ;
  assign n9386 = n8989 &  n9049 ;
  assign n9387 = n9048 &  n9386 ;
  assign n9375 = x99 | n8989 ;
  assign n9376 = x99 &  n8989 ;
  assign n9377 = ( n9375 & ~n9376 ) | ( n9375 & 1'b0 ) | ( ~n9376 & 1'b0 ) ;
  assign n9389 = ( n9032 & n9050 ) | ( n9032 & n9377 ) | ( n9050 & n9377 ) ;
  assign n9388 = n9032 | n9377 ;
  assign n9390 = ( n9387 & ~n9389 ) | ( n9387 & n9388 ) | ( ~n9389 & n9388 ) ;
  assign n9394 = n8997 &  n9049 ;
  assign n9395 = n9048 &  n9394 ;
  assign n9383 = x98 | n8997 ;
  assign n9384 = x98 &  n8997 ;
  assign n9385 = ( n9383 & ~n9384 ) | ( n9383 & 1'b0 ) | ( ~n9384 & 1'b0 ) ;
  assign n9397 = ( n9031 & n9050 ) | ( n9031 & n9385 ) | ( n9050 & n9385 ) ;
  assign n9396 = n9031 | n9385 ;
  assign n9398 = ( n9395 & ~n9397 ) | ( n9395 & n9396 ) | ( ~n9397 & n9396 ) ;
  assign n9402 = n9005 &  n9049 ;
  assign n9403 = n9048 &  n9402 ;
  assign n9391 = x97 | n9005 ;
  assign n9392 = x97 &  n9005 ;
  assign n9393 = ( n9391 & ~n9392 ) | ( n9391 & 1'b0 ) | ( ~n9392 & 1'b0 ) ;
  assign n9405 = ( n9030 & n9050 ) | ( n9030 & n9393 ) | ( n9050 & n9393 ) ;
  assign n9404 = n9030 | n9393 ;
  assign n9406 = ( n9403 & ~n9405 ) | ( n9403 & n9404 ) | ( ~n9405 & n9404 ) ;
  assign n9410 = n9013 &  n9049 ;
  assign n9411 = n9048 &  n9410 ;
  assign n9399 = x96 | n9013 ;
  assign n9400 = x96 &  n9013 ;
  assign n9401 = ( n9399 & ~n9400 ) | ( n9399 & 1'b0 ) | ( ~n9400 & 1'b0 ) ;
  assign n9413 = ( n9029 & n9050 ) | ( n9029 & n9401 ) | ( n9050 & n9401 ) ;
  assign n9412 = n9029 | n9401 ;
  assign n9414 = ( n9411 & ~n9413 ) | ( n9411 & n9412 ) | ( ~n9413 & n9412 ) ;
  assign n9415 = n9021 &  n9049 ;
  assign n9416 = n9048 &  n9415 ;
  assign n9407 = x95 | n9021 ;
  assign n9408 = x95 &  n9021 ;
  assign n9409 = ( n9407 & ~n9408 ) | ( n9407 & 1'b0 ) | ( ~n9408 & 1'b0 ) ;
  assign n9418 = ( n9028 & n9050 ) | ( n9028 & n9409 ) | ( n9050 & n9409 ) ;
  assign n9417 = n9028 | n9409 ;
  assign n9419 = ( n9416 & ~n9418 ) | ( n9416 & n9417 ) | ( ~n9418 & n9417 ) ;
  assign n9316 = n9026 &  n9049 ;
  assign n9317 = n9048 &  n9316 ;
  assign n9313 = x94 | n9026 ;
  assign n9314 = x94 &  n9026 ;
  assign n9315 = ( n9313 & ~n9314 ) | ( n9313 & 1'b0 ) | ( ~n9314 & 1'b0 ) ;
  assign n9319 = ( n9027 & n9050 ) | ( n9027 & n9315 ) | ( n9050 & n9315 ) ;
  assign n9318 = n9027 | n9315 ;
  assign n9320 = ( n9317 & ~n9319 ) | ( n9317 & n9318 ) | ( ~n9319 & n9318 ) ;
  assign n9051 = n8919 &  n9049 ;
  assign n9052 = n9048 &  n9051 ;
  assign n8920 = x93 | n8919 ;
  assign n8921 = x93 &  n8919 ;
  assign n8922 = ( n8920 & ~n8921 ) | ( n8920 & 1'b0 ) | ( ~n8921 & 1'b0 ) ;
  assign n9054 = ( n8911 & n8922 ) | ( n8911 & n9050 ) | ( n8922 & n9050 ) ;
  assign n9053 = n8911 | n8922 ;
  assign n9055 = ( n9052 & ~n9054 ) | ( n9052 & n9053 ) | ( ~n9054 & n9053 ) ;
  assign n9059 = n8662 &  n9049 ;
  assign n9060 = n9048 &  n9059 ;
  assign n8908 = x92 | n8662 ;
  assign n8909 = x92 &  n8662 ;
  assign n8910 = ( n8908 & ~n8909 ) | ( n8908 & 1'b0 ) | ( ~n8909 & 1'b0 ) ;
  assign n9061 = n8907 &  n8910 ;
  assign n9062 = ( n8907 & ~n9050 ) | ( n8907 & n8910 ) | ( ~n9050 & n8910 ) ;
  assign n9063 = ( n9060 & ~n9061 ) | ( n9060 & n9062 ) | ( ~n9061 & n9062 ) ;
  assign n9067 = n8670 &  n9049 ;
  assign n9068 = n9048 &  n9067 ;
  assign n9056 = x91 | n8670 ;
  assign n9057 = x91 &  n8670 ;
  assign n9058 = ( n9056 & ~n9057 ) | ( n9056 & 1'b0 ) | ( ~n9057 & 1'b0 ) ;
  assign n9070 = ( n8906 & n9050 ) | ( n8906 & n9058 ) | ( n9050 & n9058 ) ;
  assign n9069 = n8906 | n9058 ;
  assign n9071 = ( n9068 & ~n9070 ) | ( n9068 & n9069 ) | ( ~n9070 & n9069 ) ;
  assign n9075 = n8678 &  n9049 ;
  assign n9076 = n9048 &  n9075 ;
  assign n9064 = x90 | n8678 ;
  assign n9065 = x90 &  n8678 ;
  assign n9066 = ( n9064 & ~n9065 ) | ( n9064 & 1'b0 ) | ( ~n9065 & 1'b0 ) ;
  assign n9078 = ( n8905 & n9050 ) | ( n8905 & n9066 ) | ( n9050 & n9066 ) ;
  assign n9077 = n8905 | n9066 ;
  assign n9079 = ( n9076 & ~n9078 ) | ( n9076 & n9077 ) | ( ~n9078 & n9077 ) ;
  assign n9083 = n8686 &  n9049 ;
  assign n9084 = n9048 &  n9083 ;
  assign n9072 = x89 | n8686 ;
  assign n9073 = x89 &  n8686 ;
  assign n9074 = ( n9072 & ~n9073 ) | ( n9072 & 1'b0 ) | ( ~n9073 & 1'b0 ) ;
  assign n9086 = ( n8904 & n9050 ) | ( n8904 & n9074 ) | ( n9050 & n9074 ) ;
  assign n9085 = n8904 | n9074 ;
  assign n9087 = ( n9084 & ~n9086 ) | ( n9084 & n9085 ) | ( ~n9086 & n9085 ) ;
  assign n9091 = n8694 &  n9049 ;
  assign n9092 = n9048 &  n9091 ;
  assign n9080 = x88 | n8694 ;
  assign n9081 = x88 &  n8694 ;
  assign n9082 = ( n9080 & ~n9081 ) | ( n9080 & 1'b0 ) | ( ~n9081 & 1'b0 ) ;
  assign n9094 = ( n8903 & n9050 ) | ( n8903 & n9082 ) | ( n9050 & n9082 ) ;
  assign n9093 = n8903 | n9082 ;
  assign n9095 = ( n9092 & ~n9094 ) | ( n9092 & n9093 ) | ( ~n9094 & n9093 ) ;
  assign n9099 = n8702 &  n9049 ;
  assign n9100 = n9048 &  n9099 ;
  assign n9088 = x87 | n8702 ;
  assign n9089 = x87 &  n8702 ;
  assign n9090 = ( n9088 & ~n9089 ) | ( n9088 & 1'b0 ) | ( ~n9089 & 1'b0 ) ;
  assign n9102 = ( n8902 & n9050 ) | ( n8902 & n9090 ) | ( n9050 & n9090 ) ;
  assign n9101 = n8902 | n9090 ;
  assign n9103 = ( n9100 & ~n9102 ) | ( n9100 & n9101 ) | ( ~n9102 & n9101 ) ;
  assign n9107 = n8710 &  n9049 ;
  assign n9108 = n9048 &  n9107 ;
  assign n9096 = x86 | n8710 ;
  assign n9097 = x86 &  n8710 ;
  assign n9098 = ( n9096 & ~n9097 ) | ( n9096 & 1'b0 ) | ( ~n9097 & 1'b0 ) ;
  assign n9110 = ( n8901 & n9050 ) | ( n8901 & n9098 ) | ( n9050 & n9098 ) ;
  assign n9109 = n8901 | n9098 ;
  assign n9111 = ( n9108 & ~n9110 ) | ( n9108 & n9109 ) | ( ~n9110 & n9109 ) ;
  assign n9115 = n8718 &  n9049 ;
  assign n9116 = n9048 &  n9115 ;
  assign n9104 = x85 | n8718 ;
  assign n9105 = x85 &  n8718 ;
  assign n9106 = ( n9104 & ~n9105 ) | ( n9104 & 1'b0 ) | ( ~n9105 & 1'b0 ) ;
  assign n9118 = ( n8900 & n9050 ) | ( n8900 & n9106 ) | ( n9050 & n9106 ) ;
  assign n9117 = n8900 | n9106 ;
  assign n9119 = ( n9116 & ~n9118 ) | ( n9116 & n9117 ) | ( ~n9118 & n9117 ) ;
  assign n9123 = n8726 &  n9049 ;
  assign n9124 = n9048 &  n9123 ;
  assign n9112 = x84 | n8726 ;
  assign n9113 = x84 &  n8726 ;
  assign n9114 = ( n9112 & ~n9113 ) | ( n9112 & 1'b0 ) | ( ~n9113 & 1'b0 ) ;
  assign n9126 = ( n8899 & n9050 ) | ( n8899 & n9114 ) | ( n9050 & n9114 ) ;
  assign n9125 = n8899 | n9114 ;
  assign n9127 = ( n9124 & ~n9126 ) | ( n9124 & n9125 ) | ( ~n9126 & n9125 ) ;
  assign n9131 = n8734 &  n9049 ;
  assign n9132 = n9048 &  n9131 ;
  assign n9120 = x83 | n8734 ;
  assign n9121 = x83 &  n8734 ;
  assign n9122 = ( n9120 & ~n9121 ) | ( n9120 & 1'b0 ) | ( ~n9121 & 1'b0 ) ;
  assign n9134 = ( n8898 & n9050 ) | ( n8898 & n9122 ) | ( n9050 & n9122 ) ;
  assign n9133 = n8898 | n9122 ;
  assign n9135 = ( n9132 & ~n9134 ) | ( n9132 & n9133 ) | ( ~n9134 & n9133 ) ;
  assign n9139 = n8742 &  n9049 ;
  assign n9140 = n9048 &  n9139 ;
  assign n9128 = x82 | n8742 ;
  assign n9129 = x82 &  n8742 ;
  assign n9130 = ( n9128 & ~n9129 ) | ( n9128 & 1'b0 ) | ( ~n9129 & 1'b0 ) ;
  assign n9142 = ( n8897 & n9050 ) | ( n8897 & n9130 ) | ( n9050 & n9130 ) ;
  assign n9141 = n8897 | n9130 ;
  assign n9143 = ( n9140 & ~n9142 ) | ( n9140 & n9141 ) | ( ~n9142 & n9141 ) ;
  assign n9147 = n8750 &  n9049 ;
  assign n9148 = n9048 &  n9147 ;
  assign n9136 = x81 | n8750 ;
  assign n9137 = x81 &  n8750 ;
  assign n9138 = ( n9136 & ~n9137 ) | ( n9136 & 1'b0 ) | ( ~n9137 & 1'b0 ) ;
  assign n9150 = ( n8896 & n9050 ) | ( n8896 & n9138 ) | ( n9050 & n9138 ) ;
  assign n9149 = n8896 | n9138 ;
  assign n9151 = ( n9148 & ~n9150 ) | ( n9148 & n9149 ) | ( ~n9150 & n9149 ) ;
  assign n9155 = n8758 &  n9049 ;
  assign n9156 = n9048 &  n9155 ;
  assign n9144 = x80 | n8758 ;
  assign n9145 = x80 &  n8758 ;
  assign n9146 = ( n9144 & ~n9145 ) | ( n9144 & 1'b0 ) | ( ~n9145 & 1'b0 ) ;
  assign n9158 = ( n8895 & n9050 ) | ( n8895 & n9146 ) | ( n9050 & n9146 ) ;
  assign n9157 = n8895 | n9146 ;
  assign n9159 = ( n9156 & ~n9158 ) | ( n9156 & n9157 ) | ( ~n9158 & n9157 ) ;
  assign n9163 = n8766 &  n9049 ;
  assign n9164 = n9048 &  n9163 ;
  assign n9152 = x79 | n8766 ;
  assign n9153 = x79 &  n8766 ;
  assign n9154 = ( n9152 & ~n9153 ) | ( n9152 & 1'b0 ) | ( ~n9153 & 1'b0 ) ;
  assign n9166 = ( n8894 & n9050 ) | ( n8894 & n9154 ) | ( n9050 & n9154 ) ;
  assign n9165 = n8894 | n9154 ;
  assign n9167 = ( n9164 & ~n9166 ) | ( n9164 & n9165 ) | ( ~n9166 & n9165 ) ;
  assign n9171 = n8774 &  n9049 ;
  assign n9172 = n9048 &  n9171 ;
  assign n9160 = x78 | n8774 ;
  assign n9161 = x78 &  n8774 ;
  assign n9162 = ( n9160 & ~n9161 ) | ( n9160 & 1'b0 ) | ( ~n9161 & 1'b0 ) ;
  assign n9174 = ( n8893 & n9050 ) | ( n8893 & n9162 ) | ( n9050 & n9162 ) ;
  assign n9173 = n8893 | n9162 ;
  assign n9175 = ( n9172 & ~n9174 ) | ( n9172 & n9173 ) | ( ~n9174 & n9173 ) ;
  assign n9179 = n8782 &  n9049 ;
  assign n9180 = n9048 &  n9179 ;
  assign n9168 = x77 | n8782 ;
  assign n9169 = x77 &  n8782 ;
  assign n9170 = ( n9168 & ~n9169 ) | ( n9168 & 1'b0 ) | ( ~n9169 & 1'b0 ) ;
  assign n9182 = ( n8892 & n9050 ) | ( n8892 & n9170 ) | ( n9050 & n9170 ) ;
  assign n9181 = n8892 | n9170 ;
  assign n9183 = ( n9180 & ~n9182 ) | ( n9180 & n9181 ) | ( ~n9182 & n9181 ) ;
  assign n9187 = n8790 &  n9049 ;
  assign n9188 = n9048 &  n9187 ;
  assign n9176 = x76 | n8790 ;
  assign n9177 = x76 &  n8790 ;
  assign n9178 = ( n9176 & ~n9177 ) | ( n9176 & 1'b0 ) | ( ~n9177 & 1'b0 ) ;
  assign n9190 = ( n8891 & n9050 ) | ( n8891 & n9178 ) | ( n9050 & n9178 ) ;
  assign n9189 = n8891 | n9178 ;
  assign n9191 = ( n9188 & ~n9190 ) | ( n9188 & n9189 ) | ( ~n9190 & n9189 ) ;
  assign n9195 = n8798 &  n9049 ;
  assign n9196 = n9048 &  n9195 ;
  assign n9184 = x75 | n8798 ;
  assign n9185 = x75 &  n8798 ;
  assign n9186 = ( n9184 & ~n9185 ) | ( n9184 & 1'b0 ) | ( ~n9185 & 1'b0 ) ;
  assign n9198 = ( n8890 & n9050 ) | ( n8890 & n9186 ) | ( n9050 & n9186 ) ;
  assign n9197 = n8890 | n9186 ;
  assign n9199 = ( n9196 & ~n9198 ) | ( n9196 & n9197 ) | ( ~n9198 & n9197 ) ;
  assign n9203 = n8806 &  n9049 ;
  assign n9204 = n9048 &  n9203 ;
  assign n9192 = x74 | n8806 ;
  assign n9193 = x74 &  n8806 ;
  assign n9194 = ( n9192 & ~n9193 ) | ( n9192 & 1'b0 ) | ( ~n9193 & 1'b0 ) ;
  assign n9206 = ( n8889 & n9050 ) | ( n8889 & n9194 ) | ( n9050 & n9194 ) ;
  assign n9205 = n8889 | n9194 ;
  assign n9207 = ( n9204 & ~n9206 ) | ( n9204 & n9205 ) | ( ~n9206 & n9205 ) ;
  assign n9211 = n8814 &  n9049 ;
  assign n9212 = n9048 &  n9211 ;
  assign n9200 = x73 | n8814 ;
  assign n9201 = x73 &  n8814 ;
  assign n9202 = ( n9200 & ~n9201 ) | ( n9200 & 1'b0 ) | ( ~n9201 & 1'b0 ) ;
  assign n9214 = ( n8888 & n9050 ) | ( n8888 & n9202 ) | ( n9050 & n9202 ) ;
  assign n9213 = n8888 | n9202 ;
  assign n9215 = ( n9212 & ~n9214 ) | ( n9212 & n9213 ) | ( ~n9214 & n9213 ) ;
  assign n9219 = n8822 &  n9049 ;
  assign n9220 = n9048 &  n9219 ;
  assign n9208 = x72 | n8822 ;
  assign n9209 = x72 &  n8822 ;
  assign n9210 = ( n9208 & ~n9209 ) | ( n9208 & 1'b0 ) | ( ~n9209 & 1'b0 ) ;
  assign n9222 = ( n8887 & n9050 ) | ( n8887 & n9210 ) | ( n9050 & n9210 ) ;
  assign n9221 = n8887 | n9210 ;
  assign n9223 = ( n9220 & ~n9222 ) | ( n9220 & n9221 ) | ( ~n9222 & n9221 ) ;
  assign n9227 = n8830 &  n9049 ;
  assign n9228 = n9048 &  n9227 ;
  assign n9216 = x71 | n8830 ;
  assign n9217 = x71 &  n8830 ;
  assign n9218 = ( n9216 & ~n9217 ) | ( n9216 & 1'b0 ) | ( ~n9217 & 1'b0 ) ;
  assign n9230 = ( n8886 & n9050 ) | ( n8886 & n9218 ) | ( n9050 & n9218 ) ;
  assign n9229 = n8886 | n9218 ;
  assign n9231 = ( n9228 & ~n9230 ) | ( n9228 & n9229 ) | ( ~n9230 & n9229 ) ;
  assign n9235 = n8838 &  n9049 ;
  assign n9236 = n9048 &  n9235 ;
  assign n9224 = x70 | n8838 ;
  assign n9225 = x70 &  n8838 ;
  assign n9226 = ( n9224 & ~n9225 ) | ( n9224 & 1'b0 ) | ( ~n9225 & 1'b0 ) ;
  assign n9238 = ( n8885 & n9050 ) | ( n8885 & n9226 ) | ( n9050 & n9226 ) ;
  assign n9237 = n8885 | n9226 ;
  assign n9239 = ( n9236 & ~n9238 ) | ( n9236 & n9237 ) | ( ~n9238 & n9237 ) ;
  assign n9243 = n8846 &  n9049 ;
  assign n9244 = n9048 &  n9243 ;
  assign n9232 = x69 | n8846 ;
  assign n9233 = x69 &  n8846 ;
  assign n9234 = ( n9232 & ~n9233 ) | ( n9232 & 1'b0 ) | ( ~n9233 & 1'b0 ) ;
  assign n9246 = ( n8884 & n9050 ) | ( n8884 & n9234 ) | ( n9050 & n9234 ) ;
  assign n9245 = n8884 | n9234 ;
  assign n9247 = ( n9244 & ~n9246 ) | ( n9244 & n9245 ) | ( ~n9246 & n9245 ) ;
  assign n9251 = n8854 &  n9049 ;
  assign n9252 = n9048 &  n9251 ;
  assign n9240 = x68 | n8854 ;
  assign n9241 = x68 &  n8854 ;
  assign n9242 = ( n9240 & ~n9241 ) | ( n9240 & 1'b0 ) | ( ~n9241 & 1'b0 ) ;
  assign n9254 = ( n8883 & n9050 ) | ( n8883 & n9242 ) | ( n9050 & n9242 ) ;
  assign n9253 = n8883 | n9242 ;
  assign n9255 = ( n9252 & ~n9254 ) | ( n9252 & n9253 ) | ( ~n9254 & n9253 ) ;
  assign n9259 = n8863 &  n9049 ;
  assign n9260 = n9048 &  n9259 ;
  assign n9248 = x67 | n8863 ;
  assign n9249 = x67 &  n8863 ;
  assign n9250 = ( n9248 & ~n9249 ) | ( n9248 & 1'b0 ) | ( ~n9249 & 1'b0 ) ;
  assign n9262 = ( n8882 & n9050 ) | ( n8882 & n9250 ) | ( n9050 & n9250 ) ;
  assign n9261 = n8882 | n9250 ;
  assign n9263 = ( n9260 & ~n9262 ) | ( n9260 & n9261 ) | ( ~n9262 & n9261 ) ;
  assign n9264 = n8869 &  n9049 ;
  assign n9265 = n9048 &  n9264 ;
  assign n9256 = x66 | n8869 ;
  assign n9257 = x66 &  n8869 ;
  assign n9258 = ( n9256 & ~n9257 ) | ( n9256 & 1'b0 ) | ( ~n9257 & 1'b0 ) ;
  assign n9266 = n8881 &  n9258 ;
  assign n9267 = ( n8881 & ~n9050 ) | ( n8881 & n9258 ) | ( ~n9050 & n9258 ) ;
  assign n9268 = ( n9265 & ~n9266 ) | ( n9265 & n9267 ) | ( ~n9266 & n9267 ) ;
  assign n9269 = ( n8879 & ~x65 ) | ( n8879 & n8880 ) | ( ~x65 & n8880 ) ;
  assign n9270 = ( n8881 & ~n8880 ) | ( n8881 & n9269 ) | ( ~n8880 & n9269 ) ;
  assign n9271 = ~n9050 & n9270 ;
  assign n9272 = n8879 &  n9049 ;
  assign n9273 = n9048 &  n9272 ;
  assign n9274 = n9271 | n9273 ;
  assign n9275 = ( x64 & ~n9050 ) | ( x64 & 1'b0 ) | ( ~n9050 & 1'b0 ) ;
  assign n9276 = ( x20 & ~n9275 ) | ( x20 & 1'b0 ) | ( ~n9275 & 1'b0 ) ;
  assign n9277 = ( n8880 & ~n9050 ) | ( n8880 & 1'b0 ) | ( ~n9050 & 1'b0 ) ;
  assign n9278 = n9276 | n9277 ;
  assign n9279 = ~x19 & x64 ;
  assign n9280 = ( x65 & ~n9278 ) | ( x65 & n9279 ) | ( ~n9278 & n9279 ) ;
  assign n9281 = ( x66 & ~n9274 ) | ( x66 & n9280 ) | ( ~n9274 & n9280 ) ;
  assign n9282 = ( x67 & ~n9268 ) | ( x67 & n9281 ) | ( ~n9268 & n9281 ) ;
  assign n9283 = ( x68 & ~n9263 ) | ( x68 & n9282 ) | ( ~n9263 & n9282 ) ;
  assign n9284 = ( x69 & ~n9255 ) | ( x69 & n9283 ) | ( ~n9255 & n9283 ) ;
  assign n9285 = ( x70 & ~n9247 ) | ( x70 & n9284 ) | ( ~n9247 & n9284 ) ;
  assign n9286 = ( x71 & ~n9239 ) | ( x71 & n9285 ) | ( ~n9239 & n9285 ) ;
  assign n9287 = ( x72 & ~n9231 ) | ( x72 & n9286 ) | ( ~n9231 & n9286 ) ;
  assign n9288 = ( x73 & ~n9223 ) | ( x73 & n9287 ) | ( ~n9223 & n9287 ) ;
  assign n9289 = ( x74 & ~n9215 ) | ( x74 & n9288 ) | ( ~n9215 & n9288 ) ;
  assign n9290 = ( x75 & ~n9207 ) | ( x75 & n9289 ) | ( ~n9207 & n9289 ) ;
  assign n9291 = ( x76 & ~n9199 ) | ( x76 & n9290 ) | ( ~n9199 & n9290 ) ;
  assign n9292 = ( x77 & ~n9191 ) | ( x77 & n9291 ) | ( ~n9191 & n9291 ) ;
  assign n9293 = ( x78 & ~n9183 ) | ( x78 & n9292 ) | ( ~n9183 & n9292 ) ;
  assign n9294 = ( x79 & ~n9175 ) | ( x79 & n9293 ) | ( ~n9175 & n9293 ) ;
  assign n9295 = ( x80 & ~n9167 ) | ( x80 & n9294 ) | ( ~n9167 & n9294 ) ;
  assign n9296 = ( x81 & ~n9159 ) | ( x81 & n9295 ) | ( ~n9159 & n9295 ) ;
  assign n9297 = ( x82 & ~n9151 ) | ( x82 & n9296 ) | ( ~n9151 & n9296 ) ;
  assign n9298 = ( x83 & ~n9143 ) | ( x83 & n9297 ) | ( ~n9143 & n9297 ) ;
  assign n9299 = ( x84 & ~n9135 ) | ( x84 & n9298 ) | ( ~n9135 & n9298 ) ;
  assign n9300 = ( x85 & ~n9127 ) | ( x85 & n9299 ) | ( ~n9127 & n9299 ) ;
  assign n9301 = ( x86 & ~n9119 ) | ( x86 & n9300 ) | ( ~n9119 & n9300 ) ;
  assign n9302 = ( x87 & ~n9111 ) | ( x87 & n9301 ) | ( ~n9111 & n9301 ) ;
  assign n9303 = ( x88 & ~n9103 ) | ( x88 & n9302 ) | ( ~n9103 & n9302 ) ;
  assign n9304 = ( x89 & ~n9095 ) | ( x89 & n9303 ) | ( ~n9095 & n9303 ) ;
  assign n9305 = ( x90 & ~n9087 ) | ( x90 & n9304 ) | ( ~n9087 & n9304 ) ;
  assign n9306 = ( x91 & ~n9079 ) | ( x91 & n9305 ) | ( ~n9079 & n9305 ) ;
  assign n9307 = ( x92 & ~n9071 ) | ( x92 & n9306 ) | ( ~n9071 & n9306 ) ;
  assign n9308 = ( x93 & ~n9063 ) | ( x93 & n9307 ) | ( ~n9063 & n9307 ) ;
  assign n9312 = ( x94 & ~n9055 ) | ( x94 & n9308 ) | ( ~n9055 & n9308 ) ;
  assign n9420 = ( x95 & ~n9320 ) | ( x95 & n9312 ) | ( ~n9320 & n9312 ) ;
  assign n9421 = ( x96 & ~n9419 ) | ( x96 & n9420 ) | ( ~n9419 & n9420 ) ;
  assign n9422 = ( x97 & ~n9414 ) | ( x97 & n9421 ) | ( ~n9414 & n9421 ) ;
  assign n9423 = ( x98 & ~n9406 ) | ( x98 & n9422 ) | ( ~n9406 & n9422 ) ;
  assign n9424 = ( x99 & ~n9398 ) | ( x99 & n9423 ) | ( ~n9398 & n9423 ) ;
  assign n9425 = ( x100 & ~n9390 ) | ( x100 & n9424 ) | ( ~n9390 & n9424 ) ;
  assign n9426 = ( x101 & ~n9382 ) | ( x101 & n9425 ) | ( ~n9382 & n9425 ) ;
  assign n9427 = ( x102 & ~n9374 ) | ( x102 & n9426 ) | ( ~n9374 & n9426 ) ;
  assign n9428 = ( x103 & ~n9366 ) | ( x103 & n9427 ) | ( ~n9366 & n9427 ) ;
  assign n9429 = ( x104 & ~n9358 ) | ( x104 & n9428 ) | ( ~n9358 & n9428 ) ;
  assign n9430 = ( x105 & ~n9350 ) | ( x105 & n9429 ) | ( ~n9350 & n9429 ) ;
  assign n9431 = ( x106 & ~n9342 ) | ( x106 & n9430 ) | ( ~n9342 & n9430 ) ;
  assign n9432 = ( x107 & ~n9334 ) | ( x107 & n9431 ) | ( ~n9334 & n9431 ) ;
  assign n9440 = n425 | n427 ;
  assign n9434 = ( x107 & n9040 ) | ( x107 & n9043 ) | ( n9040 & n9043 ) ;
  assign n9433 = ( x107 & ~n9040 ) | ( x107 & n9043 ) | ( ~n9040 & n9043 ) ;
  assign n9435 = ( n9040 & ~n9434 ) | ( n9040 & n9433 ) | ( ~n9434 & n9433 ) ;
  assign n9436 = ~n9050 & n9435 ;
  assign n9437 = n8297 &  n8650 ;
  assign n9438 = n9048 &  n9437 ;
  assign n9439 = n9436 | n9438 ;
  assign n9442 = x108 &  n9439 ;
  assign n9441 = x108 | n9439 ;
  assign n9443 = ( n9440 & ~n9442 ) | ( n9440 & n9441 ) | ( ~n9442 & n9441 ) ;
  assign n9444 = n9432 | n9443 ;
  assign n9445 = ~n9439 |  n9044 ;
  assign n9465 = n9334 &  n9445 ;
  assign n9466 = n9444 &  n9465 ;
  assign n9452 = x107 | n9334 ;
  assign n9453 = x107 &  n9334 ;
  assign n9454 = ( n9452 & ~n9453 ) | ( n9452 & 1'b0 ) | ( ~n9453 & 1'b0 ) ;
  assign n9467 = n9431 &  n9454 ;
  assign n9446 = n9444 &  n9445 ;
  assign n9468 = ( n9431 & ~n9446 ) | ( n9431 & n9454 ) | ( ~n9446 & n9454 ) ;
  assign n9469 = ( n9466 & ~n9467 ) | ( n9466 & n9468 ) | ( ~n9467 & n9468 ) ;
  assign n9456 = ( x108 & n9432 ) | ( x108 & n9439 ) | ( n9432 & n9439 ) ;
  assign n9455 = ( x108 & ~n9432 ) | ( x108 & n9439 ) | ( ~n9432 & n9439 ) ;
  assign n9457 = ( n9432 & ~n9456 ) | ( n9432 & n9455 ) | ( ~n9456 & n9455 ) ;
  assign n9458 = ~n9446 & n9457 ;
  assign n9459 = n9044 &  n9439 ;
  assign n9460 = n9444 &  n9459 ;
  assign n9461 = n9458 | n9460 ;
  assign n9473 = n9342 &  n9445 ;
  assign n9474 = n9444 &  n9473 ;
  assign n9462 = x106 | n9342 ;
  assign n9463 = x106 &  n9342 ;
  assign n9464 = ( n9462 & ~n9463 ) | ( n9462 & 1'b0 ) | ( ~n9463 & 1'b0 ) ;
  assign n9475 = n9430 &  n9464 ;
  assign n9476 = ( n9430 & ~n9446 ) | ( n9430 & n9464 ) | ( ~n9446 & n9464 ) ;
  assign n9477 = ( n9474 & ~n9475 ) | ( n9474 & n9476 ) | ( ~n9475 & n9476 ) ;
  assign n9481 = n9350 &  n9445 ;
  assign n9482 = n9444 &  n9481 ;
  assign n9470 = x105 | n9350 ;
  assign n9471 = x105 &  n9350 ;
  assign n9472 = ( n9470 & ~n9471 ) | ( n9470 & 1'b0 ) | ( ~n9471 & 1'b0 ) ;
  assign n9483 = n9429 &  n9472 ;
  assign n9484 = ( n9429 & ~n9446 ) | ( n9429 & n9472 ) | ( ~n9446 & n9472 ) ;
  assign n9485 = ( n9482 & ~n9483 ) | ( n9482 & n9484 ) | ( ~n9483 & n9484 ) ;
  assign n9489 = n9358 &  n9445 ;
  assign n9490 = n9444 &  n9489 ;
  assign n9478 = x104 | n9358 ;
  assign n9479 = x104 &  n9358 ;
  assign n9480 = ( n9478 & ~n9479 ) | ( n9478 & 1'b0 ) | ( ~n9479 & 1'b0 ) ;
  assign n9491 = n9428 &  n9480 ;
  assign n9492 = ( n9428 & ~n9446 ) | ( n9428 & n9480 ) | ( ~n9446 & n9480 ) ;
  assign n9493 = ( n9490 & ~n9491 ) | ( n9490 & n9492 ) | ( ~n9491 & n9492 ) ;
  assign n9497 = n9366 &  n9445 ;
  assign n9498 = n9444 &  n9497 ;
  assign n9486 = x103 | n9366 ;
  assign n9487 = x103 &  n9366 ;
  assign n9488 = ( n9486 & ~n9487 ) | ( n9486 & 1'b0 ) | ( ~n9487 & 1'b0 ) ;
  assign n9499 = n9427 &  n9488 ;
  assign n9500 = ( n9427 & ~n9446 ) | ( n9427 & n9488 ) | ( ~n9446 & n9488 ) ;
  assign n9501 = ( n9498 & ~n9499 ) | ( n9498 & n9500 ) | ( ~n9499 & n9500 ) ;
  assign n9505 = n9374 &  n9445 ;
  assign n9506 = n9444 &  n9505 ;
  assign n9494 = x102 | n9374 ;
  assign n9495 = x102 &  n9374 ;
  assign n9496 = ( n9494 & ~n9495 ) | ( n9494 & 1'b0 ) | ( ~n9495 & 1'b0 ) ;
  assign n9508 = ( n9426 & n9446 ) | ( n9426 & n9496 ) | ( n9446 & n9496 ) ;
  assign n9507 = n9426 | n9496 ;
  assign n9509 = ( n9506 & ~n9508 ) | ( n9506 & n9507 ) | ( ~n9508 & n9507 ) ;
  assign n9513 = n9382 &  n9445 ;
  assign n9514 = n9444 &  n9513 ;
  assign n9502 = x101 | n9382 ;
  assign n9503 = x101 &  n9382 ;
  assign n9504 = ( n9502 & ~n9503 ) | ( n9502 & 1'b0 ) | ( ~n9503 & 1'b0 ) ;
  assign n9516 = ( n9425 & n9446 ) | ( n9425 & n9504 ) | ( n9446 & n9504 ) ;
  assign n9515 = n9425 | n9504 ;
  assign n9517 = ( n9514 & ~n9516 ) | ( n9514 & n9515 ) | ( ~n9516 & n9515 ) ;
  assign n9521 = n9390 &  n9445 ;
  assign n9522 = n9444 &  n9521 ;
  assign n9510 = x100 | n9390 ;
  assign n9511 = x100 &  n9390 ;
  assign n9512 = ( n9510 & ~n9511 ) | ( n9510 & 1'b0 ) | ( ~n9511 & 1'b0 ) ;
  assign n9524 = ( n9424 & n9446 ) | ( n9424 & n9512 ) | ( n9446 & n9512 ) ;
  assign n9523 = n9424 | n9512 ;
  assign n9525 = ( n9522 & ~n9524 ) | ( n9522 & n9523 ) | ( ~n9524 & n9523 ) ;
  assign n9529 = n9398 &  n9445 ;
  assign n9530 = n9444 &  n9529 ;
  assign n9518 = x99 | n9398 ;
  assign n9519 = x99 &  n9398 ;
  assign n9520 = ( n9518 & ~n9519 ) | ( n9518 & 1'b0 ) | ( ~n9519 & 1'b0 ) ;
  assign n9532 = ( n9423 & n9446 ) | ( n9423 & n9520 ) | ( n9446 & n9520 ) ;
  assign n9531 = n9423 | n9520 ;
  assign n9533 = ( n9530 & ~n9532 ) | ( n9530 & n9531 ) | ( ~n9532 & n9531 ) ;
  assign n9537 = n9406 &  n9445 ;
  assign n9538 = n9444 &  n9537 ;
  assign n9526 = x98 | n9406 ;
  assign n9527 = x98 &  n9406 ;
  assign n9528 = ( n9526 & ~n9527 ) | ( n9526 & 1'b0 ) | ( ~n9527 & 1'b0 ) ;
  assign n9540 = ( n9422 & n9446 ) | ( n9422 & n9528 ) | ( n9446 & n9528 ) ;
  assign n9539 = n9422 | n9528 ;
  assign n9541 = ( n9538 & ~n9540 ) | ( n9538 & n9539 ) | ( ~n9540 & n9539 ) ;
  assign n9545 = n9414 &  n9445 ;
  assign n9546 = n9444 &  n9545 ;
  assign n9534 = x97 | n9414 ;
  assign n9535 = x97 &  n9414 ;
  assign n9536 = ( n9534 & ~n9535 ) | ( n9534 & 1'b0 ) | ( ~n9535 & 1'b0 ) ;
  assign n9548 = ( n9421 & n9446 ) | ( n9421 & n9536 ) | ( n9446 & n9536 ) ;
  assign n9547 = n9421 | n9536 ;
  assign n9549 = ( n9546 & ~n9548 ) | ( n9546 & n9547 ) | ( ~n9548 & n9547 ) ;
  assign n9550 = n9419 &  n9445 ;
  assign n9551 = n9444 &  n9550 ;
  assign n9542 = x96 | n9419 ;
  assign n9543 = x96 &  n9419 ;
  assign n9544 = ( n9542 & ~n9543 ) | ( n9542 & 1'b0 ) | ( ~n9543 & 1'b0 ) ;
  assign n9553 = ( n9420 & n9446 ) | ( n9420 & n9544 ) | ( n9446 & n9544 ) ;
  assign n9552 = n9420 | n9544 ;
  assign n9554 = ( n9551 & ~n9553 ) | ( n9551 & n9552 ) | ( ~n9553 & n9552 ) ;
  assign n9447 = n9320 &  n9445 ;
  assign n9448 = n9444 &  n9447 ;
  assign n9321 = x95 | n9320 ;
  assign n9322 = x95 &  n9320 ;
  assign n9323 = ( n9321 & ~n9322 ) | ( n9321 & 1'b0 ) | ( ~n9322 & 1'b0 ) ;
  assign n9450 = ( n9312 & n9323 ) | ( n9312 & n9446 ) | ( n9323 & n9446 ) ;
  assign n9449 = n9312 | n9323 ;
  assign n9451 = ( n9448 & ~n9450 ) | ( n9448 & n9449 ) | ( ~n9450 & n9449 ) ;
  assign n9558 = n9055 &  n9445 ;
  assign n9559 = n9444 &  n9558 ;
  assign n9309 = x94 | n9055 ;
  assign n9310 = x94 &  n9055 ;
  assign n9311 = ( n9309 & ~n9310 ) | ( n9309 & 1'b0 ) | ( ~n9310 & 1'b0 ) ;
  assign n9560 = n9308 &  n9311 ;
  assign n9561 = ( n9308 & ~n9446 ) | ( n9308 & n9311 ) | ( ~n9446 & n9311 ) ;
  assign n9562 = ( n9559 & ~n9560 ) | ( n9559 & n9561 ) | ( ~n9560 & n9561 ) ;
  assign n9566 = n9063 &  n9445 ;
  assign n9567 = n9444 &  n9566 ;
  assign n9555 = x93 | n9063 ;
  assign n9556 = x93 &  n9063 ;
  assign n9557 = ( n9555 & ~n9556 ) | ( n9555 & 1'b0 ) | ( ~n9556 & 1'b0 ) ;
  assign n9569 = ( n9307 & n9446 ) | ( n9307 & n9557 ) | ( n9446 & n9557 ) ;
  assign n9568 = n9307 | n9557 ;
  assign n9570 = ( n9567 & ~n9569 ) | ( n9567 & n9568 ) | ( ~n9569 & n9568 ) ;
  assign n9574 = n9071 &  n9445 ;
  assign n9575 = n9444 &  n9574 ;
  assign n9563 = x92 | n9071 ;
  assign n9564 = x92 &  n9071 ;
  assign n9565 = ( n9563 & ~n9564 ) | ( n9563 & 1'b0 ) | ( ~n9564 & 1'b0 ) ;
  assign n9577 = ( n9306 & n9446 ) | ( n9306 & n9565 ) | ( n9446 & n9565 ) ;
  assign n9576 = n9306 | n9565 ;
  assign n9578 = ( n9575 & ~n9577 ) | ( n9575 & n9576 ) | ( ~n9577 & n9576 ) ;
  assign n9582 = n9079 &  n9445 ;
  assign n9583 = n9444 &  n9582 ;
  assign n9571 = x91 | n9079 ;
  assign n9572 = x91 &  n9079 ;
  assign n9573 = ( n9571 & ~n9572 ) | ( n9571 & 1'b0 ) | ( ~n9572 & 1'b0 ) ;
  assign n9585 = ( n9305 & n9446 ) | ( n9305 & n9573 ) | ( n9446 & n9573 ) ;
  assign n9584 = n9305 | n9573 ;
  assign n9586 = ( n9583 & ~n9585 ) | ( n9583 & n9584 ) | ( ~n9585 & n9584 ) ;
  assign n9590 = n9087 &  n9445 ;
  assign n9591 = n9444 &  n9590 ;
  assign n9579 = x90 | n9087 ;
  assign n9580 = x90 &  n9087 ;
  assign n9581 = ( n9579 & ~n9580 ) | ( n9579 & 1'b0 ) | ( ~n9580 & 1'b0 ) ;
  assign n9593 = ( n9304 & n9446 ) | ( n9304 & n9581 ) | ( n9446 & n9581 ) ;
  assign n9592 = n9304 | n9581 ;
  assign n9594 = ( n9591 & ~n9593 ) | ( n9591 & n9592 ) | ( ~n9593 & n9592 ) ;
  assign n9598 = n9095 &  n9445 ;
  assign n9599 = n9444 &  n9598 ;
  assign n9587 = x89 | n9095 ;
  assign n9588 = x89 &  n9095 ;
  assign n9589 = ( n9587 & ~n9588 ) | ( n9587 & 1'b0 ) | ( ~n9588 & 1'b0 ) ;
  assign n9601 = ( n9303 & n9446 ) | ( n9303 & n9589 ) | ( n9446 & n9589 ) ;
  assign n9600 = n9303 | n9589 ;
  assign n9602 = ( n9599 & ~n9601 ) | ( n9599 & n9600 ) | ( ~n9601 & n9600 ) ;
  assign n9606 = n9103 &  n9445 ;
  assign n9607 = n9444 &  n9606 ;
  assign n9595 = x88 | n9103 ;
  assign n9596 = x88 &  n9103 ;
  assign n9597 = ( n9595 & ~n9596 ) | ( n9595 & 1'b0 ) | ( ~n9596 & 1'b0 ) ;
  assign n9609 = ( n9302 & n9446 ) | ( n9302 & n9597 ) | ( n9446 & n9597 ) ;
  assign n9608 = n9302 | n9597 ;
  assign n9610 = ( n9607 & ~n9609 ) | ( n9607 & n9608 ) | ( ~n9609 & n9608 ) ;
  assign n9614 = n9111 &  n9445 ;
  assign n9615 = n9444 &  n9614 ;
  assign n9603 = x87 | n9111 ;
  assign n9604 = x87 &  n9111 ;
  assign n9605 = ( n9603 & ~n9604 ) | ( n9603 & 1'b0 ) | ( ~n9604 & 1'b0 ) ;
  assign n9617 = ( n9301 & n9446 ) | ( n9301 & n9605 ) | ( n9446 & n9605 ) ;
  assign n9616 = n9301 | n9605 ;
  assign n9618 = ( n9615 & ~n9617 ) | ( n9615 & n9616 ) | ( ~n9617 & n9616 ) ;
  assign n9622 = n9119 &  n9445 ;
  assign n9623 = n9444 &  n9622 ;
  assign n9611 = x86 | n9119 ;
  assign n9612 = x86 &  n9119 ;
  assign n9613 = ( n9611 & ~n9612 ) | ( n9611 & 1'b0 ) | ( ~n9612 & 1'b0 ) ;
  assign n9625 = ( n9300 & n9446 ) | ( n9300 & n9613 ) | ( n9446 & n9613 ) ;
  assign n9624 = n9300 | n9613 ;
  assign n9626 = ( n9623 & ~n9625 ) | ( n9623 & n9624 ) | ( ~n9625 & n9624 ) ;
  assign n9630 = n9127 &  n9445 ;
  assign n9631 = n9444 &  n9630 ;
  assign n9619 = x85 | n9127 ;
  assign n9620 = x85 &  n9127 ;
  assign n9621 = ( n9619 & ~n9620 ) | ( n9619 & 1'b0 ) | ( ~n9620 & 1'b0 ) ;
  assign n9633 = ( n9299 & n9446 ) | ( n9299 & n9621 ) | ( n9446 & n9621 ) ;
  assign n9632 = n9299 | n9621 ;
  assign n9634 = ( n9631 & ~n9633 ) | ( n9631 & n9632 ) | ( ~n9633 & n9632 ) ;
  assign n9638 = n9135 &  n9445 ;
  assign n9639 = n9444 &  n9638 ;
  assign n9627 = x84 | n9135 ;
  assign n9628 = x84 &  n9135 ;
  assign n9629 = ( n9627 & ~n9628 ) | ( n9627 & 1'b0 ) | ( ~n9628 & 1'b0 ) ;
  assign n9641 = ( n9298 & n9446 ) | ( n9298 & n9629 ) | ( n9446 & n9629 ) ;
  assign n9640 = n9298 | n9629 ;
  assign n9642 = ( n9639 & ~n9641 ) | ( n9639 & n9640 ) | ( ~n9641 & n9640 ) ;
  assign n9646 = n9143 &  n9445 ;
  assign n9647 = n9444 &  n9646 ;
  assign n9635 = x83 | n9143 ;
  assign n9636 = x83 &  n9143 ;
  assign n9637 = ( n9635 & ~n9636 ) | ( n9635 & 1'b0 ) | ( ~n9636 & 1'b0 ) ;
  assign n9649 = ( n9297 & n9446 ) | ( n9297 & n9637 ) | ( n9446 & n9637 ) ;
  assign n9648 = n9297 | n9637 ;
  assign n9650 = ( n9647 & ~n9649 ) | ( n9647 & n9648 ) | ( ~n9649 & n9648 ) ;
  assign n9654 = n9151 &  n9445 ;
  assign n9655 = n9444 &  n9654 ;
  assign n9643 = x82 | n9151 ;
  assign n9644 = x82 &  n9151 ;
  assign n9645 = ( n9643 & ~n9644 ) | ( n9643 & 1'b0 ) | ( ~n9644 & 1'b0 ) ;
  assign n9657 = ( n9296 & n9446 ) | ( n9296 & n9645 ) | ( n9446 & n9645 ) ;
  assign n9656 = n9296 | n9645 ;
  assign n9658 = ( n9655 & ~n9657 ) | ( n9655 & n9656 ) | ( ~n9657 & n9656 ) ;
  assign n9662 = n9159 &  n9445 ;
  assign n9663 = n9444 &  n9662 ;
  assign n9651 = x81 | n9159 ;
  assign n9652 = x81 &  n9159 ;
  assign n9653 = ( n9651 & ~n9652 ) | ( n9651 & 1'b0 ) | ( ~n9652 & 1'b0 ) ;
  assign n9665 = ( n9295 & n9446 ) | ( n9295 & n9653 ) | ( n9446 & n9653 ) ;
  assign n9664 = n9295 | n9653 ;
  assign n9666 = ( n9663 & ~n9665 ) | ( n9663 & n9664 ) | ( ~n9665 & n9664 ) ;
  assign n9670 = n9167 &  n9445 ;
  assign n9671 = n9444 &  n9670 ;
  assign n9659 = x80 | n9167 ;
  assign n9660 = x80 &  n9167 ;
  assign n9661 = ( n9659 & ~n9660 ) | ( n9659 & 1'b0 ) | ( ~n9660 & 1'b0 ) ;
  assign n9673 = ( n9294 & n9446 ) | ( n9294 & n9661 ) | ( n9446 & n9661 ) ;
  assign n9672 = n9294 | n9661 ;
  assign n9674 = ( n9671 & ~n9673 ) | ( n9671 & n9672 ) | ( ~n9673 & n9672 ) ;
  assign n9678 = n9175 &  n9445 ;
  assign n9679 = n9444 &  n9678 ;
  assign n9667 = x79 | n9175 ;
  assign n9668 = x79 &  n9175 ;
  assign n9669 = ( n9667 & ~n9668 ) | ( n9667 & 1'b0 ) | ( ~n9668 & 1'b0 ) ;
  assign n9681 = ( n9293 & n9446 ) | ( n9293 & n9669 ) | ( n9446 & n9669 ) ;
  assign n9680 = n9293 | n9669 ;
  assign n9682 = ( n9679 & ~n9681 ) | ( n9679 & n9680 ) | ( ~n9681 & n9680 ) ;
  assign n9686 = n9183 &  n9445 ;
  assign n9687 = n9444 &  n9686 ;
  assign n9675 = x78 | n9183 ;
  assign n9676 = x78 &  n9183 ;
  assign n9677 = ( n9675 & ~n9676 ) | ( n9675 & 1'b0 ) | ( ~n9676 & 1'b0 ) ;
  assign n9689 = ( n9292 & n9446 ) | ( n9292 & n9677 ) | ( n9446 & n9677 ) ;
  assign n9688 = n9292 | n9677 ;
  assign n9690 = ( n9687 & ~n9689 ) | ( n9687 & n9688 ) | ( ~n9689 & n9688 ) ;
  assign n9694 = n9191 &  n9445 ;
  assign n9695 = n9444 &  n9694 ;
  assign n9683 = x77 | n9191 ;
  assign n9684 = x77 &  n9191 ;
  assign n9685 = ( n9683 & ~n9684 ) | ( n9683 & 1'b0 ) | ( ~n9684 & 1'b0 ) ;
  assign n9697 = ( n9291 & n9446 ) | ( n9291 & n9685 ) | ( n9446 & n9685 ) ;
  assign n9696 = n9291 | n9685 ;
  assign n9698 = ( n9695 & ~n9697 ) | ( n9695 & n9696 ) | ( ~n9697 & n9696 ) ;
  assign n9702 = n9199 &  n9445 ;
  assign n9703 = n9444 &  n9702 ;
  assign n9691 = x76 | n9199 ;
  assign n9692 = x76 &  n9199 ;
  assign n9693 = ( n9691 & ~n9692 ) | ( n9691 & 1'b0 ) | ( ~n9692 & 1'b0 ) ;
  assign n9705 = ( n9290 & n9446 ) | ( n9290 & n9693 ) | ( n9446 & n9693 ) ;
  assign n9704 = n9290 | n9693 ;
  assign n9706 = ( n9703 & ~n9705 ) | ( n9703 & n9704 ) | ( ~n9705 & n9704 ) ;
  assign n9710 = n9207 &  n9445 ;
  assign n9711 = n9444 &  n9710 ;
  assign n9699 = x75 | n9207 ;
  assign n9700 = x75 &  n9207 ;
  assign n9701 = ( n9699 & ~n9700 ) | ( n9699 & 1'b0 ) | ( ~n9700 & 1'b0 ) ;
  assign n9713 = ( n9289 & n9446 ) | ( n9289 & n9701 ) | ( n9446 & n9701 ) ;
  assign n9712 = n9289 | n9701 ;
  assign n9714 = ( n9711 & ~n9713 ) | ( n9711 & n9712 ) | ( ~n9713 & n9712 ) ;
  assign n9718 = n9215 &  n9445 ;
  assign n9719 = n9444 &  n9718 ;
  assign n9707 = x74 | n9215 ;
  assign n9708 = x74 &  n9215 ;
  assign n9709 = ( n9707 & ~n9708 ) | ( n9707 & 1'b0 ) | ( ~n9708 & 1'b0 ) ;
  assign n9721 = ( n9288 & n9446 ) | ( n9288 & n9709 ) | ( n9446 & n9709 ) ;
  assign n9720 = n9288 | n9709 ;
  assign n9722 = ( n9719 & ~n9721 ) | ( n9719 & n9720 ) | ( ~n9721 & n9720 ) ;
  assign n9726 = n9223 &  n9445 ;
  assign n9727 = n9444 &  n9726 ;
  assign n9715 = x73 | n9223 ;
  assign n9716 = x73 &  n9223 ;
  assign n9717 = ( n9715 & ~n9716 ) | ( n9715 & 1'b0 ) | ( ~n9716 & 1'b0 ) ;
  assign n9729 = ( n9287 & n9446 ) | ( n9287 & n9717 ) | ( n9446 & n9717 ) ;
  assign n9728 = n9287 | n9717 ;
  assign n9730 = ( n9727 & ~n9729 ) | ( n9727 & n9728 ) | ( ~n9729 & n9728 ) ;
  assign n9734 = n9231 &  n9445 ;
  assign n9735 = n9444 &  n9734 ;
  assign n9723 = x72 | n9231 ;
  assign n9724 = x72 &  n9231 ;
  assign n9725 = ( n9723 & ~n9724 ) | ( n9723 & 1'b0 ) | ( ~n9724 & 1'b0 ) ;
  assign n9737 = ( n9286 & n9446 ) | ( n9286 & n9725 ) | ( n9446 & n9725 ) ;
  assign n9736 = n9286 | n9725 ;
  assign n9738 = ( n9735 & ~n9737 ) | ( n9735 & n9736 ) | ( ~n9737 & n9736 ) ;
  assign n9742 = n9239 &  n9445 ;
  assign n9743 = n9444 &  n9742 ;
  assign n9731 = x71 | n9239 ;
  assign n9732 = x71 &  n9239 ;
  assign n9733 = ( n9731 & ~n9732 ) | ( n9731 & 1'b0 ) | ( ~n9732 & 1'b0 ) ;
  assign n9745 = ( n9285 & n9446 ) | ( n9285 & n9733 ) | ( n9446 & n9733 ) ;
  assign n9744 = n9285 | n9733 ;
  assign n9746 = ( n9743 & ~n9745 ) | ( n9743 & n9744 ) | ( ~n9745 & n9744 ) ;
  assign n9750 = n9247 &  n9445 ;
  assign n9751 = n9444 &  n9750 ;
  assign n9739 = x70 | n9247 ;
  assign n9740 = x70 &  n9247 ;
  assign n9741 = ( n9739 & ~n9740 ) | ( n9739 & 1'b0 ) | ( ~n9740 & 1'b0 ) ;
  assign n9753 = ( n9284 & n9446 ) | ( n9284 & n9741 ) | ( n9446 & n9741 ) ;
  assign n9752 = n9284 | n9741 ;
  assign n9754 = ( n9751 & ~n9753 ) | ( n9751 & n9752 ) | ( ~n9753 & n9752 ) ;
  assign n9758 = n9255 &  n9445 ;
  assign n9759 = n9444 &  n9758 ;
  assign n9747 = x69 | n9255 ;
  assign n9748 = x69 &  n9255 ;
  assign n9749 = ( n9747 & ~n9748 ) | ( n9747 & 1'b0 ) | ( ~n9748 & 1'b0 ) ;
  assign n9761 = ( n9283 & n9446 ) | ( n9283 & n9749 ) | ( n9446 & n9749 ) ;
  assign n9760 = n9283 | n9749 ;
  assign n9762 = ( n9759 & ~n9761 ) | ( n9759 & n9760 ) | ( ~n9761 & n9760 ) ;
  assign n9766 = n9263 &  n9445 ;
  assign n9767 = n9444 &  n9766 ;
  assign n9755 = x68 | n9263 ;
  assign n9756 = x68 &  n9263 ;
  assign n9757 = ( n9755 & ~n9756 ) | ( n9755 & 1'b0 ) | ( ~n9756 & 1'b0 ) ;
  assign n9769 = ( n9282 & n9446 ) | ( n9282 & n9757 ) | ( n9446 & n9757 ) ;
  assign n9768 = n9282 | n9757 ;
  assign n9770 = ( n9767 & ~n9769 ) | ( n9767 & n9768 ) | ( ~n9769 & n9768 ) ;
  assign n9774 = n9268 &  n9445 ;
  assign n9775 = n9444 &  n9774 ;
  assign n9763 = x67 | n9268 ;
  assign n9764 = x67 &  n9268 ;
  assign n9765 = ( n9763 & ~n9764 ) | ( n9763 & 1'b0 ) | ( ~n9764 & 1'b0 ) ;
  assign n9777 = ( n9281 & n9446 ) | ( n9281 & n9765 ) | ( n9446 & n9765 ) ;
  assign n9776 = n9281 | n9765 ;
  assign n9778 = ( n9775 & ~n9777 ) | ( n9775 & n9776 ) | ( ~n9777 & n9776 ) ;
  assign n9779 = n9274 &  n9445 ;
  assign n9780 = n9444 &  n9779 ;
  assign n9771 = x66 | n9274 ;
  assign n9772 = x66 &  n9274 ;
  assign n9773 = ( n9771 & ~n9772 ) | ( n9771 & 1'b0 ) | ( ~n9772 & 1'b0 ) ;
  assign n9781 = n9280 &  n9773 ;
  assign n9782 = ( n9280 & ~n9446 ) | ( n9280 & n9773 ) | ( ~n9446 & n9773 ) ;
  assign n9783 = ( n9780 & ~n9781 ) | ( n9780 & n9782 ) | ( ~n9781 & n9782 ) ;
  assign n9784 = ( n9278 & ~x65 ) | ( n9278 & n9279 ) | ( ~x65 & n9279 ) ;
  assign n9785 = ( n9280 & ~n9279 ) | ( n9280 & n9784 ) | ( ~n9279 & n9784 ) ;
  assign n9786 = ~n9446 & n9785 ;
  assign n9787 = n9278 &  n9445 ;
  assign n9788 = n9444 &  n9787 ;
  assign n9789 = n9786 | n9788 ;
  assign n9790 = ( x64 & ~n9446 ) | ( x64 & 1'b0 ) | ( ~n9446 & 1'b0 ) ;
  assign n9791 = ( x19 & ~n9790 ) | ( x19 & 1'b0 ) | ( ~n9790 & 1'b0 ) ;
  assign n9792 = ( n9279 & ~n9446 ) | ( n9279 & 1'b0 ) | ( ~n9446 & 1'b0 ) ;
  assign n9793 = n9791 | n9792 ;
  assign n9794 = ~x18 & x64 ;
  assign n9795 = ( x65 & ~n9793 ) | ( x65 & n9794 ) | ( ~n9793 & n9794 ) ;
  assign n9796 = ( x66 & ~n9789 ) | ( x66 & n9795 ) | ( ~n9789 & n9795 ) ;
  assign n9797 = ( x67 & ~n9783 ) | ( x67 & n9796 ) | ( ~n9783 & n9796 ) ;
  assign n9798 = ( x68 & ~n9778 ) | ( x68 & n9797 ) | ( ~n9778 & n9797 ) ;
  assign n9799 = ( x69 & ~n9770 ) | ( x69 & n9798 ) | ( ~n9770 & n9798 ) ;
  assign n9800 = ( x70 & ~n9762 ) | ( x70 & n9799 ) | ( ~n9762 & n9799 ) ;
  assign n9801 = ( x71 & ~n9754 ) | ( x71 & n9800 ) | ( ~n9754 & n9800 ) ;
  assign n9802 = ( x72 & ~n9746 ) | ( x72 & n9801 ) | ( ~n9746 & n9801 ) ;
  assign n9803 = ( x73 & ~n9738 ) | ( x73 & n9802 ) | ( ~n9738 & n9802 ) ;
  assign n9804 = ( x74 & ~n9730 ) | ( x74 & n9803 ) | ( ~n9730 & n9803 ) ;
  assign n9805 = ( x75 & ~n9722 ) | ( x75 & n9804 ) | ( ~n9722 & n9804 ) ;
  assign n9806 = ( x76 & ~n9714 ) | ( x76 & n9805 ) | ( ~n9714 & n9805 ) ;
  assign n9807 = ( x77 & ~n9706 ) | ( x77 & n9806 ) | ( ~n9706 & n9806 ) ;
  assign n9808 = ( x78 & ~n9698 ) | ( x78 & n9807 ) | ( ~n9698 & n9807 ) ;
  assign n9809 = ( x79 & ~n9690 ) | ( x79 & n9808 ) | ( ~n9690 & n9808 ) ;
  assign n9810 = ( x80 & ~n9682 ) | ( x80 & n9809 ) | ( ~n9682 & n9809 ) ;
  assign n9811 = ( x81 & ~n9674 ) | ( x81 & n9810 ) | ( ~n9674 & n9810 ) ;
  assign n9812 = ( x82 & ~n9666 ) | ( x82 & n9811 ) | ( ~n9666 & n9811 ) ;
  assign n9813 = ( x83 & ~n9658 ) | ( x83 & n9812 ) | ( ~n9658 & n9812 ) ;
  assign n9814 = ( x84 & ~n9650 ) | ( x84 & n9813 ) | ( ~n9650 & n9813 ) ;
  assign n9815 = ( x85 & ~n9642 ) | ( x85 & n9814 ) | ( ~n9642 & n9814 ) ;
  assign n9816 = ( x86 & ~n9634 ) | ( x86 & n9815 ) | ( ~n9634 & n9815 ) ;
  assign n9817 = ( x87 & ~n9626 ) | ( x87 & n9816 ) | ( ~n9626 & n9816 ) ;
  assign n9818 = ( x88 & ~n9618 ) | ( x88 & n9817 ) | ( ~n9618 & n9817 ) ;
  assign n9819 = ( x89 & ~n9610 ) | ( x89 & n9818 ) | ( ~n9610 & n9818 ) ;
  assign n9820 = ( x90 & ~n9602 ) | ( x90 & n9819 ) | ( ~n9602 & n9819 ) ;
  assign n9821 = ( x91 & ~n9594 ) | ( x91 & n9820 ) | ( ~n9594 & n9820 ) ;
  assign n9822 = ( x92 & ~n9586 ) | ( x92 & n9821 ) | ( ~n9586 & n9821 ) ;
  assign n9823 = ( x93 & ~n9578 ) | ( x93 & n9822 ) | ( ~n9578 & n9822 ) ;
  assign n9824 = ( x94 & ~n9570 ) | ( x94 & n9823 ) | ( ~n9570 & n9823 ) ;
  assign n9825 = ( x95 & ~n9562 ) | ( x95 & n9824 ) | ( ~n9562 & n9824 ) ;
  assign n9826 = ( x96 & ~n9451 ) | ( x96 & n9825 ) | ( ~n9451 & n9825 ) ;
  assign n9827 = ( x97 & ~n9554 ) | ( x97 & n9826 ) | ( ~n9554 & n9826 ) ;
  assign n9828 = ( x98 & ~n9549 ) | ( x98 & n9827 ) | ( ~n9549 & n9827 ) ;
  assign n9829 = ( x99 & ~n9541 ) | ( x99 & n9828 ) | ( ~n9541 & n9828 ) ;
  assign n9830 = ( x100 & ~n9533 ) | ( x100 & n9829 ) | ( ~n9533 & n9829 ) ;
  assign n9831 = ( x101 & ~n9525 ) | ( x101 & n9830 ) | ( ~n9525 & n9830 ) ;
  assign n9832 = ( x102 & ~n9517 ) | ( x102 & n9831 ) | ( ~n9517 & n9831 ) ;
  assign n9833 = ( x103 & ~n9509 ) | ( x103 & n9832 ) | ( ~n9509 & n9832 ) ;
  assign n9834 = ( x104 & ~n9501 ) | ( x104 & n9833 ) | ( ~n9501 & n9833 ) ;
  assign n9835 = ( x105 & ~n9493 ) | ( x105 & n9834 ) | ( ~n9493 & n9834 ) ;
  assign n9836 = ( x106 & ~n9485 ) | ( x106 & n9835 ) | ( ~n9485 & n9835 ) ;
  assign n9837 = ( x107 & ~n9477 ) | ( x107 & n9836 ) | ( ~n9477 & n9836 ) ;
  assign n9838 = ( x108 & ~n9469 ) | ( x108 & n9837 ) | ( ~n9469 & n9837 ) ;
  assign n9839 = ( x109 & ~n9461 ) | ( x109 & n9838 ) | ( ~n9461 & n9838 ) ;
  assign n9840 = n170 | n172 ;
  assign n9841 = n160 | n9840 ;
  assign n9842 = n9839 | n9841 ;
  assign n10160 = n9469 &  n9842 ;
  assign n10164 = x108 | n9469 ;
  assign n10165 = x108 &  n9469 ;
  assign n10166 = ( n10164 & ~n10165 ) | ( n10164 & 1'b0 ) | ( ~n10165 & 1'b0 ) ;
  assign n10167 = ( n9837 & n9839 ) | ( n9837 & n10166 ) | ( n9839 & n10166 ) ;
  assign n10168 = ( n9837 & ~n9841 ) | ( n9837 & n10166 ) | ( ~n9841 & n10166 ) ;
  assign n10169 = ~n10167 & n10168 ;
  assign n10170 = n10160 | n10169 ;
  assign n10171 = n9477 &  n9842 ;
  assign n10161 = x107 | n9477 ;
  assign n10162 = x107 &  n9477 ;
  assign n10163 = ( n10161 & ~n10162 ) | ( n10161 & 1'b0 ) | ( ~n10162 & 1'b0 ) ;
  assign n10175 = ( n9836 & n9839 ) | ( n9836 & n10163 ) | ( n9839 & n10163 ) ;
  assign n10176 = ( n9836 & ~n9841 ) | ( n9836 & n10163 ) | ( ~n9841 & n10163 ) ;
  assign n10177 = ~n10175 & n10176 ;
  assign n10178 = n10171 | n10177 ;
  assign n10179 = n9485 &  n9842 ;
  assign n10172 = x106 | n9485 ;
  assign n10173 = x106 &  n9485 ;
  assign n10174 = ( n10172 & ~n10173 ) | ( n10172 & 1'b0 ) | ( ~n10173 & 1'b0 ) ;
  assign n10183 = ( n9835 & n9839 ) | ( n9835 & n10174 ) | ( n9839 & n10174 ) ;
  assign n10184 = ( n9835 & ~n9841 ) | ( n9835 & n10174 ) | ( ~n9841 & n10174 ) ;
  assign n10185 = ~n10183 & n10184 ;
  assign n10186 = n10179 | n10185 ;
  assign n10187 = n9493 &  n9842 ;
  assign n10180 = x105 | n9493 ;
  assign n10181 = x105 &  n9493 ;
  assign n10182 = ( n10180 & ~n10181 ) | ( n10180 & 1'b0 ) | ( ~n10181 & 1'b0 ) ;
  assign n10191 = ( n9834 & n9839 ) | ( n9834 & n10182 ) | ( n9839 & n10182 ) ;
  assign n10192 = ( n9834 & ~n9841 ) | ( n9834 & n10182 ) | ( ~n9841 & n10182 ) ;
  assign n10193 = ~n10191 & n10192 ;
  assign n10194 = n10187 | n10193 ;
  assign n10195 = n9501 &  n9842 ;
  assign n10188 = x104 | n9501 ;
  assign n10189 = x104 &  n9501 ;
  assign n10190 = ( n10188 & ~n10189 ) | ( n10188 & 1'b0 ) | ( ~n10189 & 1'b0 ) ;
  assign n10199 = ( n9833 & n9839 ) | ( n9833 & n10190 ) | ( n9839 & n10190 ) ;
  assign n10200 = ( n9833 & ~n9841 ) | ( n9833 & n10190 ) | ( ~n9841 & n10190 ) ;
  assign n10201 = ~n10199 & n10200 ;
  assign n10202 = n10195 | n10201 ;
  assign n10203 = n9509 &  n9842 ;
  assign n10196 = x103 | n9509 ;
  assign n10197 = x103 &  n9509 ;
  assign n10198 = ( n10196 & ~n10197 ) | ( n10196 & 1'b0 ) | ( ~n10197 & 1'b0 ) ;
  assign n10207 = ( n9832 & n9839 ) | ( n9832 & n10198 ) | ( n9839 & n10198 ) ;
  assign n10208 = ( n9832 & ~n9841 ) | ( n9832 & n10198 ) | ( ~n9841 & n10198 ) ;
  assign n10209 = ~n10207 & n10208 ;
  assign n10210 = n10203 | n10209 ;
  assign n10211 = n9517 &  n9842 ;
  assign n10204 = x102 | n9517 ;
  assign n10205 = x102 &  n9517 ;
  assign n10206 = ( n10204 & ~n10205 ) | ( n10204 & 1'b0 ) | ( ~n10205 & 1'b0 ) ;
  assign n10215 = ( n9831 & n9839 ) | ( n9831 & n10206 ) | ( n9839 & n10206 ) ;
  assign n10216 = ( n9831 & ~n9841 ) | ( n9831 & n10206 ) | ( ~n9841 & n10206 ) ;
  assign n10217 = ~n10215 & n10216 ;
  assign n10218 = n10211 | n10217 ;
  assign n10219 = n9525 &  n9842 ;
  assign n10212 = x101 | n9525 ;
  assign n10213 = x101 &  n9525 ;
  assign n10214 = ( n10212 & ~n10213 ) | ( n10212 & 1'b0 ) | ( ~n10213 & 1'b0 ) ;
  assign n10223 = ( n9830 & n9839 ) | ( n9830 & n10214 ) | ( n9839 & n10214 ) ;
  assign n10224 = ( n9830 & ~n9841 ) | ( n9830 & n10214 ) | ( ~n9841 & n10214 ) ;
  assign n10225 = ~n10223 & n10224 ;
  assign n10226 = n10219 | n10225 ;
  assign n10227 = n9533 &  n9842 ;
  assign n10220 = x100 | n9533 ;
  assign n10221 = x100 &  n9533 ;
  assign n10222 = ( n10220 & ~n10221 ) | ( n10220 & 1'b0 ) | ( ~n10221 & 1'b0 ) ;
  assign n10231 = ( n9829 & n9839 ) | ( n9829 & n10222 ) | ( n9839 & n10222 ) ;
  assign n10232 = ( n9829 & ~n9841 ) | ( n9829 & n10222 ) | ( ~n9841 & n10222 ) ;
  assign n10233 = ~n10231 & n10232 ;
  assign n10234 = n10227 | n10233 ;
  assign n10235 = n9541 &  n9842 ;
  assign n10228 = x99 | n9541 ;
  assign n10229 = x99 &  n9541 ;
  assign n10230 = ( n10228 & ~n10229 ) | ( n10228 & 1'b0 ) | ( ~n10229 & 1'b0 ) ;
  assign n10239 = ( n9828 & n9839 ) | ( n9828 & n10230 ) | ( n9839 & n10230 ) ;
  assign n10240 = ( n9828 & ~n9841 ) | ( n9828 & n10230 ) | ( ~n9841 & n10230 ) ;
  assign n10241 = ~n10239 & n10240 ;
  assign n10242 = n10235 | n10241 ;
  assign n10243 = n9549 &  n9842 ;
  assign n10236 = x98 | n9549 ;
  assign n10237 = x98 &  n9549 ;
  assign n10238 = ( n10236 & ~n10237 ) | ( n10236 & 1'b0 ) | ( ~n10237 & 1'b0 ) ;
  assign n10244 = ( n9827 & n9839 ) | ( n9827 & n10238 ) | ( n9839 & n10238 ) ;
  assign n10245 = ( n9827 & ~n9841 ) | ( n9827 & n10238 ) | ( ~n9841 & n10238 ) ;
  assign n10246 = ~n10244 & n10245 ;
  assign n10247 = n10243 | n10246 ;
  assign n10149 = n9554 &  n9842 ;
  assign n10150 = x97 | n9554 ;
  assign n10151 = x97 &  n9554 ;
  assign n10152 = ( n10150 & ~n10151 ) | ( n10150 & 1'b0 ) | ( ~n10151 & 1'b0 ) ;
  assign n10153 = ( n9826 & n9839 ) | ( n9826 & n10152 ) | ( n9839 & n10152 ) ;
  assign n10154 = ( n9826 & ~n9841 ) | ( n9826 & n10152 ) | ( ~n9841 & n10152 ) ;
  assign n10155 = ~n10153 & n10154 ;
  assign n10156 = n10149 | n10155 ;
  assign n9843 = n9451 &  n9842 ;
  assign n9847 = x96 | n9451 ;
  assign n9848 = x96 &  n9451 ;
  assign n9849 = ( n9847 & ~n9848 ) | ( n9847 & 1'b0 ) | ( ~n9848 & 1'b0 ) ;
  assign n9850 = ( n9825 & n9839 ) | ( n9825 & n9849 ) | ( n9839 & n9849 ) ;
  assign n9851 = ( n9825 & ~n9841 ) | ( n9825 & n9849 ) | ( ~n9841 & n9849 ) ;
  assign n9852 = ~n9850 & n9851 ;
  assign n9853 = n9843 | n9852 ;
  assign n9854 = n9562 &  n9842 ;
  assign n9844 = x95 | n9562 ;
  assign n9845 = x95 &  n9562 ;
  assign n9846 = ( n9844 & ~n9845 ) | ( n9844 & 1'b0 ) | ( ~n9845 & 1'b0 ) ;
  assign n9858 = ( n9824 & n9839 ) | ( n9824 & n9846 ) | ( n9839 & n9846 ) ;
  assign n9859 = ( n9824 & ~n9841 ) | ( n9824 & n9846 ) | ( ~n9841 & n9846 ) ;
  assign n9860 = ~n9858 & n9859 ;
  assign n9861 = n9854 | n9860 ;
  assign n9862 = n9570 &  n9842 ;
  assign n9855 = x94 | n9570 ;
  assign n9856 = x94 &  n9570 ;
  assign n9857 = ( n9855 & ~n9856 ) | ( n9855 & 1'b0 ) | ( ~n9856 & 1'b0 ) ;
  assign n9866 = ( n9823 & n9839 ) | ( n9823 & n9857 ) | ( n9839 & n9857 ) ;
  assign n9867 = ( n9823 & ~n9841 ) | ( n9823 & n9857 ) | ( ~n9841 & n9857 ) ;
  assign n9868 = ~n9866 & n9867 ;
  assign n9869 = n9862 | n9868 ;
  assign n9870 = n9578 &  n9842 ;
  assign n9863 = x93 | n9578 ;
  assign n9864 = x93 &  n9578 ;
  assign n9865 = ( n9863 & ~n9864 ) | ( n9863 & 1'b0 ) | ( ~n9864 & 1'b0 ) ;
  assign n9874 = ( n9822 & n9839 ) | ( n9822 & n9865 ) | ( n9839 & n9865 ) ;
  assign n9875 = ( n9822 & ~n9841 ) | ( n9822 & n9865 ) | ( ~n9841 & n9865 ) ;
  assign n9876 = ~n9874 & n9875 ;
  assign n9877 = n9870 | n9876 ;
  assign n9878 = n9586 &  n9842 ;
  assign n9871 = x92 | n9586 ;
  assign n9872 = x92 &  n9586 ;
  assign n9873 = ( n9871 & ~n9872 ) | ( n9871 & 1'b0 ) | ( ~n9872 & 1'b0 ) ;
  assign n9882 = ( n9821 & n9839 ) | ( n9821 & n9873 ) | ( n9839 & n9873 ) ;
  assign n9883 = ( n9821 & ~n9841 ) | ( n9821 & n9873 ) | ( ~n9841 & n9873 ) ;
  assign n9884 = ~n9882 & n9883 ;
  assign n9885 = n9878 | n9884 ;
  assign n9886 = n9594 &  n9842 ;
  assign n9879 = x91 | n9594 ;
  assign n9880 = x91 &  n9594 ;
  assign n9881 = ( n9879 & ~n9880 ) | ( n9879 & 1'b0 ) | ( ~n9880 & 1'b0 ) ;
  assign n9890 = ( n9820 & n9839 ) | ( n9820 & n9881 ) | ( n9839 & n9881 ) ;
  assign n9891 = ( n9820 & ~n9841 ) | ( n9820 & n9881 ) | ( ~n9841 & n9881 ) ;
  assign n9892 = ~n9890 & n9891 ;
  assign n9893 = n9886 | n9892 ;
  assign n9894 = n9602 &  n9842 ;
  assign n9887 = x90 | n9602 ;
  assign n9888 = x90 &  n9602 ;
  assign n9889 = ( n9887 & ~n9888 ) | ( n9887 & 1'b0 ) | ( ~n9888 & 1'b0 ) ;
  assign n9898 = ( n9819 & n9839 ) | ( n9819 & n9889 ) | ( n9839 & n9889 ) ;
  assign n9899 = ( n9819 & ~n9841 ) | ( n9819 & n9889 ) | ( ~n9841 & n9889 ) ;
  assign n9900 = ~n9898 & n9899 ;
  assign n9901 = n9894 | n9900 ;
  assign n9902 = n9610 &  n9842 ;
  assign n9895 = x89 | n9610 ;
  assign n9896 = x89 &  n9610 ;
  assign n9897 = ( n9895 & ~n9896 ) | ( n9895 & 1'b0 ) | ( ~n9896 & 1'b0 ) ;
  assign n9906 = ( n9818 & n9839 ) | ( n9818 & n9897 ) | ( n9839 & n9897 ) ;
  assign n9907 = ( n9818 & ~n9841 ) | ( n9818 & n9897 ) | ( ~n9841 & n9897 ) ;
  assign n9908 = ~n9906 & n9907 ;
  assign n9909 = n9902 | n9908 ;
  assign n9910 = n9618 &  n9842 ;
  assign n9903 = x88 | n9618 ;
  assign n9904 = x88 &  n9618 ;
  assign n9905 = ( n9903 & ~n9904 ) | ( n9903 & 1'b0 ) | ( ~n9904 & 1'b0 ) ;
  assign n9914 = ( n9817 & n9839 ) | ( n9817 & n9905 ) | ( n9839 & n9905 ) ;
  assign n9915 = ( n9817 & ~n9841 ) | ( n9817 & n9905 ) | ( ~n9841 & n9905 ) ;
  assign n9916 = ~n9914 & n9915 ;
  assign n9917 = n9910 | n9916 ;
  assign n9918 = n9626 &  n9842 ;
  assign n9911 = x87 | n9626 ;
  assign n9912 = x87 &  n9626 ;
  assign n9913 = ( n9911 & ~n9912 ) | ( n9911 & 1'b0 ) | ( ~n9912 & 1'b0 ) ;
  assign n9922 = ( n9816 & n9839 ) | ( n9816 & n9913 ) | ( n9839 & n9913 ) ;
  assign n9923 = ( n9816 & ~n9841 ) | ( n9816 & n9913 ) | ( ~n9841 & n9913 ) ;
  assign n9924 = ~n9922 & n9923 ;
  assign n9925 = n9918 | n9924 ;
  assign n9926 = n9634 &  n9842 ;
  assign n9919 = x86 | n9634 ;
  assign n9920 = x86 &  n9634 ;
  assign n9921 = ( n9919 & ~n9920 ) | ( n9919 & 1'b0 ) | ( ~n9920 & 1'b0 ) ;
  assign n9930 = ( n9815 & n9839 ) | ( n9815 & n9921 ) | ( n9839 & n9921 ) ;
  assign n9931 = ( n9815 & ~n9841 ) | ( n9815 & n9921 ) | ( ~n9841 & n9921 ) ;
  assign n9932 = ~n9930 & n9931 ;
  assign n9933 = n9926 | n9932 ;
  assign n9934 = n9642 &  n9842 ;
  assign n9927 = x85 | n9642 ;
  assign n9928 = x85 &  n9642 ;
  assign n9929 = ( n9927 & ~n9928 ) | ( n9927 & 1'b0 ) | ( ~n9928 & 1'b0 ) ;
  assign n9938 = ( n9814 & n9839 ) | ( n9814 & n9929 ) | ( n9839 & n9929 ) ;
  assign n9939 = ( n9814 & ~n9841 ) | ( n9814 & n9929 ) | ( ~n9841 & n9929 ) ;
  assign n9940 = ~n9938 & n9939 ;
  assign n9941 = n9934 | n9940 ;
  assign n9942 = n9650 &  n9842 ;
  assign n9935 = x84 | n9650 ;
  assign n9936 = x84 &  n9650 ;
  assign n9937 = ( n9935 & ~n9936 ) | ( n9935 & 1'b0 ) | ( ~n9936 & 1'b0 ) ;
  assign n9946 = ( n9813 & n9839 ) | ( n9813 & n9937 ) | ( n9839 & n9937 ) ;
  assign n9947 = ( n9813 & ~n9841 ) | ( n9813 & n9937 ) | ( ~n9841 & n9937 ) ;
  assign n9948 = ~n9946 & n9947 ;
  assign n9949 = n9942 | n9948 ;
  assign n9950 = n9658 &  n9842 ;
  assign n9943 = x83 | n9658 ;
  assign n9944 = x83 &  n9658 ;
  assign n9945 = ( n9943 & ~n9944 ) | ( n9943 & 1'b0 ) | ( ~n9944 & 1'b0 ) ;
  assign n9954 = ( n9812 & n9839 ) | ( n9812 & n9945 ) | ( n9839 & n9945 ) ;
  assign n9955 = ( n9812 & ~n9841 ) | ( n9812 & n9945 ) | ( ~n9841 & n9945 ) ;
  assign n9956 = ~n9954 & n9955 ;
  assign n9957 = n9950 | n9956 ;
  assign n9958 = n9666 &  n9842 ;
  assign n9951 = x82 | n9666 ;
  assign n9952 = x82 &  n9666 ;
  assign n9953 = ( n9951 & ~n9952 ) | ( n9951 & 1'b0 ) | ( ~n9952 & 1'b0 ) ;
  assign n9962 = ( n9811 & n9839 ) | ( n9811 & n9953 ) | ( n9839 & n9953 ) ;
  assign n9963 = ( n9811 & ~n9841 ) | ( n9811 & n9953 ) | ( ~n9841 & n9953 ) ;
  assign n9964 = ~n9962 & n9963 ;
  assign n9965 = n9958 | n9964 ;
  assign n9966 = n9674 &  n9842 ;
  assign n9959 = x81 | n9674 ;
  assign n9960 = x81 &  n9674 ;
  assign n9961 = ( n9959 & ~n9960 ) | ( n9959 & 1'b0 ) | ( ~n9960 & 1'b0 ) ;
  assign n9970 = ( n9810 & n9839 ) | ( n9810 & n9961 ) | ( n9839 & n9961 ) ;
  assign n9971 = ( n9810 & ~n9841 ) | ( n9810 & n9961 ) | ( ~n9841 & n9961 ) ;
  assign n9972 = ~n9970 & n9971 ;
  assign n9973 = n9966 | n9972 ;
  assign n9974 = n9682 &  n9842 ;
  assign n9967 = x80 | n9682 ;
  assign n9968 = x80 &  n9682 ;
  assign n9969 = ( n9967 & ~n9968 ) | ( n9967 & 1'b0 ) | ( ~n9968 & 1'b0 ) ;
  assign n9978 = ( n9809 & n9839 ) | ( n9809 & n9969 ) | ( n9839 & n9969 ) ;
  assign n9979 = ( n9809 & ~n9841 ) | ( n9809 & n9969 ) | ( ~n9841 & n9969 ) ;
  assign n9980 = ~n9978 & n9979 ;
  assign n9981 = n9974 | n9980 ;
  assign n9982 = n9690 &  n9842 ;
  assign n9975 = x79 | n9690 ;
  assign n9976 = x79 &  n9690 ;
  assign n9977 = ( n9975 & ~n9976 ) | ( n9975 & 1'b0 ) | ( ~n9976 & 1'b0 ) ;
  assign n9986 = ( n9808 & n9839 ) | ( n9808 & n9977 ) | ( n9839 & n9977 ) ;
  assign n9987 = ( n9808 & ~n9841 ) | ( n9808 & n9977 ) | ( ~n9841 & n9977 ) ;
  assign n9988 = ~n9986 & n9987 ;
  assign n9989 = n9982 | n9988 ;
  assign n9990 = n9698 &  n9842 ;
  assign n9983 = x78 | n9698 ;
  assign n9984 = x78 &  n9698 ;
  assign n9985 = ( n9983 & ~n9984 ) | ( n9983 & 1'b0 ) | ( ~n9984 & 1'b0 ) ;
  assign n9994 = ( n9807 & n9839 ) | ( n9807 & n9985 ) | ( n9839 & n9985 ) ;
  assign n9995 = ( n9807 & ~n9841 ) | ( n9807 & n9985 ) | ( ~n9841 & n9985 ) ;
  assign n9996 = ~n9994 & n9995 ;
  assign n9997 = n9990 | n9996 ;
  assign n9998 = n9706 &  n9842 ;
  assign n9991 = x77 | n9706 ;
  assign n9992 = x77 &  n9706 ;
  assign n9993 = ( n9991 & ~n9992 ) | ( n9991 & 1'b0 ) | ( ~n9992 & 1'b0 ) ;
  assign n10002 = ( n9806 & n9839 ) | ( n9806 & n9993 ) | ( n9839 & n9993 ) ;
  assign n10003 = ( n9806 & ~n9841 ) | ( n9806 & n9993 ) | ( ~n9841 & n9993 ) ;
  assign n10004 = ~n10002 & n10003 ;
  assign n10005 = n9998 | n10004 ;
  assign n10006 = n9714 &  n9842 ;
  assign n9999 = x76 | n9714 ;
  assign n10000 = x76 &  n9714 ;
  assign n10001 = ( n9999 & ~n10000 ) | ( n9999 & 1'b0 ) | ( ~n10000 & 1'b0 ) ;
  assign n10010 = ( n9805 & n9839 ) | ( n9805 & n10001 ) | ( n9839 & n10001 ) ;
  assign n10011 = ( n9805 & ~n9841 ) | ( n9805 & n10001 ) | ( ~n9841 & n10001 ) ;
  assign n10012 = ~n10010 & n10011 ;
  assign n10013 = n10006 | n10012 ;
  assign n10014 = n9722 &  n9842 ;
  assign n10007 = x75 | n9722 ;
  assign n10008 = x75 &  n9722 ;
  assign n10009 = ( n10007 & ~n10008 ) | ( n10007 & 1'b0 ) | ( ~n10008 & 1'b0 ) ;
  assign n10018 = ( n9804 & n9839 ) | ( n9804 & n10009 ) | ( n9839 & n10009 ) ;
  assign n10019 = ( n9804 & ~n9841 ) | ( n9804 & n10009 ) | ( ~n9841 & n10009 ) ;
  assign n10020 = ~n10018 & n10019 ;
  assign n10021 = n10014 | n10020 ;
  assign n10022 = n9730 &  n9842 ;
  assign n10015 = x74 | n9730 ;
  assign n10016 = x74 &  n9730 ;
  assign n10017 = ( n10015 & ~n10016 ) | ( n10015 & 1'b0 ) | ( ~n10016 & 1'b0 ) ;
  assign n10026 = ( n9803 & n9839 ) | ( n9803 & n10017 ) | ( n9839 & n10017 ) ;
  assign n10027 = ( n9803 & ~n9841 ) | ( n9803 & n10017 ) | ( ~n9841 & n10017 ) ;
  assign n10028 = ~n10026 & n10027 ;
  assign n10029 = n10022 | n10028 ;
  assign n10030 = n9738 &  n9842 ;
  assign n10023 = x73 | n9738 ;
  assign n10024 = x73 &  n9738 ;
  assign n10025 = ( n10023 & ~n10024 ) | ( n10023 & 1'b0 ) | ( ~n10024 & 1'b0 ) ;
  assign n10034 = ( n9802 & n9839 ) | ( n9802 & n10025 ) | ( n9839 & n10025 ) ;
  assign n10035 = ( n9802 & ~n9841 ) | ( n9802 & n10025 ) | ( ~n9841 & n10025 ) ;
  assign n10036 = ~n10034 & n10035 ;
  assign n10037 = n10030 | n10036 ;
  assign n10038 = n9746 &  n9842 ;
  assign n10031 = x72 | n9746 ;
  assign n10032 = x72 &  n9746 ;
  assign n10033 = ( n10031 & ~n10032 ) | ( n10031 & 1'b0 ) | ( ~n10032 & 1'b0 ) ;
  assign n10042 = ( n9801 & n9839 ) | ( n9801 & n10033 ) | ( n9839 & n10033 ) ;
  assign n10043 = ( n9801 & ~n9841 ) | ( n9801 & n10033 ) | ( ~n9841 & n10033 ) ;
  assign n10044 = ~n10042 & n10043 ;
  assign n10045 = n10038 | n10044 ;
  assign n10046 = n9754 &  n9842 ;
  assign n10039 = x71 | n9754 ;
  assign n10040 = x71 &  n9754 ;
  assign n10041 = ( n10039 & ~n10040 ) | ( n10039 & 1'b0 ) | ( ~n10040 & 1'b0 ) ;
  assign n10050 = ( n9800 & n9839 ) | ( n9800 & n10041 ) | ( n9839 & n10041 ) ;
  assign n10051 = ( n9800 & ~n9841 ) | ( n9800 & n10041 ) | ( ~n9841 & n10041 ) ;
  assign n10052 = ~n10050 & n10051 ;
  assign n10053 = n10046 | n10052 ;
  assign n10054 = n9762 &  n9842 ;
  assign n10047 = x70 | n9762 ;
  assign n10048 = x70 &  n9762 ;
  assign n10049 = ( n10047 & ~n10048 ) | ( n10047 & 1'b0 ) | ( ~n10048 & 1'b0 ) ;
  assign n10058 = ( n9799 & n9839 ) | ( n9799 & n10049 ) | ( n9839 & n10049 ) ;
  assign n10059 = ( n9799 & ~n9841 ) | ( n9799 & n10049 ) | ( ~n9841 & n10049 ) ;
  assign n10060 = ~n10058 & n10059 ;
  assign n10061 = n10054 | n10060 ;
  assign n10062 = n9770 &  n9842 ;
  assign n10055 = x69 | n9770 ;
  assign n10056 = x69 &  n9770 ;
  assign n10057 = ( n10055 & ~n10056 ) | ( n10055 & 1'b0 ) | ( ~n10056 & 1'b0 ) ;
  assign n10066 = ( n9798 & n9839 ) | ( n9798 & n10057 ) | ( n9839 & n10057 ) ;
  assign n10067 = ( n9798 & ~n9841 ) | ( n9798 & n10057 ) | ( ~n9841 & n10057 ) ;
  assign n10068 = ~n10066 & n10067 ;
  assign n10069 = n10062 | n10068 ;
  assign n10070 = n9778 &  n9842 ;
  assign n10063 = x68 | n9778 ;
  assign n10064 = x68 &  n9778 ;
  assign n10065 = ( n10063 & ~n10064 ) | ( n10063 & 1'b0 ) | ( ~n10064 & 1'b0 ) ;
  assign n10074 = ( n9797 & n9839 ) | ( n9797 & n10065 ) | ( n9839 & n10065 ) ;
  assign n10075 = ( n9797 & ~n9841 ) | ( n9797 & n10065 ) | ( ~n9841 & n10065 ) ;
  assign n10076 = ~n10074 & n10075 ;
  assign n10077 = n10070 | n10076 ;
  assign n10078 = n9783 &  n9842 ;
  assign n10071 = x67 | n9783 ;
  assign n10072 = x67 &  n9783 ;
  assign n10073 = ( n10071 & ~n10072 ) | ( n10071 & 1'b0 ) | ( ~n10072 & 1'b0 ) ;
  assign n10082 = ( n9796 & n9839 ) | ( n9796 & n10073 ) | ( n9839 & n10073 ) ;
  assign n10083 = ( n9796 & ~n9841 ) | ( n9796 & n10073 ) | ( ~n9841 & n10073 ) ;
  assign n10084 = ~n10082 & n10083 ;
  assign n10085 = n10078 | n10084 ;
  assign n10086 = n9789 &  n9842 ;
  assign n10079 = x66 | n9789 ;
  assign n10080 = x66 &  n9789 ;
  assign n10081 = ( n10079 & ~n10080 ) | ( n10079 & 1'b0 ) | ( ~n10080 & 1'b0 ) ;
  assign n10091 = ( n9795 & ~n9839 ) | ( n9795 & n10081 ) | ( ~n9839 & n10081 ) ;
  assign n10092 = ( n9795 & n9841 ) | ( n9795 & n10081 ) | ( n9841 & n10081 ) ;
  assign n10093 = ( n10091 & ~n10092 ) | ( n10091 & 1'b0 ) | ( ~n10092 & 1'b0 ) ;
  assign n10094 = n10086 | n10093 ;
  assign n10095 = n9793 &  n9842 ;
  assign n10087 = x65 &  n9793 ;
  assign n10088 = ( n9791 & ~x65 ) | ( n9791 & n9792 ) | ( ~x65 & n9792 ) ;
  assign n10089 = x65 | n10088 ;
  assign n10090 = ( n9794 & ~n10087 ) | ( n9794 & n10089 ) | ( ~n10087 & n10089 ) ;
  assign n10096 = ( x65 & n9793 ) | ( x65 & n9794 ) | ( n9793 & n9794 ) ;
  assign n10097 = ( n9841 & ~n10087 ) | ( n9841 & n10096 ) | ( ~n10087 & n10096 ) ;
  assign n10098 = ( n9839 & n10090 ) | ( n9839 & n10097 ) | ( n10090 & n10097 ) ;
  assign n10099 = ( n10090 & ~n10098 ) | ( n10090 & 1'b0 ) | ( ~n10098 & 1'b0 ) ;
  assign n10100 = n10095 | n10099 ;
  assign n10101 = ( x64 & ~x110 ) | ( x64 & 1'b0 ) | ( ~x110 & 1'b0 ) ;
  assign n10102 = ( n232 & ~n249 ) | ( n232 & n10101 ) | ( ~n249 & n10101 ) ;
  assign n10103 = ~n232 & n10102 ;
  assign n10104 = ~n425 & n10103 ;
  assign n10105 = n9839 &  n10104 ;
  assign n10106 = ( x18 & ~n10104 ) | ( x18 & n10105 ) | ( ~n10104 & n10105 ) ;
  assign n10107 = ~n172 & n9794 ;
  assign n10108 = ( n160 & ~n170 ) | ( n160 & n10107 ) | ( ~n170 & n10107 ) ;
  assign n10109 = ~n160 & n10108 ;
  assign n10110 = ~n9839 & n10109 ;
  assign n10111 = n10106 | n10110 ;
  assign n10112 = ~x17 & x64 ;
  assign n10113 = ( x65 & ~n10111 ) | ( x65 & n10112 ) | ( ~n10111 & n10112 ) ;
  assign n10114 = ( x66 & ~n10100 ) | ( x66 & n10113 ) | ( ~n10100 & n10113 ) ;
  assign n10115 = ( x67 & ~n10094 ) | ( x67 & n10114 ) | ( ~n10094 & n10114 ) ;
  assign n10116 = ( x68 & ~n10085 ) | ( x68 & n10115 ) | ( ~n10085 & n10115 ) ;
  assign n10117 = ( x69 & ~n10077 ) | ( x69 & n10116 ) | ( ~n10077 & n10116 ) ;
  assign n10118 = ( x70 & ~n10069 ) | ( x70 & n10117 ) | ( ~n10069 & n10117 ) ;
  assign n10119 = ( x71 & ~n10061 ) | ( x71 & n10118 ) | ( ~n10061 & n10118 ) ;
  assign n10120 = ( x72 & ~n10053 ) | ( x72 & n10119 ) | ( ~n10053 & n10119 ) ;
  assign n10121 = ( x73 & ~n10045 ) | ( x73 & n10120 ) | ( ~n10045 & n10120 ) ;
  assign n10122 = ( x74 & ~n10037 ) | ( x74 & n10121 ) | ( ~n10037 & n10121 ) ;
  assign n10123 = ( x75 & ~n10029 ) | ( x75 & n10122 ) | ( ~n10029 & n10122 ) ;
  assign n10124 = ( x76 & ~n10021 ) | ( x76 & n10123 ) | ( ~n10021 & n10123 ) ;
  assign n10125 = ( x77 & ~n10013 ) | ( x77 & n10124 ) | ( ~n10013 & n10124 ) ;
  assign n10126 = ( x78 & ~n10005 ) | ( x78 & n10125 ) | ( ~n10005 & n10125 ) ;
  assign n10127 = ( x79 & ~n9997 ) | ( x79 & n10126 ) | ( ~n9997 & n10126 ) ;
  assign n10128 = ( x80 & ~n9989 ) | ( x80 & n10127 ) | ( ~n9989 & n10127 ) ;
  assign n10129 = ( x81 & ~n9981 ) | ( x81 & n10128 ) | ( ~n9981 & n10128 ) ;
  assign n10130 = ( x82 & ~n9973 ) | ( x82 & n10129 ) | ( ~n9973 & n10129 ) ;
  assign n10131 = ( x83 & ~n9965 ) | ( x83 & n10130 ) | ( ~n9965 & n10130 ) ;
  assign n10132 = ( x84 & ~n9957 ) | ( x84 & n10131 ) | ( ~n9957 & n10131 ) ;
  assign n10133 = ( x85 & ~n9949 ) | ( x85 & n10132 ) | ( ~n9949 & n10132 ) ;
  assign n10134 = ( x86 & ~n9941 ) | ( x86 & n10133 ) | ( ~n9941 & n10133 ) ;
  assign n10135 = ( x87 & ~n9933 ) | ( x87 & n10134 ) | ( ~n9933 & n10134 ) ;
  assign n10136 = ( x88 & ~n9925 ) | ( x88 & n10135 ) | ( ~n9925 & n10135 ) ;
  assign n10137 = ( x89 & ~n9917 ) | ( x89 & n10136 ) | ( ~n9917 & n10136 ) ;
  assign n10138 = ( x90 & ~n9909 ) | ( x90 & n10137 ) | ( ~n9909 & n10137 ) ;
  assign n10139 = ( x91 & ~n9901 ) | ( x91 & n10138 ) | ( ~n9901 & n10138 ) ;
  assign n10140 = ( x92 & ~n9893 ) | ( x92 & n10139 ) | ( ~n9893 & n10139 ) ;
  assign n10141 = ( x93 & ~n9885 ) | ( x93 & n10140 ) | ( ~n9885 & n10140 ) ;
  assign n10142 = ( x94 & ~n9877 ) | ( x94 & n10141 ) | ( ~n9877 & n10141 ) ;
  assign n10143 = ( x95 & ~n9869 ) | ( x95 & n10142 ) | ( ~n9869 & n10142 ) ;
  assign n10144 = ( x96 & ~n9861 ) | ( x96 & n10143 ) | ( ~n9861 & n10143 ) ;
  assign n10148 = ( x97 & ~n9853 ) | ( x97 & n10144 ) | ( ~n9853 & n10144 ) ;
  assign n10248 = ( x98 & ~n10156 ) | ( x98 & n10148 ) | ( ~n10156 & n10148 ) ;
  assign n10249 = ( x99 & ~n10247 ) | ( x99 & n10248 ) | ( ~n10247 & n10248 ) ;
  assign n10250 = ( x100 & ~n10242 ) | ( x100 & n10249 ) | ( ~n10242 & n10249 ) ;
  assign n10251 = ( x101 & ~n10234 ) | ( x101 & n10250 ) | ( ~n10234 & n10250 ) ;
  assign n10252 = ( x102 & ~n10226 ) | ( x102 & n10251 ) | ( ~n10226 & n10251 ) ;
  assign n10253 = ( x103 & ~n10218 ) | ( x103 & n10252 ) | ( ~n10218 & n10252 ) ;
  assign n10254 = ( x104 & ~n10210 ) | ( x104 & n10253 ) | ( ~n10210 & n10253 ) ;
  assign n10255 = ( x105 & ~n10202 ) | ( x105 & n10254 ) | ( ~n10202 & n10254 ) ;
  assign n10256 = ( x106 & ~n10194 ) | ( x106 & n10255 ) | ( ~n10194 & n10255 ) ;
  assign n10257 = ( x107 & ~n10186 ) | ( x107 & n10256 ) | ( ~n10186 & n10256 ) ;
  assign n10258 = ( x108 & ~n10178 ) | ( x108 & n10257 ) | ( ~n10178 & n10257 ) ;
  assign n10259 = ( x109 & ~n10170 ) | ( x109 & n10258 ) | ( ~n10170 & n10258 ) ;
  assign n10263 = n232 | n249 ;
  assign n10264 = n425 | n10263 ;
  assign n10260 = x109 | n9838 ;
  assign n10261 = ( x109 & n9838 ) | ( x109 & n9841 ) | ( n9838 & n9841 ) ;
  assign n10262 = ( n9461 & ~n10260 ) | ( n9461 & n10261 ) | ( ~n10260 & n10261 ) ;
  assign n10266 = x110 &  n10262 ;
  assign n10265 = x110 | n10262 ;
  assign n10267 = ( n10264 & ~n10266 ) | ( n10264 & n10265 ) | ( ~n10266 & n10265 ) ;
  assign n10268 = n10259 | n10267 ;
  assign n10269 = ~n10262 |  n9841 ;
  assign n10595 = n10170 &  n10269 ;
  assign n10596 = n10268 &  n10595 ;
  assign n10592 = x109 | n10170 ;
  assign n10593 = x109 &  n10170 ;
  assign n10594 = ( n10592 & ~n10593 ) | ( n10592 & 1'b0 ) | ( ~n10593 & 1'b0 ) ;
  assign n10597 = n10258 &  n10594 ;
  assign n10270 = n10268 &  n10269 ;
  assign n10598 = ( n10258 & ~n10270 ) | ( n10258 & n10594 ) | ( ~n10270 & n10594 ) ;
  assign n10599 = ( n10596 & ~n10597 ) | ( n10596 & n10598 ) | ( ~n10597 & n10598 ) ;
  assign n10603 = n10178 &  n10269 ;
  assign n10604 = n10268 &  n10603 ;
  assign n10589 = x108 | n10178 ;
  assign n10590 = x108 &  n10178 ;
  assign n10591 = ( n10589 & ~n10590 ) | ( n10589 & 1'b0 ) | ( ~n10590 & 1'b0 ) ;
  assign n10605 = n10257 &  n10591 ;
  assign n10606 = ( n10257 & ~n10270 ) | ( n10257 & n10591 ) | ( ~n10270 & n10591 ) ;
  assign n10607 = ( n10604 & ~n10605 ) | ( n10604 & n10606 ) | ( ~n10605 & n10606 ) ;
  assign n10611 = n10186 &  n10269 ;
  assign n10612 = n10268 &  n10611 ;
  assign n10600 = x107 | n10186 ;
  assign n10601 = x107 &  n10186 ;
  assign n10602 = ( n10600 & ~n10601 ) | ( n10600 & 1'b0 ) | ( ~n10601 & 1'b0 ) ;
  assign n10613 = n10256 &  n10602 ;
  assign n10614 = ( n10256 & ~n10270 ) | ( n10256 & n10602 ) | ( ~n10270 & n10602 ) ;
  assign n10615 = ( n10612 & ~n10613 ) | ( n10612 & n10614 ) | ( ~n10613 & n10614 ) ;
  assign n10619 = n10194 &  n10269 ;
  assign n10620 = n10268 &  n10619 ;
  assign n10608 = x106 | n10194 ;
  assign n10609 = x106 &  n10194 ;
  assign n10610 = ( n10608 & ~n10609 ) | ( n10608 & 1'b0 ) | ( ~n10609 & 1'b0 ) ;
  assign n10621 = n10255 &  n10610 ;
  assign n10622 = ( n10255 & ~n10270 ) | ( n10255 & n10610 ) | ( ~n10270 & n10610 ) ;
  assign n10623 = ( n10620 & ~n10621 ) | ( n10620 & n10622 ) | ( ~n10621 & n10622 ) ;
  assign n10627 = n10202 &  n10269 ;
  assign n10628 = n10268 &  n10627 ;
  assign n10616 = x105 | n10202 ;
  assign n10617 = x105 &  n10202 ;
  assign n10618 = ( n10616 & ~n10617 ) | ( n10616 & 1'b0 ) | ( ~n10617 & 1'b0 ) ;
  assign n10629 = n10254 &  n10618 ;
  assign n10630 = ( n10254 & ~n10270 ) | ( n10254 & n10618 ) | ( ~n10270 & n10618 ) ;
  assign n10631 = ( n10628 & ~n10629 ) | ( n10628 & n10630 ) | ( ~n10629 & n10630 ) ;
  assign n10635 = n10210 &  n10269 ;
  assign n10636 = n10268 &  n10635 ;
  assign n10624 = x104 | n10210 ;
  assign n10625 = x104 &  n10210 ;
  assign n10626 = ( n10624 & ~n10625 ) | ( n10624 & 1'b0 ) | ( ~n10625 & 1'b0 ) ;
  assign n10638 = ( n10253 & n10270 ) | ( n10253 & n10626 ) | ( n10270 & n10626 ) ;
  assign n10637 = n10253 | n10626 ;
  assign n10639 = ( n10636 & ~n10638 ) | ( n10636 & n10637 ) | ( ~n10638 & n10637 ) ;
  assign n10643 = n10218 &  n10269 ;
  assign n10644 = n10268 &  n10643 ;
  assign n10632 = x103 | n10218 ;
  assign n10633 = x103 &  n10218 ;
  assign n10634 = ( n10632 & ~n10633 ) | ( n10632 & 1'b0 ) | ( ~n10633 & 1'b0 ) ;
  assign n10646 = ( n10252 & n10270 ) | ( n10252 & n10634 ) | ( n10270 & n10634 ) ;
  assign n10645 = n10252 | n10634 ;
  assign n10647 = ( n10644 & ~n10646 ) | ( n10644 & n10645 ) | ( ~n10646 & n10645 ) ;
  assign n10651 = n10226 &  n10269 ;
  assign n10652 = n10268 &  n10651 ;
  assign n10640 = x102 | n10226 ;
  assign n10641 = x102 &  n10226 ;
  assign n10642 = ( n10640 & ~n10641 ) | ( n10640 & 1'b0 ) | ( ~n10641 & 1'b0 ) ;
  assign n10654 = ( n10251 & n10270 ) | ( n10251 & n10642 ) | ( n10270 & n10642 ) ;
  assign n10653 = n10251 | n10642 ;
  assign n10655 = ( n10652 & ~n10654 ) | ( n10652 & n10653 ) | ( ~n10654 & n10653 ) ;
  assign n10659 = n10234 &  n10269 ;
  assign n10660 = n10268 &  n10659 ;
  assign n10648 = x101 | n10234 ;
  assign n10649 = x101 &  n10234 ;
  assign n10650 = ( n10648 & ~n10649 ) | ( n10648 & 1'b0 ) | ( ~n10649 & 1'b0 ) ;
  assign n10662 = ( n10250 & n10270 ) | ( n10250 & n10650 ) | ( n10270 & n10650 ) ;
  assign n10661 = n10250 | n10650 ;
  assign n10663 = ( n10660 & ~n10662 ) | ( n10660 & n10661 ) | ( ~n10662 & n10661 ) ;
  assign n10664 = n10242 &  n10269 ;
  assign n10665 = n10268 &  n10664 ;
  assign n10656 = x100 | n10242 ;
  assign n10657 = x100 &  n10242 ;
  assign n10658 = ( n10656 & ~n10657 ) | ( n10656 & 1'b0 ) | ( ~n10657 & 1'b0 ) ;
  assign n10667 = ( n10249 & n10270 ) | ( n10249 & n10658 ) | ( n10270 & n10658 ) ;
  assign n10666 = n10249 | n10658 ;
  assign n10668 = ( n10665 & ~n10667 ) | ( n10665 & n10666 ) | ( ~n10667 & n10666 ) ;
  assign n10581 = n10247 &  n10269 ;
  assign n10582 = n10268 &  n10581 ;
  assign n10578 = x99 | n10247 ;
  assign n10579 = x99 &  n10247 ;
  assign n10580 = ( n10578 & ~n10579 ) | ( n10578 & 1'b0 ) | ( ~n10579 & 1'b0 ) ;
  assign n10584 = ( n10248 & n10270 ) | ( n10248 & n10580 ) | ( n10270 & n10580 ) ;
  assign n10583 = n10248 | n10580 ;
  assign n10585 = ( n10582 & ~n10584 ) | ( n10582 & n10583 ) | ( ~n10584 & n10583 ) ;
  assign n10271 = n10156 &  n10269 ;
  assign n10272 = n10268 &  n10271 ;
  assign n10157 = x98 | n10156 ;
  assign n10158 = x98 &  n10156 ;
  assign n10159 = ( n10157 & ~n10158 ) | ( n10157 & 1'b0 ) | ( ~n10158 & 1'b0 ) ;
  assign n10274 = ( n10148 & n10159 ) | ( n10148 & n10270 ) | ( n10159 & n10270 ) ;
  assign n10273 = n10148 | n10159 ;
  assign n10275 = ( n10272 & ~n10274 ) | ( n10272 & n10273 ) | ( ~n10274 & n10273 ) ;
  assign n10279 = n9853 &  n10269 ;
  assign n10280 = n10268 &  n10279 ;
  assign n10145 = x97 | n9853 ;
  assign n10146 = x97 &  n9853 ;
  assign n10147 = ( n10145 & ~n10146 ) | ( n10145 & 1'b0 ) | ( ~n10146 & 1'b0 ) ;
  assign n10281 = n10144 &  n10147 ;
  assign n10282 = ( n10144 & ~n10270 ) | ( n10144 & n10147 ) | ( ~n10270 & n10147 ) ;
  assign n10283 = ( n10280 & ~n10281 ) | ( n10280 & n10282 ) | ( ~n10281 & n10282 ) ;
  assign n10287 = n9861 &  n10269 ;
  assign n10288 = n10268 &  n10287 ;
  assign n10276 = x96 | n9861 ;
  assign n10277 = x96 &  n9861 ;
  assign n10278 = ( n10276 & ~n10277 ) | ( n10276 & 1'b0 ) | ( ~n10277 & 1'b0 ) ;
  assign n10290 = ( n10143 & n10270 ) | ( n10143 & n10278 ) | ( n10270 & n10278 ) ;
  assign n10289 = n10143 | n10278 ;
  assign n10291 = ( n10288 & ~n10290 ) | ( n10288 & n10289 ) | ( ~n10290 & n10289 ) ;
  assign n10295 = n9869 &  n10269 ;
  assign n10296 = n10268 &  n10295 ;
  assign n10284 = x95 | n9869 ;
  assign n10285 = x95 &  n9869 ;
  assign n10286 = ( n10284 & ~n10285 ) | ( n10284 & 1'b0 ) | ( ~n10285 & 1'b0 ) ;
  assign n10298 = ( n10142 & n10270 ) | ( n10142 & n10286 ) | ( n10270 & n10286 ) ;
  assign n10297 = n10142 | n10286 ;
  assign n10299 = ( n10296 & ~n10298 ) | ( n10296 & n10297 ) | ( ~n10298 & n10297 ) ;
  assign n10303 = n9877 &  n10269 ;
  assign n10304 = n10268 &  n10303 ;
  assign n10292 = x94 | n9877 ;
  assign n10293 = x94 &  n9877 ;
  assign n10294 = ( n10292 & ~n10293 ) | ( n10292 & 1'b0 ) | ( ~n10293 & 1'b0 ) ;
  assign n10306 = ( n10141 & n10270 ) | ( n10141 & n10294 ) | ( n10270 & n10294 ) ;
  assign n10305 = n10141 | n10294 ;
  assign n10307 = ( n10304 & ~n10306 ) | ( n10304 & n10305 ) | ( ~n10306 & n10305 ) ;
  assign n10311 = n9885 &  n10269 ;
  assign n10312 = n10268 &  n10311 ;
  assign n10300 = x93 | n9885 ;
  assign n10301 = x93 &  n9885 ;
  assign n10302 = ( n10300 & ~n10301 ) | ( n10300 & 1'b0 ) | ( ~n10301 & 1'b0 ) ;
  assign n10314 = ( n10140 & n10270 ) | ( n10140 & n10302 ) | ( n10270 & n10302 ) ;
  assign n10313 = n10140 | n10302 ;
  assign n10315 = ( n10312 & ~n10314 ) | ( n10312 & n10313 ) | ( ~n10314 & n10313 ) ;
  assign n10319 = n9893 &  n10269 ;
  assign n10320 = n10268 &  n10319 ;
  assign n10308 = x92 | n9893 ;
  assign n10309 = x92 &  n9893 ;
  assign n10310 = ( n10308 & ~n10309 ) | ( n10308 & 1'b0 ) | ( ~n10309 & 1'b0 ) ;
  assign n10322 = ( n10139 & n10270 ) | ( n10139 & n10310 ) | ( n10270 & n10310 ) ;
  assign n10321 = n10139 | n10310 ;
  assign n10323 = ( n10320 & ~n10322 ) | ( n10320 & n10321 ) | ( ~n10322 & n10321 ) ;
  assign n10327 = n9901 &  n10269 ;
  assign n10328 = n10268 &  n10327 ;
  assign n10316 = x91 | n9901 ;
  assign n10317 = x91 &  n9901 ;
  assign n10318 = ( n10316 & ~n10317 ) | ( n10316 & 1'b0 ) | ( ~n10317 & 1'b0 ) ;
  assign n10330 = ( n10138 & n10270 ) | ( n10138 & n10318 ) | ( n10270 & n10318 ) ;
  assign n10329 = n10138 | n10318 ;
  assign n10331 = ( n10328 & ~n10330 ) | ( n10328 & n10329 ) | ( ~n10330 & n10329 ) ;
  assign n10335 = n9909 &  n10269 ;
  assign n10336 = n10268 &  n10335 ;
  assign n10324 = x90 | n9909 ;
  assign n10325 = x90 &  n9909 ;
  assign n10326 = ( n10324 & ~n10325 ) | ( n10324 & 1'b0 ) | ( ~n10325 & 1'b0 ) ;
  assign n10338 = ( n10137 & n10270 ) | ( n10137 & n10326 ) | ( n10270 & n10326 ) ;
  assign n10337 = n10137 | n10326 ;
  assign n10339 = ( n10336 & ~n10338 ) | ( n10336 & n10337 ) | ( ~n10338 & n10337 ) ;
  assign n10343 = n9917 &  n10269 ;
  assign n10344 = n10268 &  n10343 ;
  assign n10332 = x89 | n9917 ;
  assign n10333 = x89 &  n9917 ;
  assign n10334 = ( n10332 & ~n10333 ) | ( n10332 & 1'b0 ) | ( ~n10333 & 1'b0 ) ;
  assign n10346 = ( n10136 & n10270 ) | ( n10136 & n10334 ) | ( n10270 & n10334 ) ;
  assign n10345 = n10136 | n10334 ;
  assign n10347 = ( n10344 & ~n10346 ) | ( n10344 & n10345 ) | ( ~n10346 & n10345 ) ;
  assign n10351 = n9925 &  n10269 ;
  assign n10352 = n10268 &  n10351 ;
  assign n10340 = x88 | n9925 ;
  assign n10341 = x88 &  n9925 ;
  assign n10342 = ( n10340 & ~n10341 ) | ( n10340 & 1'b0 ) | ( ~n10341 & 1'b0 ) ;
  assign n10354 = ( n10135 & n10270 ) | ( n10135 & n10342 ) | ( n10270 & n10342 ) ;
  assign n10353 = n10135 | n10342 ;
  assign n10355 = ( n10352 & ~n10354 ) | ( n10352 & n10353 ) | ( ~n10354 & n10353 ) ;
  assign n10359 = n9933 &  n10269 ;
  assign n10360 = n10268 &  n10359 ;
  assign n10348 = x87 | n9933 ;
  assign n10349 = x87 &  n9933 ;
  assign n10350 = ( n10348 & ~n10349 ) | ( n10348 & 1'b0 ) | ( ~n10349 & 1'b0 ) ;
  assign n10362 = ( n10134 & n10270 ) | ( n10134 & n10350 ) | ( n10270 & n10350 ) ;
  assign n10361 = n10134 | n10350 ;
  assign n10363 = ( n10360 & ~n10362 ) | ( n10360 & n10361 ) | ( ~n10362 & n10361 ) ;
  assign n10367 = n9941 &  n10269 ;
  assign n10368 = n10268 &  n10367 ;
  assign n10356 = x86 | n9941 ;
  assign n10357 = x86 &  n9941 ;
  assign n10358 = ( n10356 & ~n10357 ) | ( n10356 & 1'b0 ) | ( ~n10357 & 1'b0 ) ;
  assign n10370 = ( n10133 & n10270 ) | ( n10133 & n10358 ) | ( n10270 & n10358 ) ;
  assign n10369 = n10133 | n10358 ;
  assign n10371 = ( n10368 & ~n10370 ) | ( n10368 & n10369 ) | ( ~n10370 & n10369 ) ;
  assign n10375 = n9949 &  n10269 ;
  assign n10376 = n10268 &  n10375 ;
  assign n10364 = x85 | n9949 ;
  assign n10365 = x85 &  n9949 ;
  assign n10366 = ( n10364 & ~n10365 ) | ( n10364 & 1'b0 ) | ( ~n10365 & 1'b0 ) ;
  assign n10378 = ( n10132 & n10270 ) | ( n10132 & n10366 ) | ( n10270 & n10366 ) ;
  assign n10377 = n10132 | n10366 ;
  assign n10379 = ( n10376 & ~n10378 ) | ( n10376 & n10377 ) | ( ~n10378 & n10377 ) ;
  assign n10383 = n9957 &  n10269 ;
  assign n10384 = n10268 &  n10383 ;
  assign n10372 = x84 | n9957 ;
  assign n10373 = x84 &  n9957 ;
  assign n10374 = ( n10372 & ~n10373 ) | ( n10372 & 1'b0 ) | ( ~n10373 & 1'b0 ) ;
  assign n10386 = ( n10131 & n10270 ) | ( n10131 & n10374 ) | ( n10270 & n10374 ) ;
  assign n10385 = n10131 | n10374 ;
  assign n10387 = ( n10384 & ~n10386 ) | ( n10384 & n10385 ) | ( ~n10386 & n10385 ) ;
  assign n10391 = n9965 &  n10269 ;
  assign n10392 = n10268 &  n10391 ;
  assign n10380 = x83 | n9965 ;
  assign n10381 = x83 &  n9965 ;
  assign n10382 = ( n10380 & ~n10381 ) | ( n10380 & 1'b0 ) | ( ~n10381 & 1'b0 ) ;
  assign n10394 = ( n10130 & n10270 ) | ( n10130 & n10382 ) | ( n10270 & n10382 ) ;
  assign n10393 = n10130 | n10382 ;
  assign n10395 = ( n10392 & ~n10394 ) | ( n10392 & n10393 ) | ( ~n10394 & n10393 ) ;
  assign n10399 = n9973 &  n10269 ;
  assign n10400 = n10268 &  n10399 ;
  assign n10388 = x82 | n9973 ;
  assign n10389 = x82 &  n9973 ;
  assign n10390 = ( n10388 & ~n10389 ) | ( n10388 & 1'b0 ) | ( ~n10389 & 1'b0 ) ;
  assign n10402 = ( n10129 & n10270 ) | ( n10129 & n10390 ) | ( n10270 & n10390 ) ;
  assign n10401 = n10129 | n10390 ;
  assign n10403 = ( n10400 & ~n10402 ) | ( n10400 & n10401 ) | ( ~n10402 & n10401 ) ;
  assign n10407 = n9981 &  n10269 ;
  assign n10408 = n10268 &  n10407 ;
  assign n10396 = x81 | n9981 ;
  assign n10397 = x81 &  n9981 ;
  assign n10398 = ( n10396 & ~n10397 ) | ( n10396 & 1'b0 ) | ( ~n10397 & 1'b0 ) ;
  assign n10410 = ( n10128 & n10270 ) | ( n10128 & n10398 ) | ( n10270 & n10398 ) ;
  assign n10409 = n10128 | n10398 ;
  assign n10411 = ( n10408 & ~n10410 ) | ( n10408 & n10409 ) | ( ~n10410 & n10409 ) ;
  assign n10415 = n9989 &  n10269 ;
  assign n10416 = n10268 &  n10415 ;
  assign n10404 = x80 | n9989 ;
  assign n10405 = x80 &  n9989 ;
  assign n10406 = ( n10404 & ~n10405 ) | ( n10404 & 1'b0 ) | ( ~n10405 & 1'b0 ) ;
  assign n10418 = ( n10127 & n10270 ) | ( n10127 & n10406 ) | ( n10270 & n10406 ) ;
  assign n10417 = n10127 | n10406 ;
  assign n10419 = ( n10416 & ~n10418 ) | ( n10416 & n10417 ) | ( ~n10418 & n10417 ) ;
  assign n10423 = n9997 &  n10269 ;
  assign n10424 = n10268 &  n10423 ;
  assign n10412 = x79 | n9997 ;
  assign n10413 = x79 &  n9997 ;
  assign n10414 = ( n10412 & ~n10413 ) | ( n10412 & 1'b0 ) | ( ~n10413 & 1'b0 ) ;
  assign n10426 = ( n10126 & n10270 ) | ( n10126 & n10414 ) | ( n10270 & n10414 ) ;
  assign n10425 = n10126 | n10414 ;
  assign n10427 = ( n10424 & ~n10426 ) | ( n10424 & n10425 ) | ( ~n10426 & n10425 ) ;
  assign n10431 = n10005 &  n10269 ;
  assign n10432 = n10268 &  n10431 ;
  assign n10420 = x78 | n10005 ;
  assign n10421 = x78 &  n10005 ;
  assign n10422 = ( n10420 & ~n10421 ) | ( n10420 & 1'b0 ) | ( ~n10421 & 1'b0 ) ;
  assign n10434 = ( n10125 & n10270 ) | ( n10125 & n10422 ) | ( n10270 & n10422 ) ;
  assign n10433 = n10125 | n10422 ;
  assign n10435 = ( n10432 & ~n10434 ) | ( n10432 & n10433 ) | ( ~n10434 & n10433 ) ;
  assign n10439 = n10013 &  n10269 ;
  assign n10440 = n10268 &  n10439 ;
  assign n10428 = x77 | n10013 ;
  assign n10429 = x77 &  n10013 ;
  assign n10430 = ( n10428 & ~n10429 ) | ( n10428 & 1'b0 ) | ( ~n10429 & 1'b0 ) ;
  assign n10442 = ( n10124 & n10270 ) | ( n10124 & n10430 ) | ( n10270 & n10430 ) ;
  assign n10441 = n10124 | n10430 ;
  assign n10443 = ( n10440 & ~n10442 ) | ( n10440 & n10441 ) | ( ~n10442 & n10441 ) ;
  assign n10447 = n10021 &  n10269 ;
  assign n10448 = n10268 &  n10447 ;
  assign n10436 = x76 | n10021 ;
  assign n10437 = x76 &  n10021 ;
  assign n10438 = ( n10436 & ~n10437 ) | ( n10436 & 1'b0 ) | ( ~n10437 & 1'b0 ) ;
  assign n10450 = ( n10123 & n10270 ) | ( n10123 & n10438 ) | ( n10270 & n10438 ) ;
  assign n10449 = n10123 | n10438 ;
  assign n10451 = ( n10448 & ~n10450 ) | ( n10448 & n10449 ) | ( ~n10450 & n10449 ) ;
  assign n10455 = n10029 &  n10269 ;
  assign n10456 = n10268 &  n10455 ;
  assign n10444 = x75 | n10029 ;
  assign n10445 = x75 &  n10029 ;
  assign n10446 = ( n10444 & ~n10445 ) | ( n10444 & 1'b0 ) | ( ~n10445 & 1'b0 ) ;
  assign n10458 = ( n10122 & n10270 ) | ( n10122 & n10446 ) | ( n10270 & n10446 ) ;
  assign n10457 = n10122 | n10446 ;
  assign n10459 = ( n10456 & ~n10458 ) | ( n10456 & n10457 ) | ( ~n10458 & n10457 ) ;
  assign n10463 = n10037 &  n10269 ;
  assign n10464 = n10268 &  n10463 ;
  assign n10452 = x74 | n10037 ;
  assign n10453 = x74 &  n10037 ;
  assign n10454 = ( n10452 & ~n10453 ) | ( n10452 & 1'b0 ) | ( ~n10453 & 1'b0 ) ;
  assign n10466 = ( n10121 & n10270 ) | ( n10121 & n10454 ) | ( n10270 & n10454 ) ;
  assign n10465 = n10121 | n10454 ;
  assign n10467 = ( n10464 & ~n10466 ) | ( n10464 & n10465 ) | ( ~n10466 & n10465 ) ;
  assign n10471 = n10045 &  n10269 ;
  assign n10472 = n10268 &  n10471 ;
  assign n10460 = x73 | n10045 ;
  assign n10461 = x73 &  n10045 ;
  assign n10462 = ( n10460 & ~n10461 ) | ( n10460 & 1'b0 ) | ( ~n10461 & 1'b0 ) ;
  assign n10474 = ( n10120 & n10270 ) | ( n10120 & n10462 ) | ( n10270 & n10462 ) ;
  assign n10473 = n10120 | n10462 ;
  assign n10475 = ( n10472 & ~n10474 ) | ( n10472 & n10473 ) | ( ~n10474 & n10473 ) ;
  assign n10479 = n10053 &  n10269 ;
  assign n10480 = n10268 &  n10479 ;
  assign n10468 = x72 | n10053 ;
  assign n10469 = x72 &  n10053 ;
  assign n10470 = ( n10468 & ~n10469 ) | ( n10468 & 1'b0 ) | ( ~n10469 & 1'b0 ) ;
  assign n10482 = ( n10119 & n10270 ) | ( n10119 & n10470 ) | ( n10270 & n10470 ) ;
  assign n10481 = n10119 | n10470 ;
  assign n10483 = ( n10480 & ~n10482 ) | ( n10480 & n10481 ) | ( ~n10482 & n10481 ) ;
  assign n10487 = n10061 &  n10269 ;
  assign n10488 = n10268 &  n10487 ;
  assign n10476 = x71 | n10061 ;
  assign n10477 = x71 &  n10061 ;
  assign n10478 = ( n10476 & ~n10477 ) | ( n10476 & 1'b0 ) | ( ~n10477 & 1'b0 ) ;
  assign n10490 = ( n10118 & n10270 ) | ( n10118 & n10478 ) | ( n10270 & n10478 ) ;
  assign n10489 = n10118 | n10478 ;
  assign n10491 = ( n10488 & ~n10490 ) | ( n10488 & n10489 ) | ( ~n10490 & n10489 ) ;
  assign n10495 = n10069 &  n10269 ;
  assign n10496 = n10268 &  n10495 ;
  assign n10484 = x70 | n10069 ;
  assign n10485 = x70 &  n10069 ;
  assign n10486 = ( n10484 & ~n10485 ) | ( n10484 & 1'b0 ) | ( ~n10485 & 1'b0 ) ;
  assign n10498 = ( n10117 & n10270 ) | ( n10117 & n10486 ) | ( n10270 & n10486 ) ;
  assign n10497 = n10117 | n10486 ;
  assign n10499 = ( n10496 & ~n10498 ) | ( n10496 & n10497 ) | ( ~n10498 & n10497 ) ;
  assign n10503 = n10077 &  n10269 ;
  assign n10504 = n10268 &  n10503 ;
  assign n10492 = x69 | n10077 ;
  assign n10493 = x69 &  n10077 ;
  assign n10494 = ( n10492 & ~n10493 ) | ( n10492 & 1'b0 ) | ( ~n10493 & 1'b0 ) ;
  assign n10506 = ( n10116 & n10270 ) | ( n10116 & n10494 ) | ( n10270 & n10494 ) ;
  assign n10505 = n10116 | n10494 ;
  assign n10507 = ( n10504 & ~n10506 ) | ( n10504 & n10505 ) | ( ~n10506 & n10505 ) ;
  assign n10511 = n10085 &  n10269 ;
  assign n10512 = n10268 &  n10511 ;
  assign n10500 = x68 | n10085 ;
  assign n10501 = x68 &  n10085 ;
  assign n10502 = ( n10500 & ~n10501 ) | ( n10500 & 1'b0 ) | ( ~n10501 & 1'b0 ) ;
  assign n10514 = ( n10115 & n10270 ) | ( n10115 & n10502 ) | ( n10270 & n10502 ) ;
  assign n10513 = n10115 | n10502 ;
  assign n10515 = ( n10512 & ~n10514 ) | ( n10512 & n10513 ) | ( ~n10514 & n10513 ) ;
  assign n10519 = n10094 &  n10269 ;
  assign n10520 = n10268 &  n10519 ;
  assign n10508 = x67 | n10094 ;
  assign n10509 = x67 &  n10094 ;
  assign n10510 = ( n10508 & ~n10509 ) | ( n10508 & 1'b0 ) | ( ~n10509 & 1'b0 ) ;
  assign n10522 = ( n10114 & n10270 ) | ( n10114 & n10510 ) | ( n10270 & n10510 ) ;
  assign n10521 = n10114 | n10510 ;
  assign n10523 = ( n10520 & ~n10522 ) | ( n10520 & n10521 ) | ( ~n10522 & n10521 ) ;
  assign n10524 = n10100 &  n10269 ;
  assign n10525 = n10268 &  n10524 ;
  assign n10516 = x66 | n10100 ;
  assign n10517 = x66 &  n10100 ;
  assign n10518 = ( n10516 & ~n10517 ) | ( n10516 & 1'b0 ) | ( ~n10517 & 1'b0 ) ;
  assign n10526 = n10113 &  n10518 ;
  assign n10527 = ( n10113 & ~n10270 ) | ( n10113 & n10518 ) | ( ~n10270 & n10518 ) ;
  assign n10528 = ( n10525 & ~n10526 ) | ( n10525 & n10527 ) | ( ~n10526 & n10527 ) ;
  assign n10529 = ( n10111 & ~x65 ) | ( n10111 & n10112 ) | ( ~x65 & n10112 ) ;
  assign n10530 = ( n10113 & ~n10112 ) | ( n10113 & n10529 ) | ( ~n10112 & n10529 ) ;
  assign n10531 = ~n10270 & n10530 ;
  assign n10532 = n10111 &  n10269 ;
  assign n10533 = n10268 &  n10532 ;
  assign n10534 = n10531 | n10533 ;
  assign n10535 = ( x64 & ~n10270 ) | ( x64 & 1'b0 ) | ( ~n10270 & 1'b0 ) ;
  assign n10536 = ( x17 & ~n10535 ) | ( x17 & 1'b0 ) | ( ~n10535 & 1'b0 ) ;
  assign n10537 = ( n10112 & ~n10270 ) | ( n10112 & 1'b0 ) | ( ~n10270 & 1'b0 ) ;
  assign n10538 = n10536 | n10537 ;
  assign n10539 = ~x16 & x64 ;
  assign n10540 = ( x65 & ~n10538 ) | ( x65 & n10539 ) | ( ~n10538 & n10539 ) ;
  assign n10541 = ( x66 & ~n10534 ) | ( x66 & n10540 ) | ( ~n10534 & n10540 ) ;
  assign n10542 = ( x67 & ~n10528 ) | ( x67 & n10541 ) | ( ~n10528 & n10541 ) ;
  assign n10543 = ( x68 & ~n10523 ) | ( x68 & n10542 ) | ( ~n10523 & n10542 ) ;
  assign n10544 = ( x69 & ~n10515 ) | ( x69 & n10543 ) | ( ~n10515 & n10543 ) ;
  assign n10545 = ( x70 & ~n10507 ) | ( x70 & n10544 ) | ( ~n10507 & n10544 ) ;
  assign n10546 = ( x71 & ~n10499 ) | ( x71 & n10545 ) | ( ~n10499 & n10545 ) ;
  assign n10547 = ( x72 & ~n10491 ) | ( x72 & n10546 ) | ( ~n10491 & n10546 ) ;
  assign n10548 = ( x73 & ~n10483 ) | ( x73 & n10547 ) | ( ~n10483 & n10547 ) ;
  assign n10549 = ( x74 & ~n10475 ) | ( x74 & n10548 ) | ( ~n10475 & n10548 ) ;
  assign n10550 = ( x75 & ~n10467 ) | ( x75 & n10549 ) | ( ~n10467 & n10549 ) ;
  assign n10551 = ( x76 & ~n10459 ) | ( x76 & n10550 ) | ( ~n10459 & n10550 ) ;
  assign n10552 = ( x77 & ~n10451 ) | ( x77 & n10551 ) | ( ~n10451 & n10551 ) ;
  assign n10553 = ( x78 & ~n10443 ) | ( x78 & n10552 ) | ( ~n10443 & n10552 ) ;
  assign n10554 = ( x79 & ~n10435 ) | ( x79 & n10553 ) | ( ~n10435 & n10553 ) ;
  assign n10555 = ( x80 & ~n10427 ) | ( x80 & n10554 ) | ( ~n10427 & n10554 ) ;
  assign n10556 = ( x81 & ~n10419 ) | ( x81 & n10555 ) | ( ~n10419 & n10555 ) ;
  assign n10557 = ( x82 & ~n10411 ) | ( x82 & n10556 ) | ( ~n10411 & n10556 ) ;
  assign n10558 = ( x83 & ~n10403 ) | ( x83 & n10557 ) | ( ~n10403 & n10557 ) ;
  assign n10559 = ( x84 & ~n10395 ) | ( x84 & n10558 ) | ( ~n10395 & n10558 ) ;
  assign n10560 = ( x85 & ~n10387 ) | ( x85 & n10559 ) | ( ~n10387 & n10559 ) ;
  assign n10561 = ( x86 & ~n10379 ) | ( x86 & n10560 ) | ( ~n10379 & n10560 ) ;
  assign n10562 = ( x87 & ~n10371 ) | ( x87 & n10561 ) | ( ~n10371 & n10561 ) ;
  assign n10563 = ( x88 & ~n10363 ) | ( x88 & n10562 ) | ( ~n10363 & n10562 ) ;
  assign n10564 = ( x89 & ~n10355 ) | ( x89 & n10563 ) | ( ~n10355 & n10563 ) ;
  assign n10565 = ( x90 & ~n10347 ) | ( x90 & n10564 ) | ( ~n10347 & n10564 ) ;
  assign n10566 = ( x91 & ~n10339 ) | ( x91 & n10565 ) | ( ~n10339 & n10565 ) ;
  assign n10567 = ( x92 & ~n10331 ) | ( x92 & n10566 ) | ( ~n10331 & n10566 ) ;
  assign n10568 = ( x93 & ~n10323 ) | ( x93 & n10567 ) | ( ~n10323 & n10567 ) ;
  assign n10569 = ( x94 & ~n10315 ) | ( x94 & n10568 ) | ( ~n10315 & n10568 ) ;
  assign n10570 = ( x95 & ~n10307 ) | ( x95 & n10569 ) | ( ~n10307 & n10569 ) ;
  assign n10571 = ( x96 & ~n10299 ) | ( x96 & n10570 ) | ( ~n10299 & n10570 ) ;
  assign n10572 = ( x97 & ~n10291 ) | ( x97 & n10571 ) | ( ~n10291 & n10571 ) ;
  assign n10573 = ( x98 & ~n10283 ) | ( x98 & n10572 ) | ( ~n10283 & n10572 ) ;
  assign n10577 = ( x99 & ~n10275 ) | ( x99 & n10573 ) | ( ~n10275 & n10573 ) ;
  assign n10669 = ( x100 & ~n10585 ) | ( x100 & n10577 ) | ( ~n10585 & n10577 ) ;
  assign n10670 = ( x101 & ~n10668 ) | ( x101 & n10669 ) | ( ~n10668 & n10669 ) ;
  assign n10671 = ( x102 & ~n10663 ) | ( x102 & n10670 ) | ( ~n10663 & n10670 ) ;
  assign n10672 = ( x103 & ~n10655 ) | ( x103 & n10671 ) | ( ~n10655 & n10671 ) ;
  assign n10673 = ( x104 & ~n10647 ) | ( x104 & n10672 ) | ( ~n10647 & n10672 ) ;
  assign n10674 = ( x105 & ~n10639 ) | ( x105 & n10673 ) | ( ~n10639 & n10673 ) ;
  assign n10675 = ( x106 & ~n10631 ) | ( x106 & n10674 ) | ( ~n10631 & n10674 ) ;
  assign n10676 = ( x107 & ~n10623 ) | ( x107 & n10675 ) | ( ~n10623 & n10675 ) ;
  assign n10677 = ( x108 & ~n10615 ) | ( x108 & n10676 ) | ( ~n10615 & n10676 ) ;
  assign n10678 = ( x109 & ~n10607 ) | ( x109 & n10677 ) | ( ~n10607 & n10677 ) ;
  assign n10679 = ( x110 & ~n10599 ) | ( x110 & n10678 ) | ( ~n10599 & n10678 ) ;
  assign n10681 = ( x110 & n10259 ) | ( x110 & n10262 ) | ( n10259 & n10262 ) ;
  assign n10680 = ( x110 & ~n10259 ) | ( x110 & n10262 ) | ( ~n10259 & n10262 ) ;
  assign n10682 = ( n10259 & ~n10681 ) | ( n10259 & n10680 ) | ( ~n10681 & n10680 ) ;
  assign n10683 = ~n10270 & n10682 ;
  assign n10684 = n9461 &  n9841 ;
  assign n10685 = n10268 &  n10684 ;
  assign n10686 = n10683 | n10685 ;
  assign n10687 = ~x111 & n10686 ;
  assign n10688 = ( x111 & ~n10685 ) | ( x111 & 1'b0 ) | ( ~n10685 & 1'b0 ) ;
  assign n10689 = ~n10683 & n10688 ;
  assign n10690 = n270 | n10689 ;
  assign n10691 = n10687 | n10690 ;
  assign n10692 = n10679 | n10691 ;
  assign n10693 = ~n10686 |  n10264 ;
  assign n10712 = n10599 &  n10693 ;
  assign n10713 = n10692 &  n10712 ;
  assign n10700 = x110 | n10599 ;
  assign n10701 = x110 &  n10599 ;
  assign n10702 = ( n10700 & ~n10701 ) | ( n10700 & 1'b0 ) | ( ~n10701 & 1'b0 ) ;
  assign n10714 = n10678 &  n10702 ;
  assign n10694 = n10692 &  n10693 ;
  assign n10715 = ( n10678 & ~n10694 ) | ( n10678 & n10702 ) | ( ~n10694 & n10702 ) ;
  assign n10716 = ( n10713 & ~n10714 ) | ( n10713 & n10715 ) | ( ~n10714 & n10715 ) ;
  assign n10704 = n10264 &  n10686 ;
  assign n10705 = n10692 &  n10704 ;
  assign n10703 = n10687 | n10689 ;
  assign n10707 = ( n10679 & n10694 ) | ( n10679 & n10703 ) | ( n10694 & n10703 ) ;
  assign n10706 = n10679 | n10703 ;
  assign n10708 = ( n10705 & ~n10707 ) | ( n10705 & n10706 ) | ( ~n10707 & n10706 ) ;
  assign n10720 = n10607 &  n10693 ;
  assign n10721 = n10692 &  n10720 ;
  assign n10709 = x109 | n10607 ;
  assign n10710 = x109 &  n10607 ;
  assign n10711 = ( n10709 & ~n10710 ) | ( n10709 & 1'b0 ) | ( ~n10710 & 1'b0 ) ;
  assign n10722 = n10677 &  n10711 ;
  assign n10723 = ( n10677 & ~n10694 ) | ( n10677 & n10711 ) | ( ~n10694 & n10711 ) ;
  assign n10724 = ( n10721 & ~n10722 ) | ( n10721 & n10723 ) | ( ~n10722 & n10723 ) ;
  assign n10728 = n10615 &  n10693 ;
  assign n10729 = n10692 &  n10728 ;
  assign n10717 = x108 | n10615 ;
  assign n10718 = x108 &  n10615 ;
  assign n10719 = ( n10717 & ~n10718 ) | ( n10717 & 1'b0 ) | ( ~n10718 & 1'b0 ) ;
  assign n10730 = n10676 &  n10719 ;
  assign n10731 = ( n10676 & ~n10694 ) | ( n10676 & n10719 ) | ( ~n10694 & n10719 ) ;
  assign n10732 = ( n10729 & ~n10730 ) | ( n10729 & n10731 ) | ( ~n10730 & n10731 ) ;
  assign n10736 = n10623 &  n10693 ;
  assign n10737 = n10692 &  n10736 ;
  assign n10725 = x107 | n10623 ;
  assign n10726 = x107 &  n10623 ;
  assign n10727 = ( n10725 & ~n10726 ) | ( n10725 & 1'b0 ) | ( ~n10726 & 1'b0 ) ;
  assign n10738 = n10675 &  n10727 ;
  assign n10739 = ( n10675 & ~n10694 ) | ( n10675 & n10727 ) | ( ~n10694 & n10727 ) ;
  assign n10740 = ( n10737 & ~n10738 ) | ( n10737 & n10739 ) | ( ~n10738 & n10739 ) ;
  assign n10744 = n10631 &  n10693 ;
  assign n10745 = n10692 &  n10744 ;
  assign n10733 = x106 | n10631 ;
  assign n10734 = x106 &  n10631 ;
  assign n10735 = ( n10733 & ~n10734 ) | ( n10733 & 1'b0 ) | ( ~n10734 & 1'b0 ) ;
  assign n10746 = n10674 &  n10735 ;
  assign n10747 = ( n10674 & ~n10694 ) | ( n10674 & n10735 ) | ( ~n10694 & n10735 ) ;
  assign n10748 = ( n10745 & ~n10746 ) | ( n10745 & n10747 ) | ( ~n10746 & n10747 ) ;
  assign n10752 = n10639 &  n10693 ;
  assign n10753 = n10692 &  n10752 ;
  assign n10741 = x105 | n10639 ;
  assign n10742 = x105 &  n10639 ;
  assign n10743 = ( n10741 & ~n10742 ) | ( n10741 & 1'b0 ) | ( ~n10742 & 1'b0 ) ;
  assign n10755 = ( n10673 & n10694 ) | ( n10673 & n10743 ) | ( n10694 & n10743 ) ;
  assign n10754 = n10673 | n10743 ;
  assign n10756 = ( n10753 & ~n10755 ) | ( n10753 & n10754 ) | ( ~n10755 & n10754 ) ;
  assign n10760 = n10647 &  n10693 ;
  assign n10761 = n10692 &  n10760 ;
  assign n10749 = x104 | n10647 ;
  assign n10750 = x104 &  n10647 ;
  assign n10751 = ( n10749 & ~n10750 ) | ( n10749 & 1'b0 ) | ( ~n10750 & 1'b0 ) ;
  assign n10763 = ( n10672 & n10694 ) | ( n10672 & n10751 ) | ( n10694 & n10751 ) ;
  assign n10762 = n10672 | n10751 ;
  assign n10764 = ( n10761 & ~n10763 ) | ( n10761 & n10762 ) | ( ~n10763 & n10762 ) ;
  assign n10768 = n10655 &  n10693 ;
  assign n10769 = n10692 &  n10768 ;
  assign n10757 = x103 | n10655 ;
  assign n10758 = x103 &  n10655 ;
  assign n10759 = ( n10757 & ~n10758 ) | ( n10757 & 1'b0 ) | ( ~n10758 & 1'b0 ) ;
  assign n10771 = ( n10671 & n10694 ) | ( n10671 & n10759 ) | ( n10694 & n10759 ) ;
  assign n10770 = n10671 | n10759 ;
  assign n10772 = ( n10769 & ~n10771 ) | ( n10769 & n10770 ) | ( ~n10771 & n10770 ) ;
  assign n10776 = n10663 &  n10693 ;
  assign n10777 = n10692 &  n10776 ;
  assign n10765 = x102 | n10663 ;
  assign n10766 = x102 &  n10663 ;
  assign n10767 = ( n10765 & ~n10766 ) | ( n10765 & 1'b0 ) | ( ~n10766 & 1'b0 ) ;
  assign n10779 = ( n10670 & n10694 ) | ( n10670 & n10767 ) | ( n10694 & n10767 ) ;
  assign n10778 = n10670 | n10767 ;
  assign n10780 = ( n10777 & ~n10779 ) | ( n10777 & n10778 ) | ( ~n10779 & n10778 ) ;
  assign n10781 = n10668 &  n10693 ;
  assign n10782 = n10692 &  n10781 ;
  assign n10773 = x101 | n10668 ;
  assign n10774 = x101 &  n10668 ;
  assign n10775 = ( n10773 & ~n10774 ) | ( n10773 & 1'b0 ) | ( ~n10774 & 1'b0 ) ;
  assign n10784 = ( n10669 & n10694 ) | ( n10669 & n10775 ) | ( n10694 & n10775 ) ;
  assign n10783 = n10669 | n10775 ;
  assign n10785 = ( n10782 & ~n10784 ) | ( n10782 & n10783 ) | ( ~n10784 & n10783 ) ;
  assign n10695 = n10585 &  n10693 ;
  assign n10696 = n10692 &  n10695 ;
  assign n10586 = x100 | n10585 ;
  assign n10587 = x100 &  n10585 ;
  assign n10588 = ( n10586 & ~n10587 ) | ( n10586 & 1'b0 ) | ( ~n10587 & 1'b0 ) ;
  assign n10698 = ( n10577 & n10588 ) | ( n10577 & n10694 ) | ( n10588 & n10694 ) ;
  assign n10697 = n10577 | n10588 ;
  assign n10699 = ( n10696 & ~n10698 ) | ( n10696 & n10697 ) | ( ~n10698 & n10697 ) ;
  assign n10789 = n10275 &  n10693 ;
  assign n10790 = n10692 &  n10789 ;
  assign n10574 = x99 | n10275 ;
  assign n10575 = x99 &  n10275 ;
  assign n10576 = ( n10574 & ~n10575 ) | ( n10574 & 1'b0 ) | ( ~n10575 & 1'b0 ) ;
  assign n10791 = n10573 &  n10576 ;
  assign n10792 = ( n10573 & ~n10694 ) | ( n10573 & n10576 ) | ( ~n10694 & n10576 ) ;
  assign n10793 = ( n10790 & ~n10791 ) | ( n10790 & n10792 ) | ( ~n10791 & n10792 ) ;
  assign n10797 = n10283 &  n10693 ;
  assign n10798 = n10692 &  n10797 ;
  assign n10786 = x98 | n10283 ;
  assign n10787 = x98 &  n10283 ;
  assign n10788 = ( n10786 & ~n10787 ) | ( n10786 & 1'b0 ) | ( ~n10787 & 1'b0 ) ;
  assign n10800 = ( n10572 & n10694 ) | ( n10572 & n10788 ) | ( n10694 & n10788 ) ;
  assign n10799 = n10572 | n10788 ;
  assign n10801 = ( n10798 & ~n10800 ) | ( n10798 & n10799 ) | ( ~n10800 & n10799 ) ;
  assign n10805 = n10291 &  n10693 ;
  assign n10806 = n10692 &  n10805 ;
  assign n10794 = x97 | n10291 ;
  assign n10795 = x97 &  n10291 ;
  assign n10796 = ( n10794 & ~n10795 ) | ( n10794 & 1'b0 ) | ( ~n10795 & 1'b0 ) ;
  assign n10808 = ( n10571 & n10694 ) | ( n10571 & n10796 ) | ( n10694 & n10796 ) ;
  assign n10807 = n10571 | n10796 ;
  assign n10809 = ( n10806 & ~n10808 ) | ( n10806 & n10807 ) | ( ~n10808 & n10807 ) ;
  assign n10813 = n10299 &  n10693 ;
  assign n10814 = n10692 &  n10813 ;
  assign n10802 = x96 | n10299 ;
  assign n10803 = x96 &  n10299 ;
  assign n10804 = ( n10802 & ~n10803 ) | ( n10802 & 1'b0 ) | ( ~n10803 & 1'b0 ) ;
  assign n10816 = ( n10570 & n10694 ) | ( n10570 & n10804 ) | ( n10694 & n10804 ) ;
  assign n10815 = n10570 | n10804 ;
  assign n10817 = ( n10814 & ~n10816 ) | ( n10814 & n10815 ) | ( ~n10816 & n10815 ) ;
  assign n10821 = n10307 &  n10693 ;
  assign n10822 = n10692 &  n10821 ;
  assign n10810 = x95 | n10307 ;
  assign n10811 = x95 &  n10307 ;
  assign n10812 = ( n10810 & ~n10811 ) | ( n10810 & 1'b0 ) | ( ~n10811 & 1'b0 ) ;
  assign n10824 = ( n10569 & n10694 ) | ( n10569 & n10812 ) | ( n10694 & n10812 ) ;
  assign n10823 = n10569 | n10812 ;
  assign n10825 = ( n10822 & ~n10824 ) | ( n10822 & n10823 ) | ( ~n10824 & n10823 ) ;
  assign n10829 = n10315 &  n10693 ;
  assign n10830 = n10692 &  n10829 ;
  assign n10818 = x94 | n10315 ;
  assign n10819 = x94 &  n10315 ;
  assign n10820 = ( n10818 & ~n10819 ) | ( n10818 & 1'b0 ) | ( ~n10819 & 1'b0 ) ;
  assign n10832 = ( n10568 & n10694 ) | ( n10568 & n10820 ) | ( n10694 & n10820 ) ;
  assign n10831 = n10568 | n10820 ;
  assign n10833 = ( n10830 & ~n10832 ) | ( n10830 & n10831 ) | ( ~n10832 & n10831 ) ;
  assign n10837 = n10323 &  n10693 ;
  assign n10838 = n10692 &  n10837 ;
  assign n10826 = x93 | n10323 ;
  assign n10827 = x93 &  n10323 ;
  assign n10828 = ( n10826 & ~n10827 ) | ( n10826 & 1'b0 ) | ( ~n10827 & 1'b0 ) ;
  assign n10840 = ( n10567 & n10694 ) | ( n10567 & n10828 ) | ( n10694 & n10828 ) ;
  assign n10839 = n10567 | n10828 ;
  assign n10841 = ( n10838 & ~n10840 ) | ( n10838 & n10839 ) | ( ~n10840 & n10839 ) ;
  assign n10845 = n10331 &  n10693 ;
  assign n10846 = n10692 &  n10845 ;
  assign n10834 = x92 | n10331 ;
  assign n10835 = x92 &  n10331 ;
  assign n10836 = ( n10834 & ~n10835 ) | ( n10834 & 1'b0 ) | ( ~n10835 & 1'b0 ) ;
  assign n10848 = ( n10566 & n10694 ) | ( n10566 & n10836 ) | ( n10694 & n10836 ) ;
  assign n10847 = n10566 | n10836 ;
  assign n10849 = ( n10846 & ~n10848 ) | ( n10846 & n10847 ) | ( ~n10848 & n10847 ) ;
  assign n10853 = n10339 &  n10693 ;
  assign n10854 = n10692 &  n10853 ;
  assign n10842 = x91 | n10339 ;
  assign n10843 = x91 &  n10339 ;
  assign n10844 = ( n10842 & ~n10843 ) | ( n10842 & 1'b0 ) | ( ~n10843 & 1'b0 ) ;
  assign n10856 = ( n10565 & n10694 ) | ( n10565 & n10844 ) | ( n10694 & n10844 ) ;
  assign n10855 = n10565 | n10844 ;
  assign n10857 = ( n10854 & ~n10856 ) | ( n10854 & n10855 ) | ( ~n10856 & n10855 ) ;
  assign n10861 = n10347 &  n10693 ;
  assign n10862 = n10692 &  n10861 ;
  assign n10850 = x90 | n10347 ;
  assign n10851 = x90 &  n10347 ;
  assign n10852 = ( n10850 & ~n10851 ) | ( n10850 & 1'b0 ) | ( ~n10851 & 1'b0 ) ;
  assign n10864 = ( n10564 & n10694 ) | ( n10564 & n10852 ) | ( n10694 & n10852 ) ;
  assign n10863 = n10564 | n10852 ;
  assign n10865 = ( n10862 & ~n10864 ) | ( n10862 & n10863 ) | ( ~n10864 & n10863 ) ;
  assign n10869 = n10355 &  n10693 ;
  assign n10870 = n10692 &  n10869 ;
  assign n10858 = x89 | n10355 ;
  assign n10859 = x89 &  n10355 ;
  assign n10860 = ( n10858 & ~n10859 ) | ( n10858 & 1'b0 ) | ( ~n10859 & 1'b0 ) ;
  assign n10872 = ( n10563 & n10694 ) | ( n10563 & n10860 ) | ( n10694 & n10860 ) ;
  assign n10871 = n10563 | n10860 ;
  assign n10873 = ( n10870 & ~n10872 ) | ( n10870 & n10871 ) | ( ~n10872 & n10871 ) ;
  assign n10877 = n10363 &  n10693 ;
  assign n10878 = n10692 &  n10877 ;
  assign n10866 = x88 | n10363 ;
  assign n10867 = x88 &  n10363 ;
  assign n10868 = ( n10866 & ~n10867 ) | ( n10866 & 1'b0 ) | ( ~n10867 & 1'b0 ) ;
  assign n10880 = ( n10562 & n10694 ) | ( n10562 & n10868 ) | ( n10694 & n10868 ) ;
  assign n10879 = n10562 | n10868 ;
  assign n10881 = ( n10878 & ~n10880 ) | ( n10878 & n10879 ) | ( ~n10880 & n10879 ) ;
  assign n10885 = n10371 &  n10693 ;
  assign n10886 = n10692 &  n10885 ;
  assign n10874 = x87 | n10371 ;
  assign n10875 = x87 &  n10371 ;
  assign n10876 = ( n10874 & ~n10875 ) | ( n10874 & 1'b0 ) | ( ~n10875 & 1'b0 ) ;
  assign n10888 = ( n10561 & n10694 ) | ( n10561 & n10876 ) | ( n10694 & n10876 ) ;
  assign n10887 = n10561 | n10876 ;
  assign n10889 = ( n10886 & ~n10888 ) | ( n10886 & n10887 ) | ( ~n10888 & n10887 ) ;
  assign n10893 = n10379 &  n10693 ;
  assign n10894 = n10692 &  n10893 ;
  assign n10882 = x86 | n10379 ;
  assign n10883 = x86 &  n10379 ;
  assign n10884 = ( n10882 & ~n10883 ) | ( n10882 & 1'b0 ) | ( ~n10883 & 1'b0 ) ;
  assign n10896 = ( n10560 & n10694 ) | ( n10560 & n10884 ) | ( n10694 & n10884 ) ;
  assign n10895 = n10560 | n10884 ;
  assign n10897 = ( n10894 & ~n10896 ) | ( n10894 & n10895 ) | ( ~n10896 & n10895 ) ;
  assign n10901 = n10387 &  n10693 ;
  assign n10902 = n10692 &  n10901 ;
  assign n10890 = x85 | n10387 ;
  assign n10891 = x85 &  n10387 ;
  assign n10892 = ( n10890 & ~n10891 ) | ( n10890 & 1'b0 ) | ( ~n10891 & 1'b0 ) ;
  assign n10904 = ( n10559 & n10694 ) | ( n10559 & n10892 ) | ( n10694 & n10892 ) ;
  assign n10903 = n10559 | n10892 ;
  assign n10905 = ( n10902 & ~n10904 ) | ( n10902 & n10903 ) | ( ~n10904 & n10903 ) ;
  assign n10909 = n10395 &  n10693 ;
  assign n10910 = n10692 &  n10909 ;
  assign n10898 = x84 | n10395 ;
  assign n10899 = x84 &  n10395 ;
  assign n10900 = ( n10898 & ~n10899 ) | ( n10898 & 1'b0 ) | ( ~n10899 & 1'b0 ) ;
  assign n10912 = ( n10558 & n10694 ) | ( n10558 & n10900 ) | ( n10694 & n10900 ) ;
  assign n10911 = n10558 | n10900 ;
  assign n10913 = ( n10910 & ~n10912 ) | ( n10910 & n10911 ) | ( ~n10912 & n10911 ) ;
  assign n10917 = n10403 &  n10693 ;
  assign n10918 = n10692 &  n10917 ;
  assign n10906 = x83 | n10403 ;
  assign n10907 = x83 &  n10403 ;
  assign n10908 = ( n10906 & ~n10907 ) | ( n10906 & 1'b0 ) | ( ~n10907 & 1'b0 ) ;
  assign n10920 = ( n10557 & n10694 ) | ( n10557 & n10908 ) | ( n10694 & n10908 ) ;
  assign n10919 = n10557 | n10908 ;
  assign n10921 = ( n10918 & ~n10920 ) | ( n10918 & n10919 ) | ( ~n10920 & n10919 ) ;
  assign n10925 = n10411 &  n10693 ;
  assign n10926 = n10692 &  n10925 ;
  assign n10914 = x82 | n10411 ;
  assign n10915 = x82 &  n10411 ;
  assign n10916 = ( n10914 & ~n10915 ) | ( n10914 & 1'b0 ) | ( ~n10915 & 1'b0 ) ;
  assign n10928 = ( n10556 & n10694 ) | ( n10556 & n10916 ) | ( n10694 & n10916 ) ;
  assign n10927 = n10556 | n10916 ;
  assign n10929 = ( n10926 & ~n10928 ) | ( n10926 & n10927 ) | ( ~n10928 & n10927 ) ;
  assign n10933 = n10419 &  n10693 ;
  assign n10934 = n10692 &  n10933 ;
  assign n10922 = x81 | n10419 ;
  assign n10923 = x81 &  n10419 ;
  assign n10924 = ( n10922 & ~n10923 ) | ( n10922 & 1'b0 ) | ( ~n10923 & 1'b0 ) ;
  assign n10936 = ( n10555 & n10694 ) | ( n10555 & n10924 ) | ( n10694 & n10924 ) ;
  assign n10935 = n10555 | n10924 ;
  assign n10937 = ( n10934 & ~n10936 ) | ( n10934 & n10935 ) | ( ~n10936 & n10935 ) ;
  assign n10941 = n10427 &  n10693 ;
  assign n10942 = n10692 &  n10941 ;
  assign n10930 = x80 | n10427 ;
  assign n10931 = x80 &  n10427 ;
  assign n10932 = ( n10930 & ~n10931 ) | ( n10930 & 1'b0 ) | ( ~n10931 & 1'b0 ) ;
  assign n10944 = ( n10554 & n10694 ) | ( n10554 & n10932 ) | ( n10694 & n10932 ) ;
  assign n10943 = n10554 | n10932 ;
  assign n10945 = ( n10942 & ~n10944 ) | ( n10942 & n10943 ) | ( ~n10944 & n10943 ) ;
  assign n10949 = n10435 &  n10693 ;
  assign n10950 = n10692 &  n10949 ;
  assign n10938 = x79 | n10435 ;
  assign n10939 = x79 &  n10435 ;
  assign n10940 = ( n10938 & ~n10939 ) | ( n10938 & 1'b0 ) | ( ~n10939 & 1'b0 ) ;
  assign n10952 = ( n10553 & n10694 ) | ( n10553 & n10940 ) | ( n10694 & n10940 ) ;
  assign n10951 = n10553 | n10940 ;
  assign n10953 = ( n10950 & ~n10952 ) | ( n10950 & n10951 ) | ( ~n10952 & n10951 ) ;
  assign n10957 = n10443 &  n10693 ;
  assign n10958 = n10692 &  n10957 ;
  assign n10946 = x78 | n10443 ;
  assign n10947 = x78 &  n10443 ;
  assign n10948 = ( n10946 & ~n10947 ) | ( n10946 & 1'b0 ) | ( ~n10947 & 1'b0 ) ;
  assign n10960 = ( n10552 & n10694 ) | ( n10552 & n10948 ) | ( n10694 & n10948 ) ;
  assign n10959 = n10552 | n10948 ;
  assign n10961 = ( n10958 & ~n10960 ) | ( n10958 & n10959 ) | ( ~n10960 & n10959 ) ;
  assign n10965 = n10451 &  n10693 ;
  assign n10966 = n10692 &  n10965 ;
  assign n10954 = x77 | n10451 ;
  assign n10955 = x77 &  n10451 ;
  assign n10956 = ( n10954 & ~n10955 ) | ( n10954 & 1'b0 ) | ( ~n10955 & 1'b0 ) ;
  assign n10968 = ( n10551 & n10694 ) | ( n10551 & n10956 ) | ( n10694 & n10956 ) ;
  assign n10967 = n10551 | n10956 ;
  assign n10969 = ( n10966 & ~n10968 ) | ( n10966 & n10967 ) | ( ~n10968 & n10967 ) ;
  assign n10973 = n10459 &  n10693 ;
  assign n10974 = n10692 &  n10973 ;
  assign n10962 = x76 | n10459 ;
  assign n10963 = x76 &  n10459 ;
  assign n10964 = ( n10962 & ~n10963 ) | ( n10962 & 1'b0 ) | ( ~n10963 & 1'b0 ) ;
  assign n10976 = ( n10550 & n10694 ) | ( n10550 & n10964 ) | ( n10694 & n10964 ) ;
  assign n10975 = n10550 | n10964 ;
  assign n10977 = ( n10974 & ~n10976 ) | ( n10974 & n10975 ) | ( ~n10976 & n10975 ) ;
  assign n10981 = n10467 &  n10693 ;
  assign n10982 = n10692 &  n10981 ;
  assign n10970 = x75 | n10467 ;
  assign n10971 = x75 &  n10467 ;
  assign n10972 = ( n10970 & ~n10971 ) | ( n10970 & 1'b0 ) | ( ~n10971 & 1'b0 ) ;
  assign n10984 = ( n10549 & n10694 ) | ( n10549 & n10972 ) | ( n10694 & n10972 ) ;
  assign n10983 = n10549 | n10972 ;
  assign n10985 = ( n10982 & ~n10984 ) | ( n10982 & n10983 ) | ( ~n10984 & n10983 ) ;
  assign n10989 = n10475 &  n10693 ;
  assign n10990 = n10692 &  n10989 ;
  assign n10978 = x74 | n10475 ;
  assign n10979 = x74 &  n10475 ;
  assign n10980 = ( n10978 & ~n10979 ) | ( n10978 & 1'b0 ) | ( ~n10979 & 1'b0 ) ;
  assign n10992 = ( n10548 & n10694 ) | ( n10548 & n10980 ) | ( n10694 & n10980 ) ;
  assign n10991 = n10548 | n10980 ;
  assign n10993 = ( n10990 & ~n10992 ) | ( n10990 & n10991 ) | ( ~n10992 & n10991 ) ;
  assign n10997 = n10483 &  n10693 ;
  assign n10998 = n10692 &  n10997 ;
  assign n10986 = x73 | n10483 ;
  assign n10987 = x73 &  n10483 ;
  assign n10988 = ( n10986 & ~n10987 ) | ( n10986 & 1'b0 ) | ( ~n10987 & 1'b0 ) ;
  assign n11000 = ( n10547 & n10694 ) | ( n10547 & n10988 ) | ( n10694 & n10988 ) ;
  assign n10999 = n10547 | n10988 ;
  assign n11001 = ( n10998 & ~n11000 ) | ( n10998 & n10999 ) | ( ~n11000 & n10999 ) ;
  assign n11005 = n10491 &  n10693 ;
  assign n11006 = n10692 &  n11005 ;
  assign n10994 = x72 | n10491 ;
  assign n10995 = x72 &  n10491 ;
  assign n10996 = ( n10994 & ~n10995 ) | ( n10994 & 1'b0 ) | ( ~n10995 & 1'b0 ) ;
  assign n11008 = ( n10546 & n10694 ) | ( n10546 & n10996 ) | ( n10694 & n10996 ) ;
  assign n11007 = n10546 | n10996 ;
  assign n11009 = ( n11006 & ~n11008 ) | ( n11006 & n11007 ) | ( ~n11008 & n11007 ) ;
  assign n11013 = n10499 &  n10693 ;
  assign n11014 = n10692 &  n11013 ;
  assign n11002 = x71 | n10499 ;
  assign n11003 = x71 &  n10499 ;
  assign n11004 = ( n11002 & ~n11003 ) | ( n11002 & 1'b0 ) | ( ~n11003 & 1'b0 ) ;
  assign n11016 = ( n10545 & n10694 ) | ( n10545 & n11004 ) | ( n10694 & n11004 ) ;
  assign n11015 = n10545 | n11004 ;
  assign n11017 = ( n11014 & ~n11016 ) | ( n11014 & n11015 ) | ( ~n11016 & n11015 ) ;
  assign n11021 = n10507 &  n10693 ;
  assign n11022 = n10692 &  n11021 ;
  assign n11010 = x70 | n10507 ;
  assign n11011 = x70 &  n10507 ;
  assign n11012 = ( n11010 & ~n11011 ) | ( n11010 & 1'b0 ) | ( ~n11011 & 1'b0 ) ;
  assign n11024 = ( n10544 & n10694 ) | ( n10544 & n11012 ) | ( n10694 & n11012 ) ;
  assign n11023 = n10544 | n11012 ;
  assign n11025 = ( n11022 & ~n11024 ) | ( n11022 & n11023 ) | ( ~n11024 & n11023 ) ;
  assign n11029 = n10515 &  n10693 ;
  assign n11030 = n10692 &  n11029 ;
  assign n11018 = x69 | n10515 ;
  assign n11019 = x69 &  n10515 ;
  assign n11020 = ( n11018 & ~n11019 ) | ( n11018 & 1'b0 ) | ( ~n11019 & 1'b0 ) ;
  assign n11032 = ( n10543 & n10694 ) | ( n10543 & n11020 ) | ( n10694 & n11020 ) ;
  assign n11031 = n10543 | n11020 ;
  assign n11033 = ( n11030 & ~n11032 ) | ( n11030 & n11031 ) | ( ~n11032 & n11031 ) ;
  assign n11037 = n10523 &  n10693 ;
  assign n11038 = n10692 &  n11037 ;
  assign n11026 = x68 | n10523 ;
  assign n11027 = x68 &  n10523 ;
  assign n11028 = ( n11026 & ~n11027 ) | ( n11026 & 1'b0 ) | ( ~n11027 & 1'b0 ) ;
  assign n11040 = ( n10542 & n10694 ) | ( n10542 & n11028 ) | ( n10694 & n11028 ) ;
  assign n11039 = n10542 | n11028 ;
  assign n11041 = ( n11038 & ~n11040 ) | ( n11038 & n11039 ) | ( ~n11040 & n11039 ) ;
  assign n11045 = n10528 &  n10693 ;
  assign n11046 = n10692 &  n11045 ;
  assign n11034 = x67 | n10528 ;
  assign n11035 = x67 &  n10528 ;
  assign n11036 = ( n11034 & ~n11035 ) | ( n11034 & 1'b0 ) | ( ~n11035 & 1'b0 ) ;
  assign n11048 = ( n10541 & n10694 ) | ( n10541 & n11036 ) | ( n10694 & n11036 ) ;
  assign n11047 = n10541 | n11036 ;
  assign n11049 = ( n11046 & ~n11048 ) | ( n11046 & n11047 ) | ( ~n11048 & n11047 ) ;
  assign n11050 = n10534 &  n10693 ;
  assign n11051 = n10692 &  n11050 ;
  assign n11042 = x66 | n10534 ;
  assign n11043 = x66 &  n10534 ;
  assign n11044 = ( n11042 & ~n11043 ) | ( n11042 & 1'b0 ) | ( ~n11043 & 1'b0 ) ;
  assign n11052 = n10540 &  n11044 ;
  assign n11053 = ( n10540 & ~n10694 ) | ( n10540 & n11044 ) | ( ~n10694 & n11044 ) ;
  assign n11054 = ( n11051 & ~n11052 ) | ( n11051 & n11053 ) | ( ~n11052 & n11053 ) ;
  assign n11055 = ( n10538 & ~x65 ) | ( n10538 & n10539 ) | ( ~x65 & n10539 ) ;
  assign n11056 = ( n10540 & ~n10539 ) | ( n10540 & n11055 ) | ( ~n10539 & n11055 ) ;
  assign n11057 = ~n10694 & n11056 ;
  assign n11058 = n10538 &  n10693 ;
  assign n11059 = n10692 &  n11058 ;
  assign n11060 = n11057 | n11059 ;
  assign n11061 = ( x64 & ~n10694 ) | ( x64 & 1'b0 ) | ( ~n10694 & 1'b0 ) ;
  assign n11062 = ( x16 & ~n11061 ) | ( x16 & 1'b0 ) | ( ~n11061 & 1'b0 ) ;
  assign n11063 = ( n10539 & ~n10694 ) | ( n10539 & 1'b0 ) | ( ~n10694 & 1'b0 ) ;
  assign n11064 = n11062 | n11063 ;
  assign n11065 = ~x15 & x64 ;
  assign n11066 = ( x65 & ~n11064 ) | ( x65 & n11065 ) | ( ~n11064 & n11065 ) ;
  assign n11067 = ( x66 & ~n11060 ) | ( x66 & n11066 ) | ( ~n11060 & n11066 ) ;
  assign n11068 = ( x67 & ~n11054 ) | ( x67 & n11067 ) | ( ~n11054 & n11067 ) ;
  assign n11069 = ( x68 & ~n11049 ) | ( x68 & n11068 ) | ( ~n11049 & n11068 ) ;
  assign n11070 = ( x69 & ~n11041 ) | ( x69 & n11069 ) | ( ~n11041 & n11069 ) ;
  assign n11071 = ( x70 & ~n11033 ) | ( x70 & n11070 ) | ( ~n11033 & n11070 ) ;
  assign n11072 = ( x71 & ~n11025 ) | ( x71 & n11071 ) | ( ~n11025 & n11071 ) ;
  assign n11073 = ( x72 & ~n11017 ) | ( x72 & n11072 ) | ( ~n11017 & n11072 ) ;
  assign n11074 = ( x73 & ~n11009 ) | ( x73 & n11073 ) | ( ~n11009 & n11073 ) ;
  assign n11075 = ( x74 & ~n11001 ) | ( x74 & n11074 ) | ( ~n11001 & n11074 ) ;
  assign n11076 = ( x75 & ~n10993 ) | ( x75 & n11075 ) | ( ~n10993 & n11075 ) ;
  assign n11077 = ( x76 & ~n10985 ) | ( x76 & n11076 ) | ( ~n10985 & n11076 ) ;
  assign n11078 = ( x77 & ~n10977 ) | ( x77 & n11077 ) | ( ~n10977 & n11077 ) ;
  assign n11079 = ( x78 & ~n10969 ) | ( x78 & n11078 ) | ( ~n10969 & n11078 ) ;
  assign n11080 = ( x79 & ~n10961 ) | ( x79 & n11079 ) | ( ~n10961 & n11079 ) ;
  assign n11081 = ( x80 & ~n10953 ) | ( x80 & n11080 ) | ( ~n10953 & n11080 ) ;
  assign n11082 = ( x81 & ~n10945 ) | ( x81 & n11081 ) | ( ~n10945 & n11081 ) ;
  assign n11083 = ( x82 & ~n10937 ) | ( x82 & n11082 ) | ( ~n10937 & n11082 ) ;
  assign n11084 = ( x83 & ~n10929 ) | ( x83 & n11083 ) | ( ~n10929 & n11083 ) ;
  assign n11085 = ( x84 & ~n10921 ) | ( x84 & n11084 ) | ( ~n10921 & n11084 ) ;
  assign n11086 = ( x85 & ~n10913 ) | ( x85 & n11085 ) | ( ~n10913 & n11085 ) ;
  assign n11087 = ( x86 & ~n10905 ) | ( x86 & n11086 ) | ( ~n10905 & n11086 ) ;
  assign n11088 = ( x87 & ~n10897 ) | ( x87 & n11087 ) | ( ~n10897 & n11087 ) ;
  assign n11089 = ( x88 & ~n10889 ) | ( x88 & n11088 ) | ( ~n10889 & n11088 ) ;
  assign n11090 = ( x89 & ~n10881 ) | ( x89 & n11089 ) | ( ~n10881 & n11089 ) ;
  assign n11091 = ( x90 & ~n10873 ) | ( x90 & n11090 ) | ( ~n10873 & n11090 ) ;
  assign n11092 = ( x91 & ~n10865 ) | ( x91 & n11091 ) | ( ~n10865 & n11091 ) ;
  assign n11093 = ( x92 & ~n10857 ) | ( x92 & n11092 ) | ( ~n10857 & n11092 ) ;
  assign n11094 = ( x93 & ~n10849 ) | ( x93 & n11093 ) | ( ~n10849 & n11093 ) ;
  assign n11095 = ( x94 & ~n10841 ) | ( x94 & n11094 ) | ( ~n10841 & n11094 ) ;
  assign n11096 = ( x95 & ~n10833 ) | ( x95 & n11095 ) | ( ~n10833 & n11095 ) ;
  assign n11097 = ( x96 & ~n10825 ) | ( x96 & n11096 ) | ( ~n10825 & n11096 ) ;
  assign n11098 = ( x97 & ~n10817 ) | ( x97 & n11097 ) | ( ~n10817 & n11097 ) ;
  assign n11099 = ( x98 & ~n10809 ) | ( x98 & n11098 ) | ( ~n10809 & n11098 ) ;
  assign n11100 = ( x99 & ~n10801 ) | ( x99 & n11099 ) | ( ~n10801 & n11099 ) ;
  assign n11101 = ( x100 & ~n10793 ) | ( x100 & n11100 ) | ( ~n10793 & n11100 ) ;
  assign n11102 = ( x101 & ~n10699 ) | ( x101 & n11101 ) | ( ~n10699 & n11101 ) ;
  assign n11103 = ( x102 & ~n10785 ) | ( x102 & n11102 ) | ( ~n10785 & n11102 ) ;
  assign n11104 = ( x103 & ~n10780 ) | ( x103 & n11103 ) | ( ~n10780 & n11103 ) ;
  assign n11105 = ( x104 & ~n10772 ) | ( x104 & n11104 ) | ( ~n10772 & n11104 ) ;
  assign n11106 = ( x105 & ~n10764 ) | ( x105 & n11105 ) | ( ~n10764 & n11105 ) ;
  assign n11107 = ( x106 & ~n10756 ) | ( x106 & n11106 ) | ( ~n10756 & n11106 ) ;
  assign n11108 = ( x107 & ~n10748 ) | ( x107 & n11107 ) | ( ~n10748 & n11107 ) ;
  assign n11109 = ( x108 & ~n10740 ) | ( x108 & n11108 ) | ( ~n10740 & n11108 ) ;
  assign n11110 = ( x109 & ~n10732 ) | ( x109 & n11109 ) | ( ~n10732 & n11109 ) ;
  assign n11111 = ( x110 & ~n10724 ) | ( x110 & n11110 ) | ( ~n10724 & n11110 ) ;
  assign n11112 = ( x111 & ~n10716 ) | ( x111 & n11111 ) | ( ~n10716 & n11111 ) ;
  assign n11113 = ( x112 & ~n10708 ) | ( x112 & n11112 ) | ( ~n10708 & n11112 ) ;
  assign n11114 = n240 | n11113 ;
  assign n11474 = n10716 &  n11114 ;
  assign n11478 = x111 | n10716 ;
  assign n11479 = x111 &  n10716 ;
  assign n11480 = ( n11478 & ~n11479 ) | ( n11478 & 1'b0 ) | ( ~n11479 & 1'b0 ) ;
  assign n11481 = ( n240 & n11111 ) | ( n240 & n11480 ) | ( n11111 & n11480 ) ;
  assign n11482 = ( n11111 & ~n11113 ) | ( n11111 & n11480 ) | ( ~n11113 & n11480 ) ;
  assign n11483 = ~n11481 & n11482 ;
  assign n11484 = n11474 | n11483 ;
  assign n11485 = n10724 &  n11114 ;
  assign n11475 = x110 | n10724 ;
  assign n11476 = x110 &  n10724 ;
  assign n11477 = ( n11475 & ~n11476 ) | ( n11475 & 1'b0 ) | ( ~n11476 & 1'b0 ) ;
  assign n11489 = ( n240 & n11110 ) | ( n240 & n11477 ) | ( n11110 & n11477 ) ;
  assign n11490 = ( n11110 & ~n11113 ) | ( n11110 & n11477 ) | ( ~n11113 & n11477 ) ;
  assign n11491 = ~n11489 & n11490 ;
  assign n11492 = n11485 | n11491 ;
  assign n11493 = n10732 &  n11114 ;
  assign n11486 = x109 | n10732 ;
  assign n11487 = x109 &  n10732 ;
  assign n11488 = ( n11486 & ~n11487 ) | ( n11486 & 1'b0 ) | ( ~n11487 & 1'b0 ) ;
  assign n11497 = ( n240 & n11109 ) | ( n240 & n11488 ) | ( n11109 & n11488 ) ;
  assign n11498 = ( n11109 & ~n11113 ) | ( n11109 & n11488 ) | ( ~n11113 & n11488 ) ;
  assign n11499 = ~n11497 & n11498 ;
  assign n11500 = n11493 | n11499 ;
  assign n11501 = n10740 &  n11114 ;
  assign n11494 = x108 | n10740 ;
  assign n11495 = x108 &  n10740 ;
  assign n11496 = ( n11494 & ~n11495 ) | ( n11494 & 1'b0 ) | ( ~n11495 & 1'b0 ) ;
  assign n11505 = ( n240 & n11108 ) | ( n240 & n11496 ) | ( n11108 & n11496 ) ;
  assign n11506 = ( n11108 & ~n11113 ) | ( n11108 & n11496 ) | ( ~n11113 & n11496 ) ;
  assign n11507 = ~n11505 & n11506 ;
  assign n11508 = n11501 | n11507 ;
  assign n11509 = n10748 &  n11114 ;
  assign n11502 = x107 | n10748 ;
  assign n11503 = x107 &  n10748 ;
  assign n11504 = ( n11502 & ~n11503 ) | ( n11502 & 1'b0 ) | ( ~n11503 & 1'b0 ) ;
  assign n11513 = ( n240 & n11107 ) | ( n240 & n11504 ) | ( n11107 & n11504 ) ;
  assign n11514 = ( n11107 & ~n11113 ) | ( n11107 & n11504 ) | ( ~n11113 & n11504 ) ;
  assign n11515 = ~n11513 & n11514 ;
  assign n11516 = n11509 | n11515 ;
  assign n11517 = n10756 &  n11114 ;
  assign n11510 = x106 | n10756 ;
  assign n11511 = x106 &  n10756 ;
  assign n11512 = ( n11510 & ~n11511 ) | ( n11510 & 1'b0 ) | ( ~n11511 & 1'b0 ) ;
  assign n11521 = ( n240 & n11106 ) | ( n240 & n11512 ) | ( n11106 & n11512 ) ;
  assign n11522 = ( n11106 & ~n11113 ) | ( n11106 & n11512 ) | ( ~n11113 & n11512 ) ;
  assign n11523 = ~n11521 & n11522 ;
  assign n11524 = n11517 | n11523 ;
  assign n11525 = n10764 &  n11114 ;
  assign n11518 = x105 | n10764 ;
  assign n11519 = x105 &  n10764 ;
  assign n11520 = ( n11518 & ~n11519 ) | ( n11518 & 1'b0 ) | ( ~n11519 & 1'b0 ) ;
  assign n11529 = ( n240 & n11105 ) | ( n240 & n11520 ) | ( n11105 & n11520 ) ;
  assign n11530 = ( n11105 & ~n11113 ) | ( n11105 & n11520 ) | ( ~n11113 & n11520 ) ;
  assign n11531 = ~n11529 & n11530 ;
  assign n11532 = n11525 | n11531 ;
  assign n11533 = n10772 &  n11114 ;
  assign n11526 = x104 | n10772 ;
  assign n11527 = x104 &  n10772 ;
  assign n11528 = ( n11526 & ~n11527 ) | ( n11526 & 1'b0 ) | ( ~n11527 & 1'b0 ) ;
  assign n11537 = ( n240 & n11104 ) | ( n240 & n11528 ) | ( n11104 & n11528 ) ;
  assign n11538 = ( n11104 & ~n11113 ) | ( n11104 & n11528 ) | ( ~n11113 & n11528 ) ;
  assign n11539 = ~n11537 & n11538 ;
  assign n11540 = n11533 | n11539 ;
  assign n11541 = n10780 &  n11114 ;
  assign n11534 = x103 | n10780 ;
  assign n11535 = x103 &  n10780 ;
  assign n11536 = ( n11534 & ~n11535 ) | ( n11534 & 1'b0 ) | ( ~n11535 & 1'b0 ) ;
  assign n11542 = ( n240 & n11103 ) | ( n240 & n11536 ) | ( n11103 & n11536 ) ;
  assign n11543 = ( n11103 & ~n11113 ) | ( n11103 & n11536 ) | ( ~n11113 & n11536 ) ;
  assign n11544 = ~n11542 & n11543 ;
  assign n11545 = n11541 | n11544 ;
  assign n11463 = n10785 &  n11114 ;
  assign n11464 = x102 | n10785 ;
  assign n11465 = x102 &  n10785 ;
  assign n11466 = ( n11464 & ~n11465 ) | ( n11464 & 1'b0 ) | ( ~n11465 & 1'b0 ) ;
  assign n11467 = ( n240 & n11102 ) | ( n240 & n11466 ) | ( n11102 & n11466 ) ;
  assign n11468 = ( n11102 & ~n11113 ) | ( n11102 & n11466 ) | ( ~n11113 & n11466 ) ;
  assign n11469 = ~n11467 & n11468 ;
  assign n11470 = n11463 | n11469 ;
  assign n11115 = n10699 &  n11114 ;
  assign n11119 = x101 | n10699 ;
  assign n11120 = x101 &  n10699 ;
  assign n11121 = ( n11119 & ~n11120 ) | ( n11119 & 1'b0 ) | ( ~n11120 & 1'b0 ) ;
  assign n11122 = ( n240 & n11101 ) | ( n240 & n11121 ) | ( n11101 & n11121 ) ;
  assign n11123 = ( n11101 & ~n11113 ) | ( n11101 & n11121 ) | ( ~n11113 & n11121 ) ;
  assign n11124 = ~n11122 & n11123 ;
  assign n11125 = n11115 | n11124 ;
  assign n11126 = n10793 &  n11114 ;
  assign n11116 = x100 | n10793 ;
  assign n11117 = x100 &  n10793 ;
  assign n11118 = ( n11116 & ~n11117 ) | ( n11116 & 1'b0 ) | ( ~n11117 & 1'b0 ) ;
  assign n11130 = ( n240 & n11100 ) | ( n240 & n11118 ) | ( n11100 & n11118 ) ;
  assign n11131 = ( n11100 & ~n11113 ) | ( n11100 & n11118 ) | ( ~n11113 & n11118 ) ;
  assign n11132 = ~n11130 & n11131 ;
  assign n11133 = n11126 | n11132 ;
  assign n11134 = n10801 &  n11114 ;
  assign n11127 = x99 | n10801 ;
  assign n11128 = x99 &  n10801 ;
  assign n11129 = ( n11127 & ~n11128 ) | ( n11127 & 1'b0 ) | ( ~n11128 & 1'b0 ) ;
  assign n11138 = ( n240 & n11099 ) | ( n240 & n11129 ) | ( n11099 & n11129 ) ;
  assign n11139 = ( n11099 & ~n11113 ) | ( n11099 & n11129 ) | ( ~n11113 & n11129 ) ;
  assign n11140 = ~n11138 & n11139 ;
  assign n11141 = n11134 | n11140 ;
  assign n11142 = n10809 &  n11114 ;
  assign n11135 = x98 | n10809 ;
  assign n11136 = x98 &  n10809 ;
  assign n11137 = ( n11135 & ~n11136 ) | ( n11135 & 1'b0 ) | ( ~n11136 & 1'b0 ) ;
  assign n11146 = ( n240 & n11098 ) | ( n240 & n11137 ) | ( n11098 & n11137 ) ;
  assign n11147 = ( n11098 & ~n11113 ) | ( n11098 & n11137 ) | ( ~n11113 & n11137 ) ;
  assign n11148 = ~n11146 & n11147 ;
  assign n11149 = n11142 | n11148 ;
  assign n11150 = n10817 &  n11114 ;
  assign n11143 = x97 | n10817 ;
  assign n11144 = x97 &  n10817 ;
  assign n11145 = ( n11143 & ~n11144 ) | ( n11143 & 1'b0 ) | ( ~n11144 & 1'b0 ) ;
  assign n11154 = ( n240 & n11097 ) | ( n240 & n11145 ) | ( n11097 & n11145 ) ;
  assign n11155 = ( n11097 & ~n11113 ) | ( n11097 & n11145 ) | ( ~n11113 & n11145 ) ;
  assign n11156 = ~n11154 & n11155 ;
  assign n11157 = n11150 | n11156 ;
  assign n11158 = n10825 &  n11114 ;
  assign n11151 = x96 | n10825 ;
  assign n11152 = x96 &  n10825 ;
  assign n11153 = ( n11151 & ~n11152 ) | ( n11151 & 1'b0 ) | ( ~n11152 & 1'b0 ) ;
  assign n11162 = ( n240 & n11096 ) | ( n240 & n11153 ) | ( n11096 & n11153 ) ;
  assign n11163 = ( n11096 & ~n11113 ) | ( n11096 & n11153 ) | ( ~n11113 & n11153 ) ;
  assign n11164 = ~n11162 & n11163 ;
  assign n11165 = n11158 | n11164 ;
  assign n11166 = n10833 &  n11114 ;
  assign n11159 = x95 | n10833 ;
  assign n11160 = x95 &  n10833 ;
  assign n11161 = ( n11159 & ~n11160 ) | ( n11159 & 1'b0 ) | ( ~n11160 & 1'b0 ) ;
  assign n11170 = ( n240 & n11095 ) | ( n240 & n11161 ) | ( n11095 & n11161 ) ;
  assign n11171 = ( n11095 & ~n11113 ) | ( n11095 & n11161 ) | ( ~n11113 & n11161 ) ;
  assign n11172 = ~n11170 & n11171 ;
  assign n11173 = n11166 | n11172 ;
  assign n11174 = n10841 &  n11114 ;
  assign n11167 = x94 | n10841 ;
  assign n11168 = x94 &  n10841 ;
  assign n11169 = ( n11167 & ~n11168 ) | ( n11167 & 1'b0 ) | ( ~n11168 & 1'b0 ) ;
  assign n11178 = ( n240 & n11094 ) | ( n240 & n11169 ) | ( n11094 & n11169 ) ;
  assign n11179 = ( n11094 & ~n11113 ) | ( n11094 & n11169 ) | ( ~n11113 & n11169 ) ;
  assign n11180 = ~n11178 & n11179 ;
  assign n11181 = n11174 | n11180 ;
  assign n11182 = n10849 &  n11114 ;
  assign n11175 = x93 | n10849 ;
  assign n11176 = x93 &  n10849 ;
  assign n11177 = ( n11175 & ~n11176 ) | ( n11175 & 1'b0 ) | ( ~n11176 & 1'b0 ) ;
  assign n11186 = ( n240 & n11093 ) | ( n240 & n11177 ) | ( n11093 & n11177 ) ;
  assign n11187 = ( n11093 & ~n11113 ) | ( n11093 & n11177 ) | ( ~n11113 & n11177 ) ;
  assign n11188 = ~n11186 & n11187 ;
  assign n11189 = n11182 | n11188 ;
  assign n11190 = n10857 &  n11114 ;
  assign n11183 = x92 | n10857 ;
  assign n11184 = x92 &  n10857 ;
  assign n11185 = ( n11183 & ~n11184 ) | ( n11183 & 1'b0 ) | ( ~n11184 & 1'b0 ) ;
  assign n11194 = ( n240 & n11092 ) | ( n240 & n11185 ) | ( n11092 & n11185 ) ;
  assign n11195 = ( n11092 & ~n11113 ) | ( n11092 & n11185 ) | ( ~n11113 & n11185 ) ;
  assign n11196 = ~n11194 & n11195 ;
  assign n11197 = n11190 | n11196 ;
  assign n11198 = n10865 &  n11114 ;
  assign n11191 = x91 | n10865 ;
  assign n11192 = x91 &  n10865 ;
  assign n11193 = ( n11191 & ~n11192 ) | ( n11191 & 1'b0 ) | ( ~n11192 & 1'b0 ) ;
  assign n11202 = ( n240 & n11091 ) | ( n240 & n11193 ) | ( n11091 & n11193 ) ;
  assign n11203 = ( n11091 & ~n11113 ) | ( n11091 & n11193 ) | ( ~n11113 & n11193 ) ;
  assign n11204 = ~n11202 & n11203 ;
  assign n11205 = n11198 | n11204 ;
  assign n11206 = n10873 &  n11114 ;
  assign n11199 = x90 | n10873 ;
  assign n11200 = x90 &  n10873 ;
  assign n11201 = ( n11199 & ~n11200 ) | ( n11199 & 1'b0 ) | ( ~n11200 & 1'b0 ) ;
  assign n11210 = ( n240 & n11090 ) | ( n240 & n11201 ) | ( n11090 & n11201 ) ;
  assign n11211 = ( n11090 & ~n11113 ) | ( n11090 & n11201 ) | ( ~n11113 & n11201 ) ;
  assign n11212 = ~n11210 & n11211 ;
  assign n11213 = n11206 | n11212 ;
  assign n11214 = n10881 &  n11114 ;
  assign n11207 = x89 | n10881 ;
  assign n11208 = x89 &  n10881 ;
  assign n11209 = ( n11207 & ~n11208 ) | ( n11207 & 1'b0 ) | ( ~n11208 & 1'b0 ) ;
  assign n11218 = ( n240 & n11089 ) | ( n240 & n11209 ) | ( n11089 & n11209 ) ;
  assign n11219 = ( n11089 & ~n11113 ) | ( n11089 & n11209 ) | ( ~n11113 & n11209 ) ;
  assign n11220 = ~n11218 & n11219 ;
  assign n11221 = n11214 | n11220 ;
  assign n11222 = n10889 &  n11114 ;
  assign n11215 = x88 | n10889 ;
  assign n11216 = x88 &  n10889 ;
  assign n11217 = ( n11215 & ~n11216 ) | ( n11215 & 1'b0 ) | ( ~n11216 & 1'b0 ) ;
  assign n11226 = ( n240 & n11088 ) | ( n240 & n11217 ) | ( n11088 & n11217 ) ;
  assign n11227 = ( n11088 & ~n11113 ) | ( n11088 & n11217 ) | ( ~n11113 & n11217 ) ;
  assign n11228 = ~n11226 & n11227 ;
  assign n11229 = n11222 | n11228 ;
  assign n11230 = n10897 &  n11114 ;
  assign n11223 = x87 | n10897 ;
  assign n11224 = x87 &  n10897 ;
  assign n11225 = ( n11223 & ~n11224 ) | ( n11223 & 1'b0 ) | ( ~n11224 & 1'b0 ) ;
  assign n11234 = ( n240 & n11087 ) | ( n240 & n11225 ) | ( n11087 & n11225 ) ;
  assign n11235 = ( n11087 & ~n11113 ) | ( n11087 & n11225 ) | ( ~n11113 & n11225 ) ;
  assign n11236 = ~n11234 & n11235 ;
  assign n11237 = n11230 | n11236 ;
  assign n11238 = n10905 &  n11114 ;
  assign n11231 = x86 | n10905 ;
  assign n11232 = x86 &  n10905 ;
  assign n11233 = ( n11231 & ~n11232 ) | ( n11231 & 1'b0 ) | ( ~n11232 & 1'b0 ) ;
  assign n11242 = ( n240 & n11086 ) | ( n240 & n11233 ) | ( n11086 & n11233 ) ;
  assign n11243 = ( n11086 & ~n11113 ) | ( n11086 & n11233 ) | ( ~n11113 & n11233 ) ;
  assign n11244 = ~n11242 & n11243 ;
  assign n11245 = n11238 | n11244 ;
  assign n11246 = n10913 &  n11114 ;
  assign n11239 = x85 | n10913 ;
  assign n11240 = x85 &  n10913 ;
  assign n11241 = ( n11239 & ~n11240 ) | ( n11239 & 1'b0 ) | ( ~n11240 & 1'b0 ) ;
  assign n11250 = ( n240 & n11085 ) | ( n240 & n11241 ) | ( n11085 & n11241 ) ;
  assign n11251 = ( n11085 & ~n11113 ) | ( n11085 & n11241 ) | ( ~n11113 & n11241 ) ;
  assign n11252 = ~n11250 & n11251 ;
  assign n11253 = n11246 | n11252 ;
  assign n11254 = n10921 &  n11114 ;
  assign n11247 = x84 | n10921 ;
  assign n11248 = x84 &  n10921 ;
  assign n11249 = ( n11247 & ~n11248 ) | ( n11247 & 1'b0 ) | ( ~n11248 & 1'b0 ) ;
  assign n11258 = ( n240 & n11084 ) | ( n240 & n11249 ) | ( n11084 & n11249 ) ;
  assign n11259 = ( n11084 & ~n11113 ) | ( n11084 & n11249 ) | ( ~n11113 & n11249 ) ;
  assign n11260 = ~n11258 & n11259 ;
  assign n11261 = n11254 | n11260 ;
  assign n11262 = n10929 &  n11114 ;
  assign n11255 = x83 | n10929 ;
  assign n11256 = x83 &  n10929 ;
  assign n11257 = ( n11255 & ~n11256 ) | ( n11255 & 1'b0 ) | ( ~n11256 & 1'b0 ) ;
  assign n11266 = ( n240 & n11083 ) | ( n240 & n11257 ) | ( n11083 & n11257 ) ;
  assign n11267 = ( n11083 & ~n11113 ) | ( n11083 & n11257 ) | ( ~n11113 & n11257 ) ;
  assign n11268 = ~n11266 & n11267 ;
  assign n11269 = n11262 | n11268 ;
  assign n11270 = n10937 &  n11114 ;
  assign n11263 = x82 | n10937 ;
  assign n11264 = x82 &  n10937 ;
  assign n11265 = ( n11263 & ~n11264 ) | ( n11263 & 1'b0 ) | ( ~n11264 & 1'b0 ) ;
  assign n11274 = ( n240 & n11082 ) | ( n240 & n11265 ) | ( n11082 & n11265 ) ;
  assign n11275 = ( n11082 & ~n11113 ) | ( n11082 & n11265 ) | ( ~n11113 & n11265 ) ;
  assign n11276 = ~n11274 & n11275 ;
  assign n11277 = n11270 | n11276 ;
  assign n11278 = n10945 &  n11114 ;
  assign n11271 = x81 | n10945 ;
  assign n11272 = x81 &  n10945 ;
  assign n11273 = ( n11271 & ~n11272 ) | ( n11271 & 1'b0 ) | ( ~n11272 & 1'b0 ) ;
  assign n11282 = ( n240 & n11081 ) | ( n240 & n11273 ) | ( n11081 & n11273 ) ;
  assign n11283 = ( n11081 & ~n11113 ) | ( n11081 & n11273 ) | ( ~n11113 & n11273 ) ;
  assign n11284 = ~n11282 & n11283 ;
  assign n11285 = n11278 | n11284 ;
  assign n11286 = n10953 &  n11114 ;
  assign n11279 = x80 | n10953 ;
  assign n11280 = x80 &  n10953 ;
  assign n11281 = ( n11279 & ~n11280 ) | ( n11279 & 1'b0 ) | ( ~n11280 & 1'b0 ) ;
  assign n11290 = ( n240 & n11080 ) | ( n240 & n11281 ) | ( n11080 & n11281 ) ;
  assign n11291 = ( n11080 & ~n11113 ) | ( n11080 & n11281 ) | ( ~n11113 & n11281 ) ;
  assign n11292 = ~n11290 & n11291 ;
  assign n11293 = n11286 | n11292 ;
  assign n11294 = n10961 &  n11114 ;
  assign n11287 = x79 | n10961 ;
  assign n11288 = x79 &  n10961 ;
  assign n11289 = ( n11287 & ~n11288 ) | ( n11287 & 1'b0 ) | ( ~n11288 & 1'b0 ) ;
  assign n11298 = ( n240 & n11079 ) | ( n240 & n11289 ) | ( n11079 & n11289 ) ;
  assign n11299 = ( n11079 & ~n11113 ) | ( n11079 & n11289 ) | ( ~n11113 & n11289 ) ;
  assign n11300 = ~n11298 & n11299 ;
  assign n11301 = n11294 | n11300 ;
  assign n11302 = n10969 &  n11114 ;
  assign n11295 = x78 | n10969 ;
  assign n11296 = x78 &  n10969 ;
  assign n11297 = ( n11295 & ~n11296 ) | ( n11295 & 1'b0 ) | ( ~n11296 & 1'b0 ) ;
  assign n11306 = ( n240 & n11078 ) | ( n240 & n11297 ) | ( n11078 & n11297 ) ;
  assign n11307 = ( n11078 & ~n11113 ) | ( n11078 & n11297 ) | ( ~n11113 & n11297 ) ;
  assign n11308 = ~n11306 & n11307 ;
  assign n11309 = n11302 | n11308 ;
  assign n11310 = n10977 &  n11114 ;
  assign n11303 = x77 | n10977 ;
  assign n11304 = x77 &  n10977 ;
  assign n11305 = ( n11303 & ~n11304 ) | ( n11303 & 1'b0 ) | ( ~n11304 & 1'b0 ) ;
  assign n11314 = ( n240 & n11077 ) | ( n240 & n11305 ) | ( n11077 & n11305 ) ;
  assign n11315 = ( n11077 & ~n11113 ) | ( n11077 & n11305 ) | ( ~n11113 & n11305 ) ;
  assign n11316 = ~n11314 & n11315 ;
  assign n11317 = n11310 | n11316 ;
  assign n11318 = n10985 &  n11114 ;
  assign n11311 = x76 | n10985 ;
  assign n11312 = x76 &  n10985 ;
  assign n11313 = ( n11311 & ~n11312 ) | ( n11311 & 1'b0 ) | ( ~n11312 & 1'b0 ) ;
  assign n11322 = ( n240 & n11076 ) | ( n240 & n11313 ) | ( n11076 & n11313 ) ;
  assign n11323 = ( n11076 & ~n11113 ) | ( n11076 & n11313 ) | ( ~n11113 & n11313 ) ;
  assign n11324 = ~n11322 & n11323 ;
  assign n11325 = n11318 | n11324 ;
  assign n11326 = n10993 &  n11114 ;
  assign n11319 = x75 | n10993 ;
  assign n11320 = x75 &  n10993 ;
  assign n11321 = ( n11319 & ~n11320 ) | ( n11319 & 1'b0 ) | ( ~n11320 & 1'b0 ) ;
  assign n11330 = ( n240 & n11075 ) | ( n240 & n11321 ) | ( n11075 & n11321 ) ;
  assign n11331 = ( n11075 & ~n11113 ) | ( n11075 & n11321 ) | ( ~n11113 & n11321 ) ;
  assign n11332 = ~n11330 & n11331 ;
  assign n11333 = n11326 | n11332 ;
  assign n11334 = n11001 &  n11114 ;
  assign n11327 = x74 | n11001 ;
  assign n11328 = x74 &  n11001 ;
  assign n11329 = ( n11327 & ~n11328 ) | ( n11327 & 1'b0 ) | ( ~n11328 & 1'b0 ) ;
  assign n11338 = ( n240 & n11074 ) | ( n240 & n11329 ) | ( n11074 & n11329 ) ;
  assign n11339 = ( n11074 & ~n11113 ) | ( n11074 & n11329 ) | ( ~n11113 & n11329 ) ;
  assign n11340 = ~n11338 & n11339 ;
  assign n11341 = n11334 | n11340 ;
  assign n11342 = n11009 &  n11114 ;
  assign n11335 = x73 | n11009 ;
  assign n11336 = x73 &  n11009 ;
  assign n11337 = ( n11335 & ~n11336 ) | ( n11335 & 1'b0 ) | ( ~n11336 & 1'b0 ) ;
  assign n11346 = ( n240 & n11073 ) | ( n240 & n11337 ) | ( n11073 & n11337 ) ;
  assign n11347 = ( n11073 & ~n11113 ) | ( n11073 & n11337 ) | ( ~n11113 & n11337 ) ;
  assign n11348 = ~n11346 & n11347 ;
  assign n11349 = n11342 | n11348 ;
  assign n11350 = n11017 &  n11114 ;
  assign n11343 = x72 | n11017 ;
  assign n11344 = x72 &  n11017 ;
  assign n11345 = ( n11343 & ~n11344 ) | ( n11343 & 1'b0 ) | ( ~n11344 & 1'b0 ) ;
  assign n11354 = ( n240 & n11072 ) | ( n240 & n11345 ) | ( n11072 & n11345 ) ;
  assign n11355 = ( n11072 & ~n11113 ) | ( n11072 & n11345 ) | ( ~n11113 & n11345 ) ;
  assign n11356 = ~n11354 & n11355 ;
  assign n11357 = n11350 | n11356 ;
  assign n11358 = n11025 &  n11114 ;
  assign n11351 = x71 | n11025 ;
  assign n11352 = x71 &  n11025 ;
  assign n11353 = ( n11351 & ~n11352 ) | ( n11351 & 1'b0 ) | ( ~n11352 & 1'b0 ) ;
  assign n11362 = ( n240 & n11071 ) | ( n240 & n11353 ) | ( n11071 & n11353 ) ;
  assign n11363 = ( n11071 & ~n11113 ) | ( n11071 & n11353 ) | ( ~n11113 & n11353 ) ;
  assign n11364 = ~n11362 & n11363 ;
  assign n11365 = n11358 | n11364 ;
  assign n11366 = n11033 &  n11114 ;
  assign n11359 = x70 | n11033 ;
  assign n11360 = x70 &  n11033 ;
  assign n11361 = ( n11359 & ~n11360 ) | ( n11359 & 1'b0 ) | ( ~n11360 & 1'b0 ) ;
  assign n11370 = ( n240 & n11070 ) | ( n240 & n11361 ) | ( n11070 & n11361 ) ;
  assign n11371 = ( n11070 & ~n11113 ) | ( n11070 & n11361 ) | ( ~n11113 & n11361 ) ;
  assign n11372 = ~n11370 & n11371 ;
  assign n11373 = n11366 | n11372 ;
  assign n11374 = n11041 &  n11114 ;
  assign n11367 = x69 | n11041 ;
  assign n11368 = x69 &  n11041 ;
  assign n11369 = ( n11367 & ~n11368 ) | ( n11367 & 1'b0 ) | ( ~n11368 & 1'b0 ) ;
  assign n11378 = ( n240 & n11069 ) | ( n240 & n11369 ) | ( n11069 & n11369 ) ;
  assign n11379 = ( n11069 & ~n11113 ) | ( n11069 & n11369 ) | ( ~n11113 & n11369 ) ;
  assign n11380 = ~n11378 & n11379 ;
  assign n11381 = n11374 | n11380 ;
  assign n11382 = n11049 &  n11114 ;
  assign n11375 = x68 | n11049 ;
  assign n11376 = x68 &  n11049 ;
  assign n11377 = ( n11375 & ~n11376 ) | ( n11375 & 1'b0 ) | ( ~n11376 & 1'b0 ) ;
  assign n11386 = ( n240 & n11068 ) | ( n240 & n11377 ) | ( n11068 & n11377 ) ;
  assign n11387 = ( n11068 & ~n11113 ) | ( n11068 & n11377 ) | ( ~n11113 & n11377 ) ;
  assign n11388 = ~n11386 & n11387 ;
  assign n11389 = n11382 | n11388 ;
  assign n11390 = n11054 &  n11114 ;
  assign n11383 = x67 | n11054 ;
  assign n11384 = x67 &  n11054 ;
  assign n11385 = ( n11383 & ~n11384 ) | ( n11383 & 1'b0 ) | ( ~n11384 & 1'b0 ) ;
  assign n11394 = ( n240 & n11067 ) | ( n240 & n11385 ) | ( n11067 & n11385 ) ;
  assign n11395 = ( n11067 & ~n11113 ) | ( n11067 & n11385 ) | ( ~n11113 & n11385 ) ;
  assign n11396 = ~n11394 & n11395 ;
  assign n11397 = n11390 | n11396 ;
  assign n11398 = n11060 &  n11114 ;
  assign n11391 = x66 | n11060 ;
  assign n11392 = x66 &  n11060 ;
  assign n11393 = ( n11391 & ~n11392 ) | ( n11391 & 1'b0 ) | ( ~n11392 & 1'b0 ) ;
  assign n11399 = ( n11066 & ~n240 ) | ( n11066 & n11393 ) | ( ~n240 & n11393 ) ;
  assign n11400 = ( n11066 & n11113 ) | ( n11066 & n11393 ) | ( n11113 & n11393 ) ;
  assign n11401 = ( n11399 & ~n11400 ) | ( n11399 & 1'b0 ) | ( ~n11400 & 1'b0 ) ;
  assign n11402 = n11398 | n11401 ;
  assign n11403 = n11064 &  n11114 ;
  assign n11404 = ( x65 & ~x16 ) | ( x65 & n11061 ) | ( ~x16 & n11061 ) ;
  assign n11405 = ( x16 & ~n11061 ) | ( x16 & x65 ) | ( ~n11061 & x65 ) ;
  assign n11406 = ( n11404 & ~x65 ) | ( n11404 & n11405 ) | ( ~x65 & n11405 ) ;
  assign n11407 = ( n11065 & ~n11113 ) | ( n11065 & n11406 ) | ( ~n11113 & n11406 ) ;
  assign n11408 = ( n240 & n11065 ) | ( n240 & n11406 ) | ( n11065 & n11406 ) ;
  assign n11409 = ( n11407 & ~n11408 ) | ( n11407 & 1'b0 ) | ( ~n11408 & 1'b0 ) ;
  assign n11410 = n11403 | n11409 ;
  assign n11411 = ( x64 & ~x113 ) | ( x64 & 1'b0 ) | ( ~x113 & 1'b0 ) ;
  assign n11412 = ( n158 & ~n169 ) | ( n158 & n11411 ) | ( ~n169 & n11411 ) ;
  assign n11413 = ~n158 & n11412 ;
  assign n11414 = ~n269 & n11413 ;
  assign n11415 = n11113 &  n11414 ;
  assign n11416 = ( x15 & ~n11414 ) | ( x15 & n11415 ) | ( ~n11414 & n11415 ) ;
  assign n11417 = ~n232 & n11065 ;
  assign n11418 = ~n425 & n11417 ;
  assign n11419 = ~n11113 & n11418 ;
  assign n11420 = n11416 | n11419 ;
  assign n11421 = ~x14 & x64 ;
  assign n11422 = ( x65 & ~n11420 ) | ( x65 & n11421 ) | ( ~n11420 & n11421 ) ;
  assign n11423 = ( x66 & ~n11410 ) | ( x66 & n11422 ) | ( ~n11410 & n11422 ) ;
  assign n11424 = ( x67 & ~n11402 ) | ( x67 & n11423 ) | ( ~n11402 & n11423 ) ;
  assign n11425 = ( x68 & ~n11397 ) | ( x68 & n11424 ) | ( ~n11397 & n11424 ) ;
  assign n11426 = ( x69 & ~n11389 ) | ( x69 & n11425 ) | ( ~n11389 & n11425 ) ;
  assign n11427 = ( x70 & ~n11381 ) | ( x70 & n11426 ) | ( ~n11381 & n11426 ) ;
  assign n11428 = ( x71 & ~n11373 ) | ( x71 & n11427 ) | ( ~n11373 & n11427 ) ;
  assign n11429 = ( x72 & ~n11365 ) | ( x72 & n11428 ) | ( ~n11365 & n11428 ) ;
  assign n11430 = ( x73 & ~n11357 ) | ( x73 & n11429 ) | ( ~n11357 & n11429 ) ;
  assign n11431 = ( x74 & ~n11349 ) | ( x74 & n11430 ) | ( ~n11349 & n11430 ) ;
  assign n11432 = ( x75 & ~n11341 ) | ( x75 & n11431 ) | ( ~n11341 & n11431 ) ;
  assign n11433 = ( x76 & ~n11333 ) | ( x76 & n11432 ) | ( ~n11333 & n11432 ) ;
  assign n11434 = ( x77 & ~n11325 ) | ( x77 & n11433 ) | ( ~n11325 & n11433 ) ;
  assign n11435 = ( x78 & ~n11317 ) | ( x78 & n11434 ) | ( ~n11317 & n11434 ) ;
  assign n11436 = ( x79 & ~n11309 ) | ( x79 & n11435 ) | ( ~n11309 & n11435 ) ;
  assign n11437 = ( x80 & ~n11301 ) | ( x80 & n11436 ) | ( ~n11301 & n11436 ) ;
  assign n11438 = ( x81 & ~n11293 ) | ( x81 & n11437 ) | ( ~n11293 & n11437 ) ;
  assign n11439 = ( x82 & ~n11285 ) | ( x82 & n11438 ) | ( ~n11285 & n11438 ) ;
  assign n11440 = ( x83 & ~n11277 ) | ( x83 & n11439 ) | ( ~n11277 & n11439 ) ;
  assign n11441 = ( x84 & ~n11269 ) | ( x84 & n11440 ) | ( ~n11269 & n11440 ) ;
  assign n11442 = ( x85 & ~n11261 ) | ( x85 & n11441 ) | ( ~n11261 & n11441 ) ;
  assign n11443 = ( x86 & ~n11253 ) | ( x86 & n11442 ) | ( ~n11253 & n11442 ) ;
  assign n11444 = ( x87 & ~n11245 ) | ( x87 & n11443 ) | ( ~n11245 & n11443 ) ;
  assign n11445 = ( x88 & ~n11237 ) | ( x88 & n11444 ) | ( ~n11237 & n11444 ) ;
  assign n11446 = ( x89 & ~n11229 ) | ( x89 & n11445 ) | ( ~n11229 & n11445 ) ;
  assign n11447 = ( x90 & ~n11221 ) | ( x90 & n11446 ) | ( ~n11221 & n11446 ) ;
  assign n11448 = ( x91 & ~n11213 ) | ( x91 & n11447 ) | ( ~n11213 & n11447 ) ;
  assign n11449 = ( x92 & ~n11205 ) | ( x92 & n11448 ) | ( ~n11205 & n11448 ) ;
  assign n11450 = ( x93 & ~n11197 ) | ( x93 & n11449 ) | ( ~n11197 & n11449 ) ;
  assign n11451 = ( x94 & ~n11189 ) | ( x94 & n11450 ) | ( ~n11189 & n11450 ) ;
  assign n11452 = ( x95 & ~n11181 ) | ( x95 & n11451 ) | ( ~n11181 & n11451 ) ;
  assign n11453 = ( x96 & ~n11173 ) | ( x96 & n11452 ) | ( ~n11173 & n11452 ) ;
  assign n11454 = ( x97 & ~n11165 ) | ( x97 & n11453 ) | ( ~n11165 & n11453 ) ;
  assign n11455 = ( x98 & ~n11157 ) | ( x98 & n11454 ) | ( ~n11157 & n11454 ) ;
  assign n11456 = ( x99 & ~n11149 ) | ( x99 & n11455 ) | ( ~n11149 & n11455 ) ;
  assign n11457 = ( x100 & ~n11141 ) | ( x100 & n11456 ) | ( ~n11141 & n11456 ) ;
  assign n11458 = ( x101 & ~n11133 ) | ( x101 & n11457 ) | ( ~n11133 & n11457 ) ;
  assign n11462 = ( x102 & ~n11125 ) | ( x102 & n11458 ) | ( ~n11125 & n11458 ) ;
  assign n11546 = ( x103 & ~n11470 ) | ( x103 & n11462 ) | ( ~n11470 & n11462 ) ;
  assign n11547 = ( x104 & ~n11545 ) | ( x104 & n11546 ) | ( ~n11545 & n11546 ) ;
  assign n11548 = ( x105 & ~n11540 ) | ( x105 & n11547 ) | ( ~n11540 & n11547 ) ;
  assign n11549 = ( x106 & ~n11532 ) | ( x106 & n11548 ) | ( ~n11532 & n11548 ) ;
  assign n11550 = ( x107 & ~n11524 ) | ( x107 & n11549 ) | ( ~n11524 & n11549 ) ;
  assign n11551 = ( x108 & ~n11516 ) | ( x108 & n11550 ) | ( ~n11516 & n11550 ) ;
  assign n11552 = ( x109 & ~n11508 ) | ( x109 & n11551 ) | ( ~n11508 & n11551 ) ;
  assign n11553 = ( x110 & ~n11500 ) | ( x110 & n11552 ) | ( ~n11500 & n11552 ) ;
  assign n11554 = ( x111 & ~n11492 ) | ( x111 & n11553 ) | ( ~n11492 & n11553 ) ;
  assign n11555 = ( x112 & ~n11484 ) | ( x112 & n11554 ) | ( ~n11484 & n11554 ) ;
  assign n11559 = n158 | n169 ;
  assign n11560 = n269 | n11559 ;
  assign n11557 = ( x112 & ~n240 ) | ( x112 & n11112 ) | ( ~n240 & n11112 ) ;
  assign n11556 = x112 &  n11112 ;
  assign n11558 = ( n10708 & ~n11557 ) | ( n10708 & n11556 ) | ( ~n11557 & n11556 ) ;
  assign n11562 = x113 &  n11558 ;
  assign n11561 = x113 | n11558 ;
  assign n11563 = ( n11560 & ~n11562 ) | ( n11560 & n11561 ) | ( ~n11562 & n11561 ) ;
  assign n11564 = n11555 | n11563 ;
  assign n11565 = ~n11558 |  n240 ;
  assign n11936 = n11484 &  n11565 ;
  assign n11937 = n11564 &  n11936 ;
  assign n11933 = x112 | n11484 ;
  assign n11934 = x112 &  n11484 ;
  assign n11935 = ( n11933 & ~n11934 ) | ( n11933 & 1'b0 ) | ( ~n11934 & 1'b0 ) ;
  assign n11938 = n11554 &  n11935 ;
  assign n11566 = n11564 &  n11565 ;
  assign n11939 = ( n11554 & ~n11566 ) | ( n11554 & n11935 ) | ( ~n11566 & n11935 ) ;
  assign n11940 = ( n11937 & ~n11938 ) | ( n11937 & n11939 ) | ( ~n11938 & n11939 ) ;
  assign n11944 = n11492 &  n11565 ;
  assign n11945 = n11564 &  n11944 ;
  assign n11930 = x111 | n11492 ;
  assign n11931 = x111 &  n11492 ;
  assign n11932 = ( n11930 & ~n11931 ) | ( n11930 & 1'b0 ) | ( ~n11931 & 1'b0 ) ;
  assign n11946 = n11553 &  n11932 ;
  assign n11947 = ( n11553 & ~n11566 ) | ( n11553 & n11932 ) | ( ~n11566 & n11932 ) ;
  assign n11948 = ( n11945 & ~n11946 ) | ( n11945 & n11947 ) | ( ~n11946 & n11947 ) ;
  assign n11952 = n11500 &  n11565 ;
  assign n11953 = n11564 &  n11952 ;
  assign n11941 = x110 | n11500 ;
  assign n11942 = x110 &  n11500 ;
  assign n11943 = ( n11941 & ~n11942 ) | ( n11941 & 1'b0 ) | ( ~n11942 & 1'b0 ) ;
  assign n11954 = n11552 &  n11943 ;
  assign n11955 = ( n11552 & ~n11566 ) | ( n11552 & n11943 ) | ( ~n11566 & n11943 ) ;
  assign n11956 = ( n11953 & ~n11954 ) | ( n11953 & n11955 ) | ( ~n11954 & n11955 ) ;
  assign n11960 = n11508 &  n11565 ;
  assign n11961 = n11564 &  n11960 ;
  assign n11949 = x109 | n11508 ;
  assign n11950 = x109 &  n11508 ;
  assign n11951 = ( n11949 & ~n11950 ) | ( n11949 & 1'b0 ) | ( ~n11950 & 1'b0 ) ;
  assign n11962 = n11551 &  n11951 ;
  assign n11963 = ( n11551 & ~n11566 ) | ( n11551 & n11951 ) | ( ~n11566 & n11951 ) ;
  assign n11964 = ( n11961 & ~n11962 ) | ( n11961 & n11963 ) | ( ~n11962 & n11963 ) ;
  assign n11968 = n11516 &  n11565 ;
  assign n11969 = n11564 &  n11968 ;
  assign n11957 = x108 | n11516 ;
  assign n11958 = x108 &  n11516 ;
  assign n11959 = ( n11957 & ~n11958 ) | ( n11957 & 1'b0 ) | ( ~n11958 & 1'b0 ) ;
  assign n11970 = n11550 &  n11959 ;
  assign n11971 = ( n11550 & ~n11566 ) | ( n11550 & n11959 ) | ( ~n11566 & n11959 ) ;
  assign n11972 = ( n11969 & ~n11970 ) | ( n11969 & n11971 ) | ( ~n11970 & n11971 ) ;
  assign n11976 = n11524 &  n11565 ;
  assign n11977 = n11564 &  n11976 ;
  assign n11965 = x107 | n11524 ;
  assign n11966 = x107 &  n11524 ;
  assign n11967 = ( n11965 & ~n11966 ) | ( n11965 & 1'b0 ) | ( ~n11966 & 1'b0 ) ;
  assign n11979 = ( n11549 & n11566 ) | ( n11549 & n11967 ) | ( n11566 & n11967 ) ;
  assign n11978 = n11549 | n11967 ;
  assign n11980 = ( n11977 & ~n11979 ) | ( n11977 & n11978 ) | ( ~n11979 & n11978 ) ;
  assign n11984 = n11532 &  n11565 ;
  assign n11985 = n11564 &  n11984 ;
  assign n11973 = x106 | n11532 ;
  assign n11974 = x106 &  n11532 ;
  assign n11975 = ( n11973 & ~n11974 ) | ( n11973 & 1'b0 ) | ( ~n11974 & 1'b0 ) ;
  assign n11987 = ( n11548 & n11566 ) | ( n11548 & n11975 ) | ( n11566 & n11975 ) ;
  assign n11986 = n11548 | n11975 ;
  assign n11988 = ( n11985 & ~n11987 ) | ( n11985 & n11986 ) | ( ~n11987 & n11986 ) ;
  assign n11989 = n11540 &  n11565 ;
  assign n11990 = n11564 &  n11989 ;
  assign n11981 = x105 | n11540 ;
  assign n11982 = x105 &  n11540 ;
  assign n11983 = ( n11981 & ~n11982 ) | ( n11981 & 1'b0 ) | ( ~n11982 & 1'b0 ) ;
  assign n11992 = ( n11547 & n11566 ) | ( n11547 & n11983 ) | ( n11566 & n11983 ) ;
  assign n11991 = n11547 | n11983 ;
  assign n11993 = ( n11990 & ~n11992 ) | ( n11990 & n11991 ) | ( ~n11992 & n11991 ) ;
  assign n11922 = n11545 &  n11565 ;
  assign n11923 = n11564 &  n11922 ;
  assign n11919 = x104 | n11545 ;
  assign n11920 = x104 &  n11545 ;
  assign n11921 = ( n11919 & ~n11920 ) | ( n11919 & 1'b0 ) | ( ~n11920 & 1'b0 ) ;
  assign n11925 = ( n11546 & n11566 ) | ( n11546 & n11921 ) | ( n11566 & n11921 ) ;
  assign n11924 = n11546 | n11921 ;
  assign n11926 = ( n11923 & ~n11925 ) | ( n11923 & n11924 ) | ( ~n11925 & n11924 ) ;
  assign n11567 = n11470 &  n11565 ;
  assign n11568 = n11564 &  n11567 ;
  assign n11471 = x103 | n11470 ;
  assign n11472 = x103 &  n11470 ;
  assign n11473 = ( n11471 & ~n11472 ) | ( n11471 & 1'b0 ) | ( ~n11472 & 1'b0 ) ;
  assign n11570 = ( n11462 & n11473 ) | ( n11462 & n11566 ) | ( n11473 & n11566 ) ;
  assign n11569 = n11462 | n11473 ;
  assign n11571 = ( n11568 & ~n11570 ) | ( n11568 & n11569 ) | ( ~n11570 & n11569 ) ;
  assign n11575 = n11125 &  n11565 ;
  assign n11576 = n11564 &  n11575 ;
  assign n11459 = x102 | n11125 ;
  assign n11460 = x102 &  n11125 ;
  assign n11461 = ( n11459 & ~n11460 ) | ( n11459 & 1'b0 ) | ( ~n11460 & 1'b0 ) ;
  assign n11577 = n11458 &  n11461 ;
  assign n11578 = ( n11458 & ~n11566 ) | ( n11458 & n11461 ) | ( ~n11566 & n11461 ) ;
  assign n11579 = ( n11576 & ~n11577 ) | ( n11576 & n11578 ) | ( ~n11577 & n11578 ) ;
  assign n11583 = n11133 &  n11565 ;
  assign n11584 = n11564 &  n11583 ;
  assign n11572 = x101 | n11133 ;
  assign n11573 = x101 &  n11133 ;
  assign n11574 = ( n11572 & ~n11573 ) | ( n11572 & 1'b0 ) | ( ~n11573 & 1'b0 ) ;
  assign n11586 = ( n11457 & n11566 ) | ( n11457 & n11574 ) | ( n11566 & n11574 ) ;
  assign n11585 = n11457 | n11574 ;
  assign n11587 = ( n11584 & ~n11586 ) | ( n11584 & n11585 ) | ( ~n11586 & n11585 ) ;
  assign n11591 = n11141 &  n11565 ;
  assign n11592 = n11564 &  n11591 ;
  assign n11580 = x100 | n11141 ;
  assign n11581 = x100 &  n11141 ;
  assign n11582 = ( n11580 & ~n11581 ) | ( n11580 & 1'b0 ) | ( ~n11581 & 1'b0 ) ;
  assign n11594 = ( n11456 & n11566 ) | ( n11456 & n11582 ) | ( n11566 & n11582 ) ;
  assign n11593 = n11456 | n11582 ;
  assign n11595 = ( n11592 & ~n11594 ) | ( n11592 & n11593 ) | ( ~n11594 & n11593 ) ;
  assign n11599 = n11149 &  n11565 ;
  assign n11600 = n11564 &  n11599 ;
  assign n11588 = x99 | n11149 ;
  assign n11589 = x99 &  n11149 ;
  assign n11590 = ( n11588 & ~n11589 ) | ( n11588 & 1'b0 ) | ( ~n11589 & 1'b0 ) ;
  assign n11602 = ( n11455 & n11566 ) | ( n11455 & n11590 ) | ( n11566 & n11590 ) ;
  assign n11601 = n11455 | n11590 ;
  assign n11603 = ( n11600 & ~n11602 ) | ( n11600 & n11601 ) | ( ~n11602 & n11601 ) ;
  assign n11607 = n11157 &  n11565 ;
  assign n11608 = n11564 &  n11607 ;
  assign n11596 = x98 | n11157 ;
  assign n11597 = x98 &  n11157 ;
  assign n11598 = ( n11596 & ~n11597 ) | ( n11596 & 1'b0 ) | ( ~n11597 & 1'b0 ) ;
  assign n11610 = ( n11454 & n11566 ) | ( n11454 & n11598 ) | ( n11566 & n11598 ) ;
  assign n11609 = n11454 | n11598 ;
  assign n11611 = ( n11608 & ~n11610 ) | ( n11608 & n11609 ) | ( ~n11610 & n11609 ) ;
  assign n11615 = n11165 &  n11565 ;
  assign n11616 = n11564 &  n11615 ;
  assign n11604 = x97 | n11165 ;
  assign n11605 = x97 &  n11165 ;
  assign n11606 = ( n11604 & ~n11605 ) | ( n11604 & 1'b0 ) | ( ~n11605 & 1'b0 ) ;
  assign n11618 = ( n11453 & n11566 ) | ( n11453 & n11606 ) | ( n11566 & n11606 ) ;
  assign n11617 = n11453 | n11606 ;
  assign n11619 = ( n11616 & ~n11618 ) | ( n11616 & n11617 ) | ( ~n11618 & n11617 ) ;
  assign n11623 = n11173 &  n11565 ;
  assign n11624 = n11564 &  n11623 ;
  assign n11612 = x96 | n11173 ;
  assign n11613 = x96 &  n11173 ;
  assign n11614 = ( n11612 & ~n11613 ) | ( n11612 & 1'b0 ) | ( ~n11613 & 1'b0 ) ;
  assign n11626 = ( n11452 & n11566 ) | ( n11452 & n11614 ) | ( n11566 & n11614 ) ;
  assign n11625 = n11452 | n11614 ;
  assign n11627 = ( n11624 & ~n11626 ) | ( n11624 & n11625 ) | ( ~n11626 & n11625 ) ;
  assign n11631 = n11181 &  n11565 ;
  assign n11632 = n11564 &  n11631 ;
  assign n11620 = x95 | n11181 ;
  assign n11621 = x95 &  n11181 ;
  assign n11622 = ( n11620 & ~n11621 ) | ( n11620 & 1'b0 ) | ( ~n11621 & 1'b0 ) ;
  assign n11634 = ( n11451 & n11566 ) | ( n11451 & n11622 ) | ( n11566 & n11622 ) ;
  assign n11633 = n11451 | n11622 ;
  assign n11635 = ( n11632 & ~n11634 ) | ( n11632 & n11633 ) | ( ~n11634 & n11633 ) ;
  assign n11639 = n11189 &  n11565 ;
  assign n11640 = n11564 &  n11639 ;
  assign n11628 = x94 | n11189 ;
  assign n11629 = x94 &  n11189 ;
  assign n11630 = ( n11628 & ~n11629 ) | ( n11628 & 1'b0 ) | ( ~n11629 & 1'b0 ) ;
  assign n11642 = ( n11450 & n11566 ) | ( n11450 & n11630 ) | ( n11566 & n11630 ) ;
  assign n11641 = n11450 | n11630 ;
  assign n11643 = ( n11640 & ~n11642 ) | ( n11640 & n11641 ) | ( ~n11642 & n11641 ) ;
  assign n11647 = n11197 &  n11565 ;
  assign n11648 = n11564 &  n11647 ;
  assign n11636 = x93 | n11197 ;
  assign n11637 = x93 &  n11197 ;
  assign n11638 = ( n11636 & ~n11637 ) | ( n11636 & 1'b0 ) | ( ~n11637 & 1'b0 ) ;
  assign n11650 = ( n11449 & n11566 ) | ( n11449 & n11638 ) | ( n11566 & n11638 ) ;
  assign n11649 = n11449 | n11638 ;
  assign n11651 = ( n11648 & ~n11650 ) | ( n11648 & n11649 ) | ( ~n11650 & n11649 ) ;
  assign n11655 = n11205 &  n11565 ;
  assign n11656 = n11564 &  n11655 ;
  assign n11644 = x92 | n11205 ;
  assign n11645 = x92 &  n11205 ;
  assign n11646 = ( n11644 & ~n11645 ) | ( n11644 & 1'b0 ) | ( ~n11645 & 1'b0 ) ;
  assign n11658 = ( n11448 & n11566 ) | ( n11448 & n11646 ) | ( n11566 & n11646 ) ;
  assign n11657 = n11448 | n11646 ;
  assign n11659 = ( n11656 & ~n11658 ) | ( n11656 & n11657 ) | ( ~n11658 & n11657 ) ;
  assign n11663 = n11213 &  n11565 ;
  assign n11664 = n11564 &  n11663 ;
  assign n11652 = x91 | n11213 ;
  assign n11653 = x91 &  n11213 ;
  assign n11654 = ( n11652 & ~n11653 ) | ( n11652 & 1'b0 ) | ( ~n11653 & 1'b0 ) ;
  assign n11666 = ( n11447 & n11566 ) | ( n11447 & n11654 ) | ( n11566 & n11654 ) ;
  assign n11665 = n11447 | n11654 ;
  assign n11667 = ( n11664 & ~n11666 ) | ( n11664 & n11665 ) | ( ~n11666 & n11665 ) ;
  assign n11671 = n11221 &  n11565 ;
  assign n11672 = n11564 &  n11671 ;
  assign n11660 = x90 | n11221 ;
  assign n11661 = x90 &  n11221 ;
  assign n11662 = ( n11660 & ~n11661 ) | ( n11660 & 1'b0 ) | ( ~n11661 & 1'b0 ) ;
  assign n11674 = ( n11446 & n11566 ) | ( n11446 & n11662 ) | ( n11566 & n11662 ) ;
  assign n11673 = n11446 | n11662 ;
  assign n11675 = ( n11672 & ~n11674 ) | ( n11672 & n11673 ) | ( ~n11674 & n11673 ) ;
  assign n11679 = n11229 &  n11565 ;
  assign n11680 = n11564 &  n11679 ;
  assign n11668 = x89 | n11229 ;
  assign n11669 = x89 &  n11229 ;
  assign n11670 = ( n11668 & ~n11669 ) | ( n11668 & 1'b0 ) | ( ~n11669 & 1'b0 ) ;
  assign n11682 = ( n11445 & n11566 ) | ( n11445 & n11670 ) | ( n11566 & n11670 ) ;
  assign n11681 = n11445 | n11670 ;
  assign n11683 = ( n11680 & ~n11682 ) | ( n11680 & n11681 ) | ( ~n11682 & n11681 ) ;
  assign n11687 = n11237 &  n11565 ;
  assign n11688 = n11564 &  n11687 ;
  assign n11676 = x88 | n11237 ;
  assign n11677 = x88 &  n11237 ;
  assign n11678 = ( n11676 & ~n11677 ) | ( n11676 & 1'b0 ) | ( ~n11677 & 1'b0 ) ;
  assign n11690 = ( n11444 & n11566 ) | ( n11444 & n11678 ) | ( n11566 & n11678 ) ;
  assign n11689 = n11444 | n11678 ;
  assign n11691 = ( n11688 & ~n11690 ) | ( n11688 & n11689 ) | ( ~n11690 & n11689 ) ;
  assign n11695 = n11245 &  n11565 ;
  assign n11696 = n11564 &  n11695 ;
  assign n11684 = x87 | n11245 ;
  assign n11685 = x87 &  n11245 ;
  assign n11686 = ( n11684 & ~n11685 ) | ( n11684 & 1'b0 ) | ( ~n11685 & 1'b0 ) ;
  assign n11698 = ( n11443 & n11566 ) | ( n11443 & n11686 ) | ( n11566 & n11686 ) ;
  assign n11697 = n11443 | n11686 ;
  assign n11699 = ( n11696 & ~n11698 ) | ( n11696 & n11697 ) | ( ~n11698 & n11697 ) ;
  assign n11703 = n11253 &  n11565 ;
  assign n11704 = n11564 &  n11703 ;
  assign n11692 = x86 | n11253 ;
  assign n11693 = x86 &  n11253 ;
  assign n11694 = ( n11692 & ~n11693 ) | ( n11692 & 1'b0 ) | ( ~n11693 & 1'b0 ) ;
  assign n11706 = ( n11442 & n11566 ) | ( n11442 & n11694 ) | ( n11566 & n11694 ) ;
  assign n11705 = n11442 | n11694 ;
  assign n11707 = ( n11704 & ~n11706 ) | ( n11704 & n11705 ) | ( ~n11706 & n11705 ) ;
  assign n11711 = n11261 &  n11565 ;
  assign n11712 = n11564 &  n11711 ;
  assign n11700 = x85 | n11261 ;
  assign n11701 = x85 &  n11261 ;
  assign n11702 = ( n11700 & ~n11701 ) | ( n11700 & 1'b0 ) | ( ~n11701 & 1'b0 ) ;
  assign n11714 = ( n11441 & n11566 ) | ( n11441 & n11702 ) | ( n11566 & n11702 ) ;
  assign n11713 = n11441 | n11702 ;
  assign n11715 = ( n11712 & ~n11714 ) | ( n11712 & n11713 ) | ( ~n11714 & n11713 ) ;
  assign n11719 = n11269 &  n11565 ;
  assign n11720 = n11564 &  n11719 ;
  assign n11708 = x84 | n11269 ;
  assign n11709 = x84 &  n11269 ;
  assign n11710 = ( n11708 & ~n11709 ) | ( n11708 & 1'b0 ) | ( ~n11709 & 1'b0 ) ;
  assign n11722 = ( n11440 & n11566 ) | ( n11440 & n11710 ) | ( n11566 & n11710 ) ;
  assign n11721 = n11440 | n11710 ;
  assign n11723 = ( n11720 & ~n11722 ) | ( n11720 & n11721 ) | ( ~n11722 & n11721 ) ;
  assign n11727 = n11277 &  n11565 ;
  assign n11728 = n11564 &  n11727 ;
  assign n11716 = x83 | n11277 ;
  assign n11717 = x83 &  n11277 ;
  assign n11718 = ( n11716 & ~n11717 ) | ( n11716 & 1'b0 ) | ( ~n11717 & 1'b0 ) ;
  assign n11730 = ( n11439 & n11566 ) | ( n11439 & n11718 ) | ( n11566 & n11718 ) ;
  assign n11729 = n11439 | n11718 ;
  assign n11731 = ( n11728 & ~n11730 ) | ( n11728 & n11729 ) | ( ~n11730 & n11729 ) ;
  assign n11735 = n11285 &  n11565 ;
  assign n11736 = n11564 &  n11735 ;
  assign n11724 = x82 | n11285 ;
  assign n11725 = x82 &  n11285 ;
  assign n11726 = ( n11724 & ~n11725 ) | ( n11724 & 1'b0 ) | ( ~n11725 & 1'b0 ) ;
  assign n11738 = ( n11438 & n11566 ) | ( n11438 & n11726 ) | ( n11566 & n11726 ) ;
  assign n11737 = n11438 | n11726 ;
  assign n11739 = ( n11736 & ~n11738 ) | ( n11736 & n11737 ) | ( ~n11738 & n11737 ) ;
  assign n11743 = n11293 &  n11565 ;
  assign n11744 = n11564 &  n11743 ;
  assign n11732 = x81 | n11293 ;
  assign n11733 = x81 &  n11293 ;
  assign n11734 = ( n11732 & ~n11733 ) | ( n11732 & 1'b0 ) | ( ~n11733 & 1'b0 ) ;
  assign n11746 = ( n11437 & n11566 ) | ( n11437 & n11734 ) | ( n11566 & n11734 ) ;
  assign n11745 = n11437 | n11734 ;
  assign n11747 = ( n11744 & ~n11746 ) | ( n11744 & n11745 ) | ( ~n11746 & n11745 ) ;
  assign n11751 = n11301 &  n11565 ;
  assign n11752 = n11564 &  n11751 ;
  assign n11740 = x80 | n11301 ;
  assign n11741 = x80 &  n11301 ;
  assign n11742 = ( n11740 & ~n11741 ) | ( n11740 & 1'b0 ) | ( ~n11741 & 1'b0 ) ;
  assign n11754 = ( n11436 & n11566 ) | ( n11436 & n11742 ) | ( n11566 & n11742 ) ;
  assign n11753 = n11436 | n11742 ;
  assign n11755 = ( n11752 & ~n11754 ) | ( n11752 & n11753 ) | ( ~n11754 & n11753 ) ;
  assign n11759 = n11309 &  n11565 ;
  assign n11760 = n11564 &  n11759 ;
  assign n11748 = x79 | n11309 ;
  assign n11749 = x79 &  n11309 ;
  assign n11750 = ( n11748 & ~n11749 ) | ( n11748 & 1'b0 ) | ( ~n11749 & 1'b0 ) ;
  assign n11762 = ( n11435 & n11566 ) | ( n11435 & n11750 ) | ( n11566 & n11750 ) ;
  assign n11761 = n11435 | n11750 ;
  assign n11763 = ( n11760 & ~n11762 ) | ( n11760 & n11761 ) | ( ~n11762 & n11761 ) ;
  assign n11767 = n11317 &  n11565 ;
  assign n11768 = n11564 &  n11767 ;
  assign n11756 = x78 | n11317 ;
  assign n11757 = x78 &  n11317 ;
  assign n11758 = ( n11756 & ~n11757 ) | ( n11756 & 1'b0 ) | ( ~n11757 & 1'b0 ) ;
  assign n11770 = ( n11434 & n11566 ) | ( n11434 & n11758 ) | ( n11566 & n11758 ) ;
  assign n11769 = n11434 | n11758 ;
  assign n11771 = ( n11768 & ~n11770 ) | ( n11768 & n11769 ) | ( ~n11770 & n11769 ) ;
  assign n11775 = n11325 &  n11565 ;
  assign n11776 = n11564 &  n11775 ;
  assign n11764 = x77 | n11325 ;
  assign n11765 = x77 &  n11325 ;
  assign n11766 = ( n11764 & ~n11765 ) | ( n11764 & 1'b0 ) | ( ~n11765 & 1'b0 ) ;
  assign n11778 = ( n11433 & n11566 ) | ( n11433 & n11766 ) | ( n11566 & n11766 ) ;
  assign n11777 = n11433 | n11766 ;
  assign n11779 = ( n11776 & ~n11778 ) | ( n11776 & n11777 ) | ( ~n11778 & n11777 ) ;
  assign n11783 = n11333 &  n11565 ;
  assign n11784 = n11564 &  n11783 ;
  assign n11772 = x76 | n11333 ;
  assign n11773 = x76 &  n11333 ;
  assign n11774 = ( n11772 & ~n11773 ) | ( n11772 & 1'b0 ) | ( ~n11773 & 1'b0 ) ;
  assign n11786 = ( n11432 & n11566 ) | ( n11432 & n11774 ) | ( n11566 & n11774 ) ;
  assign n11785 = n11432 | n11774 ;
  assign n11787 = ( n11784 & ~n11786 ) | ( n11784 & n11785 ) | ( ~n11786 & n11785 ) ;
  assign n11791 = n11341 &  n11565 ;
  assign n11792 = n11564 &  n11791 ;
  assign n11780 = x75 | n11341 ;
  assign n11781 = x75 &  n11341 ;
  assign n11782 = ( n11780 & ~n11781 ) | ( n11780 & 1'b0 ) | ( ~n11781 & 1'b0 ) ;
  assign n11794 = ( n11431 & n11566 ) | ( n11431 & n11782 ) | ( n11566 & n11782 ) ;
  assign n11793 = n11431 | n11782 ;
  assign n11795 = ( n11792 & ~n11794 ) | ( n11792 & n11793 ) | ( ~n11794 & n11793 ) ;
  assign n11799 = n11349 &  n11565 ;
  assign n11800 = n11564 &  n11799 ;
  assign n11788 = x74 | n11349 ;
  assign n11789 = x74 &  n11349 ;
  assign n11790 = ( n11788 & ~n11789 ) | ( n11788 & 1'b0 ) | ( ~n11789 & 1'b0 ) ;
  assign n11802 = ( n11430 & n11566 ) | ( n11430 & n11790 ) | ( n11566 & n11790 ) ;
  assign n11801 = n11430 | n11790 ;
  assign n11803 = ( n11800 & ~n11802 ) | ( n11800 & n11801 ) | ( ~n11802 & n11801 ) ;
  assign n11807 = n11357 &  n11565 ;
  assign n11808 = n11564 &  n11807 ;
  assign n11796 = x73 | n11357 ;
  assign n11797 = x73 &  n11357 ;
  assign n11798 = ( n11796 & ~n11797 ) | ( n11796 & 1'b0 ) | ( ~n11797 & 1'b0 ) ;
  assign n11810 = ( n11429 & n11566 ) | ( n11429 & n11798 ) | ( n11566 & n11798 ) ;
  assign n11809 = n11429 | n11798 ;
  assign n11811 = ( n11808 & ~n11810 ) | ( n11808 & n11809 ) | ( ~n11810 & n11809 ) ;
  assign n11815 = n11365 &  n11565 ;
  assign n11816 = n11564 &  n11815 ;
  assign n11804 = x72 | n11365 ;
  assign n11805 = x72 &  n11365 ;
  assign n11806 = ( n11804 & ~n11805 ) | ( n11804 & 1'b0 ) | ( ~n11805 & 1'b0 ) ;
  assign n11818 = ( n11428 & n11566 ) | ( n11428 & n11806 ) | ( n11566 & n11806 ) ;
  assign n11817 = n11428 | n11806 ;
  assign n11819 = ( n11816 & ~n11818 ) | ( n11816 & n11817 ) | ( ~n11818 & n11817 ) ;
  assign n11823 = n11373 &  n11565 ;
  assign n11824 = n11564 &  n11823 ;
  assign n11812 = x71 | n11373 ;
  assign n11813 = x71 &  n11373 ;
  assign n11814 = ( n11812 & ~n11813 ) | ( n11812 & 1'b0 ) | ( ~n11813 & 1'b0 ) ;
  assign n11826 = ( n11427 & n11566 ) | ( n11427 & n11814 ) | ( n11566 & n11814 ) ;
  assign n11825 = n11427 | n11814 ;
  assign n11827 = ( n11824 & ~n11826 ) | ( n11824 & n11825 ) | ( ~n11826 & n11825 ) ;
  assign n11831 = n11381 &  n11565 ;
  assign n11832 = n11564 &  n11831 ;
  assign n11820 = x70 | n11381 ;
  assign n11821 = x70 &  n11381 ;
  assign n11822 = ( n11820 & ~n11821 ) | ( n11820 & 1'b0 ) | ( ~n11821 & 1'b0 ) ;
  assign n11834 = ( n11426 & n11566 ) | ( n11426 & n11822 ) | ( n11566 & n11822 ) ;
  assign n11833 = n11426 | n11822 ;
  assign n11835 = ( n11832 & ~n11834 ) | ( n11832 & n11833 ) | ( ~n11834 & n11833 ) ;
  assign n11839 = n11389 &  n11565 ;
  assign n11840 = n11564 &  n11839 ;
  assign n11828 = x69 | n11389 ;
  assign n11829 = x69 &  n11389 ;
  assign n11830 = ( n11828 & ~n11829 ) | ( n11828 & 1'b0 ) | ( ~n11829 & 1'b0 ) ;
  assign n11842 = ( n11425 & n11566 ) | ( n11425 & n11830 ) | ( n11566 & n11830 ) ;
  assign n11841 = n11425 | n11830 ;
  assign n11843 = ( n11840 & ~n11842 ) | ( n11840 & n11841 ) | ( ~n11842 & n11841 ) ;
  assign n11847 = n11397 &  n11565 ;
  assign n11848 = n11564 &  n11847 ;
  assign n11836 = x68 | n11397 ;
  assign n11837 = x68 &  n11397 ;
  assign n11838 = ( n11836 & ~n11837 ) | ( n11836 & 1'b0 ) | ( ~n11837 & 1'b0 ) ;
  assign n11850 = ( n11424 & n11566 ) | ( n11424 & n11838 ) | ( n11566 & n11838 ) ;
  assign n11849 = n11424 | n11838 ;
  assign n11851 = ( n11848 & ~n11850 ) | ( n11848 & n11849 ) | ( ~n11850 & n11849 ) ;
  assign n11855 = n11402 &  n11565 ;
  assign n11856 = n11564 &  n11855 ;
  assign n11844 = x67 | n11402 ;
  assign n11845 = x67 &  n11402 ;
  assign n11846 = ( n11844 & ~n11845 ) | ( n11844 & 1'b0 ) | ( ~n11845 & 1'b0 ) ;
  assign n11858 = ( n11423 & n11566 ) | ( n11423 & n11846 ) | ( n11566 & n11846 ) ;
  assign n11857 = n11423 | n11846 ;
  assign n11859 = ( n11856 & ~n11858 ) | ( n11856 & n11857 ) | ( ~n11858 & n11857 ) ;
  assign n11860 = n11410 &  n11565 ;
  assign n11861 = n11564 &  n11860 ;
  assign n11852 = x66 | n11410 ;
  assign n11853 = x66 &  n11410 ;
  assign n11854 = ( n11852 & ~n11853 ) | ( n11852 & 1'b0 ) | ( ~n11853 & 1'b0 ) ;
  assign n11862 = n11422 &  n11854 ;
  assign n11863 = ( n11422 & ~n11566 ) | ( n11422 & n11854 ) | ( ~n11566 & n11854 ) ;
  assign n11864 = ( n11861 & ~n11862 ) | ( n11861 & n11863 ) | ( ~n11862 & n11863 ) ;
  assign n11865 = ( n11420 & ~x65 ) | ( n11420 & n11421 ) | ( ~x65 & n11421 ) ;
  assign n11866 = ( n11422 & ~n11421 ) | ( n11422 & n11865 ) | ( ~n11421 & n11865 ) ;
  assign n11867 = ~n11566 & n11866 ;
  assign n11868 = n11420 &  n11565 ;
  assign n11869 = n11564 &  n11868 ;
  assign n11870 = n11867 | n11869 ;
  assign n11871 = ( x64 & ~n11566 ) | ( x64 & 1'b0 ) | ( ~n11566 & 1'b0 ) ;
  assign n11872 = ( x14 & ~n11871 ) | ( x14 & 1'b0 ) | ( ~n11871 & 1'b0 ) ;
  assign n11873 = ( n11421 & ~n11566 ) | ( n11421 & 1'b0 ) | ( ~n11566 & 1'b0 ) ;
  assign n11874 = n11872 | n11873 ;
  assign n11875 = ~x13 & x64 ;
  assign n11876 = ( x65 & ~n11874 ) | ( x65 & n11875 ) | ( ~n11874 & n11875 ) ;
  assign n11877 = ( x66 & ~n11870 ) | ( x66 & n11876 ) | ( ~n11870 & n11876 ) ;
  assign n11878 = ( x67 & ~n11864 ) | ( x67 & n11877 ) | ( ~n11864 & n11877 ) ;
  assign n11879 = ( x68 & ~n11859 ) | ( x68 & n11878 ) | ( ~n11859 & n11878 ) ;
  assign n11880 = ( x69 & ~n11851 ) | ( x69 & n11879 ) | ( ~n11851 & n11879 ) ;
  assign n11881 = ( x70 & ~n11843 ) | ( x70 & n11880 ) | ( ~n11843 & n11880 ) ;
  assign n11882 = ( x71 & ~n11835 ) | ( x71 & n11881 ) | ( ~n11835 & n11881 ) ;
  assign n11883 = ( x72 & ~n11827 ) | ( x72 & n11882 ) | ( ~n11827 & n11882 ) ;
  assign n11884 = ( x73 & ~n11819 ) | ( x73 & n11883 ) | ( ~n11819 & n11883 ) ;
  assign n11885 = ( x74 & ~n11811 ) | ( x74 & n11884 ) | ( ~n11811 & n11884 ) ;
  assign n11886 = ( x75 & ~n11803 ) | ( x75 & n11885 ) | ( ~n11803 & n11885 ) ;
  assign n11887 = ( x76 & ~n11795 ) | ( x76 & n11886 ) | ( ~n11795 & n11886 ) ;
  assign n11888 = ( x77 & ~n11787 ) | ( x77 & n11887 ) | ( ~n11787 & n11887 ) ;
  assign n11889 = ( x78 & ~n11779 ) | ( x78 & n11888 ) | ( ~n11779 & n11888 ) ;
  assign n11890 = ( x79 & ~n11771 ) | ( x79 & n11889 ) | ( ~n11771 & n11889 ) ;
  assign n11891 = ( x80 & ~n11763 ) | ( x80 & n11890 ) | ( ~n11763 & n11890 ) ;
  assign n11892 = ( x81 & ~n11755 ) | ( x81 & n11891 ) | ( ~n11755 & n11891 ) ;
  assign n11893 = ( x82 & ~n11747 ) | ( x82 & n11892 ) | ( ~n11747 & n11892 ) ;
  assign n11894 = ( x83 & ~n11739 ) | ( x83 & n11893 ) | ( ~n11739 & n11893 ) ;
  assign n11895 = ( x84 & ~n11731 ) | ( x84 & n11894 ) | ( ~n11731 & n11894 ) ;
  assign n11896 = ( x85 & ~n11723 ) | ( x85 & n11895 ) | ( ~n11723 & n11895 ) ;
  assign n11897 = ( x86 & ~n11715 ) | ( x86 & n11896 ) | ( ~n11715 & n11896 ) ;
  assign n11898 = ( x87 & ~n11707 ) | ( x87 & n11897 ) | ( ~n11707 & n11897 ) ;
  assign n11899 = ( x88 & ~n11699 ) | ( x88 & n11898 ) | ( ~n11699 & n11898 ) ;
  assign n11900 = ( x89 & ~n11691 ) | ( x89 & n11899 ) | ( ~n11691 & n11899 ) ;
  assign n11901 = ( x90 & ~n11683 ) | ( x90 & n11900 ) | ( ~n11683 & n11900 ) ;
  assign n11902 = ( x91 & ~n11675 ) | ( x91 & n11901 ) | ( ~n11675 & n11901 ) ;
  assign n11903 = ( x92 & ~n11667 ) | ( x92 & n11902 ) | ( ~n11667 & n11902 ) ;
  assign n11904 = ( x93 & ~n11659 ) | ( x93 & n11903 ) | ( ~n11659 & n11903 ) ;
  assign n11905 = ( x94 & ~n11651 ) | ( x94 & n11904 ) | ( ~n11651 & n11904 ) ;
  assign n11906 = ( x95 & ~n11643 ) | ( x95 & n11905 ) | ( ~n11643 & n11905 ) ;
  assign n11907 = ( x96 & ~n11635 ) | ( x96 & n11906 ) | ( ~n11635 & n11906 ) ;
  assign n11908 = ( x97 & ~n11627 ) | ( x97 & n11907 ) | ( ~n11627 & n11907 ) ;
  assign n11909 = ( x98 & ~n11619 ) | ( x98 & n11908 ) | ( ~n11619 & n11908 ) ;
  assign n11910 = ( x99 & ~n11611 ) | ( x99 & n11909 ) | ( ~n11611 & n11909 ) ;
  assign n11911 = ( x100 & ~n11603 ) | ( x100 & n11910 ) | ( ~n11603 & n11910 ) ;
  assign n11912 = ( x101 & ~n11595 ) | ( x101 & n11911 ) | ( ~n11595 & n11911 ) ;
  assign n11913 = ( x102 & ~n11587 ) | ( x102 & n11912 ) | ( ~n11587 & n11912 ) ;
  assign n11914 = ( x103 & ~n11579 ) | ( x103 & n11913 ) | ( ~n11579 & n11913 ) ;
  assign n11918 = ( x104 & ~n11571 ) | ( x104 & n11914 ) | ( ~n11571 & n11914 ) ;
  assign n11994 = ( x105 & ~n11926 ) | ( x105 & n11918 ) | ( ~n11926 & n11918 ) ;
  assign n11995 = ( x106 & ~n11993 ) | ( x106 & n11994 ) | ( ~n11993 & n11994 ) ;
  assign n11996 = ( x107 & ~n11988 ) | ( x107 & n11995 ) | ( ~n11988 & n11995 ) ;
  assign n11997 = ( x108 & ~n11980 ) | ( x108 & n11996 ) | ( ~n11980 & n11996 ) ;
  assign n11998 = ( x109 & ~n11972 ) | ( x109 & n11997 ) | ( ~n11972 & n11997 ) ;
  assign n11999 = ( x110 & ~n11964 ) | ( x110 & n11998 ) | ( ~n11964 & n11998 ) ;
  assign n12000 = ( x111 & ~n11956 ) | ( x111 & n11999 ) | ( ~n11956 & n11999 ) ;
  assign n12001 = ( x112 & ~n11948 ) | ( x112 & n12000 ) | ( ~n11948 & n12000 ) ;
  assign n12002 = ( x113 & ~n11940 ) | ( x113 & n12001 ) | ( ~n11940 & n12001 ) ;
  assign n12010 = n229 | n231 ;
  assign n12011 = n239 | n12010 ;
  assign n12004 = ( x113 & n11555 ) | ( x113 & n11558 ) | ( n11555 & n11558 ) ;
  assign n12003 = ( x113 & ~n11555 ) | ( x113 & n11558 ) | ( ~n11555 & n11558 ) ;
  assign n12005 = ( n11555 & ~n12004 ) | ( n11555 & n12003 ) | ( ~n12004 & n12003 ) ;
  assign n12006 = ~n11566 & n12005 ;
  assign n12007 = n240 &  n10708 ;
  assign n12008 = n11564 &  n12007 ;
  assign n12009 = n12006 | n12008 ;
  assign n12013 = x114 &  n12009 ;
  assign n12012 = x114 | n12009 ;
  assign n12014 = ( n12011 & ~n12013 ) | ( n12011 & n12012 ) | ( ~n12013 & n12012 ) ;
  assign n12015 = n12002 | n12014 ;
  assign n12016 = ~n12009 |  n11560 ;
  assign n12036 = n11940 &  n12016 ;
  assign n12037 = n12015 &  n12036 ;
  assign n12023 = x113 | n11940 ;
  assign n12024 = x113 &  n11940 ;
  assign n12025 = ( n12023 & ~n12024 ) | ( n12023 & 1'b0 ) | ( ~n12024 & 1'b0 ) ;
  assign n12038 = n12001 &  n12025 ;
  assign n12017 = n12015 &  n12016 ;
  assign n12039 = ( n12001 & ~n12017 ) | ( n12001 & n12025 ) | ( ~n12017 & n12025 ) ;
  assign n12040 = ( n12037 & ~n12038 ) | ( n12037 & n12039 ) | ( ~n12038 & n12039 ) ;
  assign n12027 = ( x114 & n12002 ) | ( x114 & n12009 ) | ( n12002 & n12009 ) ;
  assign n12026 = ( x114 & ~n12002 ) | ( x114 & n12009 ) | ( ~n12002 & n12009 ) ;
  assign n12028 = ( n12002 & ~n12027 ) | ( n12002 & n12026 ) | ( ~n12027 & n12026 ) ;
  assign n12029 = ~n12017 & n12028 ;
  assign n12030 = n11560 &  n12009 ;
  assign n12031 = n12015 &  n12030 ;
  assign n12032 = n12029 | n12031 ;
  assign n12044 = n11948 &  n12016 ;
  assign n12045 = n12015 &  n12044 ;
  assign n12033 = x112 | n11948 ;
  assign n12034 = x112 &  n11948 ;
  assign n12035 = ( n12033 & ~n12034 ) | ( n12033 & 1'b0 ) | ( ~n12034 & 1'b0 ) ;
  assign n12046 = n12000 &  n12035 ;
  assign n12047 = ( n12000 & ~n12017 ) | ( n12000 & n12035 ) | ( ~n12017 & n12035 ) ;
  assign n12048 = ( n12045 & ~n12046 ) | ( n12045 & n12047 ) | ( ~n12046 & n12047 ) ;
  assign n12052 = n11956 &  n12016 ;
  assign n12053 = n12015 &  n12052 ;
  assign n12041 = x111 | n11956 ;
  assign n12042 = x111 &  n11956 ;
  assign n12043 = ( n12041 & ~n12042 ) | ( n12041 & 1'b0 ) | ( ~n12042 & 1'b0 ) ;
  assign n12054 = n11999 &  n12043 ;
  assign n12055 = ( n11999 & ~n12017 ) | ( n11999 & n12043 ) | ( ~n12017 & n12043 ) ;
  assign n12056 = ( n12053 & ~n12054 ) | ( n12053 & n12055 ) | ( ~n12054 & n12055 ) ;
  assign n12060 = n11964 &  n12016 ;
  assign n12061 = n12015 &  n12060 ;
  assign n12049 = x110 | n11964 ;
  assign n12050 = x110 &  n11964 ;
  assign n12051 = ( n12049 & ~n12050 ) | ( n12049 & 1'b0 ) | ( ~n12050 & 1'b0 ) ;
  assign n12062 = n11998 &  n12051 ;
  assign n12063 = ( n11998 & ~n12017 ) | ( n11998 & n12051 ) | ( ~n12017 & n12051 ) ;
  assign n12064 = ( n12061 & ~n12062 ) | ( n12061 & n12063 ) | ( ~n12062 & n12063 ) ;
  assign n12068 = n11972 &  n12016 ;
  assign n12069 = n12015 &  n12068 ;
  assign n12057 = x109 | n11972 ;
  assign n12058 = x109 &  n11972 ;
  assign n12059 = ( n12057 & ~n12058 ) | ( n12057 & 1'b0 ) | ( ~n12058 & 1'b0 ) ;
  assign n12070 = n11997 &  n12059 ;
  assign n12071 = ( n11997 & ~n12017 ) | ( n11997 & n12059 ) | ( ~n12017 & n12059 ) ;
  assign n12072 = ( n12069 & ~n12070 ) | ( n12069 & n12071 ) | ( ~n12070 & n12071 ) ;
  assign n12076 = n11980 &  n12016 ;
  assign n12077 = n12015 &  n12076 ;
  assign n12065 = x108 | n11980 ;
  assign n12066 = x108 &  n11980 ;
  assign n12067 = ( n12065 & ~n12066 ) | ( n12065 & 1'b0 ) | ( ~n12066 & 1'b0 ) ;
  assign n12079 = ( n11996 & n12017 ) | ( n11996 & n12067 ) | ( n12017 & n12067 ) ;
  assign n12078 = n11996 | n12067 ;
  assign n12080 = ( n12077 & ~n12079 ) | ( n12077 & n12078 ) | ( ~n12079 & n12078 ) ;
  assign n12084 = n11988 &  n12016 ;
  assign n12085 = n12015 &  n12084 ;
  assign n12073 = x107 | n11988 ;
  assign n12074 = x107 &  n11988 ;
  assign n12075 = ( n12073 & ~n12074 ) | ( n12073 & 1'b0 ) | ( ~n12074 & 1'b0 ) ;
  assign n12087 = ( n11995 & n12017 ) | ( n11995 & n12075 ) | ( n12017 & n12075 ) ;
  assign n12086 = n11995 | n12075 ;
  assign n12088 = ( n12085 & ~n12087 ) | ( n12085 & n12086 ) | ( ~n12087 & n12086 ) ;
  assign n12089 = n11993 &  n12016 ;
  assign n12090 = n12015 &  n12089 ;
  assign n12081 = x106 | n11993 ;
  assign n12082 = x106 &  n11993 ;
  assign n12083 = ( n12081 & ~n12082 ) | ( n12081 & 1'b0 ) | ( ~n12082 & 1'b0 ) ;
  assign n12092 = ( n11994 & n12017 ) | ( n11994 & n12083 ) | ( n12017 & n12083 ) ;
  assign n12091 = n11994 | n12083 ;
  assign n12093 = ( n12090 & ~n12092 ) | ( n12090 & n12091 ) | ( ~n12092 & n12091 ) ;
  assign n12018 = n11926 &  n12016 ;
  assign n12019 = n12015 &  n12018 ;
  assign n11927 = x105 | n11926 ;
  assign n11928 = x105 &  n11926 ;
  assign n11929 = ( n11927 & ~n11928 ) | ( n11927 & 1'b0 ) | ( ~n11928 & 1'b0 ) ;
  assign n12021 = ( n11918 & n11929 ) | ( n11918 & n12017 ) | ( n11929 & n12017 ) ;
  assign n12020 = n11918 | n11929 ;
  assign n12022 = ( n12019 & ~n12021 ) | ( n12019 & n12020 ) | ( ~n12021 & n12020 ) ;
  assign n12097 = n11571 &  n12016 ;
  assign n12098 = n12015 &  n12097 ;
  assign n11915 = x104 | n11571 ;
  assign n11916 = x104 &  n11571 ;
  assign n11917 = ( n11915 & ~n11916 ) | ( n11915 & 1'b0 ) | ( ~n11916 & 1'b0 ) ;
  assign n12099 = n11914 &  n11917 ;
  assign n12100 = ( n11914 & ~n12017 ) | ( n11914 & n11917 ) | ( ~n12017 & n11917 ) ;
  assign n12101 = ( n12098 & ~n12099 ) | ( n12098 & n12100 ) | ( ~n12099 & n12100 ) ;
  assign n12105 = n11579 &  n12016 ;
  assign n12106 = n12015 &  n12105 ;
  assign n12094 = x103 | n11579 ;
  assign n12095 = x103 &  n11579 ;
  assign n12096 = ( n12094 & ~n12095 ) | ( n12094 & 1'b0 ) | ( ~n12095 & 1'b0 ) ;
  assign n12108 = ( n11913 & n12017 ) | ( n11913 & n12096 ) | ( n12017 & n12096 ) ;
  assign n12107 = n11913 | n12096 ;
  assign n12109 = ( n12106 & ~n12108 ) | ( n12106 & n12107 ) | ( ~n12108 & n12107 ) ;
  assign n12113 = n11587 &  n12016 ;
  assign n12114 = n12015 &  n12113 ;
  assign n12102 = x102 | n11587 ;
  assign n12103 = x102 &  n11587 ;
  assign n12104 = ( n12102 & ~n12103 ) | ( n12102 & 1'b0 ) | ( ~n12103 & 1'b0 ) ;
  assign n12116 = ( n11912 & n12017 ) | ( n11912 & n12104 ) | ( n12017 & n12104 ) ;
  assign n12115 = n11912 | n12104 ;
  assign n12117 = ( n12114 & ~n12116 ) | ( n12114 & n12115 ) | ( ~n12116 & n12115 ) ;
  assign n12121 = n11595 &  n12016 ;
  assign n12122 = n12015 &  n12121 ;
  assign n12110 = x101 | n11595 ;
  assign n12111 = x101 &  n11595 ;
  assign n12112 = ( n12110 & ~n12111 ) | ( n12110 & 1'b0 ) | ( ~n12111 & 1'b0 ) ;
  assign n12124 = ( n11911 & n12017 ) | ( n11911 & n12112 ) | ( n12017 & n12112 ) ;
  assign n12123 = n11911 | n12112 ;
  assign n12125 = ( n12122 & ~n12124 ) | ( n12122 & n12123 ) | ( ~n12124 & n12123 ) ;
  assign n12129 = n11603 &  n12016 ;
  assign n12130 = n12015 &  n12129 ;
  assign n12118 = x100 | n11603 ;
  assign n12119 = x100 &  n11603 ;
  assign n12120 = ( n12118 & ~n12119 ) | ( n12118 & 1'b0 ) | ( ~n12119 & 1'b0 ) ;
  assign n12132 = ( n11910 & n12017 ) | ( n11910 & n12120 ) | ( n12017 & n12120 ) ;
  assign n12131 = n11910 | n12120 ;
  assign n12133 = ( n12130 & ~n12132 ) | ( n12130 & n12131 ) | ( ~n12132 & n12131 ) ;
  assign n12137 = n11611 &  n12016 ;
  assign n12138 = n12015 &  n12137 ;
  assign n12126 = x99 | n11611 ;
  assign n12127 = x99 &  n11611 ;
  assign n12128 = ( n12126 & ~n12127 ) | ( n12126 & 1'b0 ) | ( ~n12127 & 1'b0 ) ;
  assign n12140 = ( n11909 & n12017 ) | ( n11909 & n12128 ) | ( n12017 & n12128 ) ;
  assign n12139 = n11909 | n12128 ;
  assign n12141 = ( n12138 & ~n12140 ) | ( n12138 & n12139 ) | ( ~n12140 & n12139 ) ;
  assign n12145 = n11619 &  n12016 ;
  assign n12146 = n12015 &  n12145 ;
  assign n12134 = x98 | n11619 ;
  assign n12135 = x98 &  n11619 ;
  assign n12136 = ( n12134 & ~n12135 ) | ( n12134 & 1'b0 ) | ( ~n12135 & 1'b0 ) ;
  assign n12148 = ( n11908 & n12017 ) | ( n11908 & n12136 ) | ( n12017 & n12136 ) ;
  assign n12147 = n11908 | n12136 ;
  assign n12149 = ( n12146 & ~n12148 ) | ( n12146 & n12147 ) | ( ~n12148 & n12147 ) ;
  assign n12153 = n11627 &  n12016 ;
  assign n12154 = n12015 &  n12153 ;
  assign n12142 = x97 | n11627 ;
  assign n12143 = x97 &  n11627 ;
  assign n12144 = ( n12142 & ~n12143 ) | ( n12142 & 1'b0 ) | ( ~n12143 & 1'b0 ) ;
  assign n12156 = ( n11907 & n12017 ) | ( n11907 & n12144 ) | ( n12017 & n12144 ) ;
  assign n12155 = n11907 | n12144 ;
  assign n12157 = ( n12154 & ~n12156 ) | ( n12154 & n12155 ) | ( ~n12156 & n12155 ) ;
  assign n12161 = n11635 &  n12016 ;
  assign n12162 = n12015 &  n12161 ;
  assign n12150 = x96 | n11635 ;
  assign n12151 = x96 &  n11635 ;
  assign n12152 = ( n12150 & ~n12151 ) | ( n12150 & 1'b0 ) | ( ~n12151 & 1'b0 ) ;
  assign n12164 = ( n11906 & n12017 ) | ( n11906 & n12152 ) | ( n12017 & n12152 ) ;
  assign n12163 = n11906 | n12152 ;
  assign n12165 = ( n12162 & ~n12164 ) | ( n12162 & n12163 ) | ( ~n12164 & n12163 ) ;
  assign n12169 = n11643 &  n12016 ;
  assign n12170 = n12015 &  n12169 ;
  assign n12158 = x95 | n11643 ;
  assign n12159 = x95 &  n11643 ;
  assign n12160 = ( n12158 & ~n12159 ) | ( n12158 & 1'b0 ) | ( ~n12159 & 1'b0 ) ;
  assign n12172 = ( n11905 & n12017 ) | ( n11905 & n12160 ) | ( n12017 & n12160 ) ;
  assign n12171 = n11905 | n12160 ;
  assign n12173 = ( n12170 & ~n12172 ) | ( n12170 & n12171 ) | ( ~n12172 & n12171 ) ;
  assign n12177 = n11651 &  n12016 ;
  assign n12178 = n12015 &  n12177 ;
  assign n12166 = x94 | n11651 ;
  assign n12167 = x94 &  n11651 ;
  assign n12168 = ( n12166 & ~n12167 ) | ( n12166 & 1'b0 ) | ( ~n12167 & 1'b0 ) ;
  assign n12180 = ( n11904 & n12017 ) | ( n11904 & n12168 ) | ( n12017 & n12168 ) ;
  assign n12179 = n11904 | n12168 ;
  assign n12181 = ( n12178 & ~n12180 ) | ( n12178 & n12179 ) | ( ~n12180 & n12179 ) ;
  assign n12185 = n11659 &  n12016 ;
  assign n12186 = n12015 &  n12185 ;
  assign n12174 = x93 | n11659 ;
  assign n12175 = x93 &  n11659 ;
  assign n12176 = ( n12174 & ~n12175 ) | ( n12174 & 1'b0 ) | ( ~n12175 & 1'b0 ) ;
  assign n12188 = ( n11903 & n12017 ) | ( n11903 & n12176 ) | ( n12017 & n12176 ) ;
  assign n12187 = n11903 | n12176 ;
  assign n12189 = ( n12186 & ~n12188 ) | ( n12186 & n12187 ) | ( ~n12188 & n12187 ) ;
  assign n12193 = n11667 &  n12016 ;
  assign n12194 = n12015 &  n12193 ;
  assign n12182 = x92 | n11667 ;
  assign n12183 = x92 &  n11667 ;
  assign n12184 = ( n12182 & ~n12183 ) | ( n12182 & 1'b0 ) | ( ~n12183 & 1'b0 ) ;
  assign n12196 = ( n11902 & n12017 ) | ( n11902 & n12184 ) | ( n12017 & n12184 ) ;
  assign n12195 = n11902 | n12184 ;
  assign n12197 = ( n12194 & ~n12196 ) | ( n12194 & n12195 ) | ( ~n12196 & n12195 ) ;
  assign n12201 = n11675 &  n12016 ;
  assign n12202 = n12015 &  n12201 ;
  assign n12190 = x91 | n11675 ;
  assign n12191 = x91 &  n11675 ;
  assign n12192 = ( n12190 & ~n12191 ) | ( n12190 & 1'b0 ) | ( ~n12191 & 1'b0 ) ;
  assign n12204 = ( n11901 & n12017 ) | ( n11901 & n12192 ) | ( n12017 & n12192 ) ;
  assign n12203 = n11901 | n12192 ;
  assign n12205 = ( n12202 & ~n12204 ) | ( n12202 & n12203 ) | ( ~n12204 & n12203 ) ;
  assign n12209 = n11683 &  n12016 ;
  assign n12210 = n12015 &  n12209 ;
  assign n12198 = x90 | n11683 ;
  assign n12199 = x90 &  n11683 ;
  assign n12200 = ( n12198 & ~n12199 ) | ( n12198 & 1'b0 ) | ( ~n12199 & 1'b0 ) ;
  assign n12212 = ( n11900 & n12017 ) | ( n11900 & n12200 ) | ( n12017 & n12200 ) ;
  assign n12211 = n11900 | n12200 ;
  assign n12213 = ( n12210 & ~n12212 ) | ( n12210 & n12211 ) | ( ~n12212 & n12211 ) ;
  assign n12217 = n11691 &  n12016 ;
  assign n12218 = n12015 &  n12217 ;
  assign n12206 = x89 | n11691 ;
  assign n12207 = x89 &  n11691 ;
  assign n12208 = ( n12206 & ~n12207 ) | ( n12206 & 1'b0 ) | ( ~n12207 & 1'b0 ) ;
  assign n12220 = ( n11899 & n12017 ) | ( n11899 & n12208 ) | ( n12017 & n12208 ) ;
  assign n12219 = n11899 | n12208 ;
  assign n12221 = ( n12218 & ~n12220 ) | ( n12218 & n12219 ) | ( ~n12220 & n12219 ) ;
  assign n12225 = n11699 &  n12016 ;
  assign n12226 = n12015 &  n12225 ;
  assign n12214 = x88 | n11699 ;
  assign n12215 = x88 &  n11699 ;
  assign n12216 = ( n12214 & ~n12215 ) | ( n12214 & 1'b0 ) | ( ~n12215 & 1'b0 ) ;
  assign n12228 = ( n11898 & n12017 ) | ( n11898 & n12216 ) | ( n12017 & n12216 ) ;
  assign n12227 = n11898 | n12216 ;
  assign n12229 = ( n12226 & ~n12228 ) | ( n12226 & n12227 ) | ( ~n12228 & n12227 ) ;
  assign n12233 = n11707 &  n12016 ;
  assign n12234 = n12015 &  n12233 ;
  assign n12222 = x87 | n11707 ;
  assign n12223 = x87 &  n11707 ;
  assign n12224 = ( n12222 & ~n12223 ) | ( n12222 & 1'b0 ) | ( ~n12223 & 1'b0 ) ;
  assign n12236 = ( n11897 & n12017 ) | ( n11897 & n12224 ) | ( n12017 & n12224 ) ;
  assign n12235 = n11897 | n12224 ;
  assign n12237 = ( n12234 & ~n12236 ) | ( n12234 & n12235 ) | ( ~n12236 & n12235 ) ;
  assign n12241 = n11715 &  n12016 ;
  assign n12242 = n12015 &  n12241 ;
  assign n12230 = x86 | n11715 ;
  assign n12231 = x86 &  n11715 ;
  assign n12232 = ( n12230 & ~n12231 ) | ( n12230 & 1'b0 ) | ( ~n12231 & 1'b0 ) ;
  assign n12244 = ( n11896 & n12017 ) | ( n11896 & n12232 ) | ( n12017 & n12232 ) ;
  assign n12243 = n11896 | n12232 ;
  assign n12245 = ( n12242 & ~n12244 ) | ( n12242 & n12243 ) | ( ~n12244 & n12243 ) ;
  assign n12249 = n11723 &  n12016 ;
  assign n12250 = n12015 &  n12249 ;
  assign n12238 = x85 | n11723 ;
  assign n12239 = x85 &  n11723 ;
  assign n12240 = ( n12238 & ~n12239 ) | ( n12238 & 1'b0 ) | ( ~n12239 & 1'b0 ) ;
  assign n12252 = ( n11895 & n12017 ) | ( n11895 & n12240 ) | ( n12017 & n12240 ) ;
  assign n12251 = n11895 | n12240 ;
  assign n12253 = ( n12250 & ~n12252 ) | ( n12250 & n12251 ) | ( ~n12252 & n12251 ) ;
  assign n12257 = n11731 &  n12016 ;
  assign n12258 = n12015 &  n12257 ;
  assign n12246 = x84 | n11731 ;
  assign n12247 = x84 &  n11731 ;
  assign n12248 = ( n12246 & ~n12247 ) | ( n12246 & 1'b0 ) | ( ~n12247 & 1'b0 ) ;
  assign n12260 = ( n11894 & n12017 ) | ( n11894 & n12248 ) | ( n12017 & n12248 ) ;
  assign n12259 = n11894 | n12248 ;
  assign n12261 = ( n12258 & ~n12260 ) | ( n12258 & n12259 ) | ( ~n12260 & n12259 ) ;
  assign n12265 = n11739 &  n12016 ;
  assign n12266 = n12015 &  n12265 ;
  assign n12254 = x83 | n11739 ;
  assign n12255 = x83 &  n11739 ;
  assign n12256 = ( n12254 & ~n12255 ) | ( n12254 & 1'b0 ) | ( ~n12255 & 1'b0 ) ;
  assign n12268 = ( n11893 & n12017 ) | ( n11893 & n12256 ) | ( n12017 & n12256 ) ;
  assign n12267 = n11893 | n12256 ;
  assign n12269 = ( n12266 & ~n12268 ) | ( n12266 & n12267 ) | ( ~n12268 & n12267 ) ;
  assign n12273 = n11747 &  n12016 ;
  assign n12274 = n12015 &  n12273 ;
  assign n12262 = x82 | n11747 ;
  assign n12263 = x82 &  n11747 ;
  assign n12264 = ( n12262 & ~n12263 ) | ( n12262 & 1'b0 ) | ( ~n12263 & 1'b0 ) ;
  assign n12276 = ( n11892 & n12017 ) | ( n11892 & n12264 ) | ( n12017 & n12264 ) ;
  assign n12275 = n11892 | n12264 ;
  assign n12277 = ( n12274 & ~n12276 ) | ( n12274 & n12275 ) | ( ~n12276 & n12275 ) ;
  assign n12281 = n11755 &  n12016 ;
  assign n12282 = n12015 &  n12281 ;
  assign n12270 = x81 | n11755 ;
  assign n12271 = x81 &  n11755 ;
  assign n12272 = ( n12270 & ~n12271 ) | ( n12270 & 1'b0 ) | ( ~n12271 & 1'b0 ) ;
  assign n12284 = ( n11891 & n12017 ) | ( n11891 & n12272 ) | ( n12017 & n12272 ) ;
  assign n12283 = n11891 | n12272 ;
  assign n12285 = ( n12282 & ~n12284 ) | ( n12282 & n12283 ) | ( ~n12284 & n12283 ) ;
  assign n12289 = n11763 &  n12016 ;
  assign n12290 = n12015 &  n12289 ;
  assign n12278 = x80 | n11763 ;
  assign n12279 = x80 &  n11763 ;
  assign n12280 = ( n12278 & ~n12279 ) | ( n12278 & 1'b0 ) | ( ~n12279 & 1'b0 ) ;
  assign n12292 = ( n11890 & n12017 ) | ( n11890 & n12280 ) | ( n12017 & n12280 ) ;
  assign n12291 = n11890 | n12280 ;
  assign n12293 = ( n12290 & ~n12292 ) | ( n12290 & n12291 ) | ( ~n12292 & n12291 ) ;
  assign n12297 = n11771 &  n12016 ;
  assign n12298 = n12015 &  n12297 ;
  assign n12286 = x79 | n11771 ;
  assign n12287 = x79 &  n11771 ;
  assign n12288 = ( n12286 & ~n12287 ) | ( n12286 & 1'b0 ) | ( ~n12287 & 1'b0 ) ;
  assign n12300 = ( n11889 & n12017 ) | ( n11889 & n12288 ) | ( n12017 & n12288 ) ;
  assign n12299 = n11889 | n12288 ;
  assign n12301 = ( n12298 & ~n12300 ) | ( n12298 & n12299 ) | ( ~n12300 & n12299 ) ;
  assign n12305 = n11779 &  n12016 ;
  assign n12306 = n12015 &  n12305 ;
  assign n12294 = x78 | n11779 ;
  assign n12295 = x78 &  n11779 ;
  assign n12296 = ( n12294 & ~n12295 ) | ( n12294 & 1'b0 ) | ( ~n12295 & 1'b0 ) ;
  assign n12308 = ( n11888 & n12017 ) | ( n11888 & n12296 ) | ( n12017 & n12296 ) ;
  assign n12307 = n11888 | n12296 ;
  assign n12309 = ( n12306 & ~n12308 ) | ( n12306 & n12307 ) | ( ~n12308 & n12307 ) ;
  assign n12313 = n11787 &  n12016 ;
  assign n12314 = n12015 &  n12313 ;
  assign n12302 = x77 | n11787 ;
  assign n12303 = x77 &  n11787 ;
  assign n12304 = ( n12302 & ~n12303 ) | ( n12302 & 1'b0 ) | ( ~n12303 & 1'b0 ) ;
  assign n12316 = ( n11887 & n12017 ) | ( n11887 & n12304 ) | ( n12017 & n12304 ) ;
  assign n12315 = n11887 | n12304 ;
  assign n12317 = ( n12314 & ~n12316 ) | ( n12314 & n12315 ) | ( ~n12316 & n12315 ) ;
  assign n12321 = n11795 &  n12016 ;
  assign n12322 = n12015 &  n12321 ;
  assign n12310 = x76 | n11795 ;
  assign n12311 = x76 &  n11795 ;
  assign n12312 = ( n12310 & ~n12311 ) | ( n12310 & 1'b0 ) | ( ~n12311 & 1'b0 ) ;
  assign n12324 = ( n11886 & n12017 ) | ( n11886 & n12312 ) | ( n12017 & n12312 ) ;
  assign n12323 = n11886 | n12312 ;
  assign n12325 = ( n12322 & ~n12324 ) | ( n12322 & n12323 ) | ( ~n12324 & n12323 ) ;
  assign n12329 = n11803 &  n12016 ;
  assign n12330 = n12015 &  n12329 ;
  assign n12318 = x75 | n11803 ;
  assign n12319 = x75 &  n11803 ;
  assign n12320 = ( n12318 & ~n12319 ) | ( n12318 & 1'b0 ) | ( ~n12319 & 1'b0 ) ;
  assign n12332 = ( n11885 & n12017 ) | ( n11885 & n12320 ) | ( n12017 & n12320 ) ;
  assign n12331 = n11885 | n12320 ;
  assign n12333 = ( n12330 & ~n12332 ) | ( n12330 & n12331 ) | ( ~n12332 & n12331 ) ;
  assign n12337 = n11811 &  n12016 ;
  assign n12338 = n12015 &  n12337 ;
  assign n12326 = x74 | n11811 ;
  assign n12327 = x74 &  n11811 ;
  assign n12328 = ( n12326 & ~n12327 ) | ( n12326 & 1'b0 ) | ( ~n12327 & 1'b0 ) ;
  assign n12340 = ( n11884 & n12017 ) | ( n11884 & n12328 ) | ( n12017 & n12328 ) ;
  assign n12339 = n11884 | n12328 ;
  assign n12341 = ( n12338 & ~n12340 ) | ( n12338 & n12339 ) | ( ~n12340 & n12339 ) ;
  assign n12345 = n11819 &  n12016 ;
  assign n12346 = n12015 &  n12345 ;
  assign n12334 = x73 | n11819 ;
  assign n12335 = x73 &  n11819 ;
  assign n12336 = ( n12334 & ~n12335 ) | ( n12334 & 1'b0 ) | ( ~n12335 & 1'b0 ) ;
  assign n12348 = ( n11883 & n12017 ) | ( n11883 & n12336 ) | ( n12017 & n12336 ) ;
  assign n12347 = n11883 | n12336 ;
  assign n12349 = ( n12346 & ~n12348 ) | ( n12346 & n12347 ) | ( ~n12348 & n12347 ) ;
  assign n12353 = n11827 &  n12016 ;
  assign n12354 = n12015 &  n12353 ;
  assign n12342 = x72 | n11827 ;
  assign n12343 = x72 &  n11827 ;
  assign n12344 = ( n12342 & ~n12343 ) | ( n12342 & 1'b0 ) | ( ~n12343 & 1'b0 ) ;
  assign n12356 = ( n11882 & n12017 ) | ( n11882 & n12344 ) | ( n12017 & n12344 ) ;
  assign n12355 = n11882 | n12344 ;
  assign n12357 = ( n12354 & ~n12356 ) | ( n12354 & n12355 ) | ( ~n12356 & n12355 ) ;
  assign n12361 = n11835 &  n12016 ;
  assign n12362 = n12015 &  n12361 ;
  assign n12350 = x71 | n11835 ;
  assign n12351 = x71 &  n11835 ;
  assign n12352 = ( n12350 & ~n12351 ) | ( n12350 & 1'b0 ) | ( ~n12351 & 1'b0 ) ;
  assign n12364 = ( n11881 & n12017 ) | ( n11881 & n12352 ) | ( n12017 & n12352 ) ;
  assign n12363 = n11881 | n12352 ;
  assign n12365 = ( n12362 & ~n12364 ) | ( n12362 & n12363 ) | ( ~n12364 & n12363 ) ;
  assign n12369 = n11843 &  n12016 ;
  assign n12370 = n12015 &  n12369 ;
  assign n12358 = x70 | n11843 ;
  assign n12359 = x70 &  n11843 ;
  assign n12360 = ( n12358 & ~n12359 ) | ( n12358 & 1'b0 ) | ( ~n12359 & 1'b0 ) ;
  assign n12372 = ( n11880 & n12017 ) | ( n11880 & n12360 ) | ( n12017 & n12360 ) ;
  assign n12371 = n11880 | n12360 ;
  assign n12373 = ( n12370 & ~n12372 ) | ( n12370 & n12371 ) | ( ~n12372 & n12371 ) ;
  assign n12377 = n11851 &  n12016 ;
  assign n12378 = n12015 &  n12377 ;
  assign n12366 = x69 | n11851 ;
  assign n12367 = x69 &  n11851 ;
  assign n12368 = ( n12366 & ~n12367 ) | ( n12366 & 1'b0 ) | ( ~n12367 & 1'b0 ) ;
  assign n12380 = ( n11879 & n12017 ) | ( n11879 & n12368 ) | ( n12017 & n12368 ) ;
  assign n12379 = n11879 | n12368 ;
  assign n12381 = ( n12378 & ~n12380 ) | ( n12378 & n12379 ) | ( ~n12380 & n12379 ) ;
  assign n12385 = n11859 &  n12016 ;
  assign n12386 = n12015 &  n12385 ;
  assign n12374 = x68 | n11859 ;
  assign n12375 = x68 &  n11859 ;
  assign n12376 = ( n12374 & ~n12375 ) | ( n12374 & 1'b0 ) | ( ~n12375 & 1'b0 ) ;
  assign n12388 = ( n11878 & n12017 ) | ( n11878 & n12376 ) | ( n12017 & n12376 ) ;
  assign n12387 = n11878 | n12376 ;
  assign n12389 = ( n12386 & ~n12388 ) | ( n12386 & n12387 ) | ( ~n12388 & n12387 ) ;
  assign n12393 = n11864 &  n12016 ;
  assign n12394 = n12015 &  n12393 ;
  assign n12382 = x67 | n11864 ;
  assign n12383 = x67 &  n11864 ;
  assign n12384 = ( n12382 & ~n12383 ) | ( n12382 & 1'b0 ) | ( ~n12383 & 1'b0 ) ;
  assign n12396 = ( n11877 & n12017 ) | ( n11877 & n12384 ) | ( n12017 & n12384 ) ;
  assign n12395 = n11877 | n12384 ;
  assign n12397 = ( n12394 & ~n12396 ) | ( n12394 & n12395 ) | ( ~n12396 & n12395 ) ;
  assign n12398 = n11870 &  n12016 ;
  assign n12399 = n12015 &  n12398 ;
  assign n12390 = x66 | n11870 ;
  assign n12391 = x66 &  n11870 ;
  assign n12392 = ( n12390 & ~n12391 ) | ( n12390 & 1'b0 ) | ( ~n12391 & 1'b0 ) ;
  assign n12400 = n11876 &  n12392 ;
  assign n12401 = ( n11876 & ~n12017 ) | ( n11876 & n12392 ) | ( ~n12017 & n12392 ) ;
  assign n12402 = ( n12399 & ~n12400 ) | ( n12399 & n12401 ) | ( ~n12400 & n12401 ) ;
  assign n12403 = ( n11874 & ~x65 ) | ( n11874 & n11875 ) | ( ~x65 & n11875 ) ;
  assign n12404 = ( n11876 & ~n11875 ) | ( n11876 & n12403 ) | ( ~n11875 & n12403 ) ;
  assign n12405 = ~n12017 & n12404 ;
  assign n12406 = n11874 &  n12016 ;
  assign n12407 = n12015 &  n12406 ;
  assign n12408 = n12405 | n12407 ;
  assign n12409 = ( x64 & ~n12017 ) | ( x64 & 1'b0 ) | ( ~n12017 & 1'b0 ) ;
  assign n12410 = ( x13 & ~n12409 ) | ( x13 & 1'b0 ) | ( ~n12409 & 1'b0 ) ;
  assign n12411 = ( n11875 & ~n12017 ) | ( n11875 & 1'b0 ) | ( ~n12017 & 1'b0 ) ;
  assign n12412 = n12410 | n12411 ;
  assign n12413 = ~x12 & x64 ;
  assign n12414 = ( x65 & ~n12412 ) | ( x65 & n12413 ) | ( ~n12412 & n12413 ) ;
  assign n12415 = ( x66 & ~n12408 ) | ( x66 & n12414 ) | ( ~n12408 & n12414 ) ;
  assign n12416 = ( x67 & ~n12402 ) | ( x67 & n12415 ) | ( ~n12402 & n12415 ) ;
  assign n12417 = ( x68 & ~n12397 ) | ( x68 & n12416 ) | ( ~n12397 & n12416 ) ;
  assign n12418 = ( x69 & ~n12389 ) | ( x69 & n12417 ) | ( ~n12389 & n12417 ) ;
  assign n12419 = ( x70 & ~n12381 ) | ( x70 & n12418 ) | ( ~n12381 & n12418 ) ;
  assign n12420 = ( x71 & ~n12373 ) | ( x71 & n12419 ) | ( ~n12373 & n12419 ) ;
  assign n12421 = ( x72 & ~n12365 ) | ( x72 & n12420 ) | ( ~n12365 & n12420 ) ;
  assign n12422 = ( x73 & ~n12357 ) | ( x73 & n12421 ) | ( ~n12357 & n12421 ) ;
  assign n12423 = ( x74 & ~n12349 ) | ( x74 & n12422 ) | ( ~n12349 & n12422 ) ;
  assign n12424 = ( x75 & ~n12341 ) | ( x75 & n12423 ) | ( ~n12341 & n12423 ) ;
  assign n12425 = ( x76 & ~n12333 ) | ( x76 & n12424 ) | ( ~n12333 & n12424 ) ;
  assign n12426 = ( x77 & ~n12325 ) | ( x77 & n12425 ) | ( ~n12325 & n12425 ) ;
  assign n12427 = ( x78 & ~n12317 ) | ( x78 & n12426 ) | ( ~n12317 & n12426 ) ;
  assign n12428 = ( x79 & ~n12309 ) | ( x79 & n12427 ) | ( ~n12309 & n12427 ) ;
  assign n12429 = ( x80 & ~n12301 ) | ( x80 & n12428 ) | ( ~n12301 & n12428 ) ;
  assign n12430 = ( x81 & ~n12293 ) | ( x81 & n12429 ) | ( ~n12293 & n12429 ) ;
  assign n12431 = ( x82 & ~n12285 ) | ( x82 & n12430 ) | ( ~n12285 & n12430 ) ;
  assign n12432 = ( x83 & ~n12277 ) | ( x83 & n12431 ) | ( ~n12277 & n12431 ) ;
  assign n12433 = ( x84 & ~n12269 ) | ( x84 & n12432 ) | ( ~n12269 & n12432 ) ;
  assign n12434 = ( x85 & ~n12261 ) | ( x85 & n12433 ) | ( ~n12261 & n12433 ) ;
  assign n12435 = ( x86 & ~n12253 ) | ( x86 & n12434 ) | ( ~n12253 & n12434 ) ;
  assign n12436 = ( x87 & ~n12245 ) | ( x87 & n12435 ) | ( ~n12245 & n12435 ) ;
  assign n12437 = ( x88 & ~n12237 ) | ( x88 & n12436 ) | ( ~n12237 & n12436 ) ;
  assign n12438 = ( x89 & ~n12229 ) | ( x89 & n12437 ) | ( ~n12229 & n12437 ) ;
  assign n12439 = ( x90 & ~n12221 ) | ( x90 & n12438 ) | ( ~n12221 & n12438 ) ;
  assign n12440 = ( x91 & ~n12213 ) | ( x91 & n12439 ) | ( ~n12213 & n12439 ) ;
  assign n12441 = ( x92 & ~n12205 ) | ( x92 & n12440 ) | ( ~n12205 & n12440 ) ;
  assign n12442 = ( x93 & ~n12197 ) | ( x93 & n12441 ) | ( ~n12197 & n12441 ) ;
  assign n12443 = ( x94 & ~n12189 ) | ( x94 & n12442 ) | ( ~n12189 & n12442 ) ;
  assign n12444 = ( x95 & ~n12181 ) | ( x95 & n12443 ) | ( ~n12181 & n12443 ) ;
  assign n12445 = ( x96 & ~n12173 ) | ( x96 & n12444 ) | ( ~n12173 & n12444 ) ;
  assign n12446 = ( x97 & ~n12165 ) | ( x97 & n12445 ) | ( ~n12165 & n12445 ) ;
  assign n12447 = ( x98 & ~n12157 ) | ( x98 & n12446 ) | ( ~n12157 & n12446 ) ;
  assign n12448 = ( x99 & ~n12149 ) | ( x99 & n12447 ) | ( ~n12149 & n12447 ) ;
  assign n12449 = ( x100 & ~n12141 ) | ( x100 & n12448 ) | ( ~n12141 & n12448 ) ;
  assign n12450 = ( x101 & ~n12133 ) | ( x101 & n12449 ) | ( ~n12133 & n12449 ) ;
  assign n12451 = ( x102 & ~n12125 ) | ( x102 & n12450 ) | ( ~n12125 & n12450 ) ;
  assign n12452 = ( x103 & ~n12117 ) | ( x103 & n12451 ) | ( ~n12117 & n12451 ) ;
  assign n12453 = ( x104 & ~n12109 ) | ( x104 & n12452 ) | ( ~n12109 & n12452 ) ;
  assign n12454 = ( x105 & ~n12101 ) | ( x105 & n12453 ) | ( ~n12101 & n12453 ) ;
  assign n12455 = ( x106 & ~n12022 ) | ( x106 & n12454 ) | ( ~n12022 & n12454 ) ;
  assign n12456 = ( x107 & ~n12093 ) | ( x107 & n12455 ) | ( ~n12093 & n12455 ) ;
  assign n12457 = ( x108 & ~n12088 ) | ( x108 & n12456 ) | ( ~n12088 & n12456 ) ;
  assign n12458 = ( x109 & ~n12080 ) | ( x109 & n12457 ) | ( ~n12080 & n12457 ) ;
  assign n12459 = ( x110 & ~n12072 ) | ( x110 & n12458 ) | ( ~n12072 & n12458 ) ;
  assign n12460 = ( x111 & ~n12064 ) | ( x111 & n12459 ) | ( ~n12064 & n12459 ) ;
  assign n12461 = ( x112 & ~n12056 ) | ( x112 & n12460 ) | ( ~n12056 & n12460 ) ;
  assign n12462 = ( x113 & ~n12048 ) | ( x113 & n12461 ) | ( ~n12048 & n12461 ) ;
  assign n12463 = ( x114 & ~n12040 ) | ( x114 & n12462 ) | ( ~n12040 & n12462 ) ;
  assign n12464 = ( x115 & ~n12032 ) | ( x115 & n12463 ) | ( ~n12032 & n12463 ) ;
  assign n12465 = n160 | n12464 ;
  assign n12869 = n12040 &  n12465 ;
  assign n12873 = x114 | n12040 ;
  assign n12874 = x114 &  n12040 ;
  assign n12875 = ( n12873 & ~n12874 ) | ( n12873 & 1'b0 ) | ( ~n12874 & 1'b0 ) ;
  assign n12876 = ( n160 & n12462 ) | ( n160 & n12875 ) | ( n12462 & n12875 ) ;
  assign n12877 = ( n12462 & ~n12464 ) | ( n12462 & n12875 ) | ( ~n12464 & n12875 ) ;
  assign n12878 = ~n12876 & n12877 ;
  assign n12879 = n12869 | n12878 ;
  assign n12880 = n12048 &  n12465 ;
  assign n12870 = x113 | n12048 ;
  assign n12871 = x113 &  n12048 ;
  assign n12872 = ( n12870 & ~n12871 ) | ( n12870 & 1'b0 ) | ( ~n12871 & 1'b0 ) ;
  assign n12884 = ( n160 & n12461 ) | ( n160 & n12872 ) | ( n12461 & n12872 ) ;
  assign n12885 = ( n12461 & ~n12464 ) | ( n12461 & n12872 ) | ( ~n12464 & n12872 ) ;
  assign n12886 = ~n12884 & n12885 ;
  assign n12887 = n12880 | n12886 ;
  assign n12888 = n12056 &  n12465 ;
  assign n12881 = x112 | n12056 ;
  assign n12882 = x112 &  n12056 ;
  assign n12883 = ( n12881 & ~n12882 ) | ( n12881 & 1'b0 ) | ( ~n12882 & 1'b0 ) ;
  assign n12892 = ( n160 & n12460 ) | ( n160 & n12883 ) | ( n12460 & n12883 ) ;
  assign n12893 = ( n12460 & ~n12464 ) | ( n12460 & n12883 ) | ( ~n12464 & n12883 ) ;
  assign n12894 = ~n12892 & n12893 ;
  assign n12895 = n12888 | n12894 ;
  assign n12896 = n12064 &  n12465 ;
  assign n12889 = x111 | n12064 ;
  assign n12890 = x111 &  n12064 ;
  assign n12891 = ( n12889 & ~n12890 ) | ( n12889 & 1'b0 ) | ( ~n12890 & 1'b0 ) ;
  assign n12900 = ( n160 & n12459 ) | ( n160 & n12891 ) | ( n12459 & n12891 ) ;
  assign n12901 = ( n12459 & ~n12464 ) | ( n12459 & n12891 ) | ( ~n12464 & n12891 ) ;
  assign n12902 = ~n12900 & n12901 ;
  assign n12903 = n12896 | n12902 ;
  assign n12904 = n12072 &  n12465 ;
  assign n12897 = x110 | n12072 ;
  assign n12898 = x110 &  n12072 ;
  assign n12899 = ( n12897 & ~n12898 ) | ( n12897 & 1'b0 ) | ( ~n12898 & 1'b0 ) ;
  assign n12908 = ( n160 & n12458 ) | ( n160 & n12899 ) | ( n12458 & n12899 ) ;
  assign n12909 = ( n12458 & ~n12464 ) | ( n12458 & n12899 ) | ( ~n12464 & n12899 ) ;
  assign n12910 = ~n12908 & n12909 ;
  assign n12911 = n12904 | n12910 ;
  assign n12912 = n12080 &  n12465 ;
  assign n12905 = x109 | n12080 ;
  assign n12906 = x109 &  n12080 ;
  assign n12907 = ( n12905 & ~n12906 ) | ( n12905 & 1'b0 ) | ( ~n12906 & 1'b0 ) ;
  assign n12916 = ( n160 & n12457 ) | ( n160 & n12907 ) | ( n12457 & n12907 ) ;
  assign n12917 = ( n12457 & ~n12464 ) | ( n12457 & n12907 ) | ( ~n12464 & n12907 ) ;
  assign n12918 = ~n12916 & n12917 ;
  assign n12919 = n12912 | n12918 ;
  assign n12920 = n12088 &  n12465 ;
  assign n12913 = x108 | n12088 ;
  assign n12914 = x108 &  n12088 ;
  assign n12915 = ( n12913 & ~n12914 ) | ( n12913 & 1'b0 ) | ( ~n12914 & 1'b0 ) ;
  assign n12921 = ( n160 & n12456 ) | ( n160 & n12915 ) | ( n12456 & n12915 ) ;
  assign n12922 = ( n12456 & ~n12464 ) | ( n12456 & n12915 ) | ( ~n12464 & n12915 ) ;
  assign n12923 = ~n12921 & n12922 ;
  assign n12924 = n12920 | n12923 ;
  assign n12858 = n12093 &  n12465 ;
  assign n12859 = x107 | n12093 ;
  assign n12860 = x107 &  n12093 ;
  assign n12861 = ( n12859 & ~n12860 ) | ( n12859 & 1'b0 ) | ( ~n12860 & 1'b0 ) ;
  assign n12862 = ( n160 & n12455 ) | ( n160 & n12861 ) | ( n12455 & n12861 ) ;
  assign n12863 = ( n12455 & ~n12464 ) | ( n12455 & n12861 ) | ( ~n12464 & n12861 ) ;
  assign n12864 = ~n12862 & n12863 ;
  assign n12865 = n12858 | n12864 ;
  assign n12466 = n12022 &  n12465 ;
  assign n12470 = x106 | n12022 ;
  assign n12471 = x106 &  n12022 ;
  assign n12472 = ( n12470 & ~n12471 ) | ( n12470 & 1'b0 ) | ( ~n12471 & 1'b0 ) ;
  assign n12473 = ( n160 & n12454 ) | ( n160 & n12472 ) | ( n12454 & n12472 ) ;
  assign n12474 = ( n12454 & ~n12464 ) | ( n12454 & n12472 ) | ( ~n12464 & n12472 ) ;
  assign n12475 = ~n12473 & n12474 ;
  assign n12476 = n12466 | n12475 ;
  assign n12477 = n12101 &  n12465 ;
  assign n12467 = x105 | n12101 ;
  assign n12468 = x105 &  n12101 ;
  assign n12469 = ( n12467 & ~n12468 ) | ( n12467 & 1'b0 ) | ( ~n12468 & 1'b0 ) ;
  assign n12481 = ( n160 & n12453 ) | ( n160 & n12469 ) | ( n12453 & n12469 ) ;
  assign n12482 = ( n12453 & ~n12464 ) | ( n12453 & n12469 ) | ( ~n12464 & n12469 ) ;
  assign n12483 = ~n12481 & n12482 ;
  assign n12484 = n12477 | n12483 ;
  assign n12485 = n12109 &  n12465 ;
  assign n12478 = x104 | n12109 ;
  assign n12479 = x104 &  n12109 ;
  assign n12480 = ( n12478 & ~n12479 ) | ( n12478 & 1'b0 ) | ( ~n12479 & 1'b0 ) ;
  assign n12489 = ( n160 & n12452 ) | ( n160 & n12480 ) | ( n12452 & n12480 ) ;
  assign n12490 = ( n12452 & ~n12464 ) | ( n12452 & n12480 ) | ( ~n12464 & n12480 ) ;
  assign n12491 = ~n12489 & n12490 ;
  assign n12492 = n12485 | n12491 ;
  assign n12493 = n12117 &  n12465 ;
  assign n12486 = x103 | n12117 ;
  assign n12487 = x103 &  n12117 ;
  assign n12488 = ( n12486 & ~n12487 ) | ( n12486 & 1'b0 ) | ( ~n12487 & 1'b0 ) ;
  assign n12497 = ( n160 & n12451 ) | ( n160 & n12488 ) | ( n12451 & n12488 ) ;
  assign n12498 = ( n12451 & ~n12464 ) | ( n12451 & n12488 ) | ( ~n12464 & n12488 ) ;
  assign n12499 = ~n12497 & n12498 ;
  assign n12500 = n12493 | n12499 ;
  assign n12501 = n12125 &  n12465 ;
  assign n12494 = x102 | n12125 ;
  assign n12495 = x102 &  n12125 ;
  assign n12496 = ( n12494 & ~n12495 ) | ( n12494 & 1'b0 ) | ( ~n12495 & 1'b0 ) ;
  assign n12505 = ( n160 & n12450 ) | ( n160 & n12496 ) | ( n12450 & n12496 ) ;
  assign n12506 = ( n12450 & ~n12464 ) | ( n12450 & n12496 ) | ( ~n12464 & n12496 ) ;
  assign n12507 = ~n12505 & n12506 ;
  assign n12508 = n12501 | n12507 ;
  assign n12509 = n12133 &  n12465 ;
  assign n12502 = x101 | n12133 ;
  assign n12503 = x101 &  n12133 ;
  assign n12504 = ( n12502 & ~n12503 ) | ( n12502 & 1'b0 ) | ( ~n12503 & 1'b0 ) ;
  assign n12513 = ( n160 & n12449 ) | ( n160 & n12504 ) | ( n12449 & n12504 ) ;
  assign n12514 = ( n12449 & ~n12464 ) | ( n12449 & n12504 ) | ( ~n12464 & n12504 ) ;
  assign n12515 = ~n12513 & n12514 ;
  assign n12516 = n12509 | n12515 ;
  assign n12517 = n12141 &  n12465 ;
  assign n12510 = x100 | n12141 ;
  assign n12511 = x100 &  n12141 ;
  assign n12512 = ( n12510 & ~n12511 ) | ( n12510 & 1'b0 ) | ( ~n12511 & 1'b0 ) ;
  assign n12521 = ( n160 & n12448 ) | ( n160 & n12512 ) | ( n12448 & n12512 ) ;
  assign n12522 = ( n12448 & ~n12464 ) | ( n12448 & n12512 ) | ( ~n12464 & n12512 ) ;
  assign n12523 = ~n12521 & n12522 ;
  assign n12524 = n12517 | n12523 ;
  assign n12525 = n12149 &  n12465 ;
  assign n12518 = x99 | n12149 ;
  assign n12519 = x99 &  n12149 ;
  assign n12520 = ( n12518 & ~n12519 ) | ( n12518 & 1'b0 ) | ( ~n12519 & 1'b0 ) ;
  assign n12529 = ( n160 & n12447 ) | ( n160 & n12520 ) | ( n12447 & n12520 ) ;
  assign n12530 = ( n12447 & ~n12464 ) | ( n12447 & n12520 ) | ( ~n12464 & n12520 ) ;
  assign n12531 = ~n12529 & n12530 ;
  assign n12532 = n12525 | n12531 ;
  assign n12533 = n12157 &  n12465 ;
  assign n12526 = x98 | n12157 ;
  assign n12527 = x98 &  n12157 ;
  assign n12528 = ( n12526 & ~n12527 ) | ( n12526 & 1'b0 ) | ( ~n12527 & 1'b0 ) ;
  assign n12537 = ( n160 & n12446 ) | ( n160 & n12528 ) | ( n12446 & n12528 ) ;
  assign n12538 = ( n12446 & ~n12464 ) | ( n12446 & n12528 ) | ( ~n12464 & n12528 ) ;
  assign n12539 = ~n12537 & n12538 ;
  assign n12540 = n12533 | n12539 ;
  assign n12541 = n12165 &  n12465 ;
  assign n12534 = x97 | n12165 ;
  assign n12535 = x97 &  n12165 ;
  assign n12536 = ( n12534 & ~n12535 ) | ( n12534 & 1'b0 ) | ( ~n12535 & 1'b0 ) ;
  assign n12545 = ( n160 & n12445 ) | ( n160 & n12536 ) | ( n12445 & n12536 ) ;
  assign n12546 = ( n12445 & ~n12464 ) | ( n12445 & n12536 ) | ( ~n12464 & n12536 ) ;
  assign n12547 = ~n12545 & n12546 ;
  assign n12548 = n12541 | n12547 ;
  assign n12549 = n12173 &  n12465 ;
  assign n12542 = x96 | n12173 ;
  assign n12543 = x96 &  n12173 ;
  assign n12544 = ( n12542 & ~n12543 ) | ( n12542 & 1'b0 ) | ( ~n12543 & 1'b0 ) ;
  assign n12553 = ( n160 & n12444 ) | ( n160 & n12544 ) | ( n12444 & n12544 ) ;
  assign n12554 = ( n12444 & ~n12464 ) | ( n12444 & n12544 ) | ( ~n12464 & n12544 ) ;
  assign n12555 = ~n12553 & n12554 ;
  assign n12556 = n12549 | n12555 ;
  assign n12557 = n12181 &  n12465 ;
  assign n12550 = x95 | n12181 ;
  assign n12551 = x95 &  n12181 ;
  assign n12552 = ( n12550 & ~n12551 ) | ( n12550 & 1'b0 ) | ( ~n12551 & 1'b0 ) ;
  assign n12561 = ( n160 & n12443 ) | ( n160 & n12552 ) | ( n12443 & n12552 ) ;
  assign n12562 = ( n12443 & ~n12464 ) | ( n12443 & n12552 ) | ( ~n12464 & n12552 ) ;
  assign n12563 = ~n12561 & n12562 ;
  assign n12564 = n12557 | n12563 ;
  assign n12565 = n12189 &  n12465 ;
  assign n12558 = x94 | n12189 ;
  assign n12559 = x94 &  n12189 ;
  assign n12560 = ( n12558 & ~n12559 ) | ( n12558 & 1'b0 ) | ( ~n12559 & 1'b0 ) ;
  assign n12569 = ( n160 & n12442 ) | ( n160 & n12560 ) | ( n12442 & n12560 ) ;
  assign n12570 = ( n12442 & ~n12464 ) | ( n12442 & n12560 ) | ( ~n12464 & n12560 ) ;
  assign n12571 = ~n12569 & n12570 ;
  assign n12572 = n12565 | n12571 ;
  assign n12573 = n12197 &  n12465 ;
  assign n12566 = x93 | n12197 ;
  assign n12567 = x93 &  n12197 ;
  assign n12568 = ( n12566 & ~n12567 ) | ( n12566 & 1'b0 ) | ( ~n12567 & 1'b0 ) ;
  assign n12577 = ( n160 & n12441 ) | ( n160 & n12568 ) | ( n12441 & n12568 ) ;
  assign n12578 = ( n12441 & ~n12464 ) | ( n12441 & n12568 ) | ( ~n12464 & n12568 ) ;
  assign n12579 = ~n12577 & n12578 ;
  assign n12580 = n12573 | n12579 ;
  assign n12581 = n12205 &  n12465 ;
  assign n12574 = x92 | n12205 ;
  assign n12575 = x92 &  n12205 ;
  assign n12576 = ( n12574 & ~n12575 ) | ( n12574 & 1'b0 ) | ( ~n12575 & 1'b0 ) ;
  assign n12585 = ( n160 & n12440 ) | ( n160 & n12576 ) | ( n12440 & n12576 ) ;
  assign n12586 = ( n12440 & ~n12464 ) | ( n12440 & n12576 ) | ( ~n12464 & n12576 ) ;
  assign n12587 = ~n12585 & n12586 ;
  assign n12588 = n12581 | n12587 ;
  assign n12589 = n12213 &  n12465 ;
  assign n12582 = x91 | n12213 ;
  assign n12583 = x91 &  n12213 ;
  assign n12584 = ( n12582 & ~n12583 ) | ( n12582 & 1'b0 ) | ( ~n12583 & 1'b0 ) ;
  assign n12593 = ( n160 & n12439 ) | ( n160 & n12584 ) | ( n12439 & n12584 ) ;
  assign n12594 = ( n12439 & ~n12464 ) | ( n12439 & n12584 ) | ( ~n12464 & n12584 ) ;
  assign n12595 = ~n12593 & n12594 ;
  assign n12596 = n12589 | n12595 ;
  assign n12597 = n12221 &  n12465 ;
  assign n12590 = x90 | n12221 ;
  assign n12591 = x90 &  n12221 ;
  assign n12592 = ( n12590 & ~n12591 ) | ( n12590 & 1'b0 ) | ( ~n12591 & 1'b0 ) ;
  assign n12601 = ( n160 & n12438 ) | ( n160 & n12592 ) | ( n12438 & n12592 ) ;
  assign n12602 = ( n12438 & ~n12464 ) | ( n12438 & n12592 ) | ( ~n12464 & n12592 ) ;
  assign n12603 = ~n12601 & n12602 ;
  assign n12604 = n12597 | n12603 ;
  assign n12605 = n12229 &  n12465 ;
  assign n12598 = x89 | n12229 ;
  assign n12599 = x89 &  n12229 ;
  assign n12600 = ( n12598 & ~n12599 ) | ( n12598 & 1'b0 ) | ( ~n12599 & 1'b0 ) ;
  assign n12609 = ( n160 & n12437 ) | ( n160 & n12600 ) | ( n12437 & n12600 ) ;
  assign n12610 = ( n12437 & ~n12464 ) | ( n12437 & n12600 ) | ( ~n12464 & n12600 ) ;
  assign n12611 = ~n12609 & n12610 ;
  assign n12612 = n12605 | n12611 ;
  assign n12613 = n12237 &  n12465 ;
  assign n12606 = x88 | n12237 ;
  assign n12607 = x88 &  n12237 ;
  assign n12608 = ( n12606 & ~n12607 ) | ( n12606 & 1'b0 ) | ( ~n12607 & 1'b0 ) ;
  assign n12617 = ( n160 & n12436 ) | ( n160 & n12608 ) | ( n12436 & n12608 ) ;
  assign n12618 = ( n12436 & ~n12464 ) | ( n12436 & n12608 ) | ( ~n12464 & n12608 ) ;
  assign n12619 = ~n12617 & n12618 ;
  assign n12620 = n12613 | n12619 ;
  assign n12621 = n12245 &  n12465 ;
  assign n12614 = x87 | n12245 ;
  assign n12615 = x87 &  n12245 ;
  assign n12616 = ( n12614 & ~n12615 ) | ( n12614 & 1'b0 ) | ( ~n12615 & 1'b0 ) ;
  assign n12625 = ( n160 & n12435 ) | ( n160 & n12616 ) | ( n12435 & n12616 ) ;
  assign n12626 = ( n12435 & ~n12464 ) | ( n12435 & n12616 ) | ( ~n12464 & n12616 ) ;
  assign n12627 = ~n12625 & n12626 ;
  assign n12628 = n12621 | n12627 ;
  assign n12629 = n12253 &  n12465 ;
  assign n12622 = x86 | n12253 ;
  assign n12623 = x86 &  n12253 ;
  assign n12624 = ( n12622 & ~n12623 ) | ( n12622 & 1'b0 ) | ( ~n12623 & 1'b0 ) ;
  assign n12633 = ( n160 & n12434 ) | ( n160 & n12624 ) | ( n12434 & n12624 ) ;
  assign n12634 = ( n12434 & ~n12464 ) | ( n12434 & n12624 ) | ( ~n12464 & n12624 ) ;
  assign n12635 = ~n12633 & n12634 ;
  assign n12636 = n12629 | n12635 ;
  assign n12637 = n12261 &  n12465 ;
  assign n12630 = x85 | n12261 ;
  assign n12631 = x85 &  n12261 ;
  assign n12632 = ( n12630 & ~n12631 ) | ( n12630 & 1'b0 ) | ( ~n12631 & 1'b0 ) ;
  assign n12641 = ( n160 & n12433 ) | ( n160 & n12632 ) | ( n12433 & n12632 ) ;
  assign n12642 = ( n12433 & ~n12464 ) | ( n12433 & n12632 ) | ( ~n12464 & n12632 ) ;
  assign n12643 = ~n12641 & n12642 ;
  assign n12644 = n12637 | n12643 ;
  assign n12645 = n12269 &  n12465 ;
  assign n12638 = x84 | n12269 ;
  assign n12639 = x84 &  n12269 ;
  assign n12640 = ( n12638 & ~n12639 ) | ( n12638 & 1'b0 ) | ( ~n12639 & 1'b0 ) ;
  assign n12649 = ( n160 & n12432 ) | ( n160 & n12640 ) | ( n12432 & n12640 ) ;
  assign n12650 = ( n12432 & ~n12464 ) | ( n12432 & n12640 ) | ( ~n12464 & n12640 ) ;
  assign n12651 = ~n12649 & n12650 ;
  assign n12652 = n12645 | n12651 ;
  assign n12653 = n12277 &  n12465 ;
  assign n12646 = x83 | n12277 ;
  assign n12647 = x83 &  n12277 ;
  assign n12648 = ( n12646 & ~n12647 ) | ( n12646 & 1'b0 ) | ( ~n12647 & 1'b0 ) ;
  assign n12657 = ( n160 & n12431 ) | ( n160 & n12648 ) | ( n12431 & n12648 ) ;
  assign n12658 = ( n12431 & ~n12464 ) | ( n12431 & n12648 ) | ( ~n12464 & n12648 ) ;
  assign n12659 = ~n12657 & n12658 ;
  assign n12660 = n12653 | n12659 ;
  assign n12661 = n12285 &  n12465 ;
  assign n12654 = x82 | n12285 ;
  assign n12655 = x82 &  n12285 ;
  assign n12656 = ( n12654 & ~n12655 ) | ( n12654 & 1'b0 ) | ( ~n12655 & 1'b0 ) ;
  assign n12665 = ( n160 & n12430 ) | ( n160 & n12656 ) | ( n12430 & n12656 ) ;
  assign n12666 = ( n12430 & ~n12464 ) | ( n12430 & n12656 ) | ( ~n12464 & n12656 ) ;
  assign n12667 = ~n12665 & n12666 ;
  assign n12668 = n12661 | n12667 ;
  assign n12669 = n12293 &  n12465 ;
  assign n12662 = x81 | n12293 ;
  assign n12663 = x81 &  n12293 ;
  assign n12664 = ( n12662 & ~n12663 ) | ( n12662 & 1'b0 ) | ( ~n12663 & 1'b0 ) ;
  assign n12673 = ( n160 & n12429 ) | ( n160 & n12664 ) | ( n12429 & n12664 ) ;
  assign n12674 = ( n12429 & ~n12464 ) | ( n12429 & n12664 ) | ( ~n12464 & n12664 ) ;
  assign n12675 = ~n12673 & n12674 ;
  assign n12676 = n12669 | n12675 ;
  assign n12677 = n12301 &  n12465 ;
  assign n12670 = x80 | n12301 ;
  assign n12671 = x80 &  n12301 ;
  assign n12672 = ( n12670 & ~n12671 ) | ( n12670 & 1'b0 ) | ( ~n12671 & 1'b0 ) ;
  assign n12681 = ( n160 & n12428 ) | ( n160 & n12672 ) | ( n12428 & n12672 ) ;
  assign n12682 = ( n12428 & ~n12464 ) | ( n12428 & n12672 ) | ( ~n12464 & n12672 ) ;
  assign n12683 = ~n12681 & n12682 ;
  assign n12684 = n12677 | n12683 ;
  assign n12685 = n12309 &  n12465 ;
  assign n12678 = x79 | n12309 ;
  assign n12679 = x79 &  n12309 ;
  assign n12680 = ( n12678 & ~n12679 ) | ( n12678 & 1'b0 ) | ( ~n12679 & 1'b0 ) ;
  assign n12689 = ( n160 & n12427 ) | ( n160 & n12680 ) | ( n12427 & n12680 ) ;
  assign n12690 = ( n12427 & ~n12464 ) | ( n12427 & n12680 ) | ( ~n12464 & n12680 ) ;
  assign n12691 = ~n12689 & n12690 ;
  assign n12692 = n12685 | n12691 ;
  assign n12693 = n12317 &  n12465 ;
  assign n12686 = x78 | n12317 ;
  assign n12687 = x78 &  n12317 ;
  assign n12688 = ( n12686 & ~n12687 ) | ( n12686 & 1'b0 ) | ( ~n12687 & 1'b0 ) ;
  assign n12697 = ( n160 & n12426 ) | ( n160 & n12688 ) | ( n12426 & n12688 ) ;
  assign n12698 = ( n12426 & ~n12464 ) | ( n12426 & n12688 ) | ( ~n12464 & n12688 ) ;
  assign n12699 = ~n12697 & n12698 ;
  assign n12700 = n12693 | n12699 ;
  assign n12701 = n12325 &  n12465 ;
  assign n12694 = x77 | n12325 ;
  assign n12695 = x77 &  n12325 ;
  assign n12696 = ( n12694 & ~n12695 ) | ( n12694 & 1'b0 ) | ( ~n12695 & 1'b0 ) ;
  assign n12705 = ( n160 & n12425 ) | ( n160 & n12696 ) | ( n12425 & n12696 ) ;
  assign n12706 = ( n12425 & ~n12464 ) | ( n12425 & n12696 ) | ( ~n12464 & n12696 ) ;
  assign n12707 = ~n12705 & n12706 ;
  assign n12708 = n12701 | n12707 ;
  assign n12709 = n12333 &  n12465 ;
  assign n12702 = x76 | n12333 ;
  assign n12703 = x76 &  n12333 ;
  assign n12704 = ( n12702 & ~n12703 ) | ( n12702 & 1'b0 ) | ( ~n12703 & 1'b0 ) ;
  assign n12713 = ( n160 & n12424 ) | ( n160 & n12704 ) | ( n12424 & n12704 ) ;
  assign n12714 = ( n12424 & ~n12464 ) | ( n12424 & n12704 ) | ( ~n12464 & n12704 ) ;
  assign n12715 = ~n12713 & n12714 ;
  assign n12716 = n12709 | n12715 ;
  assign n12717 = n12341 &  n12465 ;
  assign n12710 = x75 | n12341 ;
  assign n12711 = x75 &  n12341 ;
  assign n12712 = ( n12710 & ~n12711 ) | ( n12710 & 1'b0 ) | ( ~n12711 & 1'b0 ) ;
  assign n12721 = ( n160 & n12423 ) | ( n160 & n12712 ) | ( n12423 & n12712 ) ;
  assign n12722 = ( n12423 & ~n12464 ) | ( n12423 & n12712 ) | ( ~n12464 & n12712 ) ;
  assign n12723 = ~n12721 & n12722 ;
  assign n12724 = n12717 | n12723 ;
  assign n12725 = n12349 &  n12465 ;
  assign n12718 = x74 | n12349 ;
  assign n12719 = x74 &  n12349 ;
  assign n12720 = ( n12718 & ~n12719 ) | ( n12718 & 1'b0 ) | ( ~n12719 & 1'b0 ) ;
  assign n12729 = ( n160 & n12422 ) | ( n160 & n12720 ) | ( n12422 & n12720 ) ;
  assign n12730 = ( n12422 & ~n12464 ) | ( n12422 & n12720 ) | ( ~n12464 & n12720 ) ;
  assign n12731 = ~n12729 & n12730 ;
  assign n12732 = n12725 | n12731 ;
  assign n12733 = n12357 &  n12465 ;
  assign n12726 = x73 | n12357 ;
  assign n12727 = x73 &  n12357 ;
  assign n12728 = ( n12726 & ~n12727 ) | ( n12726 & 1'b0 ) | ( ~n12727 & 1'b0 ) ;
  assign n12737 = ( n160 & n12421 ) | ( n160 & n12728 ) | ( n12421 & n12728 ) ;
  assign n12738 = ( n12421 & ~n12464 ) | ( n12421 & n12728 ) | ( ~n12464 & n12728 ) ;
  assign n12739 = ~n12737 & n12738 ;
  assign n12740 = n12733 | n12739 ;
  assign n12741 = n12365 &  n12465 ;
  assign n12734 = x72 | n12365 ;
  assign n12735 = x72 &  n12365 ;
  assign n12736 = ( n12734 & ~n12735 ) | ( n12734 & 1'b0 ) | ( ~n12735 & 1'b0 ) ;
  assign n12745 = ( n160 & n12420 ) | ( n160 & n12736 ) | ( n12420 & n12736 ) ;
  assign n12746 = ( n12420 & ~n12464 ) | ( n12420 & n12736 ) | ( ~n12464 & n12736 ) ;
  assign n12747 = ~n12745 & n12746 ;
  assign n12748 = n12741 | n12747 ;
  assign n12749 = n12373 &  n12465 ;
  assign n12742 = x71 | n12373 ;
  assign n12743 = x71 &  n12373 ;
  assign n12744 = ( n12742 & ~n12743 ) | ( n12742 & 1'b0 ) | ( ~n12743 & 1'b0 ) ;
  assign n12753 = ( n160 & n12419 ) | ( n160 & n12744 ) | ( n12419 & n12744 ) ;
  assign n12754 = ( n12419 & ~n12464 ) | ( n12419 & n12744 ) | ( ~n12464 & n12744 ) ;
  assign n12755 = ~n12753 & n12754 ;
  assign n12756 = n12749 | n12755 ;
  assign n12757 = n12381 &  n12465 ;
  assign n12750 = x70 | n12381 ;
  assign n12751 = x70 &  n12381 ;
  assign n12752 = ( n12750 & ~n12751 ) | ( n12750 & 1'b0 ) | ( ~n12751 & 1'b0 ) ;
  assign n12761 = ( n160 & n12418 ) | ( n160 & n12752 ) | ( n12418 & n12752 ) ;
  assign n12762 = ( n12418 & ~n12464 ) | ( n12418 & n12752 ) | ( ~n12464 & n12752 ) ;
  assign n12763 = ~n12761 & n12762 ;
  assign n12764 = n12757 | n12763 ;
  assign n12765 = n12389 &  n12465 ;
  assign n12758 = x69 | n12389 ;
  assign n12759 = x69 &  n12389 ;
  assign n12760 = ( n12758 & ~n12759 ) | ( n12758 & 1'b0 ) | ( ~n12759 & 1'b0 ) ;
  assign n12769 = ( n160 & n12417 ) | ( n160 & n12760 ) | ( n12417 & n12760 ) ;
  assign n12770 = ( n12417 & ~n12464 ) | ( n12417 & n12760 ) | ( ~n12464 & n12760 ) ;
  assign n12771 = ~n12769 & n12770 ;
  assign n12772 = n12765 | n12771 ;
  assign n12773 = n12397 &  n12465 ;
  assign n12766 = x68 | n12397 ;
  assign n12767 = x68 &  n12397 ;
  assign n12768 = ( n12766 & ~n12767 ) | ( n12766 & 1'b0 ) | ( ~n12767 & 1'b0 ) ;
  assign n12777 = ( n160 & n12416 ) | ( n160 & n12768 ) | ( n12416 & n12768 ) ;
  assign n12778 = ( n12416 & ~n12464 ) | ( n12416 & n12768 ) | ( ~n12464 & n12768 ) ;
  assign n12779 = ~n12777 & n12778 ;
  assign n12780 = n12773 | n12779 ;
  assign n12781 = n12402 &  n12465 ;
  assign n12774 = x67 | n12402 ;
  assign n12775 = x67 &  n12402 ;
  assign n12776 = ( n12774 & ~n12775 ) | ( n12774 & 1'b0 ) | ( ~n12775 & 1'b0 ) ;
  assign n12785 = ( n160 & n12415 ) | ( n160 & n12776 ) | ( n12415 & n12776 ) ;
  assign n12786 = ( n12415 & ~n12464 ) | ( n12415 & n12776 ) | ( ~n12464 & n12776 ) ;
  assign n12787 = ~n12785 & n12786 ;
  assign n12788 = n12781 | n12787 ;
  assign n12789 = n12408 &  n12465 ;
  assign n12782 = x66 | n12408 ;
  assign n12783 = x66 &  n12408 ;
  assign n12784 = ( n12782 & ~n12783 ) | ( n12782 & 1'b0 ) | ( ~n12783 & 1'b0 ) ;
  assign n12790 = ( n12414 & ~n160 ) | ( n12414 & n12784 ) | ( ~n160 & n12784 ) ;
  assign n12791 = ( n12414 & n12464 ) | ( n12414 & n12784 ) | ( n12464 & n12784 ) ;
  assign n12792 = ( n12790 & ~n12791 ) | ( n12790 & 1'b0 ) | ( ~n12791 & 1'b0 ) ;
  assign n12793 = n12789 | n12792 ;
  assign n12794 = n12412 &  n12465 ;
  assign n12795 = ( x65 & ~x13 ) | ( x65 & n12409 ) | ( ~x13 & n12409 ) ;
  assign n12796 = ( x13 & ~n12409 ) | ( x13 & x65 ) | ( ~n12409 & x65 ) ;
  assign n12797 = ( n12795 & ~x65 ) | ( n12795 & n12796 ) | ( ~x65 & n12796 ) ;
  assign n12798 = ( n12413 & ~n12464 ) | ( n12413 & n12797 ) | ( ~n12464 & n12797 ) ;
  assign n12799 = ( n160 & n12413 ) | ( n160 & n12797 ) | ( n12413 & n12797 ) ;
  assign n12800 = ( n12798 & ~n12799 ) | ( n12798 & 1'b0 ) | ( ~n12799 & 1'b0 ) ;
  assign n12801 = n12794 | n12800 ;
  assign n12802 = ( x64 & ~x116 ) | ( x64 & 1'b0 ) | ( ~x116 & 1'b0 ) ;
  assign n12803 = ( n229 & ~n239 ) | ( n229 & n12802 ) | ( ~n239 & n12802 ) ;
  assign n12804 = ~n229 & n12803 ;
  assign n12805 = n12464 &  n12804 ;
  assign n12806 = ( x12 & ~n12804 ) | ( x12 & n12805 ) | ( ~n12804 & n12805 ) ;
  assign n12807 = ~n158 & n12413 ;
  assign n12808 = ~n269 & n12807 ;
  assign n12809 = ~n12464 & n12808 ;
  assign n12810 = n12806 | n12809 ;
  assign n12811 = ~x11 & x64 ;
  assign n12812 = ( x65 & ~n12810 ) | ( x65 & n12811 ) | ( ~n12810 & n12811 ) ;
  assign n12813 = ( x66 & ~n12801 ) | ( x66 & n12812 ) | ( ~n12801 & n12812 ) ;
  assign n12814 = ( x67 & ~n12793 ) | ( x67 & n12813 ) | ( ~n12793 & n12813 ) ;
  assign n12815 = ( x68 & ~n12788 ) | ( x68 & n12814 ) | ( ~n12788 & n12814 ) ;
  assign n12816 = ( x69 & ~n12780 ) | ( x69 & n12815 ) | ( ~n12780 & n12815 ) ;
  assign n12817 = ( x70 & ~n12772 ) | ( x70 & n12816 ) | ( ~n12772 & n12816 ) ;
  assign n12818 = ( x71 & ~n12764 ) | ( x71 & n12817 ) | ( ~n12764 & n12817 ) ;
  assign n12819 = ( x72 & ~n12756 ) | ( x72 & n12818 ) | ( ~n12756 & n12818 ) ;
  assign n12820 = ( x73 & ~n12748 ) | ( x73 & n12819 ) | ( ~n12748 & n12819 ) ;
  assign n12821 = ( x74 & ~n12740 ) | ( x74 & n12820 ) | ( ~n12740 & n12820 ) ;
  assign n12822 = ( x75 & ~n12732 ) | ( x75 & n12821 ) | ( ~n12732 & n12821 ) ;
  assign n12823 = ( x76 & ~n12724 ) | ( x76 & n12822 ) | ( ~n12724 & n12822 ) ;
  assign n12824 = ( x77 & ~n12716 ) | ( x77 & n12823 ) | ( ~n12716 & n12823 ) ;
  assign n12825 = ( x78 & ~n12708 ) | ( x78 & n12824 ) | ( ~n12708 & n12824 ) ;
  assign n12826 = ( x79 & ~n12700 ) | ( x79 & n12825 ) | ( ~n12700 & n12825 ) ;
  assign n12827 = ( x80 & ~n12692 ) | ( x80 & n12826 ) | ( ~n12692 & n12826 ) ;
  assign n12828 = ( x81 & ~n12684 ) | ( x81 & n12827 ) | ( ~n12684 & n12827 ) ;
  assign n12829 = ( x82 & ~n12676 ) | ( x82 & n12828 ) | ( ~n12676 & n12828 ) ;
  assign n12830 = ( x83 & ~n12668 ) | ( x83 & n12829 ) | ( ~n12668 & n12829 ) ;
  assign n12831 = ( x84 & ~n12660 ) | ( x84 & n12830 ) | ( ~n12660 & n12830 ) ;
  assign n12832 = ( x85 & ~n12652 ) | ( x85 & n12831 ) | ( ~n12652 & n12831 ) ;
  assign n12833 = ( x86 & ~n12644 ) | ( x86 & n12832 ) | ( ~n12644 & n12832 ) ;
  assign n12834 = ( x87 & ~n12636 ) | ( x87 & n12833 ) | ( ~n12636 & n12833 ) ;
  assign n12835 = ( x88 & ~n12628 ) | ( x88 & n12834 ) | ( ~n12628 & n12834 ) ;
  assign n12836 = ( x89 & ~n12620 ) | ( x89 & n12835 ) | ( ~n12620 & n12835 ) ;
  assign n12837 = ( x90 & ~n12612 ) | ( x90 & n12836 ) | ( ~n12612 & n12836 ) ;
  assign n12838 = ( x91 & ~n12604 ) | ( x91 & n12837 ) | ( ~n12604 & n12837 ) ;
  assign n12839 = ( x92 & ~n12596 ) | ( x92 & n12838 ) | ( ~n12596 & n12838 ) ;
  assign n12840 = ( x93 & ~n12588 ) | ( x93 & n12839 ) | ( ~n12588 & n12839 ) ;
  assign n12841 = ( x94 & ~n12580 ) | ( x94 & n12840 ) | ( ~n12580 & n12840 ) ;
  assign n12842 = ( x95 & ~n12572 ) | ( x95 & n12841 ) | ( ~n12572 & n12841 ) ;
  assign n12843 = ( x96 & ~n12564 ) | ( x96 & n12842 ) | ( ~n12564 & n12842 ) ;
  assign n12844 = ( x97 & ~n12556 ) | ( x97 & n12843 ) | ( ~n12556 & n12843 ) ;
  assign n12845 = ( x98 & ~n12548 ) | ( x98 & n12844 ) | ( ~n12548 & n12844 ) ;
  assign n12846 = ( x99 & ~n12540 ) | ( x99 & n12845 ) | ( ~n12540 & n12845 ) ;
  assign n12847 = ( x100 & ~n12532 ) | ( x100 & n12846 ) | ( ~n12532 & n12846 ) ;
  assign n12848 = ( x101 & ~n12524 ) | ( x101 & n12847 ) | ( ~n12524 & n12847 ) ;
  assign n12849 = ( x102 & ~n12516 ) | ( x102 & n12848 ) | ( ~n12516 & n12848 ) ;
  assign n12850 = ( x103 & ~n12508 ) | ( x103 & n12849 ) | ( ~n12508 & n12849 ) ;
  assign n12851 = ( x104 & ~n12500 ) | ( x104 & n12850 ) | ( ~n12500 & n12850 ) ;
  assign n12852 = ( x105 & ~n12492 ) | ( x105 & n12851 ) | ( ~n12492 & n12851 ) ;
  assign n12853 = ( x106 & ~n12484 ) | ( x106 & n12852 ) | ( ~n12484 & n12852 ) ;
  assign n12857 = ( x107 & ~n12476 ) | ( x107 & n12853 ) | ( ~n12476 & n12853 ) ;
  assign n12925 = ( x108 & ~n12865 ) | ( x108 & n12857 ) | ( ~n12865 & n12857 ) ;
  assign n12926 = ( x109 & ~n12924 ) | ( x109 & n12925 ) | ( ~n12924 & n12925 ) ;
  assign n12927 = ( x110 & ~n12919 ) | ( x110 & n12926 ) | ( ~n12919 & n12926 ) ;
  assign n12928 = ( x111 & ~n12911 ) | ( x111 & n12927 ) | ( ~n12911 & n12927 ) ;
  assign n12929 = ( x112 & ~n12903 ) | ( x112 & n12928 ) | ( ~n12903 & n12928 ) ;
  assign n12930 = ( x113 & ~n12895 ) | ( x113 & n12929 ) | ( ~n12895 & n12929 ) ;
  assign n12931 = ( x114 & ~n12887 ) | ( x114 & n12930 ) | ( ~n12887 & n12930 ) ;
  assign n12932 = ( x115 & ~n12879 ) | ( x115 & n12931 ) | ( ~n12879 & n12931 ) ;
  assign n12933 = n12032 &  n12465 ;
  assign n12934 = ( n160 & n12032 ) | ( n160 & n12463 ) | ( n12032 & n12463 ) ;
  assign n12935 = ( x115 & ~n12934 ) | ( x115 & n12032 ) | ( ~n12934 & n12032 ) ;
  assign n12936 = ~x115 & n12935 ;
  assign n12937 = n12933 | n12936 ;
  assign n12938 = ~x116 & n12937 ;
  assign n12939 = ( x116 & ~n12933 ) | ( x116 & 1'b0 ) | ( ~n12933 & 1'b0 ) ;
  assign n12940 = ~n12936 & n12939 ;
  assign n12941 = n425 | n12940 ;
  assign n12942 = n12938 | n12941 ;
  assign n12943 = n12932 | n12942 ;
  assign n12944 = ~n12937 |  n160 ;
  assign n13360 = n12879 &  n12944 ;
  assign n13361 = n12943 &  n13360 ;
  assign n13357 = x115 | n12879 ;
  assign n13358 = x115 &  n12879 ;
  assign n13359 = ( n13357 & ~n13358 ) | ( n13357 & 1'b0 ) | ( ~n13358 & 1'b0 ) ;
  assign n13362 = n12931 &  n13359 ;
  assign n12945 = n12943 &  n12944 ;
  assign n13363 = ( n12931 & ~n12945 ) | ( n12931 & n13359 ) | ( ~n12945 & n13359 ) ;
  assign n13364 = ( n13361 & ~n13362 ) | ( n13361 & n13363 ) | ( ~n13362 & n13363 ) ;
  assign n13368 = n12887 &  n12944 ;
  assign n13369 = n12943 &  n13368 ;
  assign n13354 = x114 | n12887 ;
  assign n13355 = x114 &  n12887 ;
  assign n13356 = ( n13354 & ~n13355 ) | ( n13354 & 1'b0 ) | ( ~n13355 & 1'b0 ) ;
  assign n13370 = n12930 &  n13356 ;
  assign n13371 = ( n12930 & ~n12945 ) | ( n12930 & n13356 ) | ( ~n12945 & n13356 ) ;
  assign n13372 = ( n13369 & ~n13370 ) | ( n13369 & n13371 ) | ( ~n13370 & n13371 ) ;
  assign n13376 = n12895 &  n12944 ;
  assign n13377 = n12943 &  n13376 ;
  assign n13365 = x113 | n12895 ;
  assign n13366 = x113 &  n12895 ;
  assign n13367 = ( n13365 & ~n13366 ) | ( n13365 & 1'b0 ) | ( ~n13366 & 1'b0 ) ;
  assign n13378 = n12929 &  n13367 ;
  assign n13379 = ( n12929 & ~n12945 ) | ( n12929 & n13367 ) | ( ~n12945 & n13367 ) ;
  assign n13380 = ( n13377 & ~n13378 ) | ( n13377 & n13379 ) | ( ~n13378 & n13379 ) ;
  assign n13384 = n12903 &  n12944 ;
  assign n13385 = n12943 &  n13384 ;
  assign n13373 = x112 | n12903 ;
  assign n13374 = x112 &  n12903 ;
  assign n13375 = ( n13373 & ~n13374 ) | ( n13373 & 1'b0 ) | ( ~n13374 & 1'b0 ) ;
  assign n13386 = n12928 &  n13375 ;
  assign n13387 = ( n12928 & ~n12945 ) | ( n12928 & n13375 ) | ( ~n12945 & n13375 ) ;
  assign n13388 = ( n13385 & ~n13386 ) | ( n13385 & n13387 ) | ( ~n13386 & n13387 ) ;
  assign n13392 = n12911 &  n12944 ;
  assign n13393 = n12943 &  n13392 ;
  assign n13381 = x111 | n12911 ;
  assign n13382 = x111 &  n12911 ;
  assign n13383 = ( n13381 & ~n13382 ) | ( n13381 & 1'b0 ) | ( ~n13382 & 1'b0 ) ;
  assign n13394 = n12927 &  n13383 ;
  assign n13395 = ( n12927 & ~n12945 ) | ( n12927 & n13383 ) | ( ~n12945 & n13383 ) ;
  assign n13396 = ( n13393 & ~n13394 ) | ( n13393 & n13395 ) | ( ~n13394 & n13395 ) ;
  assign n13397 = n12919 &  n12944 ;
  assign n13398 = n12943 &  n13397 ;
  assign n13389 = x110 | n12919 ;
  assign n13390 = x110 &  n12919 ;
  assign n13391 = ( n13389 & ~n13390 ) | ( n13389 & 1'b0 ) | ( ~n13390 & 1'b0 ) ;
  assign n13400 = ( n12926 & n12945 ) | ( n12926 & n13391 ) | ( n12945 & n13391 ) ;
  assign n13399 = n12926 | n13391 ;
  assign n13401 = ( n13398 & ~n13400 ) | ( n13398 & n13399 ) | ( ~n13400 & n13399 ) ;
  assign n13346 = n12924 &  n12944 ;
  assign n13347 = n12943 &  n13346 ;
  assign n13343 = x109 | n12924 ;
  assign n13344 = x109 &  n12924 ;
  assign n13345 = ( n13343 & ~n13344 ) | ( n13343 & 1'b0 ) | ( ~n13344 & 1'b0 ) ;
  assign n13349 = ( n12925 & n12945 ) | ( n12925 & n13345 ) | ( n12945 & n13345 ) ;
  assign n13348 = n12925 | n13345 ;
  assign n13350 = ( n13347 & ~n13349 ) | ( n13347 & n13348 ) | ( ~n13349 & n13348 ) ;
  assign n12946 = n12865 &  n12944 ;
  assign n12947 = n12943 &  n12946 ;
  assign n12866 = x108 | n12865 ;
  assign n12867 = x108 &  n12865 ;
  assign n12868 = ( n12866 & ~n12867 ) | ( n12866 & 1'b0 ) | ( ~n12867 & 1'b0 ) ;
  assign n12949 = ( n12857 & n12868 ) | ( n12857 & n12945 ) | ( n12868 & n12945 ) ;
  assign n12948 = n12857 | n12868 ;
  assign n12950 = ( n12947 & ~n12949 ) | ( n12947 & n12948 ) | ( ~n12949 & n12948 ) ;
  assign n12954 = n12476 &  n12944 ;
  assign n12955 = n12943 &  n12954 ;
  assign n12854 = x107 | n12476 ;
  assign n12855 = x107 &  n12476 ;
  assign n12856 = ( n12854 & ~n12855 ) | ( n12854 & 1'b0 ) | ( ~n12855 & 1'b0 ) ;
  assign n12956 = n12853 &  n12856 ;
  assign n12957 = ( n12853 & ~n12945 ) | ( n12853 & n12856 ) | ( ~n12945 & n12856 ) ;
  assign n12958 = ( n12955 & ~n12956 ) | ( n12955 & n12957 ) | ( ~n12956 & n12957 ) ;
  assign n12962 = n12484 &  n12944 ;
  assign n12963 = n12943 &  n12962 ;
  assign n12951 = x106 | n12484 ;
  assign n12952 = x106 &  n12484 ;
  assign n12953 = ( n12951 & ~n12952 ) | ( n12951 & 1'b0 ) | ( ~n12952 & 1'b0 ) ;
  assign n12965 = ( n12852 & n12945 ) | ( n12852 & n12953 ) | ( n12945 & n12953 ) ;
  assign n12964 = n12852 | n12953 ;
  assign n12966 = ( n12963 & ~n12965 ) | ( n12963 & n12964 ) | ( ~n12965 & n12964 ) ;
  assign n12970 = n12492 &  n12944 ;
  assign n12971 = n12943 &  n12970 ;
  assign n12959 = x105 | n12492 ;
  assign n12960 = x105 &  n12492 ;
  assign n12961 = ( n12959 & ~n12960 ) | ( n12959 & 1'b0 ) | ( ~n12960 & 1'b0 ) ;
  assign n12973 = ( n12851 & n12945 ) | ( n12851 & n12961 ) | ( n12945 & n12961 ) ;
  assign n12972 = n12851 | n12961 ;
  assign n12974 = ( n12971 & ~n12973 ) | ( n12971 & n12972 ) | ( ~n12973 & n12972 ) ;
  assign n12978 = n12500 &  n12944 ;
  assign n12979 = n12943 &  n12978 ;
  assign n12967 = x104 | n12500 ;
  assign n12968 = x104 &  n12500 ;
  assign n12969 = ( n12967 & ~n12968 ) | ( n12967 & 1'b0 ) | ( ~n12968 & 1'b0 ) ;
  assign n12981 = ( n12850 & n12945 ) | ( n12850 & n12969 ) | ( n12945 & n12969 ) ;
  assign n12980 = n12850 | n12969 ;
  assign n12982 = ( n12979 & ~n12981 ) | ( n12979 & n12980 ) | ( ~n12981 & n12980 ) ;
  assign n12986 = n12508 &  n12944 ;
  assign n12987 = n12943 &  n12986 ;
  assign n12975 = x103 | n12508 ;
  assign n12976 = x103 &  n12508 ;
  assign n12977 = ( n12975 & ~n12976 ) | ( n12975 & 1'b0 ) | ( ~n12976 & 1'b0 ) ;
  assign n12989 = ( n12849 & n12945 ) | ( n12849 & n12977 ) | ( n12945 & n12977 ) ;
  assign n12988 = n12849 | n12977 ;
  assign n12990 = ( n12987 & ~n12989 ) | ( n12987 & n12988 ) | ( ~n12989 & n12988 ) ;
  assign n12994 = n12516 &  n12944 ;
  assign n12995 = n12943 &  n12994 ;
  assign n12983 = x102 | n12516 ;
  assign n12984 = x102 &  n12516 ;
  assign n12985 = ( n12983 & ~n12984 ) | ( n12983 & 1'b0 ) | ( ~n12984 & 1'b0 ) ;
  assign n12997 = ( n12848 & n12945 ) | ( n12848 & n12985 ) | ( n12945 & n12985 ) ;
  assign n12996 = n12848 | n12985 ;
  assign n12998 = ( n12995 & ~n12997 ) | ( n12995 & n12996 ) | ( ~n12997 & n12996 ) ;
  assign n13002 = n12524 &  n12944 ;
  assign n13003 = n12943 &  n13002 ;
  assign n12991 = x101 | n12524 ;
  assign n12992 = x101 &  n12524 ;
  assign n12993 = ( n12991 & ~n12992 ) | ( n12991 & 1'b0 ) | ( ~n12992 & 1'b0 ) ;
  assign n13005 = ( n12847 & n12945 ) | ( n12847 & n12993 ) | ( n12945 & n12993 ) ;
  assign n13004 = n12847 | n12993 ;
  assign n13006 = ( n13003 & ~n13005 ) | ( n13003 & n13004 ) | ( ~n13005 & n13004 ) ;
  assign n13010 = n12532 &  n12944 ;
  assign n13011 = n12943 &  n13010 ;
  assign n12999 = x100 | n12532 ;
  assign n13000 = x100 &  n12532 ;
  assign n13001 = ( n12999 & ~n13000 ) | ( n12999 & 1'b0 ) | ( ~n13000 & 1'b0 ) ;
  assign n13013 = ( n12846 & n12945 ) | ( n12846 & n13001 ) | ( n12945 & n13001 ) ;
  assign n13012 = n12846 | n13001 ;
  assign n13014 = ( n13011 & ~n13013 ) | ( n13011 & n13012 ) | ( ~n13013 & n13012 ) ;
  assign n13018 = n12540 &  n12944 ;
  assign n13019 = n12943 &  n13018 ;
  assign n13007 = x99 | n12540 ;
  assign n13008 = x99 &  n12540 ;
  assign n13009 = ( n13007 & ~n13008 ) | ( n13007 & 1'b0 ) | ( ~n13008 & 1'b0 ) ;
  assign n13021 = ( n12845 & n12945 ) | ( n12845 & n13009 ) | ( n12945 & n13009 ) ;
  assign n13020 = n12845 | n13009 ;
  assign n13022 = ( n13019 & ~n13021 ) | ( n13019 & n13020 ) | ( ~n13021 & n13020 ) ;
  assign n13026 = n12548 &  n12944 ;
  assign n13027 = n12943 &  n13026 ;
  assign n13015 = x98 | n12548 ;
  assign n13016 = x98 &  n12548 ;
  assign n13017 = ( n13015 & ~n13016 ) | ( n13015 & 1'b0 ) | ( ~n13016 & 1'b0 ) ;
  assign n13029 = ( n12844 & n12945 ) | ( n12844 & n13017 ) | ( n12945 & n13017 ) ;
  assign n13028 = n12844 | n13017 ;
  assign n13030 = ( n13027 & ~n13029 ) | ( n13027 & n13028 ) | ( ~n13029 & n13028 ) ;
  assign n13034 = n12556 &  n12944 ;
  assign n13035 = n12943 &  n13034 ;
  assign n13023 = x97 | n12556 ;
  assign n13024 = x97 &  n12556 ;
  assign n13025 = ( n13023 & ~n13024 ) | ( n13023 & 1'b0 ) | ( ~n13024 & 1'b0 ) ;
  assign n13037 = ( n12843 & n12945 ) | ( n12843 & n13025 ) | ( n12945 & n13025 ) ;
  assign n13036 = n12843 | n13025 ;
  assign n13038 = ( n13035 & ~n13037 ) | ( n13035 & n13036 ) | ( ~n13037 & n13036 ) ;
  assign n13042 = n12564 &  n12944 ;
  assign n13043 = n12943 &  n13042 ;
  assign n13031 = x96 | n12564 ;
  assign n13032 = x96 &  n12564 ;
  assign n13033 = ( n13031 & ~n13032 ) | ( n13031 & 1'b0 ) | ( ~n13032 & 1'b0 ) ;
  assign n13045 = ( n12842 & n12945 ) | ( n12842 & n13033 ) | ( n12945 & n13033 ) ;
  assign n13044 = n12842 | n13033 ;
  assign n13046 = ( n13043 & ~n13045 ) | ( n13043 & n13044 ) | ( ~n13045 & n13044 ) ;
  assign n13050 = n12572 &  n12944 ;
  assign n13051 = n12943 &  n13050 ;
  assign n13039 = x95 | n12572 ;
  assign n13040 = x95 &  n12572 ;
  assign n13041 = ( n13039 & ~n13040 ) | ( n13039 & 1'b0 ) | ( ~n13040 & 1'b0 ) ;
  assign n13053 = ( n12841 & n12945 ) | ( n12841 & n13041 ) | ( n12945 & n13041 ) ;
  assign n13052 = n12841 | n13041 ;
  assign n13054 = ( n13051 & ~n13053 ) | ( n13051 & n13052 ) | ( ~n13053 & n13052 ) ;
  assign n13058 = n12580 &  n12944 ;
  assign n13059 = n12943 &  n13058 ;
  assign n13047 = x94 | n12580 ;
  assign n13048 = x94 &  n12580 ;
  assign n13049 = ( n13047 & ~n13048 ) | ( n13047 & 1'b0 ) | ( ~n13048 & 1'b0 ) ;
  assign n13061 = ( n12840 & n12945 ) | ( n12840 & n13049 ) | ( n12945 & n13049 ) ;
  assign n13060 = n12840 | n13049 ;
  assign n13062 = ( n13059 & ~n13061 ) | ( n13059 & n13060 ) | ( ~n13061 & n13060 ) ;
  assign n13066 = n12588 &  n12944 ;
  assign n13067 = n12943 &  n13066 ;
  assign n13055 = x93 | n12588 ;
  assign n13056 = x93 &  n12588 ;
  assign n13057 = ( n13055 & ~n13056 ) | ( n13055 & 1'b0 ) | ( ~n13056 & 1'b0 ) ;
  assign n13069 = ( n12839 & n12945 ) | ( n12839 & n13057 ) | ( n12945 & n13057 ) ;
  assign n13068 = n12839 | n13057 ;
  assign n13070 = ( n13067 & ~n13069 ) | ( n13067 & n13068 ) | ( ~n13069 & n13068 ) ;
  assign n13074 = n12596 &  n12944 ;
  assign n13075 = n12943 &  n13074 ;
  assign n13063 = x92 | n12596 ;
  assign n13064 = x92 &  n12596 ;
  assign n13065 = ( n13063 & ~n13064 ) | ( n13063 & 1'b0 ) | ( ~n13064 & 1'b0 ) ;
  assign n13077 = ( n12838 & n12945 ) | ( n12838 & n13065 ) | ( n12945 & n13065 ) ;
  assign n13076 = n12838 | n13065 ;
  assign n13078 = ( n13075 & ~n13077 ) | ( n13075 & n13076 ) | ( ~n13077 & n13076 ) ;
  assign n13082 = n12604 &  n12944 ;
  assign n13083 = n12943 &  n13082 ;
  assign n13071 = x91 | n12604 ;
  assign n13072 = x91 &  n12604 ;
  assign n13073 = ( n13071 & ~n13072 ) | ( n13071 & 1'b0 ) | ( ~n13072 & 1'b0 ) ;
  assign n13085 = ( n12837 & n12945 ) | ( n12837 & n13073 ) | ( n12945 & n13073 ) ;
  assign n13084 = n12837 | n13073 ;
  assign n13086 = ( n13083 & ~n13085 ) | ( n13083 & n13084 ) | ( ~n13085 & n13084 ) ;
  assign n13090 = n12612 &  n12944 ;
  assign n13091 = n12943 &  n13090 ;
  assign n13079 = x90 | n12612 ;
  assign n13080 = x90 &  n12612 ;
  assign n13081 = ( n13079 & ~n13080 ) | ( n13079 & 1'b0 ) | ( ~n13080 & 1'b0 ) ;
  assign n13093 = ( n12836 & n12945 ) | ( n12836 & n13081 ) | ( n12945 & n13081 ) ;
  assign n13092 = n12836 | n13081 ;
  assign n13094 = ( n13091 & ~n13093 ) | ( n13091 & n13092 ) | ( ~n13093 & n13092 ) ;
  assign n13098 = n12620 &  n12944 ;
  assign n13099 = n12943 &  n13098 ;
  assign n13087 = x89 | n12620 ;
  assign n13088 = x89 &  n12620 ;
  assign n13089 = ( n13087 & ~n13088 ) | ( n13087 & 1'b0 ) | ( ~n13088 & 1'b0 ) ;
  assign n13101 = ( n12835 & n12945 ) | ( n12835 & n13089 ) | ( n12945 & n13089 ) ;
  assign n13100 = n12835 | n13089 ;
  assign n13102 = ( n13099 & ~n13101 ) | ( n13099 & n13100 ) | ( ~n13101 & n13100 ) ;
  assign n13106 = n12628 &  n12944 ;
  assign n13107 = n12943 &  n13106 ;
  assign n13095 = x88 | n12628 ;
  assign n13096 = x88 &  n12628 ;
  assign n13097 = ( n13095 & ~n13096 ) | ( n13095 & 1'b0 ) | ( ~n13096 & 1'b0 ) ;
  assign n13109 = ( n12834 & n12945 ) | ( n12834 & n13097 ) | ( n12945 & n13097 ) ;
  assign n13108 = n12834 | n13097 ;
  assign n13110 = ( n13107 & ~n13109 ) | ( n13107 & n13108 ) | ( ~n13109 & n13108 ) ;
  assign n13114 = n12636 &  n12944 ;
  assign n13115 = n12943 &  n13114 ;
  assign n13103 = x87 | n12636 ;
  assign n13104 = x87 &  n12636 ;
  assign n13105 = ( n13103 & ~n13104 ) | ( n13103 & 1'b0 ) | ( ~n13104 & 1'b0 ) ;
  assign n13117 = ( n12833 & n12945 ) | ( n12833 & n13105 ) | ( n12945 & n13105 ) ;
  assign n13116 = n12833 | n13105 ;
  assign n13118 = ( n13115 & ~n13117 ) | ( n13115 & n13116 ) | ( ~n13117 & n13116 ) ;
  assign n13122 = n12644 &  n12944 ;
  assign n13123 = n12943 &  n13122 ;
  assign n13111 = x86 | n12644 ;
  assign n13112 = x86 &  n12644 ;
  assign n13113 = ( n13111 & ~n13112 ) | ( n13111 & 1'b0 ) | ( ~n13112 & 1'b0 ) ;
  assign n13125 = ( n12832 & n12945 ) | ( n12832 & n13113 ) | ( n12945 & n13113 ) ;
  assign n13124 = n12832 | n13113 ;
  assign n13126 = ( n13123 & ~n13125 ) | ( n13123 & n13124 ) | ( ~n13125 & n13124 ) ;
  assign n13130 = n12652 &  n12944 ;
  assign n13131 = n12943 &  n13130 ;
  assign n13119 = x85 | n12652 ;
  assign n13120 = x85 &  n12652 ;
  assign n13121 = ( n13119 & ~n13120 ) | ( n13119 & 1'b0 ) | ( ~n13120 & 1'b0 ) ;
  assign n13133 = ( n12831 & n12945 ) | ( n12831 & n13121 ) | ( n12945 & n13121 ) ;
  assign n13132 = n12831 | n13121 ;
  assign n13134 = ( n13131 & ~n13133 ) | ( n13131 & n13132 ) | ( ~n13133 & n13132 ) ;
  assign n13138 = n12660 &  n12944 ;
  assign n13139 = n12943 &  n13138 ;
  assign n13127 = x84 | n12660 ;
  assign n13128 = x84 &  n12660 ;
  assign n13129 = ( n13127 & ~n13128 ) | ( n13127 & 1'b0 ) | ( ~n13128 & 1'b0 ) ;
  assign n13141 = ( n12830 & n12945 ) | ( n12830 & n13129 ) | ( n12945 & n13129 ) ;
  assign n13140 = n12830 | n13129 ;
  assign n13142 = ( n13139 & ~n13141 ) | ( n13139 & n13140 ) | ( ~n13141 & n13140 ) ;
  assign n13146 = n12668 &  n12944 ;
  assign n13147 = n12943 &  n13146 ;
  assign n13135 = x83 | n12668 ;
  assign n13136 = x83 &  n12668 ;
  assign n13137 = ( n13135 & ~n13136 ) | ( n13135 & 1'b0 ) | ( ~n13136 & 1'b0 ) ;
  assign n13149 = ( n12829 & n12945 ) | ( n12829 & n13137 ) | ( n12945 & n13137 ) ;
  assign n13148 = n12829 | n13137 ;
  assign n13150 = ( n13147 & ~n13149 ) | ( n13147 & n13148 ) | ( ~n13149 & n13148 ) ;
  assign n13154 = n12676 &  n12944 ;
  assign n13155 = n12943 &  n13154 ;
  assign n13143 = x82 | n12676 ;
  assign n13144 = x82 &  n12676 ;
  assign n13145 = ( n13143 & ~n13144 ) | ( n13143 & 1'b0 ) | ( ~n13144 & 1'b0 ) ;
  assign n13157 = ( n12828 & n12945 ) | ( n12828 & n13145 ) | ( n12945 & n13145 ) ;
  assign n13156 = n12828 | n13145 ;
  assign n13158 = ( n13155 & ~n13157 ) | ( n13155 & n13156 ) | ( ~n13157 & n13156 ) ;
  assign n13162 = n12684 &  n12944 ;
  assign n13163 = n12943 &  n13162 ;
  assign n13151 = x81 | n12684 ;
  assign n13152 = x81 &  n12684 ;
  assign n13153 = ( n13151 & ~n13152 ) | ( n13151 & 1'b0 ) | ( ~n13152 & 1'b0 ) ;
  assign n13165 = ( n12827 & n12945 ) | ( n12827 & n13153 ) | ( n12945 & n13153 ) ;
  assign n13164 = n12827 | n13153 ;
  assign n13166 = ( n13163 & ~n13165 ) | ( n13163 & n13164 ) | ( ~n13165 & n13164 ) ;
  assign n13170 = n12692 &  n12944 ;
  assign n13171 = n12943 &  n13170 ;
  assign n13159 = x80 | n12692 ;
  assign n13160 = x80 &  n12692 ;
  assign n13161 = ( n13159 & ~n13160 ) | ( n13159 & 1'b0 ) | ( ~n13160 & 1'b0 ) ;
  assign n13173 = ( n12826 & n12945 ) | ( n12826 & n13161 ) | ( n12945 & n13161 ) ;
  assign n13172 = n12826 | n13161 ;
  assign n13174 = ( n13171 & ~n13173 ) | ( n13171 & n13172 ) | ( ~n13173 & n13172 ) ;
  assign n13178 = n12700 &  n12944 ;
  assign n13179 = n12943 &  n13178 ;
  assign n13167 = x79 | n12700 ;
  assign n13168 = x79 &  n12700 ;
  assign n13169 = ( n13167 & ~n13168 ) | ( n13167 & 1'b0 ) | ( ~n13168 & 1'b0 ) ;
  assign n13181 = ( n12825 & n12945 ) | ( n12825 & n13169 ) | ( n12945 & n13169 ) ;
  assign n13180 = n12825 | n13169 ;
  assign n13182 = ( n13179 & ~n13181 ) | ( n13179 & n13180 ) | ( ~n13181 & n13180 ) ;
  assign n13186 = n12708 &  n12944 ;
  assign n13187 = n12943 &  n13186 ;
  assign n13175 = x78 | n12708 ;
  assign n13176 = x78 &  n12708 ;
  assign n13177 = ( n13175 & ~n13176 ) | ( n13175 & 1'b0 ) | ( ~n13176 & 1'b0 ) ;
  assign n13189 = ( n12824 & n12945 ) | ( n12824 & n13177 ) | ( n12945 & n13177 ) ;
  assign n13188 = n12824 | n13177 ;
  assign n13190 = ( n13187 & ~n13189 ) | ( n13187 & n13188 ) | ( ~n13189 & n13188 ) ;
  assign n13194 = n12716 &  n12944 ;
  assign n13195 = n12943 &  n13194 ;
  assign n13183 = x77 | n12716 ;
  assign n13184 = x77 &  n12716 ;
  assign n13185 = ( n13183 & ~n13184 ) | ( n13183 & 1'b0 ) | ( ~n13184 & 1'b0 ) ;
  assign n13197 = ( n12823 & n12945 ) | ( n12823 & n13185 ) | ( n12945 & n13185 ) ;
  assign n13196 = n12823 | n13185 ;
  assign n13198 = ( n13195 & ~n13197 ) | ( n13195 & n13196 ) | ( ~n13197 & n13196 ) ;
  assign n13202 = n12724 &  n12944 ;
  assign n13203 = n12943 &  n13202 ;
  assign n13191 = x76 | n12724 ;
  assign n13192 = x76 &  n12724 ;
  assign n13193 = ( n13191 & ~n13192 ) | ( n13191 & 1'b0 ) | ( ~n13192 & 1'b0 ) ;
  assign n13205 = ( n12822 & n12945 ) | ( n12822 & n13193 ) | ( n12945 & n13193 ) ;
  assign n13204 = n12822 | n13193 ;
  assign n13206 = ( n13203 & ~n13205 ) | ( n13203 & n13204 ) | ( ~n13205 & n13204 ) ;
  assign n13210 = n12732 &  n12944 ;
  assign n13211 = n12943 &  n13210 ;
  assign n13199 = x75 | n12732 ;
  assign n13200 = x75 &  n12732 ;
  assign n13201 = ( n13199 & ~n13200 ) | ( n13199 & 1'b0 ) | ( ~n13200 & 1'b0 ) ;
  assign n13213 = ( n12821 & n12945 ) | ( n12821 & n13201 ) | ( n12945 & n13201 ) ;
  assign n13212 = n12821 | n13201 ;
  assign n13214 = ( n13211 & ~n13213 ) | ( n13211 & n13212 ) | ( ~n13213 & n13212 ) ;
  assign n13218 = n12740 &  n12944 ;
  assign n13219 = n12943 &  n13218 ;
  assign n13207 = x74 | n12740 ;
  assign n13208 = x74 &  n12740 ;
  assign n13209 = ( n13207 & ~n13208 ) | ( n13207 & 1'b0 ) | ( ~n13208 & 1'b0 ) ;
  assign n13221 = ( n12820 & n12945 ) | ( n12820 & n13209 ) | ( n12945 & n13209 ) ;
  assign n13220 = n12820 | n13209 ;
  assign n13222 = ( n13219 & ~n13221 ) | ( n13219 & n13220 ) | ( ~n13221 & n13220 ) ;
  assign n13226 = n12748 &  n12944 ;
  assign n13227 = n12943 &  n13226 ;
  assign n13215 = x73 | n12748 ;
  assign n13216 = x73 &  n12748 ;
  assign n13217 = ( n13215 & ~n13216 ) | ( n13215 & 1'b0 ) | ( ~n13216 & 1'b0 ) ;
  assign n13229 = ( n12819 & n12945 ) | ( n12819 & n13217 ) | ( n12945 & n13217 ) ;
  assign n13228 = n12819 | n13217 ;
  assign n13230 = ( n13227 & ~n13229 ) | ( n13227 & n13228 ) | ( ~n13229 & n13228 ) ;
  assign n13234 = n12756 &  n12944 ;
  assign n13235 = n12943 &  n13234 ;
  assign n13223 = x72 | n12756 ;
  assign n13224 = x72 &  n12756 ;
  assign n13225 = ( n13223 & ~n13224 ) | ( n13223 & 1'b0 ) | ( ~n13224 & 1'b0 ) ;
  assign n13237 = ( n12818 & n12945 ) | ( n12818 & n13225 ) | ( n12945 & n13225 ) ;
  assign n13236 = n12818 | n13225 ;
  assign n13238 = ( n13235 & ~n13237 ) | ( n13235 & n13236 ) | ( ~n13237 & n13236 ) ;
  assign n13242 = n12764 &  n12944 ;
  assign n13243 = n12943 &  n13242 ;
  assign n13231 = x71 | n12764 ;
  assign n13232 = x71 &  n12764 ;
  assign n13233 = ( n13231 & ~n13232 ) | ( n13231 & 1'b0 ) | ( ~n13232 & 1'b0 ) ;
  assign n13245 = ( n12817 & n12945 ) | ( n12817 & n13233 ) | ( n12945 & n13233 ) ;
  assign n13244 = n12817 | n13233 ;
  assign n13246 = ( n13243 & ~n13245 ) | ( n13243 & n13244 ) | ( ~n13245 & n13244 ) ;
  assign n13250 = n12772 &  n12944 ;
  assign n13251 = n12943 &  n13250 ;
  assign n13239 = x70 | n12772 ;
  assign n13240 = x70 &  n12772 ;
  assign n13241 = ( n13239 & ~n13240 ) | ( n13239 & 1'b0 ) | ( ~n13240 & 1'b0 ) ;
  assign n13253 = ( n12816 & n12945 ) | ( n12816 & n13241 ) | ( n12945 & n13241 ) ;
  assign n13252 = n12816 | n13241 ;
  assign n13254 = ( n13251 & ~n13253 ) | ( n13251 & n13252 ) | ( ~n13253 & n13252 ) ;
  assign n13258 = n12780 &  n12944 ;
  assign n13259 = n12943 &  n13258 ;
  assign n13247 = x69 | n12780 ;
  assign n13248 = x69 &  n12780 ;
  assign n13249 = ( n13247 & ~n13248 ) | ( n13247 & 1'b0 ) | ( ~n13248 & 1'b0 ) ;
  assign n13261 = ( n12815 & n12945 ) | ( n12815 & n13249 ) | ( n12945 & n13249 ) ;
  assign n13260 = n12815 | n13249 ;
  assign n13262 = ( n13259 & ~n13261 ) | ( n13259 & n13260 ) | ( ~n13261 & n13260 ) ;
  assign n13266 = n12788 &  n12944 ;
  assign n13267 = n12943 &  n13266 ;
  assign n13255 = x68 | n12788 ;
  assign n13256 = x68 &  n12788 ;
  assign n13257 = ( n13255 & ~n13256 ) | ( n13255 & 1'b0 ) | ( ~n13256 & 1'b0 ) ;
  assign n13269 = ( n12814 & n12945 ) | ( n12814 & n13257 ) | ( n12945 & n13257 ) ;
  assign n13268 = n12814 | n13257 ;
  assign n13270 = ( n13267 & ~n13269 ) | ( n13267 & n13268 ) | ( ~n13269 & n13268 ) ;
  assign n13274 = n12793 &  n12944 ;
  assign n13275 = n12943 &  n13274 ;
  assign n13263 = x67 | n12793 ;
  assign n13264 = x67 &  n12793 ;
  assign n13265 = ( n13263 & ~n13264 ) | ( n13263 & 1'b0 ) | ( ~n13264 & 1'b0 ) ;
  assign n13277 = ( n12813 & n12945 ) | ( n12813 & n13265 ) | ( n12945 & n13265 ) ;
  assign n13276 = n12813 | n13265 ;
  assign n13278 = ( n13275 & ~n13277 ) | ( n13275 & n13276 ) | ( ~n13277 & n13276 ) ;
  assign n13279 = n12801 &  n12944 ;
  assign n13280 = n12943 &  n13279 ;
  assign n13271 = x66 | n12801 ;
  assign n13272 = x66 &  n12801 ;
  assign n13273 = ( n13271 & ~n13272 ) | ( n13271 & 1'b0 ) | ( ~n13272 & 1'b0 ) ;
  assign n13281 = n12812 &  n13273 ;
  assign n13282 = ( n12812 & ~n12945 ) | ( n12812 & n13273 ) | ( ~n12945 & n13273 ) ;
  assign n13283 = ( n13280 & ~n13281 ) | ( n13280 & n13282 ) | ( ~n13281 & n13282 ) ;
  assign n13284 = ( n12810 & ~x65 ) | ( n12810 & n12811 ) | ( ~x65 & n12811 ) ;
  assign n13285 = ( n12812 & ~n12811 ) | ( n12812 & n13284 ) | ( ~n12811 & n13284 ) ;
  assign n13286 = ~n12945 & n13285 ;
  assign n13287 = n12810 &  n12944 ;
  assign n13288 = n12943 &  n13287 ;
  assign n13289 = n13286 | n13288 ;
  assign n13290 = ( x64 & ~n12945 ) | ( x64 & 1'b0 ) | ( ~n12945 & 1'b0 ) ;
  assign n13291 = ( x11 & ~n13290 ) | ( x11 & 1'b0 ) | ( ~n13290 & 1'b0 ) ;
  assign n13292 = ( n12811 & ~n12945 ) | ( n12811 & 1'b0 ) | ( ~n12945 & 1'b0 ) ;
  assign n13293 = n13291 | n13292 ;
  assign n13294 = ~x10 & x64 ;
  assign n13295 = ( x65 & ~n13293 ) | ( x65 & n13294 ) | ( ~n13293 & n13294 ) ;
  assign n13296 = ( x66 & ~n13289 ) | ( x66 & n13295 ) | ( ~n13289 & n13295 ) ;
  assign n13297 = ( x67 & ~n13283 ) | ( x67 & n13296 ) | ( ~n13283 & n13296 ) ;
  assign n13298 = ( x68 & ~n13278 ) | ( x68 & n13297 ) | ( ~n13278 & n13297 ) ;
  assign n13299 = ( x69 & ~n13270 ) | ( x69 & n13298 ) | ( ~n13270 & n13298 ) ;
  assign n13300 = ( x70 & ~n13262 ) | ( x70 & n13299 ) | ( ~n13262 & n13299 ) ;
  assign n13301 = ( x71 & ~n13254 ) | ( x71 & n13300 ) | ( ~n13254 & n13300 ) ;
  assign n13302 = ( x72 & ~n13246 ) | ( x72 & n13301 ) | ( ~n13246 & n13301 ) ;
  assign n13303 = ( x73 & ~n13238 ) | ( x73 & n13302 ) | ( ~n13238 & n13302 ) ;
  assign n13304 = ( x74 & ~n13230 ) | ( x74 & n13303 ) | ( ~n13230 & n13303 ) ;
  assign n13305 = ( x75 & ~n13222 ) | ( x75 & n13304 ) | ( ~n13222 & n13304 ) ;
  assign n13306 = ( x76 & ~n13214 ) | ( x76 & n13305 ) | ( ~n13214 & n13305 ) ;
  assign n13307 = ( x77 & ~n13206 ) | ( x77 & n13306 ) | ( ~n13206 & n13306 ) ;
  assign n13308 = ( x78 & ~n13198 ) | ( x78 & n13307 ) | ( ~n13198 & n13307 ) ;
  assign n13309 = ( x79 & ~n13190 ) | ( x79 & n13308 ) | ( ~n13190 & n13308 ) ;
  assign n13310 = ( x80 & ~n13182 ) | ( x80 & n13309 ) | ( ~n13182 & n13309 ) ;
  assign n13311 = ( x81 & ~n13174 ) | ( x81 & n13310 ) | ( ~n13174 & n13310 ) ;
  assign n13312 = ( x82 & ~n13166 ) | ( x82 & n13311 ) | ( ~n13166 & n13311 ) ;
  assign n13313 = ( x83 & ~n13158 ) | ( x83 & n13312 ) | ( ~n13158 & n13312 ) ;
  assign n13314 = ( x84 & ~n13150 ) | ( x84 & n13313 ) | ( ~n13150 & n13313 ) ;
  assign n13315 = ( x85 & ~n13142 ) | ( x85 & n13314 ) | ( ~n13142 & n13314 ) ;
  assign n13316 = ( x86 & ~n13134 ) | ( x86 & n13315 ) | ( ~n13134 & n13315 ) ;
  assign n13317 = ( x87 & ~n13126 ) | ( x87 & n13316 ) | ( ~n13126 & n13316 ) ;
  assign n13318 = ( x88 & ~n13118 ) | ( x88 & n13317 ) | ( ~n13118 & n13317 ) ;
  assign n13319 = ( x89 & ~n13110 ) | ( x89 & n13318 ) | ( ~n13110 & n13318 ) ;
  assign n13320 = ( x90 & ~n13102 ) | ( x90 & n13319 ) | ( ~n13102 & n13319 ) ;
  assign n13321 = ( x91 & ~n13094 ) | ( x91 & n13320 ) | ( ~n13094 & n13320 ) ;
  assign n13322 = ( x92 & ~n13086 ) | ( x92 & n13321 ) | ( ~n13086 & n13321 ) ;
  assign n13323 = ( x93 & ~n13078 ) | ( x93 & n13322 ) | ( ~n13078 & n13322 ) ;
  assign n13324 = ( x94 & ~n13070 ) | ( x94 & n13323 ) | ( ~n13070 & n13323 ) ;
  assign n13325 = ( x95 & ~n13062 ) | ( x95 & n13324 ) | ( ~n13062 & n13324 ) ;
  assign n13326 = ( x96 & ~n13054 ) | ( x96 & n13325 ) | ( ~n13054 & n13325 ) ;
  assign n13327 = ( x97 & ~n13046 ) | ( x97 & n13326 ) | ( ~n13046 & n13326 ) ;
  assign n13328 = ( x98 & ~n13038 ) | ( x98 & n13327 ) | ( ~n13038 & n13327 ) ;
  assign n13329 = ( x99 & ~n13030 ) | ( x99 & n13328 ) | ( ~n13030 & n13328 ) ;
  assign n13330 = ( x100 & ~n13022 ) | ( x100 & n13329 ) | ( ~n13022 & n13329 ) ;
  assign n13331 = ( x101 & ~n13014 ) | ( x101 & n13330 ) | ( ~n13014 & n13330 ) ;
  assign n13332 = ( x102 & ~n13006 ) | ( x102 & n13331 ) | ( ~n13006 & n13331 ) ;
  assign n13333 = ( x103 & ~n12998 ) | ( x103 & n13332 ) | ( ~n12998 & n13332 ) ;
  assign n13334 = ( x104 & ~n12990 ) | ( x104 & n13333 ) | ( ~n12990 & n13333 ) ;
  assign n13335 = ( x105 & ~n12982 ) | ( x105 & n13334 ) | ( ~n12982 & n13334 ) ;
  assign n13336 = ( x106 & ~n12974 ) | ( x106 & n13335 ) | ( ~n12974 & n13335 ) ;
  assign n13337 = ( x107 & ~n12966 ) | ( x107 & n13336 ) | ( ~n12966 & n13336 ) ;
  assign n13338 = ( x108 & ~n12958 ) | ( x108 & n13337 ) | ( ~n12958 & n13337 ) ;
  assign n13342 = ( x109 & ~n12950 ) | ( x109 & n13338 ) | ( ~n12950 & n13338 ) ;
  assign n13402 = ( x110 & ~n13350 ) | ( x110 & n13342 ) | ( ~n13350 & n13342 ) ;
  assign n13403 = ( x111 & ~n13401 ) | ( x111 & n13402 ) | ( ~n13401 & n13402 ) ;
  assign n13404 = ( x112 & ~n13396 ) | ( x112 & n13403 ) | ( ~n13396 & n13403 ) ;
  assign n13405 = ( x113 & ~n13388 ) | ( x113 & n13404 ) | ( ~n13388 & n13404 ) ;
  assign n13406 = ( x114 & ~n13380 ) | ( x114 & n13405 ) | ( ~n13380 & n13405 ) ;
  assign n13407 = ( x115 & ~n13372 ) | ( x115 & n13406 ) | ( ~n13372 & n13406 ) ;
  assign n13408 = ( x116 & ~n13364 ) | ( x116 & n13407 ) | ( ~n13364 & n13407 ) ;
  assign n13415 = n155 | n157 ;
  assign n13416 = n152 | n13415 ;
  assign n13410 = n160 &  n12032 ;
  assign n13411 = n12943 &  n13410 ;
  assign n13409 = n12938 | n12940 ;
  assign n13413 = ( n12932 & n12945 ) | ( n12932 & n13409 ) | ( n12945 & n13409 ) ;
  assign n13412 = n12932 | n13409 ;
  assign n13414 = ( n13411 & ~n13413 ) | ( n13411 & n13412 ) | ( ~n13413 & n13412 ) ;
  assign n13418 = x117 &  n13414 ;
  assign n13417 = x117 | n13414 ;
  assign n13419 = ( n13416 & ~n13418 ) | ( n13416 & n13417 ) | ( ~n13418 & n13417 ) ;
  assign n13420 = n13408 | n13419 ;
  assign n13421 = ~n13414 |  n425 ;
  assign n13441 = n13364 &  n13421 ;
  assign n13442 = n13420 &  n13441 ;
  assign n13428 = x116 | n13364 ;
  assign n13429 = x116 &  n13364 ;
  assign n13430 = ( n13428 & ~n13429 ) | ( n13428 & 1'b0 ) | ( ~n13429 & 1'b0 ) ;
  assign n13443 = n13407 &  n13430 ;
  assign n13422 = n13420 &  n13421 ;
  assign n13444 = ( n13407 & ~n13422 ) | ( n13407 & n13430 ) | ( ~n13422 & n13430 ) ;
  assign n13445 = ( n13442 & ~n13443 ) | ( n13442 & n13444 ) | ( ~n13443 & n13444 ) ;
  assign n13432 = ( x117 & n13408 ) | ( x117 & n13414 ) | ( n13408 & n13414 ) ;
  assign n13431 = ( x117 & ~n13408 ) | ( x117 & n13414 ) | ( ~n13408 & n13414 ) ;
  assign n13433 = ( n13408 & ~n13432 ) | ( n13408 & n13431 ) | ( ~n13432 & n13431 ) ;
  assign n13434 = ~n13422 & n13433 ;
  assign n13435 = n425 &  n13414 ;
  assign n13436 = n13420 &  n13435 ;
  assign n13437 = n13434 | n13436 ;
  assign n13449 = n13372 &  n13421 ;
  assign n13450 = n13420 &  n13449 ;
  assign n13438 = x115 | n13372 ;
  assign n13439 = x115 &  n13372 ;
  assign n13440 = ( n13438 & ~n13439 ) | ( n13438 & 1'b0 ) | ( ~n13439 & 1'b0 ) ;
  assign n13451 = n13406 &  n13440 ;
  assign n13452 = ( n13406 & ~n13422 ) | ( n13406 & n13440 ) | ( ~n13422 & n13440 ) ;
  assign n13453 = ( n13450 & ~n13451 ) | ( n13450 & n13452 ) | ( ~n13451 & n13452 ) ;
  assign n13457 = n13380 &  n13421 ;
  assign n13458 = n13420 &  n13457 ;
  assign n13446 = x114 | n13380 ;
  assign n13447 = x114 &  n13380 ;
  assign n13448 = ( n13446 & ~n13447 ) | ( n13446 & 1'b0 ) | ( ~n13447 & 1'b0 ) ;
  assign n13459 = n13405 &  n13448 ;
  assign n13460 = ( n13405 & ~n13422 ) | ( n13405 & n13448 ) | ( ~n13422 & n13448 ) ;
  assign n13461 = ( n13458 & ~n13459 ) | ( n13458 & n13460 ) | ( ~n13459 & n13460 ) ;
  assign n13465 = n13388 &  n13421 ;
  assign n13466 = n13420 &  n13465 ;
  assign n13454 = x113 | n13388 ;
  assign n13455 = x113 &  n13388 ;
  assign n13456 = ( n13454 & ~n13455 ) | ( n13454 & 1'b0 ) | ( ~n13455 & 1'b0 ) ;
  assign n13467 = n13404 &  n13456 ;
  assign n13468 = ( n13404 & ~n13422 ) | ( n13404 & n13456 ) | ( ~n13422 & n13456 ) ;
  assign n13469 = ( n13466 & ~n13467 ) | ( n13466 & n13468 ) | ( ~n13467 & n13468 ) ;
  assign n13473 = n13396 &  n13421 ;
  assign n13474 = n13420 &  n13473 ;
  assign n13462 = x112 | n13396 ;
  assign n13463 = x112 &  n13396 ;
  assign n13464 = ( n13462 & ~n13463 ) | ( n13462 & 1'b0 ) | ( ~n13463 & 1'b0 ) ;
  assign n13475 = n13403 &  n13464 ;
  assign n13476 = ( n13403 & ~n13422 ) | ( n13403 & n13464 ) | ( ~n13422 & n13464 ) ;
  assign n13477 = ( n13474 & ~n13475 ) | ( n13474 & n13476 ) | ( ~n13475 & n13476 ) ;
  assign n13478 = n13401 &  n13421 ;
  assign n13479 = n13420 &  n13478 ;
  assign n13470 = x111 | n13401 ;
  assign n13471 = x111 &  n13401 ;
  assign n13472 = ( n13470 & ~n13471 ) | ( n13470 & 1'b0 ) | ( ~n13471 & 1'b0 ) ;
  assign n13481 = ( n13402 & n13422 ) | ( n13402 & n13472 ) | ( n13422 & n13472 ) ;
  assign n13480 = n13402 | n13472 ;
  assign n13482 = ( n13479 & ~n13481 ) | ( n13479 & n13480 ) | ( ~n13481 & n13480 ) ;
  assign n13423 = n13350 &  n13421 ;
  assign n13424 = n13420 &  n13423 ;
  assign n13351 = x110 | n13350 ;
  assign n13352 = x110 &  n13350 ;
  assign n13353 = ( n13351 & ~n13352 ) | ( n13351 & 1'b0 ) | ( ~n13352 & 1'b0 ) ;
  assign n13426 = ( n13342 & n13353 ) | ( n13342 & n13422 ) | ( n13353 & n13422 ) ;
  assign n13425 = n13342 | n13353 ;
  assign n13427 = ( n13424 & ~n13426 ) | ( n13424 & n13425 ) | ( ~n13426 & n13425 ) ;
  assign n13486 = n12950 &  n13421 ;
  assign n13487 = n13420 &  n13486 ;
  assign n13339 = x109 | n12950 ;
  assign n13340 = x109 &  n12950 ;
  assign n13341 = ( n13339 & ~n13340 ) | ( n13339 & 1'b0 ) | ( ~n13340 & 1'b0 ) ;
  assign n13488 = n13338 &  n13341 ;
  assign n13489 = ( n13338 & ~n13422 ) | ( n13338 & n13341 ) | ( ~n13422 & n13341 ) ;
  assign n13490 = ( n13487 & ~n13488 ) | ( n13487 & n13489 ) | ( ~n13488 & n13489 ) ;
  assign n13494 = n12958 &  n13421 ;
  assign n13495 = n13420 &  n13494 ;
  assign n13483 = x108 | n12958 ;
  assign n13484 = x108 &  n12958 ;
  assign n13485 = ( n13483 & ~n13484 ) | ( n13483 & 1'b0 ) | ( ~n13484 & 1'b0 ) ;
  assign n13497 = ( n13337 & n13422 ) | ( n13337 & n13485 ) | ( n13422 & n13485 ) ;
  assign n13496 = n13337 | n13485 ;
  assign n13498 = ( n13495 & ~n13497 ) | ( n13495 & n13496 ) | ( ~n13497 & n13496 ) ;
  assign n13502 = n12966 &  n13421 ;
  assign n13503 = n13420 &  n13502 ;
  assign n13491 = x107 | n12966 ;
  assign n13492 = x107 &  n12966 ;
  assign n13493 = ( n13491 & ~n13492 ) | ( n13491 & 1'b0 ) | ( ~n13492 & 1'b0 ) ;
  assign n13505 = ( n13336 & n13422 ) | ( n13336 & n13493 ) | ( n13422 & n13493 ) ;
  assign n13504 = n13336 | n13493 ;
  assign n13506 = ( n13503 & ~n13505 ) | ( n13503 & n13504 ) | ( ~n13505 & n13504 ) ;
  assign n13510 = n12974 &  n13421 ;
  assign n13511 = n13420 &  n13510 ;
  assign n13499 = x106 | n12974 ;
  assign n13500 = x106 &  n12974 ;
  assign n13501 = ( n13499 & ~n13500 ) | ( n13499 & 1'b0 ) | ( ~n13500 & 1'b0 ) ;
  assign n13513 = ( n13335 & n13422 ) | ( n13335 & n13501 ) | ( n13422 & n13501 ) ;
  assign n13512 = n13335 | n13501 ;
  assign n13514 = ( n13511 & ~n13513 ) | ( n13511 & n13512 ) | ( ~n13513 & n13512 ) ;
  assign n13518 = n12982 &  n13421 ;
  assign n13519 = n13420 &  n13518 ;
  assign n13507 = x105 | n12982 ;
  assign n13508 = x105 &  n12982 ;
  assign n13509 = ( n13507 & ~n13508 ) | ( n13507 & 1'b0 ) | ( ~n13508 & 1'b0 ) ;
  assign n13521 = ( n13334 & n13422 ) | ( n13334 & n13509 ) | ( n13422 & n13509 ) ;
  assign n13520 = n13334 | n13509 ;
  assign n13522 = ( n13519 & ~n13521 ) | ( n13519 & n13520 ) | ( ~n13521 & n13520 ) ;
  assign n13526 = n12990 &  n13421 ;
  assign n13527 = n13420 &  n13526 ;
  assign n13515 = x104 | n12990 ;
  assign n13516 = x104 &  n12990 ;
  assign n13517 = ( n13515 & ~n13516 ) | ( n13515 & 1'b0 ) | ( ~n13516 & 1'b0 ) ;
  assign n13529 = ( n13333 & n13422 ) | ( n13333 & n13517 ) | ( n13422 & n13517 ) ;
  assign n13528 = n13333 | n13517 ;
  assign n13530 = ( n13527 & ~n13529 ) | ( n13527 & n13528 ) | ( ~n13529 & n13528 ) ;
  assign n13534 = n12998 &  n13421 ;
  assign n13535 = n13420 &  n13534 ;
  assign n13523 = x103 | n12998 ;
  assign n13524 = x103 &  n12998 ;
  assign n13525 = ( n13523 & ~n13524 ) | ( n13523 & 1'b0 ) | ( ~n13524 & 1'b0 ) ;
  assign n13537 = ( n13332 & n13422 ) | ( n13332 & n13525 ) | ( n13422 & n13525 ) ;
  assign n13536 = n13332 | n13525 ;
  assign n13538 = ( n13535 & ~n13537 ) | ( n13535 & n13536 ) | ( ~n13537 & n13536 ) ;
  assign n13542 = n13006 &  n13421 ;
  assign n13543 = n13420 &  n13542 ;
  assign n13531 = x102 | n13006 ;
  assign n13532 = x102 &  n13006 ;
  assign n13533 = ( n13531 & ~n13532 ) | ( n13531 & 1'b0 ) | ( ~n13532 & 1'b0 ) ;
  assign n13545 = ( n13331 & n13422 ) | ( n13331 & n13533 ) | ( n13422 & n13533 ) ;
  assign n13544 = n13331 | n13533 ;
  assign n13546 = ( n13543 & ~n13545 ) | ( n13543 & n13544 ) | ( ~n13545 & n13544 ) ;
  assign n13550 = n13014 &  n13421 ;
  assign n13551 = n13420 &  n13550 ;
  assign n13539 = x101 | n13014 ;
  assign n13540 = x101 &  n13014 ;
  assign n13541 = ( n13539 & ~n13540 ) | ( n13539 & 1'b0 ) | ( ~n13540 & 1'b0 ) ;
  assign n13553 = ( n13330 & n13422 ) | ( n13330 & n13541 ) | ( n13422 & n13541 ) ;
  assign n13552 = n13330 | n13541 ;
  assign n13554 = ( n13551 & ~n13553 ) | ( n13551 & n13552 ) | ( ~n13553 & n13552 ) ;
  assign n13558 = n13022 &  n13421 ;
  assign n13559 = n13420 &  n13558 ;
  assign n13547 = x100 | n13022 ;
  assign n13548 = x100 &  n13022 ;
  assign n13549 = ( n13547 & ~n13548 ) | ( n13547 & 1'b0 ) | ( ~n13548 & 1'b0 ) ;
  assign n13561 = ( n13329 & n13422 ) | ( n13329 & n13549 ) | ( n13422 & n13549 ) ;
  assign n13560 = n13329 | n13549 ;
  assign n13562 = ( n13559 & ~n13561 ) | ( n13559 & n13560 ) | ( ~n13561 & n13560 ) ;
  assign n13566 = n13030 &  n13421 ;
  assign n13567 = n13420 &  n13566 ;
  assign n13555 = x99 | n13030 ;
  assign n13556 = x99 &  n13030 ;
  assign n13557 = ( n13555 & ~n13556 ) | ( n13555 & 1'b0 ) | ( ~n13556 & 1'b0 ) ;
  assign n13569 = ( n13328 & n13422 ) | ( n13328 & n13557 ) | ( n13422 & n13557 ) ;
  assign n13568 = n13328 | n13557 ;
  assign n13570 = ( n13567 & ~n13569 ) | ( n13567 & n13568 ) | ( ~n13569 & n13568 ) ;
  assign n13574 = n13038 &  n13421 ;
  assign n13575 = n13420 &  n13574 ;
  assign n13563 = x98 | n13038 ;
  assign n13564 = x98 &  n13038 ;
  assign n13565 = ( n13563 & ~n13564 ) | ( n13563 & 1'b0 ) | ( ~n13564 & 1'b0 ) ;
  assign n13577 = ( n13327 & n13422 ) | ( n13327 & n13565 ) | ( n13422 & n13565 ) ;
  assign n13576 = n13327 | n13565 ;
  assign n13578 = ( n13575 & ~n13577 ) | ( n13575 & n13576 ) | ( ~n13577 & n13576 ) ;
  assign n13582 = n13046 &  n13421 ;
  assign n13583 = n13420 &  n13582 ;
  assign n13571 = x97 | n13046 ;
  assign n13572 = x97 &  n13046 ;
  assign n13573 = ( n13571 & ~n13572 ) | ( n13571 & 1'b0 ) | ( ~n13572 & 1'b0 ) ;
  assign n13585 = ( n13326 & n13422 ) | ( n13326 & n13573 ) | ( n13422 & n13573 ) ;
  assign n13584 = n13326 | n13573 ;
  assign n13586 = ( n13583 & ~n13585 ) | ( n13583 & n13584 ) | ( ~n13585 & n13584 ) ;
  assign n13590 = n13054 &  n13421 ;
  assign n13591 = n13420 &  n13590 ;
  assign n13579 = x96 | n13054 ;
  assign n13580 = x96 &  n13054 ;
  assign n13581 = ( n13579 & ~n13580 ) | ( n13579 & 1'b0 ) | ( ~n13580 & 1'b0 ) ;
  assign n13593 = ( n13325 & n13422 ) | ( n13325 & n13581 ) | ( n13422 & n13581 ) ;
  assign n13592 = n13325 | n13581 ;
  assign n13594 = ( n13591 & ~n13593 ) | ( n13591 & n13592 ) | ( ~n13593 & n13592 ) ;
  assign n13598 = n13062 &  n13421 ;
  assign n13599 = n13420 &  n13598 ;
  assign n13587 = x95 | n13062 ;
  assign n13588 = x95 &  n13062 ;
  assign n13589 = ( n13587 & ~n13588 ) | ( n13587 & 1'b0 ) | ( ~n13588 & 1'b0 ) ;
  assign n13601 = ( n13324 & n13422 ) | ( n13324 & n13589 ) | ( n13422 & n13589 ) ;
  assign n13600 = n13324 | n13589 ;
  assign n13602 = ( n13599 & ~n13601 ) | ( n13599 & n13600 ) | ( ~n13601 & n13600 ) ;
  assign n13606 = n13070 &  n13421 ;
  assign n13607 = n13420 &  n13606 ;
  assign n13595 = x94 | n13070 ;
  assign n13596 = x94 &  n13070 ;
  assign n13597 = ( n13595 & ~n13596 ) | ( n13595 & 1'b0 ) | ( ~n13596 & 1'b0 ) ;
  assign n13609 = ( n13323 & n13422 ) | ( n13323 & n13597 ) | ( n13422 & n13597 ) ;
  assign n13608 = n13323 | n13597 ;
  assign n13610 = ( n13607 & ~n13609 ) | ( n13607 & n13608 ) | ( ~n13609 & n13608 ) ;
  assign n13614 = n13078 &  n13421 ;
  assign n13615 = n13420 &  n13614 ;
  assign n13603 = x93 | n13078 ;
  assign n13604 = x93 &  n13078 ;
  assign n13605 = ( n13603 & ~n13604 ) | ( n13603 & 1'b0 ) | ( ~n13604 & 1'b0 ) ;
  assign n13617 = ( n13322 & n13422 ) | ( n13322 & n13605 ) | ( n13422 & n13605 ) ;
  assign n13616 = n13322 | n13605 ;
  assign n13618 = ( n13615 & ~n13617 ) | ( n13615 & n13616 ) | ( ~n13617 & n13616 ) ;
  assign n13622 = n13086 &  n13421 ;
  assign n13623 = n13420 &  n13622 ;
  assign n13611 = x92 | n13086 ;
  assign n13612 = x92 &  n13086 ;
  assign n13613 = ( n13611 & ~n13612 ) | ( n13611 & 1'b0 ) | ( ~n13612 & 1'b0 ) ;
  assign n13625 = ( n13321 & n13422 ) | ( n13321 & n13613 ) | ( n13422 & n13613 ) ;
  assign n13624 = n13321 | n13613 ;
  assign n13626 = ( n13623 & ~n13625 ) | ( n13623 & n13624 ) | ( ~n13625 & n13624 ) ;
  assign n13630 = n13094 &  n13421 ;
  assign n13631 = n13420 &  n13630 ;
  assign n13619 = x91 | n13094 ;
  assign n13620 = x91 &  n13094 ;
  assign n13621 = ( n13619 & ~n13620 ) | ( n13619 & 1'b0 ) | ( ~n13620 & 1'b0 ) ;
  assign n13633 = ( n13320 & n13422 ) | ( n13320 & n13621 ) | ( n13422 & n13621 ) ;
  assign n13632 = n13320 | n13621 ;
  assign n13634 = ( n13631 & ~n13633 ) | ( n13631 & n13632 ) | ( ~n13633 & n13632 ) ;
  assign n13638 = n13102 &  n13421 ;
  assign n13639 = n13420 &  n13638 ;
  assign n13627 = x90 | n13102 ;
  assign n13628 = x90 &  n13102 ;
  assign n13629 = ( n13627 & ~n13628 ) | ( n13627 & 1'b0 ) | ( ~n13628 & 1'b0 ) ;
  assign n13641 = ( n13319 & n13422 ) | ( n13319 & n13629 ) | ( n13422 & n13629 ) ;
  assign n13640 = n13319 | n13629 ;
  assign n13642 = ( n13639 & ~n13641 ) | ( n13639 & n13640 ) | ( ~n13641 & n13640 ) ;
  assign n13646 = n13110 &  n13421 ;
  assign n13647 = n13420 &  n13646 ;
  assign n13635 = x89 | n13110 ;
  assign n13636 = x89 &  n13110 ;
  assign n13637 = ( n13635 & ~n13636 ) | ( n13635 & 1'b0 ) | ( ~n13636 & 1'b0 ) ;
  assign n13649 = ( n13318 & n13422 ) | ( n13318 & n13637 ) | ( n13422 & n13637 ) ;
  assign n13648 = n13318 | n13637 ;
  assign n13650 = ( n13647 & ~n13649 ) | ( n13647 & n13648 ) | ( ~n13649 & n13648 ) ;
  assign n13654 = n13118 &  n13421 ;
  assign n13655 = n13420 &  n13654 ;
  assign n13643 = x88 | n13118 ;
  assign n13644 = x88 &  n13118 ;
  assign n13645 = ( n13643 & ~n13644 ) | ( n13643 & 1'b0 ) | ( ~n13644 & 1'b0 ) ;
  assign n13657 = ( n13317 & n13422 ) | ( n13317 & n13645 ) | ( n13422 & n13645 ) ;
  assign n13656 = n13317 | n13645 ;
  assign n13658 = ( n13655 & ~n13657 ) | ( n13655 & n13656 ) | ( ~n13657 & n13656 ) ;
  assign n13662 = n13126 &  n13421 ;
  assign n13663 = n13420 &  n13662 ;
  assign n13651 = x87 | n13126 ;
  assign n13652 = x87 &  n13126 ;
  assign n13653 = ( n13651 & ~n13652 ) | ( n13651 & 1'b0 ) | ( ~n13652 & 1'b0 ) ;
  assign n13665 = ( n13316 & n13422 ) | ( n13316 & n13653 ) | ( n13422 & n13653 ) ;
  assign n13664 = n13316 | n13653 ;
  assign n13666 = ( n13663 & ~n13665 ) | ( n13663 & n13664 ) | ( ~n13665 & n13664 ) ;
  assign n13670 = n13134 &  n13421 ;
  assign n13671 = n13420 &  n13670 ;
  assign n13659 = x86 | n13134 ;
  assign n13660 = x86 &  n13134 ;
  assign n13661 = ( n13659 & ~n13660 ) | ( n13659 & 1'b0 ) | ( ~n13660 & 1'b0 ) ;
  assign n13673 = ( n13315 & n13422 ) | ( n13315 & n13661 ) | ( n13422 & n13661 ) ;
  assign n13672 = n13315 | n13661 ;
  assign n13674 = ( n13671 & ~n13673 ) | ( n13671 & n13672 ) | ( ~n13673 & n13672 ) ;
  assign n13678 = n13142 &  n13421 ;
  assign n13679 = n13420 &  n13678 ;
  assign n13667 = x85 | n13142 ;
  assign n13668 = x85 &  n13142 ;
  assign n13669 = ( n13667 & ~n13668 ) | ( n13667 & 1'b0 ) | ( ~n13668 & 1'b0 ) ;
  assign n13681 = ( n13314 & n13422 ) | ( n13314 & n13669 ) | ( n13422 & n13669 ) ;
  assign n13680 = n13314 | n13669 ;
  assign n13682 = ( n13679 & ~n13681 ) | ( n13679 & n13680 ) | ( ~n13681 & n13680 ) ;
  assign n13686 = n13150 &  n13421 ;
  assign n13687 = n13420 &  n13686 ;
  assign n13675 = x84 | n13150 ;
  assign n13676 = x84 &  n13150 ;
  assign n13677 = ( n13675 & ~n13676 ) | ( n13675 & 1'b0 ) | ( ~n13676 & 1'b0 ) ;
  assign n13689 = ( n13313 & n13422 ) | ( n13313 & n13677 ) | ( n13422 & n13677 ) ;
  assign n13688 = n13313 | n13677 ;
  assign n13690 = ( n13687 & ~n13689 ) | ( n13687 & n13688 ) | ( ~n13689 & n13688 ) ;
  assign n13694 = n13158 &  n13421 ;
  assign n13695 = n13420 &  n13694 ;
  assign n13683 = x83 | n13158 ;
  assign n13684 = x83 &  n13158 ;
  assign n13685 = ( n13683 & ~n13684 ) | ( n13683 & 1'b0 ) | ( ~n13684 & 1'b0 ) ;
  assign n13697 = ( n13312 & n13422 ) | ( n13312 & n13685 ) | ( n13422 & n13685 ) ;
  assign n13696 = n13312 | n13685 ;
  assign n13698 = ( n13695 & ~n13697 ) | ( n13695 & n13696 ) | ( ~n13697 & n13696 ) ;
  assign n13702 = n13166 &  n13421 ;
  assign n13703 = n13420 &  n13702 ;
  assign n13691 = x82 | n13166 ;
  assign n13692 = x82 &  n13166 ;
  assign n13693 = ( n13691 & ~n13692 ) | ( n13691 & 1'b0 ) | ( ~n13692 & 1'b0 ) ;
  assign n13705 = ( n13311 & n13422 ) | ( n13311 & n13693 ) | ( n13422 & n13693 ) ;
  assign n13704 = n13311 | n13693 ;
  assign n13706 = ( n13703 & ~n13705 ) | ( n13703 & n13704 ) | ( ~n13705 & n13704 ) ;
  assign n13710 = n13174 &  n13421 ;
  assign n13711 = n13420 &  n13710 ;
  assign n13699 = x81 | n13174 ;
  assign n13700 = x81 &  n13174 ;
  assign n13701 = ( n13699 & ~n13700 ) | ( n13699 & 1'b0 ) | ( ~n13700 & 1'b0 ) ;
  assign n13713 = ( n13310 & n13422 ) | ( n13310 & n13701 ) | ( n13422 & n13701 ) ;
  assign n13712 = n13310 | n13701 ;
  assign n13714 = ( n13711 & ~n13713 ) | ( n13711 & n13712 ) | ( ~n13713 & n13712 ) ;
  assign n13718 = n13182 &  n13421 ;
  assign n13719 = n13420 &  n13718 ;
  assign n13707 = x80 | n13182 ;
  assign n13708 = x80 &  n13182 ;
  assign n13709 = ( n13707 & ~n13708 ) | ( n13707 & 1'b0 ) | ( ~n13708 & 1'b0 ) ;
  assign n13721 = ( n13309 & n13422 ) | ( n13309 & n13709 ) | ( n13422 & n13709 ) ;
  assign n13720 = n13309 | n13709 ;
  assign n13722 = ( n13719 & ~n13721 ) | ( n13719 & n13720 ) | ( ~n13721 & n13720 ) ;
  assign n13726 = n13190 &  n13421 ;
  assign n13727 = n13420 &  n13726 ;
  assign n13715 = x79 | n13190 ;
  assign n13716 = x79 &  n13190 ;
  assign n13717 = ( n13715 & ~n13716 ) | ( n13715 & 1'b0 ) | ( ~n13716 & 1'b0 ) ;
  assign n13729 = ( n13308 & n13422 ) | ( n13308 & n13717 ) | ( n13422 & n13717 ) ;
  assign n13728 = n13308 | n13717 ;
  assign n13730 = ( n13727 & ~n13729 ) | ( n13727 & n13728 ) | ( ~n13729 & n13728 ) ;
  assign n13734 = n13198 &  n13421 ;
  assign n13735 = n13420 &  n13734 ;
  assign n13723 = x78 | n13198 ;
  assign n13724 = x78 &  n13198 ;
  assign n13725 = ( n13723 & ~n13724 ) | ( n13723 & 1'b0 ) | ( ~n13724 & 1'b0 ) ;
  assign n13737 = ( n13307 & n13422 ) | ( n13307 & n13725 ) | ( n13422 & n13725 ) ;
  assign n13736 = n13307 | n13725 ;
  assign n13738 = ( n13735 & ~n13737 ) | ( n13735 & n13736 ) | ( ~n13737 & n13736 ) ;
  assign n13742 = n13206 &  n13421 ;
  assign n13743 = n13420 &  n13742 ;
  assign n13731 = x77 | n13206 ;
  assign n13732 = x77 &  n13206 ;
  assign n13733 = ( n13731 & ~n13732 ) | ( n13731 & 1'b0 ) | ( ~n13732 & 1'b0 ) ;
  assign n13745 = ( n13306 & n13422 ) | ( n13306 & n13733 ) | ( n13422 & n13733 ) ;
  assign n13744 = n13306 | n13733 ;
  assign n13746 = ( n13743 & ~n13745 ) | ( n13743 & n13744 ) | ( ~n13745 & n13744 ) ;
  assign n13750 = n13214 &  n13421 ;
  assign n13751 = n13420 &  n13750 ;
  assign n13739 = x76 | n13214 ;
  assign n13740 = x76 &  n13214 ;
  assign n13741 = ( n13739 & ~n13740 ) | ( n13739 & 1'b0 ) | ( ~n13740 & 1'b0 ) ;
  assign n13753 = ( n13305 & n13422 ) | ( n13305 & n13741 ) | ( n13422 & n13741 ) ;
  assign n13752 = n13305 | n13741 ;
  assign n13754 = ( n13751 & ~n13753 ) | ( n13751 & n13752 ) | ( ~n13753 & n13752 ) ;
  assign n13758 = n13222 &  n13421 ;
  assign n13759 = n13420 &  n13758 ;
  assign n13747 = x75 | n13222 ;
  assign n13748 = x75 &  n13222 ;
  assign n13749 = ( n13747 & ~n13748 ) | ( n13747 & 1'b0 ) | ( ~n13748 & 1'b0 ) ;
  assign n13761 = ( n13304 & n13422 ) | ( n13304 & n13749 ) | ( n13422 & n13749 ) ;
  assign n13760 = n13304 | n13749 ;
  assign n13762 = ( n13759 & ~n13761 ) | ( n13759 & n13760 ) | ( ~n13761 & n13760 ) ;
  assign n13766 = n13230 &  n13421 ;
  assign n13767 = n13420 &  n13766 ;
  assign n13755 = x74 | n13230 ;
  assign n13756 = x74 &  n13230 ;
  assign n13757 = ( n13755 & ~n13756 ) | ( n13755 & 1'b0 ) | ( ~n13756 & 1'b0 ) ;
  assign n13769 = ( n13303 & n13422 ) | ( n13303 & n13757 ) | ( n13422 & n13757 ) ;
  assign n13768 = n13303 | n13757 ;
  assign n13770 = ( n13767 & ~n13769 ) | ( n13767 & n13768 ) | ( ~n13769 & n13768 ) ;
  assign n13774 = n13238 &  n13421 ;
  assign n13775 = n13420 &  n13774 ;
  assign n13763 = x73 | n13238 ;
  assign n13764 = x73 &  n13238 ;
  assign n13765 = ( n13763 & ~n13764 ) | ( n13763 & 1'b0 ) | ( ~n13764 & 1'b0 ) ;
  assign n13777 = ( n13302 & n13422 ) | ( n13302 & n13765 ) | ( n13422 & n13765 ) ;
  assign n13776 = n13302 | n13765 ;
  assign n13778 = ( n13775 & ~n13777 ) | ( n13775 & n13776 ) | ( ~n13777 & n13776 ) ;
  assign n13782 = n13246 &  n13421 ;
  assign n13783 = n13420 &  n13782 ;
  assign n13771 = x72 | n13246 ;
  assign n13772 = x72 &  n13246 ;
  assign n13773 = ( n13771 & ~n13772 ) | ( n13771 & 1'b0 ) | ( ~n13772 & 1'b0 ) ;
  assign n13785 = ( n13301 & n13422 ) | ( n13301 & n13773 ) | ( n13422 & n13773 ) ;
  assign n13784 = n13301 | n13773 ;
  assign n13786 = ( n13783 & ~n13785 ) | ( n13783 & n13784 ) | ( ~n13785 & n13784 ) ;
  assign n13790 = n13254 &  n13421 ;
  assign n13791 = n13420 &  n13790 ;
  assign n13779 = x71 | n13254 ;
  assign n13780 = x71 &  n13254 ;
  assign n13781 = ( n13779 & ~n13780 ) | ( n13779 & 1'b0 ) | ( ~n13780 & 1'b0 ) ;
  assign n13793 = ( n13300 & n13422 ) | ( n13300 & n13781 ) | ( n13422 & n13781 ) ;
  assign n13792 = n13300 | n13781 ;
  assign n13794 = ( n13791 & ~n13793 ) | ( n13791 & n13792 ) | ( ~n13793 & n13792 ) ;
  assign n13798 = n13262 &  n13421 ;
  assign n13799 = n13420 &  n13798 ;
  assign n13787 = x70 | n13262 ;
  assign n13788 = x70 &  n13262 ;
  assign n13789 = ( n13787 & ~n13788 ) | ( n13787 & 1'b0 ) | ( ~n13788 & 1'b0 ) ;
  assign n13801 = ( n13299 & n13422 ) | ( n13299 & n13789 ) | ( n13422 & n13789 ) ;
  assign n13800 = n13299 | n13789 ;
  assign n13802 = ( n13799 & ~n13801 ) | ( n13799 & n13800 ) | ( ~n13801 & n13800 ) ;
  assign n13806 = n13270 &  n13421 ;
  assign n13807 = n13420 &  n13806 ;
  assign n13795 = x69 | n13270 ;
  assign n13796 = x69 &  n13270 ;
  assign n13797 = ( n13795 & ~n13796 ) | ( n13795 & 1'b0 ) | ( ~n13796 & 1'b0 ) ;
  assign n13809 = ( n13298 & n13422 ) | ( n13298 & n13797 ) | ( n13422 & n13797 ) ;
  assign n13808 = n13298 | n13797 ;
  assign n13810 = ( n13807 & ~n13809 ) | ( n13807 & n13808 ) | ( ~n13809 & n13808 ) ;
  assign n13814 = n13278 &  n13421 ;
  assign n13815 = n13420 &  n13814 ;
  assign n13803 = x68 | n13278 ;
  assign n13804 = x68 &  n13278 ;
  assign n13805 = ( n13803 & ~n13804 ) | ( n13803 & 1'b0 ) | ( ~n13804 & 1'b0 ) ;
  assign n13817 = ( n13297 & n13422 ) | ( n13297 & n13805 ) | ( n13422 & n13805 ) ;
  assign n13816 = n13297 | n13805 ;
  assign n13818 = ( n13815 & ~n13817 ) | ( n13815 & n13816 ) | ( ~n13817 & n13816 ) ;
  assign n13822 = n13283 &  n13421 ;
  assign n13823 = n13420 &  n13822 ;
  assign n13811 = x67 | n13283 ;
  assign n13812 = x67 &  n13283 ;
  assign n13813 = ( n13811 & ~n13812 ) | ( n13811 & 1'b0 ) | ( ~n13812 & 1'b0 ) ;
  assign n13825 = ( n13296 & n13422 ) | ( n13296 & n13813 ) | ( n13422 & n13813 ) ;
  assign n13824 = n13296 | n13813 ;
  assign n13826 = ( n13823 & ~n13825 ) | ( n13823 & n13824 ) | ( ~n13825 & n13824 ) ;
  assign n13827 = n13289 &  n13421 ;
  assign n13828 = n13420 &  n13827 ;
  assign n13819 = x66 | n13289 ;
  assign n13820 = x66 &  n13289 ;
  assign n13821 = ( n13819 & ~n13820 ) | ( n13819 & 1'b0 ) | ( ~n13820 & 1'b0 ) ;
  assign n13829 = n13295 &  n13821 ;
  assign n13830 = ( n13295 & ~n13422 ) | ( n13295 & n13821 ) | ( ~n13422 & n13821 ) ;
  assign n13831 = ( n13828 & ~n13829 ) | ( n13828 & n13830 ) | ( ~n13829 & n13830 ) ;
  assign n13832 = ( n13293 & ~x65 ) | ( n13293 & n13294 ) | ( ~x65 & n13294 ) ;
  assign n13833 = ( n13295 & ~n13294 ) | ( n13295 & n13832 ) | ( ~n13294 & n13832 ) ;
  assign n13834 = ~n13422 & n13833 ;
  assign n13835 = n13293 &  n13421 ;
  assign n13836 = n13420 &  n13835 ;
  assign n13837 = n13834 | n13836 ;
  assign n13838 = ( x64 & ~n13422 ) | ( x64 & 1'b0 ) | ( ~n13422 & 1'b0 ) ;
  assign n13839 = ( x10 & ~n13838 ) | ( x10 & 1'b0 ) | ( ~n13838 & 1'b0 ) ;
  assign n13840 = ( n13294 & ~n13422 ) | ( n13294 & 1'b0 ) | ( ~n13422 & 1'b0 ) ;
  assign n13841 = n13839 | n13840 ;
  assign n13842 = ~x9 & x64 ;
  assign n13843 = ( x65 & ~n13841 ) | ( x65 & n13842 ) | ( ~n13841 & n13842 ) ;
  assign n13844 = ( x66 & ~n13837 ) | ( x66 & n13843 ) | ( ~n13837 & n13843 ) ;
  assign n13845 = ( x67 & ~n13831 ) | ( x67 & n13844 ) | ( ~n13831 & n13844 ) ;
  assign n13846 = ( x68 & ~n13826 ) | ( x68 & n13845 ) | ( ~n13826 & n13845 ) ;
  assign n13847 = ( x69 & ~n13818 ) | ( x69 & n13846 ) | ( ~n13818 & n13846 ) ;
  assign n13848 = ( x70 & ~n13810 ) | ( x70 & n13847 ) | ( ~n13810 & n13847 ) ;
  assign n13849 = ( x71 & ~n13802 ) | ( x71 & n13848 ) | ( ~n13802 & n13848 ) ;
  assign n13850 = ( x72 & ~n13794 ) | ( x72 & n13849 ) | ( ~n13794 & n13849 ) ;
  assign n13851 = ( x73 & ~n13786 ) | ( x73 & n13850 ) | ( ~n13786 & n13850 ) ;
  assign n13852 = ( x74 & ~n13778 ) | ( x74 & n13851 ) | ( ~n13778 & n13851 ) ;
  assign n13853 = ( x75 & ~n13770 ) | ( x75 & n13852 ) | ( ~n13770 & n13852 ) ;
  assign n13854 = ( x76 & ~n13762 ) | ( x76 & n13853 ) | ( ~n13762 & n13853 ) ;
  assign n13855 = ( x77 & ~n13754 ) | ( x77 & n13854 ) | ( ~n13754 & n13854 ) ;
  assign n13856 = ( x78 & ~n13746 ) | ( x78 & n13855 ) | ( ~n13746 & n13855 ) ;
  assign n13857 = ( x79 & ~n13738 ) | ( x79 & n13856 ) | ( ~n13738 & n13856 ) ;
  assign n13858 = ( x80 & ~n13730 ) | ( x80 & n13857 ) | ( ~n13730 & n13857 ) ;
  assign n13859 = ( x81 & ~n13722 ) | ( x81 & n13858 ) | ( ~n13722 & n13858 ) ;
  assign n13860 = ( x82 & ~n13714 ) | ( x82 & n13859 ) | ( ~n13714 & n13859 ) ;
  assign n13861 = ( x83 & ~n13706 ) | ( x83 & n13860 ) | ( ~n13706 & n13860 ) ;
  assign n13862 = ( x84 & ~n13698 ) | ( x84 & n13861 ) | ( ~n13698 & n13861 ) ;
  assign n13863 = ( x85 & ~n13690 ) | ( x85 & n13862 ) | ( ~n13690 & n13862 ) ;
  assign n13864 = ( x86 & ~n13682 ) | ( x86 & n13863 ) | ( ~n13682 & n13863 ) ;
  assign n13865 = ( x87 & ~n13674 ) | ( x87 & n13864 ) | ( ~n13674 & n13864 ) ;
  assign n13866 = ( x88 & ~n13666 ) | ( x88 & n13865 ) | ( ~n13666 & n13865 ) ;
  assign n13867 = ( x89 & ~n13658 ) | ( x89 & n13866 ) | ( ~n13658 & n13866 ) ;
  assign n13868 = ( x90 & ~n13650 ) | ( x90 & n13867 ) | ( ~n13650 & n13867 ) ;
  assign n13869 = ( x91 & ~n13642 ) | ( x91 & n13868 ) | ( ~n13642 & n13868 ) ;
  assign n13870 = ( x92 & ~n13634 ) | ( x92 & n13869 ) | ( ~n13634 & n13869 ) ;
  assign n13871 = ( x93 & ~n13626 ) | ( x93 & n13870 ) | ( ~n13626 & n13870 ) ;
  assign n13872 = ( x94 & ~n13618 ) | ( x94 & n13871 ) | ( ~n13618 & n13871 ) ;
  assign n13873 = ( x95 & ~n13610 ) | ( x95 & n13872 ) | ( ~n13610 & n13872 ) ;
  assign n13874 = ( x96 & ~n13602 ) | ( x96 & n13873 ) | ( ~n13602 & n13873 ) ;
  assign n13875 = ( x97 & ~n13594 ) | ( x97 & n13874 ) | ( ~n13594 & n13874 ) ;
  assign n13876 = ( x98 & ~n13586 ) | ( x98 & n13875 ) | ( ~n13586 & n13875 ) ;
  assign n13877 = ( x99 & ~n13578 ) | ( x99 & n13876 ) | ( ~n13578 & n13876 ) ;
  assign n13878 = ( x100 & ~n13570 ) | ( x100 & n13877 ) | ( ~n13570 & n13877 ) ;
  assign n13879 = ( x101 & ~n13562 ) | ( x101 & n13878 ) | ( ~n13562 & n13878 ) ;
  assign n13880 = ( x102 & ~n13554 ) | ( x102 & n13879 ) | ( ~n13554 & n13879 ) ;
  assign n13881 = ( x103 & ~n13546 ) | ( x103 & n13880 ) | ( ~n13546 & n13880 ) ;
  assign n13882 = ( x104 & ~n13538 ) | ( x104 & n13881 ) | ( ~n13538 & n13881 ) ;
  assign n13883 = ( x105 & ~n13530 ) | ( x105 & n13882 ) | ( ~n13530 & n13882 ) ;
  assign n13884 = ( x106 & ~n13522 ) | ( x106 & n13883 ) | ( ~n13522 & n13883 ) ;
  assign n13885 = ( x107 & ~n13514 ) | ( x107 & n13884 ) | ( ~n13514 & n13884 ) ;
  assign n13886 = ( x108 & ~n13506 ) | ( x108 & n13885 ) | ( ~n13506 & n13885 ) ;
  assign n13887 = ( x109 & ~n13498 ) | ( x109 & n13886 ) | ( ~n13498 & n13886 ) ;
  assign n13888 = ( x110 & ~n13490 ) | ( x110 & n13887 ) | ( ~n13490 & n13887 ) ;
  assign n13889 = ( x111 & ~n13427 ) | ( x111 & n13888 ) | ( ~n13427 & n13888 ) ;
  assign n13890 = ( x112 & ~n13482 ) | ( x112 & n13889 ) | ( ~n13482 & n13889 ) ;
  assign n13891 = ( x113 & ~n13477 ) | ( x113 & n13890 ) | ( ~n13477 & n13890 ) ;
  assign n13892 = ( x114 & ~n13469 ) | ( x114 & n13891 ) | ( ~n13469 & n13891 ) ;
  assign n13893 = ( x115 & ~n13461 ) | ( x115 & n13892 ) | ( ~n13461 & n13892 ) ;
  assign n13894 = ( x116 & ~n13453 ) | ( x116 & n13893 ) | ( ~n13453 & n13893 ) ;
  assign n13895 = ( x117 & ~n13445 ) | ( x117 & n13894 ) | ( ~n13445 & n13894 ) ;
  assign n13896 = ( x118 & ~n13437 ) | ( x118 & n13895 ) | ( ~n13437 & n13895 ) ;
  assign n13897 = n228 | n238 ;
  assign n13898 = n235 | n13897 ;
  assign n13899 = n13896 | n13898 ;
  assign n14351 = n13445 &  n13899 ;
  assign n14355 = x117 | n13445 ;
  assign n14356 = x117 &  n13445 ;
  assign n14357 = ( n14355 & ~n14356 ) | ( n14355 & 1'b0 ) | ( ~n14356 & 1'b0 ) ;
  assign n14358 = ( n13894 & n13896 ) | ( n13894 & n14357 ) | ( n13896 & n14357 ) ;
  assign n14359 = ( n13894 & ~n13898 ) | ( n13894 & n14357 ) | ( ~n13898 & n14357 ) ;
  assign n14360 = ~n14358 & n14359 ;
  assign n14361 = n14351 | n14360 ;
  assign n14362 = n13453 &  n13899 ;
  assign n14352 = x116 | n13453 ;
  assign n14353 = x116 &  n13453 ;
  assign n14354 = ( n14352 & ~n14353 ) | ( n14352 & 1'b0 ) | ( ~n14353 & 1'b0 ) ;
  assign n14366 = ( n13893 & n13896 ) | ( n13893 & n14354 ) | ( n13896 & n14354 ) ;
  assign n14367 = ( n13893 & ~n13898 ) | ( n13893 & n14354 ) | ( ~n13898 & n14354 ) ;
  assign n14368 = ~n14366 & n14367 ;
  assign n14369 = n14362 | n14368 ;
  assign n14370 = n13461 &  n13899 ;
  assign n14363 = x115 | n13461 ;
  assign n14364 = x115 &  n13461 ;
  assign n14365 = ( n14363 & ~n14364 ) | ( n14363 & 1'b0 ) | ( ~n14364 & 1'b0 ) ;
  assign n14374 = ( n13892 & n13896 ) | ( n13892 & n14365 ) | ( n13896 & n14365 ) ;
  assign n14375 = ( n13892 & ~n13898 ) | ( n13892 & n14365 ) | ( ~n13898 & n14365 ) ;
  assign n14376 = ~n14374 & n14375 ;
  assign n14377 = n14370 | n14376 ;
  assign n14378 = n13469 &  n13899 ;
  assign n14371 = x114 | n13469 ;
  assign n14372 = x114 &  n13469 ;
  assign n14373 = ( n14371 & ~n14372 ) | ( n14371 & 1'b0 ) | ( ~n14372 & 1'b0 ) ;
  assign n14382 = ( n13891 & n13896 ) | ( n13891 & n14373 ) | ( n13896 & n14373 ) ;
  assign n14383 = ( n13891 & ~n13898 ) | ( n13891 & n14373 ) | ( ~n13898 & n14373 ) ;
  assign n14384 = ~n14382 & n14383 ;
  assign n14385 = n14378 | n14384 ;
  assign n14386 = n13477 &  n13899 ;
  assign n14379 = x113 | n13477 ;
  assign n14380 = x113 &  n13477 ;
  assign n14381 = ( n14379 & ~n14380 ) | ( n14379 & 1'b0 ) | ( ~n14380 & 1'b0 ) ;
  assign n14387 = ( n13890 & n13896 ) | ( n13890 & n14381 ) | ( n13896 & n14381 ) ;
  assign n14388 = ( n13890 & ~n13898 ) | ( n13890 & n14381 ) | ( ~n13898 & n14381 ) ;
  assign n14389 = ~n14387 & n14388 ;
  assign n14390 = n14386 | n14389 ;
  assign n14340 = n13482 &  n13899 ;
  assign n14341 = x112 | n13482 ;
  assign n14342 = x112 &  n13482 ;
  assign n14343 = ( n14341 & ~n14342 ) | ( n14341 & 1'b0 ) | ( ~n14342 & 1'b0 ) ;
  assign n14344 = ( n13889 & n13896 ) | ( n13889 & n14343 ) | ( n13896 & n14343 ) ;
  assign n14345 = ( n13889 & ~n13898 ) | ( n13889 & n14343 ) | ( ~n13898 & n14343 ) ;
  assign n14346 = ~n14344 & n14345 ;
  assign n14347 = n14340 | n14346 ;
  assign n13900 = n13427 &  n13899 ;
  assign n13904 = x111 | n13427 ;
  assign n13905 = x111 &  n13427 ;
  assign n13906 = ( n13904 & ~n13905 ) | ( n13904 & 1'b0 ) | ( ~n13905 & 1'b0 ) ;
  assign n13907 = ( n13888 & n13896 ) | ( n13888 & n13906 ) | ( n13896 & n13906 ) ;
  assign n13908 = ( n13888 & ~n13898 ) | ( n13888 & n13906 ) | ( ~n13898 & n13906 ) ;
  assign n13909 = ~n13907 & n13908 ;
  assign n13910 = n13900 | n13909 ;
  assign n13911 = n13490 &  n13899 ;
  assign n13901 = x110 | n13490 ;
  assign n13902 = x110 &  n13490 ;
  assign n13903 = ( n13901 & ~n13902 ) | ( n13901 & 1'b0 ) | ( ~n13902 & 1'b0 ) ;
  assign n13915 = ( n13887 & n13896 ) | ( n13887 & n13903 ) | ( n13896 & n13903 ) ;
  assign n13916 = ( n13887 & ~n13898 ) | ( n13887 & n13903 ) | ( ~n13898 & n13903 ) ;
  assign n13917 = ~n13915 & n13916 ;
  assign n13918 = n13911 | n13917 ;
  assign n13919 = n13498 &  n13899 ;
  assign n13912 = x109 | n13498 ;
  assign n13913 = x109 &  n13498 ;
  assign n13914 = ( n13912 & ~n13913 ) | ( n13912 & 1'b0 ) | ( ~n13913 & 1'b0 ) ;
  assign n13923 = ( n13886 & n13896 ) | ( n13886 & n13914 ) | ( n13896 & n13914 ) ;
  assign n13924 = ( n13886 & ~n13898 ) | ( n13886 & n13914 ) | ( ~n13898 & n13914 ) ;
  assign n13925 = ~n13923 & n13924 ;
  assign n13926 = n13919 | n13925 ;
  assign n13927 = n13506 &  n13899 ;
  assign n13920 = x108 | n13506 ;
  assign n13921 = x108 &  n13506 ;
  assign n13922 = ( n13920 & ~n13921 ) | ( n13920 & 1'b0 ) | ( ~n13921 & 1'b0 ) ;
  assign n13931 = ( n13885 & n13896 ) | ( n13885 & n13922 ) | ( n13896 & n13922 ) ;
  assign n13932 = ( n13885 & ~n13898 ) | ( n13885 & n13922 ) | ( ~n13898 & n13922 ) ;
  assign n13933 = ~n13931 & n13932 ;
  assign n13934 = n13927 | n13933 ;
  assign n13935 = n13514 &  n13899 ;
  assign n13928 = x107 | n13514 ;
  assign n13929 = x107 &  n13514 ;
  assign n13930 = ( n13928 & ~n13929 ) | ( n13928 & 1'b0 ) | ( ~n13929 & 1'b0 ) ;
  assign n13939 = ( n13884 & n13896 ) | ( n13884 & n13930 ) | ( n13896 & n13930 ) ;
  assign n13940 = ( n13884 & ~n13898 ) | ( n13884 & n13930 ) | ( ~n13898 & n13930 ) ;
  assign n13941 = ~n13939 & n13940 ;
  assign n13942 = n13935 | n13941 ;
  assign n13943 = n13522 &  n13899 ;
  assign n13936 = x106 | n13522 ;
  assign n13937 = x106 &  n13522 ;
  assign n13938 = ( n13936 & ~n13937 ) | ( n13936 & 1'b0 ) | ( ~n13937 & 1'b0 ) ;
  assign n13947 = ( n13883 & n13896 ) | ( n13883 & n13938 ) | ( n13896 & n13938 ) ;
  assign n13948 = ( n13883 & ~n13898 ) | ( n13883 & n13938 ) | ( ~n13898 & n13938 ) ;
  assign n13949 = ~n13947 & n13948 ;
  assign n13950 = n13943 | n13949 ;
  assign n13951 = n13530 &  n13899 ;
  assign n13944 = x105 | n13530 ;
  assign n13945 = x105 &  n13530 ;
  assign n13946 = ( n13944 & ~n13945 ) | ( n13944 & 1'b0 ) | ( ~n13945 & 1'b0 ) ;
  assign n13955 = ( n13882 & n13896 ) | ( n13882 & n13946 ) | ( n13896 & n13946 ) ;
  assign n13956 = ( n13882 & ~n13898 ) | ( n13882 & n13946 ) | ( ~n13898 & n13946 ) ;
  assign n13957 = ~n13955 & n13956 ;
  assign n13958 = n13951 | n13957 ;
  assign n13959 = n13538 &  n13899 ;
  assign n13952 = x104 | n13538 ;
  assign n13953 = x104 &  n13538 ;
  assign n13954 = ( n13952 & ~n13953 ) | ( n13952 & 1'b0 ) | ( ~n13953 & 1'b0 ) ;
  assign n13963 = ( n13881 & n13896 ) | ( n13881 & n13954 ) | ( n13896 & n13954 ) ;
  assign n13964 = ( n13881 & ~n13898 ) | ( n13881 & n13954 ) | ( ~n13898 & n13954 ) ;
  assign n13965 = ~n13963 & n13964 ;
  assign n13966 = n13959 | n13965 ;
  assign n13967 = n13546 &  n13899 ;
  assign n13960 = x103 | n13546 ;
  assign n13961 = x103 &  n13546 ;
  assign n13962 = ( n13960 & ~n13961 ) | ( n13960 & 1'b0 ) | ( ~n13961 & 1'b0 ) ;
  assign n13971 = ( n13880 & n13896 ) | ( n13880 & n13962 ) | ( n13896 & n13962 ) ;
  assign n13972 = ( n13880 & ~n13898 ) | ( n13880 & n13962 ) | ( ~n13898 & n13962 ) ;
  assign n13973 = ~n13971 & n13972 ;
  assign n13974 = n13967 | n13973 ;
  assign n13975 = n13554 &  n13899 ;
  assign n13968 = x102 | n13554 ;
  assign n13969 = x102 &  n13554 ;
  assign n13970 = ( n13968 & ~n13969 ) | ( n13968 & 1'b0 ) | ( ~n13969 & 1'b0 ) ;
  assign n13979 = ( n13879 & n13896 ) | ( n13879 & n13970 ) | ( n13896 & n13970 ) ;
  assign n13980 = ( n13879 & ~n13898 ) | ( n13879 & n13970 ) | ( ~n13898 & n13970 ) ;
  assign n13981 = ~n13979 & n13980 ;
  assign n13982 = n13975 | n13981 ;
  assign n13983 = n13562 &  n13899 ;
  assign n13976 = x101 | n13562 ;
  assign n13977 = x101 &  n13562 ;
  assign n13978 = ( n13976 & ~n13977 ) | ( n13976 & 1'b0 ) | ( ~n13977 & 1'b0 ) ;
  assign n13987 = ( n13878 & n13896 ) | ( n13878 & n13978 ) | ( n13896 & n13978 ) ;
  assign n13988 = ( n13878 & ~n13898 ) | ( n13878 & n13978 ) | ( ~n13898 & n13978 ) ;
  assign n13989 = ~n13987 & n13988 ;
  assign n13990 = n13983 | n13989 ;
  assign n13991 = n13570 &  n13899 ;
  assign n13984 = x100 | n13570 ;
  assign n13985 = x100 &  n13570 ;
  assign n13986 = ( n13984 & ~n13985 ) | ( n13984 & 1'b0 ) | ( ~n13985 & 1'b0 ) ;
  assign n13995 = ( n13877 & n13896 ) | ( n13877 & n13986 ) | ( n13896 & n13986 ) ;
  assign n13996 = ( n13877 & ~n13898 ) | ( n13877 & n13986 ) | ( ~n13898 & n13986 ) ;
  assign n13997 = ~n13995 & n13996 ;
  assign n13998 = n13991 | n13997 ;
  assign n13999 = n13578 &  n13899 ;
  assign n13992 = x99 | n13578 ;
  assign n13993 = x99 &  n13578 ;
  assign n13994 = ( n13992 & ~n13993 ) | ( n13992 & 1'b0 ) | ( ~n13993 & 1'b0 ) ;
  assign n14003 = ( n13876 & n13896 ) | ( n13876 & n13994 ) | ( n13896 & n13994 ) ;
  assign n14004 = ( n13876 & ~n13898 ) | ( n13876 & n13994 ) | ( ~n13898 & n13994 ) ;
  assign n14005 = ~n14003 & n14004 ;
  assign n14006 = n13999 | n14005 ;
  assign n14007 = n13586 &  n13899 ;
  assign n14000 = x98 | n13586 ;
  assign n14001 = x98 &  n13586 ;
  assign n14002 = ( n14000 & ~n14001 ) | ( n14000 & 1'b0 ) | ( ~n14001 & 1'b0 ) ;
  assign n14011 = ( n13875 & n13896 ) | ( n13875 & n14002 ) | ( n13896 & n14002 ) ;
  assign n14012 = ( n13875 & ~n13898 ) | ( n13875 & n14002 ) | ( ~n13898 & n14002 ) ;
  assign n14013 = ~n14011 & n14012 ;
  assign n14014 = n14007 | n14013 ;
  assign n14015 = n13594 &  n13899 ;
  assign n14008 = x97 | n13594 ;
  assign n14009 = x97 &  n13594 ;
  assign n14010 = ( n14008 & ~n14009 ) | ( n14008 & 1'b0 ) | ( ~n14009 & 1'b0 ) ;
  assign n14019 = ( n13874 & n13896 ) | ( n13874 & n14010 ) | ( n13896 & n14010 ) ;
  assign n14020 = ( n13874 & ~n13898 ) | ( n13874 & n14010 ) | ( ~n13898 & n14010 ) ;
  assign n14021 = ~n14019 & n14020 ;
  assign n14022 = n14015 | n14021 ;
  assign n14023 = n13602 &  n13899 ;
  assign n14016 = x96 | n13602 ;
  assign n14017 = x96 &  n13602 ;
  assign n14018 = ( n14016 & ~n14017 ) | ( n14016 & 1'b0 ) | ( ~n14017 & 1'b0 ) ;
  assign n14027 = ( n13873 & n13896 ) | ( n13873 & n14018 ) | ( n13896 & n14018 ) ;
  assign n14028 = ( n13873 & ~n13898 ) | ( n13873 & n14018 ) | ( ~n13898 & n14018 ) ;
  assign n14029 = ~n14027 & n14028 ;
  assign n14030 = n14023 | n14029 ;
  assign n14031 = n13610 &  n13899 ;
  assign n14024 = x95 | n13610 ;
  assign n14025 = x95 &  n13610 ;
  assign n14026 = ( n14024 & ~n14025 ) | ( n14024 & 1'b0 ) | ( ~n14025 & 1'b0 ) ;
  assign n14035 = ( n13872 & n13896 ) | ( n13872 & n14026 ) | ( n13896 & n14026 ) ;
  assign n14036 = ( n13872 & ~n13898 ) | ( n13872 & n14026 ) | ( ~n13898 & n14026 ) ;
  assign n14037 = ~n14035 & n14036 ;
  assign n14038 = n14031 | n14037 ;
  assign n14039 = n13618 &  n13899 ;
  assign n14032 = x94 | n13618 ;
  assign n14033 = x94 &  n13618 ;
  assign n14034 = ( n14032 & ~n14033 ) | ( n14032 & 1'b0 ) | ( ~n14033 & 1'b0 ) ;
  assign n14043 = ( n13871 & n13896 ) | ( n13871 & n14034 ) | ( n13896 & n14034 ) ;
  assign n14044 = ( n13871 & ~n13898 ) | ( n13871 & n14034 ) | ( ~n13898 & n14034 ) ;
  assign n14045 = ~n14043 & n14044 ;
  assign n14046 = n14039 | n14045 ;
  assign n14047 = n13626 &  n13899 ;
  assign n14040 = x93 | n13626 ;
  assign n14041 = x93 &  n13626 ;
  assign n14042 = ( n14040 & ~n14041 ) | ( n14040 & 1'b0 ) | ( ~n14041 & 1'b0 ) ;
  assign n14051 = ( n13870 & n13896 ) | ( n13870 & n14042 ) | ( n13896 & n14042 ) ;
  assign n14052 = ( n13870 & ~n13898 ) | ( n13870 & n14042 ) | ( ~n13898 & n14042 ) ;
  assign n14053 = ~n14051 & n14052 ;
  assign n14054 = n14047 | n14053 ;
  assign n14055 = n13634 &  n13899 ;
  assign n14048 = x92 | n13634 ;
  assign n14049 = x92 &  n13634 ;
  assign n14050 = ( n14048 & ~n14049 ) | ( n14048 & 1'b0 ) | ( ~n14049 & 1'b0 ) ;
  assign n14059 = ( n13869 & n13896 ) | ( n13869 & n14050 ) | ( n13896 & n14050 ) ;
  assign n14060 = ( n13869 & ~n13898 ) | ( n13869 & n14050 ) | ( ~n13898 & n14050 ) ;
  assign n14061 = ~n14059 & n14060 ;
  assign n14062 = n14055 | n14061 ;
  assign n14063 = n13642 &  n13899 ;
  assign n14056 = x91 | n13642 ;
  assign n14057 = x91 &  n13642 ;
  assign n14058 = ( n14056 & ~n14057 ) | ( n14056 & 1'b0 ) | ( ~n14057 & 1'b0 ) ;
  assign n14067 = ( n13868 & n13896 ) | ( n13868 & n14058 ) | ( n13896 & n14058 ) ;
  assign n14068 = ( n13868 & ~n13898 ) | ( n13868 & n14058 ) | ( ~n13898 & n14058 ) ;
  assign n14069 = ~n14067 & n14068 ;
  assign n14070 = n14063 | n14069 ;
  assign n14071 = n13650 &  n13899 ;
  assign n14064 = x90 | n13650 ;
  assign n14065 = x90 &  n13650 ;
  assign n14066 = ( n14064 & ~n14065 ) | ( n14064 & 1'b0 ) | ( ~n14065 & 1'b0 ) ;
  assign n14075 = ( n13867 & n13896 ) | ( n13867 & n14066 ) | ( n13896 & n14066 ) ;
  assign n14076 = ( n13867 & ~n13898 ) | ( n13867 & n14066 ) | ( ~n13898 & n14066 ) ;
  assign n14077 = ~n14075 & n14076 ;
  assign n14078 = n14071 | n14077 ;
  assign n14079 = n13658 &  n13899 ;
  assign n14072 = x89 | n13658 ;
  assign n14073 = x89 &  n13658 ;
  assign n14074 = ( n14072 & ~n14073 ) | ( n14072 & 1'b0 ) | ( ~n14073 & 1'b0 ) ;
  assign n14083 = ( n13866 & n13896 ) | ( n13866 & n14074 ) | ( n13896 & n14074 ) ;
  assign n14084 = ( n13866 & ~n13898 ) | ( n13866 & n14074 ) | ( ~n13898 & n14074 ) ;
  assign n14085 = ~n14083 & n14084 ;
  assign n14086 = n14079 | n14085 ;
  assign n14087 = n13666 &  n13899 ;
  assign n14080 = x88 | n13666 ;
  assign n14081 = x88 &  n13666 ;
  assign n14082 = ( n14080 & ~n14081 ) | ( n14080 & 1'b0 ) | ( ~n14081 & 1'b0 ) ;
  assign n14091 = ( n13865 & n13896 ) | ( n13865 & n14082 ) | ( n13896 & n14082 ) ;
  assign n14092 = ( n13865 & ~n13898 ) | ( n13865 & n14082 ) | ( ~n13898 & n14082 ) ;
  assign n14093 = ~n14091 & n14092 ;
  assign n14094 = n14087 | n14093 ;
  assign n14095 = n13674 &  n13899 ;
  assign n14088 = x87 | n13674 ;
  assign n14089 = x87 &  n13674 ;
  assign n14090 = ( n14088 & ~n14089 ) | ( n14088 & 1'b0 ) | ( ~n14089 & 1'b0 ) ;
  assign n14099 = ( n13864 & n13896 ) | ( n13864 & n14090 ) | ( n13896 & n14090 ) ;
  assign n14100 = ( n13864 & ~n13898 ) | ( n13864 & n14090 ) | ( ~n13898 & n14090 ) ;
  assign n14101 = ~n14099 & n14100 ;
  assign n14102 = n14095 | n14101 ;
  assign n14103 = n13682 &  n13899 ;
  assign n14096 = x86 | n13682 ;
  assign n14097 = x86 &  n13682 ;
  assign n14098 = ( n14096 & ~n14097 ) | ( n14096 & 1'b0 ) | ( ~n14097 & 1'b0 ) ;
  assign n14107 = ( n13863 & n13896 ) | ( n13863 & n14098 ) | ( n13896 & n14098 ) ;
  assign n14108 = ( n13863 & ~n13898 ) | ( n13863 & n14098 ) | ( ~n13898 & n14098 ) ;
  assign n14109 = ~n14107 & n14108 ;
  assign n14110 = n14103 | n14109 ;
  assign n14111 = n13690 &  n13899 ;
  assign n14104 = x85 | n13690 ;
  assign n14105 = x85 &  n13690 ;
  assign n14106 = ( n14104 & ~n14105 ) | ( n14104 & 1'b0 ) | ( ~n14105 & 1'b0 ) ;
  assign n14115 = ( n13862 & n13896 ) | ( n13862 & n14106 ) | ( n13896 & n14106 ) ;
  assign n14116 = ( n13862 & ~n13898 ) | ( n13862 & n14106 ) | ( ~n13898 & n14106 ) ;
  assign n14117 = ~n14115 & n14116 ;
  assign n14118 = n14111 | n14117 ;
  assign n14119 = n13698 &  n13899 ;
  assign n14112 = x84 | n13698 ;
  assign n14113 = x84 &  n13698 ;
  assign n14114 = ( n14112 & ~n14113 ) | ( n14112 & 1'b0 ) | ( ~n14113 & 1'b0 ) ;
  assign n14123 = ( n13861 & n13896 ) | ( n13861 & n14114 ) | ( n13896 & n14114 ) ;
  assign n14124 = ( n13861 & ~n13898 ) | ( n13861 & n14114 ) | ( ~n13898 & n14114 ) ;
  assign n14125 = ~n14123 & n14124 ;
  assign n14126 = n14119 | n14125 ;
  assign n14127 = n13706 &  n13899 ;
  assign n14120 = x83 | n13706 ;
  assign n14121 = x83 &  n13706 ;
  assign n14122 = ( n14120 & ~n14121 ) | ( n14120 & 1'b0 ) | ( ~n14121 & 1'b0 ) ;
  assign n14131 = ( n13860 & n13896 ) | ( n13860 & n14122 ) | ( n13896 & n14122 ) ;
  assign n14132 = ( n13860 & ~n13898 ) | ( n13860 & n14122 ) | ( ~n13898 & n14122 ) ;
  assign n14133 = ~n14131 & n14132 ;
  assign n14134 = n14127 | n14133 ;
  assign n14135 = n13714 &  n13899 ;
  assign n14128 = x82 | n13714 ;
  assign n14129 = x82 &  n13714 ;
  assign n14130 = ( n14128 & ~n14129 ) | ( n14128 & 1'b0 ) | ( ~n14129 & 1'b0 ) ;
  assign n14139 = ( n13859 & n13896 ) | ( n13859 & n14130 ) | ( n13896 & n14130 ) ;
  assign n14140 = ( n13859 & ~n13898 ) | ( n13859 & n14130 ) | ( ~n13898 & n14130 ) ;
  assign n14141 = ~n14139 & n14140 ;
  assign n14142 = n14135 | n14141 ;
  assign n14143 = n13722 &  n13899 ;
  assign n14136 = x81 | n13722 ;
  assign n14137 = x81 &  n13722 ;
  assign n14138 = ( n14136 & ~n14137 ) | ( n14136 & 1'b0 ) | ( ~n14137 & 1'b0 ) ;
  assign n14147 = ( n13858 & n13896 ) | ( n13858 & n14138 ) | ( n13896 & n14138 ) ;
  assign n14148 = ( n13858 & ~n13898 ) | ( n13858 & n14138 ) | ( ~n13898 & n14138 ) ;
  assign n14149 = ~n14147 & n14148 ;
  assign n14150 = n14143 | n14149 ;
  assign n14151 = n13730 &  n13899 ;
  assign n14144 = x80 | n13730 ;
  assign n14145 = x80 &  n13730 ;
  assign n14146 = ( n14144 & ~n14145 ) | ( n14144 & 1'b0 ) | ( ~n14145 & 1'b0 ) ;
  assign n14155 = ( n13857 & n13896 ) | ( n13857 & n14146 ) | ( n13896 & n14146 ) ;
  assign n14156 = ( n13857 & ~n13898 ) | ( n13857 & n14146 ) | ( ~n13898 & n14146 ) ;
  assign n14157 = ~n14155 & n14156 ;
  assign n14158 = n14151 | n14157 ;
  assign n14159 = n13738 &  n13899 ;
  assign n14152 = x79 | n13738 ;
  assign n14153 = x79 &  n13738 ;
  assign n14154 = ( n14152 & ~n14153 ) | ( n14152 & 1'b0 ) | ( ~n14153 & 1'b0 ) ;
  assign n14163 = ( n13856 & n13896 ) | ( n13856 & n14154 ) | ( n13896 & n14154 ) ;
  assign n14164 = ( n13856 & ~n13898 ) | ( n13856 & n14154 ) | ( ~n13898 & n14154 ) ;
  assign n14165 = ~n14163 & n14164 ;
  assign n14166 = n14159 | n14165 ;
  assign n14167 = n13746 &  n13899 ;
  assign n14160 = x78 | n13746 ;
  assign n14161 = x78 &  n13746 ;
  assign n14162 = ( n14160 & ~n14161 ) | ( n14160 & 1'b0 ) | ( ~n14161 & 1'b0 ) ;
  assign n14171 = ( n13855 & n13896 ) | ( n13855 & n14162 ) | ( n13896 & n14162 ) ;
  assign n14172 = ( n13855 & ~n13898 ) | ( n13855 & n14162 ) | ( ~n13898 & n14162 ) ;
  assign n14173 = ~n14171 & n14172 ;
  assign n14174 = n14167 | n14173 ;
  assign n14175 = n13754 &  n13899 ;
  assign n14168 = x77 | n13754 ;
  assign n14169 = x77 &  n13754 ;
  assign n14170 = ( n14168 & ~n14169 ) | ( n14168 & 1'b0 ) | ( ~n14169 & 1'b0 ) ;
  assign n14179 = ( n13854 & n13896 ) | ( n13854 & n14170 ) | ( n13896 & n14170 ) ;
  assign n14180 = ( n13854 & ~n13898 ) | ( n13854 & n14170 ) | ( ~n13898 & n14170 ) ;
  assign n14181 = ~n14179 & n14180 ;
  assign n14182 = n14175 | n14181 ;
  assign n14183 = n13762 &  n13899 ;
  assign n14176 = x76 | n13762 ;
  assign n14177 = x76 &  n13762 ;
  assign n14178 = ( n14176 & ~n14177 ) | ( n14176 & 1'b0 ) | ( ~n14177 & 1'b0 ) ;
  assign n14187 = ( n13853 & n13896 ) | ( n13853 & n14178 ) | ( n13896 & n14178 ) ;
  assign n14188 = ( n13853 & ~n13898 ) | ( n13853 & n14178 ) | ( ~n13898 & n14178 ) ;
  assign n14189 = ~n14187 & n14188 ;
  assign n14190 = n14183 | n14189 ;
  assign n14191 = n13770 &  n13899 ;
  assign n14184 = x75 | n13770 ;
  assign n14185 = x75 &  n13770 ;
  assign n14186 = ( n14184 & ~n14185 ) | ( n14184 & 1'b0 ) | ( ~n14185 & 1'b0 ) ;
  assign n14195 = ( n13852 & n13896 ) | ( n13852 & n14186 ) | ( n13896 & n14186 ) ;
  assign n14196 = ( n13852 & ~n13898 ) | ( n13852 & n14186 ) | ( ~n13898 & n14186 ) ;
  assign n14197 = ~n14195 & n14196 ;
  assign n14198 = n14191 | n14197 ;
  assign n14199 = n13778 &  n13899 ;
  assign n14192 = x74 | n13778 ;
  assign n14193 = x74 &  n13778 ;
  assign n14194 = ( n14192 & ~n14193 ) | ( n14192 & 1'b0 ) | ( ~n14193 & 1'b0 ) ;
  assign n14203 = ( n13851 & n13896 ) | ( n13851 & n14194 ) | ( n13896 & n14194 ) ;
  assign n14204 = ( n13851 & ~n13898 ) | ( n13851 & n14194 ) | ( ~n13898 & n14194 ) ;
  assign n14205 = ~n14203 & n14204 ;
  assign n14206 = n14199 | n14205 ;
  assign n14207 = n13786 &  n13899 ;
  assign n14200 = x73 | n13786 ;
  assign n14201 = x73 &  n13786 ;
  assign n14202 = ( n14200 & ~n14201 ) | ( n14200 & 1'b0 ) | ( ~n14201 & 1'b0 ) ;
  assign n14211 = ( n13850 & n13896 ) | ( n13850 & n14202 ) | ( n13896 & n14202 ) ;
  assign n14212 = ( n13850 & ~n13898 ) | ( n13850 & n14202 ) | ( ~n13898 & n14202 ) ;
  assign n14213 = ~n14211 & n14212 ;
  assign n14214 = n14207 | n14213 ;
  assign n14215 = n13794 &  n13899 ;
  assign n14208 = x72 | n13794 ;
  assign n14209 = x72 &  n13794 ;
  assign n14210 = ( n14208 & ~n14209 ) | ( n14208 & 1'b0 ) | ( ~n14209 & 1'b0 ) ;
  assign n14219 = ( n13849 & n13896 ) | ( n13849 & n14210 ) | ( n13896 & n14210 ) ;
  assign n14220 = ( n13849 & ~n13898 ) | ( n13849 & n14210 ) | ( ~n13898 & n14210 ) ;
  assign n14221 = ~n14219 & n14220 ;
  assign n14222 = n14215 | n14221 ;
  assign n14223 = n13802 &  n13899 ;
  assign n14216 = x71 | n13802 ;
  assign n14217 = x71 &  n13802 ;
  assign n14218 = ( n14216 & ~n14217 ) | ( n14216 & 1'b0 ) | ( ~n14217 & 1'b0 ) ;
  assign n14227 = ( n13848 & n13896 ) | ( n13848 & n14218 ) | ( n13896 & n14218 ) ;
  assign n14228 = ( n13848 & ~n13898 ) | ( n13848 & n14218 ) | ( ~n13898 & n14218 ) ;
  assign n14229 = ~n14227 & n14228 ;
  assign n14230 = n14223 | n14229 ;
  assign n14231 = n13810 &  n13899 ;
  assign n14224 = x70 | n13810 ;
  assign n14225 = x70 &  n13810 ;
  assign n14226 = ( n14224 & ~n14225 ) | ( n14224 & 1'b0 ) | ( ~n14225 & 1'b0 ) ;
  assign n14235 = ( n13847 & n13896 ) | ( n13847 & n14226 ) | ( n13896 & n14226 ) ;
  assign n14236 = ( n13847 & ~n13898 ) | ( n13847 & n14226 ) | ( ~n13898 & n14226 ) ;
  assign n14237 = ~n14235 & n14236 ;
  assign n14238 = n14231 | n14237 ;
  assign n14239 = n13818 &  n13899 ;
  assign n14232 = x69 | n13818 ;
  assign n14233 = x69 &  n13818 ;
  assign n14234 = ( n14232 & ~n14233 ) | ( n14232 & 1'b0 ) | ( ~n14233 & 1'b0 ) ;
  assign n14243 = ( n13846 & n13896 ) | ( n13846 & n14234 ) | ( n13896 & n14234 ) ;
  assign n14244 = ( n13846 & ~n13898 ) | ( n13846 & n14234 ) | ( ~n13898 & n14234 ) ;
  assign n14245 = ~n14243 & n14244 ;
  assign n14246 = n14239 | n14245 ;
  assign n14247 = n13826 &  n13899 ;
  assign n14240 = x68 | n13826 ;
  assign n14241 = x68 &  n13826 ;
  assign n14242 = ( n14240 & ~n14241 ) | ( n14240 & 1'b0 ) | ( ~n14241 & 1'b0 ) ;
  assign n14251 = ( n13845 & n13896 ) | ( n13845 & n14242 ) | ( n13896 & n14242 ) ;
  assign n14252 = ( n13845 & ~n13898 ) | ( n13845 & n14242 ) | ( ~n13898 & n14242 ) ;
  assign n14253 = ~n14251 & n14252 ;
  assign n14254 = n14247 | n14253 ;
  assign n14255 = n13831 &  n13899 ;
  assign n14248 = x67 | n13831 ;
  assign n14249 = x67 &  n13831 ;
  assign n14250 = ( n14248 & ~n14249 ) | ( n14248 & 1'b0 ) | ( ~n14249 & 1'b0 ) ;
  assign n14259 = ( n13844 & n13896 ) | ( n13844 & n14250 ) | ( n13896 & n14250 ) ;
  assign n14260 = ( n13844 & ~n13898 ) | ( n13844 & n14250 ) | ( ~n13898 & n14250 ) ;
  assign n14261 = ~n14259 & n14260 ;
  assign n14262 = n14255 | n14261 ;
  assign n14263 = n13837 &  n13899 ;
  assign n14256 = x66 | n13837 ;
  assign n14257 = x66 &  n13837 ;
  assign n14258 = ( n14256 & ~n14257 ) | ( n14256 & 1'b0 ) | ( ~n14257 & 1'b0 ) ;
  assign n14268 = ( n13843 & ~n13896 ) | ( n13843 & n14258 ) | ( ~n13896 & n14258 ) ;
  assign n14269 = ( n13843 & n13898 ) | ( n13843 & n14258 ) | ( n13898 & n14258 ) ;
  assign n14270 = ( n14268 & ~n14269 ) | ( n14268 & 1'b0 ) | ( ~n14269 & 1'b0 ) ;
  assign n14271 = n14263 | n14270 ;
  assign n14272 = n13841 &  n13899 ;
  assign n14264 = x65 &  n13841 ;
  assign n14265 = ( n13839 & ~x65 ) | ( n13839 & n13840 ) | ( ~x65 & n13840 ) ;
  assign n14266 = x65 | n14265 ;
  assign n14267 = ( n13842 & ~n14264 ) | ( n13842 & n14266 ) | ( ~n14264 & n14266 ) ;
  assign n14273 = ( x65 & n13841 ) | ( x65 & n13842 ) | ( n13841 & n13842 ) ;
  assign n14274 = ( n13898 & ~n14264 ) | ( n13898 & n14273 ) | ( ~n14264 & n14273 ) ;
  assign n14275 = ( n13896 & n14267 ) | ( n13896 & n14274 ) | ( n14267 & n14274 ) ;
  assign n14276 = ( n14267 & ~n14275 ) | ( n14267 & 1'b0 ) | ( ~n14275 & 1'b0 ) ;
  assign n14277 = n14272 | n14276 ;
  assign n14278 = ( x64 & ~x119 ) | ( x64 & 1'b0 ) | ( ~x119 & 1'b0 ) ;
  assign n14279 = ( n152 & ~n155 ) | ( n152 & n14278 ) | ( ~n155 & n14278 ) ;
  assign n14280 = ~n152 & n14279 ;
  assign n14281 = n13896 &  n14280 ;
  assign n14282 = ( x9 & ~n14280 ) | ( x9 & n14281 ) | ( ~n14280 & n14281 ) ;
  assign n14283 = ~n228 & n13842 ;
  assign n14284 = ( n235 & ~n238 ) | ( n235 & n14283 ) | ( ~n238 & n14283 ) ;
  assign n14285 = ~n235 & n14284 ;
  assign n14286 = ~n13896 & n14285 ;
  assign n14287 = n14282 | n14286 ;
  assign n14288 = ~x8 & x64 ;
  assign n14289 = ( x65 & ~n14287 ) | ( x65 & n14288 ) | ( ~n14287 & n14288 ) ;
  assign n14290 = ( x66 & ~n14277 ) | ( x66 & n14289 ) | ( ~n14277 & n14289 ) ;
  assign n14291 = ( x67 & ~n14271 ) | ( x67 & n14290 ) | ( ~n14271 & n14290 ) ;
  assign n14292 = ( x68 & ~n14262 ) | ( x68 & n14291 ) | ( ~n14262 & n14291 ) ;
  assign n14293 = ( x69 & ~n14254 ) | ( x69 & n14292 ) | ( ~n14254 & n14292 ) ;
  assign n14294 = ( x70 & ~n14246 ) | ( x70 & n14293 ) | ( ~n14246 & n14293 ) ;
  assign n14295 = ( x71 & ~n14238 ) | ( x71 & n14294 ) | ( ~n14238 & n14294 ) ;
  assign n14296 = ( x72 & ~n14230 ) | ( x72 & n14295 ) | ( ~n14230 & n14295 ) ;
  assign n14297 = ( x73 & ~n14222 ) | ( x73 & n14296 ) | ( ~n14222 & n14296 ) ;
  assign n14298 = ( x74 & ~n14214 ) | ( x74 & n14297 ) | ( ~n14214 & n14297 ) ;
  assign n14299 = ( x75 & ~n14206 ) | ( x75 & n14298 ) | ( ~n14206 & n14298 ) ;
  assign n14300 = ( x76 & ~n14198 ) | ( x76 & n14299 ) | ( ~n14198 & n14299 ) ;
  assign n14301 = ( x77 & ~n14190 ) | ( x77 & n14300 ) | ( ~n14190 & n14300 ) ;
  assign n14302 = ( x78 & ~n14182 ) | ( x78 & n14301 ) | ( ~n14182 & n14301 ) ;
  assign n14303 = ( x79 & ~n14174 ) | ( x79 & n14302 ) | ( ~n14174 & n14302 ) ;
  assign n14304 = ( x80 & ~n14166 ) | ( x80 & n14303 ) | ( ~n14166 & n14303 ) ;
  assign n14305 = ( x81 & ~n14158 ) | ( x81 & n14304 ) | ( ~n14158 & n14304 ) ;
  assign n14306 = ( x82 & ~n14150 ) | ( x82 & n14305 ) | ( ~n14150 & n14305 ) ;
  assign n14307 = ( x83 & ~n14142 ) | ( x83 & n14306 ) | ( ~n14142 & n14306 ) ;
  assign n14308 = ( x84 & ~n14134 ) | ( x84 & n14307 ) | ( ~n14134 & n14307 ) ;
  assign n14309 = ( x85 & ~n14126 ) | ( x85 & n14308 ) | ( ~n14126 & n14308 ) ;
  assign n14310 = ( x86 & ~n14118 ) | ( x86 & n14309 ) | ( ~n14118 & n14309 ) ;
  assign n14311 = ( x87 & ~n14110 ) | ( x87 & n14310 ) | ( ~n14110 & n14310 ) ;
  assign n14312 = ( x88 & ~n14102 ) | ( x88 & n14311 ) | ( ~n14102 & n14311 ) ;
  assign n14313 = ( x89 & ~n14094 ) | ( x89 & n14312 ) | ( ~n14094 & n14312 ) ;
  assign n14314 = ( x90 & ~n14086 ) | ( x90 & n14313 ) | ( ~n14086 & n14313 ) ;
  assign n14315 = ( x91 & ~n14078 ) | ( x91 & n14314 ) | ( ~n14078 & n14314 ) ;
  assign n14316 = ( x92 & ~n14070 ) | ( x92 & n14315 ) | ( ~n14070 & n14315 ) ;
  assign n14317 = ( x93 & ~n14062 ) | ( x93 & n14316 ) | ( ~n14062 & n14316 ) ;
  assign n14318 = ( x94 & ~n14054 ) | ( x94 & n14317 ) | ( ~n14054 & n14317 ) ;
  assign n14319 = ( x95 & ~n14046 ) | ( x95 & n14318 ) | ( ~n14046 & n14318 ) ;
  assign n14320 = ( x96 & ~n14038 ) | ( x96 & n14319 ) | ( ~n14038 & n14319 ) ;
  assign n14321 = ( x97 & ~n14030 ) | ( x97 & n14320 ) | ( ~n14030 & n14320 ) ;
  assign n14322 = ( x98 & ~n14022 ) | ( x98 & n14321 ) | ( ~n14022 & n14321 ) ;
  assign n14323 = ( x99 & ~n14014 ) | ( x99 & n14322 ) | ( ~n14014 & n14322 ) ;
  assign n14324 = ( x100 & ~n14006 ) | ( x100 & n14323 ) | ( ~n14006 & n14323 ) ;
  assign n14325 = ( x101 & ~n13998 ) | ( x101 & n14324 ) | ( ~n13998 & n14324 ) ;
  assign n14326 = ( x102 & ~n13990 ) | ( x102 & n14325 ) | ( ~n13990 & n14325 ) ;
  assign n14327 = ( x103 & ~n13982 ) | ( x103 & n14326 ) | ( ~n13982 & n14326 ) ;
  assign n14328 = ( x104 & ~n13974 ) | ( x104 & n14327 ) | ( ~n13974 & n14327 ) ;
  assign n14329 = ( x105 & ~n13966 ) | ( x105 & n14328 ) | ( ~n13966 & n14328 ) ;
  assign n14330 = ( x106 & ~n13958 ) | ( x106 & n14329 ) | ( ~n13958 & n14329 ) ;
  assign n14331 = ( x107 & ~n13950 ) | ( x107 & n14330 ) | ( ~n13950 & n14330 ) ;
  assign n14332 = ( x108 & ~n13942 ) | ( x108 & n14331 ) | ( ~n13942 & n14331 ) ;
  assign n14333 = ( x109 & ~n13934 ) | ( x109 & n14332 ) | ( ~n13934 & n14332 ) ;
  assign n14334 = ( x110 & ~n13926 ) | ( x110 & n14333 ) | ( ~n13926 & n14333 ) ;
  assign n14335 = ( x111 & ~n13918 ) | ( x111 & n14334 ) | ( ~n13918 & n14334 ) ;
  assign n14339 = ( x112 & ~n13910 ) | ( x112 & n14335 ) | ( ~n13910 & n14335 ) ;
  assign n14391 = ( x113 & ~n14347 ) | ( x113 & n14339 ) | ( ~n14347 & n14339 ) ;
  assign n14392 = ( x114 & ~n14390 ) | ( x114 & n14391 ) | ( ~n14390 & n14391 ) ;
  assign n14393 = ( x115 & ~n14385 ) | ( x115 & n14392 ) | ( ~n14385 & n14392 ) ;
  assign n14394 = ( x116 & ~n14377 ) | ( x116 & n14393 ) | ( ~n14377 & n14393 ) ;
  assign n14395 = ( x117 & ~n14369 ) | ( x117 & n14394 ) | ( ~n14369 & n14394 ) ;
  assign n14396 = ( x118 & ~n14361 ) | ( x118 & n14395 ) | ( ~n14361 & n14395 ) ;
  assign n14397 = n13437 &  n13899 ;
  assign n14398 = ( n13437 & ~n13898 ) | ( n13437 & n13895 ) | ( ~n13898 & n13895 ) ;
  assign n14399 = ( x118 & ~n13895 ) | ( x118 & n14398 ) | ( ~n13895 & n14398 ) ;
  assign n14400 = ~x118 & n14399 ;
  assign n14401 = n14397 | n14400 ;
  assign n14402 = ~x119 & n14401 ;
  assign n14403 = ( x119 & ~n14397 ) | ( x119 & 1'b0 ) | ( ~n14397 & 1'b0 ) ;
  assign n14404 = ~n14400 & n14403 ;
  assign n14405 = n269 | n14404 ;
  assign n14406 = n14402 | n14405 ;
  assign n14407 = n14396 | n14406 ;
  assign n14408 = ~n14401 |  n13898 ;
  assign n14869 = n14361 &  n14408 ;
  assign n14870 = n14407 &  n14869 ;
  assign n14866 = x118 | n14361 ;
  assign n14867 = x118 &  n14361 ;
  assign n14868 = ( n14866 & ~n14867 ) | ( n14866 & 1'b0 ) | ( ~n14867 & 1'b0 ) ;
  assign n14871 = n14395 &  n14868 ;
  assign n14409 = n14407 &  n14408 ;
  assign n14872 = ( n14395 & ~n14409 ) | ( n14395 & n14868 ) | ( ~n14409 & n14868 ) ;
  assign n14873 = ( n14870 & ~n14871 ) | ( n14870 & n14872 ) | ( ~n14871 & n14872 ) ;
  assign n14877 = n14369 &  n14408 ;
  assign n14878 = n14407 &  n14877 ;
  assign n14863 = x117 | n14369 ;
  assign n14864 = x117 &  n14369 ;
  assign n14865 = ( n14863 & ~n14864 ) | ( n14863 & 1'b0 ) | ( ~n14864 & 1'b0 ) ;
  assign n14879 = n14394 &  n14865 ;
  assign n14880 = ( n14394 & ~n14409 ) | ( n14394 & n14865 ) | ( ~n14409 & n14865 ) ;
  assign n14881 = ( n14878 & ~n14879 ) | ( n14878 & n14880 ) | ( ~n14879 & n14880 ) ;
  assign n14885 = n14377 &  n14408 ;
  assign n14886 = n14407 &  n14885 ;
  assign n14874 = x116 | n14377 ;
  assign n14875 = x116 &  n14377 ;
  assign n14876 = ( n14874 & ~n14875 ) | ( n14874 & 1'b0 ) | ( ~n14875 & 1'b0 ) ;
  assign n14887 = n14393 &  n14876 ;
  assign n14888 = ( n14393 & ~n14409 ) | ( n14393 & n14876 ) | ( ~n14409 & n14876 ) ;
  assign n14889 = ( n14886 & ~n14887 ) | ( n14886 & n14888 ) | ( ~n14887 & n14888 ) ;
  assign n14890 = n14385 &  n14408 ;
  assign n14891 = n14407 &  n14890 ;
  assign n14882 = x115 | n14385 ;
  assign n14883 = x115 &  n14385 ;
  assign n14884 = ( n14882 & ~n14883 ) | ( n14882 & 1'b0 ) | ( ~n14883 & 1'b0 ) ;
  assign n14892 = n14392 &  n14884 ;
  assign n14893 = ( n14392 & ~n14409 ) | ( n14392 & n14884 ) | ( ~n14409 & n14884 ) ;
  assign n14894 = ( n14891 & ~n14892 ) | ( n14891 & n14893 ) | ( ~n14892 & n14893 ) ;
  assign n14855 = n14390 &  n14408 ;
  assign n14856 = n14407 &  n14855 ;
  assign n14852 = x114 | n14390 ;
  assign n14853 = x114 &  n14390 ;
  assign n14854 = ( n14852 & ~n14853 ) | ( n14852 & 1'b0 ) | ( ~n14853 & 1'b0 ) ;
  assign n14857 = n14391 &  n14854 ;
  assign n14858 = ( n14391 & ~n14409 ) | ( n14391 & n14854 ) | ( ~n14409 & n14854 ) ;
  assign n14859 = ( n14856 & ~n14857 ) | ( n14856 & n14858 ) | ( ~n14857 & n14858 ) ;
  assign n14410 = n14347 &  n14408 ;
  assign n14411 = n14407 &  n14410 ;
  assign n14348 = x113 | n14347 ;
  assign n14349 = x113 &  n14347 ;
  assign n14350 = ( n14348 & ~n14349 ) | ( n14348 & 1'b0 ) | ( ~n14349 & 1'b0 ) ;
  assign n14413 = ( n14339 & n14350 ) | ( n14339 & n14409 ) | ( n14350 & n14409 ) ;
  assign n14412 = n14339 | n14350 ;
  assign n14414 = ( n14411 & ~n14413 ) | ( n14411 & n14412 ) | ( ~n14413 & n14412 ) ;
  assign n14418 = n13910 &  n14408 ;
  assign n14419 = n14407 &  n14418 ;
  assign n14336 = x112 | n13910 ;
  assign n14337 = x112 &  n13910 ;
  assign n14338 = ( n14336 & ~n14337 ) | ( n14336 & 1'b0 ) | ( ~n14337 & 1'b0 ) ;
  assign n14420 = n14335 &  n14338 ;
  assign n14421 = ( n14335 & ~n14409 ) | ( n14335 & n14338 ) | ( ~n14409 & n14338 ) ;
  assign n14422 = ( n14419 & ~n14420 ) | ( n14419 & n14421 ) | ( ~n14420 & n14421 ) ;
  assign n14426 = n13918 &  n14408 ;
  assign n14427 = n14407 &  n14426 ;
  assign n14415 = x111 | n13918 ;
  assign n14416 = x111 &  n13918 ;
  assign n14417 = ( n14415 & ~n14416 ) | ( n14415 & 1'b0 ) | ( ~n14416 & 1'b0 ) ;
  assign n14429 = ( n14334 & n14409 ) | ( n14334 & n14417 ) | ( n14409 & n14417 ) ;
  assign n14428 = n14334 | n14417 ;
  assign n14430 = ( n14427 & ~n14429 ) | ( n14427 & n14428 ) | ( ~n14429 & n14428 ) ;
  assign n14434 = n13926 &  n14408 ;
  assign n14435 = n14407 &  n14434 ;
  assign n14423 = x110 | n13926 ;
  assign n14424 = x110 &  n13926 ;
  assign n14425 = ( n14423 & ~n14424 ) | ( n14423 & 1'b0 ) | ( ~n14424 & 1'b0 ) ;
  assign n14437 = ( n14333 & n14409 ) | ( n14333 & n14425 ) | ( n14409 & n14425 ) ;
  assign n14436 = n14333 | n14425 ;
  assign n14438 = ( n14435 & ~n14437 ) | ( n14435 & n14436 ) | ( ~n14437 & n14436 ) ;
  assign n14442 = n13934 &  n14408 ;
  assign n14443 = n14407 &  n14442 ;
  assign n14431 = x109 | n13934 ;
  assign n14432 = x109 &  n13934 ;
  assign n14433 = ( n14431 & ~n14432 ) | ( n14431 & 1'b0 ) | ( ~n14432 & 1'b0 ) ;
  assign n14445 = ( n14332 & n14409 ) | ( n14332 & n14433 ) | ( n14409 & n14433 ) ;
  assign n14444 = n14332 | n14433 ;
  assign n14446 = ( n14443 & ~n14445 ) | ( n14443 & n14444 ) | ( ~n14445 & n14444 ) ;
  assign n14450 = n13942 &  n14408 ;
  assign n14451 = n14407 &  n14450 ;
  assign n14439 = x108 | n13942 ;
  assign n14440 = x108 &  n13942 ;
  assign n14441 = ( n14439 & ~n14440 ) | ( n14439 & 1'b0 ) | ( ~n14440 & 1'b0 ) ;
  assign n14453 = ( n14331 & n14409 ) | ( n14331 & n14441 ) | ( n14409 & n14441 ) ;
  assign n14452 = n14331 | n14441 ;
  assign n14454 = ( n14451 & ~n14453 ) | ( n14451 & n14452 ) | ( ~n14453 & n14452 ) ;
  assign n14458 = n13950 &  n14408 ;
  assign n14459 = n14407 &  n14458 ;
  assign n14447 = x107 | n13950 ;
  assign n14448 = x107 &  n13950 ;
  assign n14449 = ( n14447 & ~n14448 ) | ( n14447 & 1'b0 ) | ( ~n14448 & 1'b0 ) ;
  assign n14461 = ( n14330 & n14409 ) | ( n14330 & n14449 ) | ( n14409 & n14449 ) ;
  assign n14460 = n14330 | n14449 ;
  assign n14462 = ( n14459 & ~n14461 ) | ( n14459 & n14460 ) | ( ~n14461 & n14460 ) ;
  assign n14466 = n13958 &  n14408 ;
  assign n14467 = n14407 &  n14466 ;
  assign n14455 = x106 | n13958 ;
  assign n14456 = x106 &  n13958 ;
  assign n14457 = ( n14455 & ~n14456 ) | ( n14455 & 1'b0 ) | ( ~n14456 & 1'b0 ) ;
  assign n14469 = ( n14329 & n14409 ) | ( n14329 & n14457 ) | ( n14409 & n14457 ) ;
  assign n14468 = n14329 | n14457 ;
  assign n14470 = ( n14467 & ~n14469 ) | ( n14467 & n14468 ) | ( ~n14469 & n14468 ) ;
  assign n14474 = n13966 &  n14408 ;
  assign n14475 = n14407 &  n14474 ;
  assign n14463 = x105 | n13966 ;
  assign n14464 = x105 &  n13966 ;
  assign n14465 = ( n14463 & ~n14464 ) | ( n14463 & 1'b0 ) | ( ~n14464 & 1'b0 ) ;
  assign n14477 = ( n14328 & n14409 ) | ( n14328 & n14465 ) | ( n14409 & n14465 ) ;
  assign n14476 = n14328 | n14465 ;
  assign n14478 = ( n14475 & ~n14477 ) | ( n14475 & n14476 ) | ( ~n14477 & n14476 ) ;
  assign n14482 = n13974 &  n14408 ;
  assign n14483 = n14407 &  n14482 ;
  assign n14471 = x104 | n13974 ;
  assign n14472 = x104 &  n13974 ;
  assign n14473 = ( n14471 & ~n14472 ) | ( n14471 & 1'b0 ) | ( ~n14472 & 1'b0 ) ;
  assign n14485 = ( n14327 & n14409 ) | ( n14327 & n14473 ) | ( n14409 & n14473 ) ;
  assign n14484 = n14327 | n14473 ;
  assign n14486 = ( n14483 & ~n14485 ) | ( n14483 & n14484 ) | ( ~n14485 & n14484 ) ;
  assign n14490 = n13982 &  n14408 ;
  assign n14491 = n14407 &  n14490 ;
  assign n14479 = x103 | n13982 ;
  assign n14480 = x103 &  n13982 ;
  assign n14481 = ( n14479 & ~n14480 ) | ( n14479 & 1'b0 ) | ( ~n14480 & 1'b0 ) ;
  assign n14493 = ( n14326 & n14409 ) | ( n14326 & n14481 ) | ( n14409 & n14481 ) ;
  assign n14492 = n14326 | n14481 ;
  assign n14494 = ( n14491 & ~n14493 ) | ( n14491 & n14492 ) | ( ~n14493 & n14492 ) ;
  assign n14498 = n13990 &  n14408 ;
  assign n14499 = n14407 &  n14498 ;
  assign n14487 = x102 | n13990 ;
  assign n14488 = x102 &  n13990 ;
  assign n14489 = ( n14487 & ~n14488 ) | ( n14487 & 1'b0 ) | ( ~n14488 & 1'b0 ) ;
  assign n14501 = ( n14325 & n14409 ) | ( n14325 & n14489 ) | ( n14409 & n14489 ) ;
  assign n14500 = n14325 | n14489 ;
  assign n14502 = ( n14499 & ~n14501 ) | ( n14499 & n14500 ) | ( ~n14501 & n14500 ) ;
  assign n14506 = n13998 &  n14408 ;
  assign n14507 = n14407 &  n14506 ;
  assign n14495 = x101 | n13998 ;
  assign n14496 = x101 &  n13998 ;
  assign n14497 = ( n14495 & ~n14496 ) | ( n14495 & 1'b0 ) | ( ~n14496 & 1'b0 ) ;
  assign n14509 = ( n14324 & n14409 ) | ( n14324 & n14497 ) | ( n14409 & n14497 ) ;
  assign n14508 = n14324 | n14497 ;
  assign n14510 = ( n14507 & ~n14509 ) | ( n14507 & n14508 ) | ( ~n14509 & n14508 ) ;
  assign n14514 = n14006 &  n14408 ;
  assign n14515 = n14407 &  n14514 ;
  assign n14503 = x100 | n14006 ;
  assign n14504 = x100 &  n14006 ;
  assign n14505 = ( n14503 & ~n14504 ) | ( n14503 & 1'b0 ) | ( ~n14504 & 1'b0 ) ;
  assign n14517 = ( n14323 & n14409 ) | ( n14323 & n14505 ) | ( n14409 & n14505 ) ;
  assign n14516 = n14323 | n14505 ;
  assign n14518 = ( n14515 & ~n14517 ) | ( n14515 & n14516 ) | ( ~n14517 & n14516 ) ;
  assign n14522 = n14014 &  n14408 ;
  assign n14523 = n14407 &  n14522 ;
  assign n14511 = x99 | n14014 ;
  assign n14512 = x99 &  n14014 ;
  assign n14513 = ( n14511 & ~n14512 ) | ( n14511 & 1'b0 ) | ( ~n14512 & 1'b0 ) ;
  assign n14525 = ( n14322 & n14409 ) | ( n14322 & n14513 ) | ( n14409 & n14513 ) ;
  assign n14524 = n14322 | n14513 ;
  assign n14526 = ( n14523 & ~n14525 ) | ( n14523 & n14524 ) | ( ~n14525 & n14524 ) ;
  assign n14530 = n14022 &  n14408 ;
  assign n14531 = n14407 &  n14530 ;
  assign n14519 = x98 | n14022 ;
  assign n14520 = x98 &  n14022 ;
  assign n14521 = ( n14519 & ~n14520 ) | ( n14519 & 1'b0 ) | ( ~n14520 & 1'b0 ) ;
  assign n14533 = ( n14321 & n14409 ) | ( n14321 & n14521 ) | ( n14409 & n14521 ) ;
  assign n14532 = n14321 | n14521 ;
  assign n14534 = ( n14531 & ~n14533 ) | ( n14531 & n14532 ) | ( ~n14533 & n14532 ) ;
  assign n14538 = n14030 &  n14408 ;
  assign n14539 = n14407 &  n14538 ;
  assign n14527 = x97 | n14030 ;
  assign n14528 = x97 &  n14030 ;
  assign n14529 = ( n14527 & ~n14528 ) | ( n14527 & 1'b0 ) | ( ~n14528 & 1'b0 ) ;
  assign n14541 = ( n14320 & n14409 ) | ( n14320 & n14529 ) | ( n14409 & n14529 ) ;
  assign n14540 = n14320 | n14529 ;
  assign n14542 = ( n14539 & ~n14541 ) | ( n14539 & n14540 ) | ( ~n14541 & n14540 ) ;
  assign n14546 = n14038 &  n14408 ;
  assign n14547 = n14407 &  n14546 ;
  assign n14535 = x96 | n14038 ;
  assign n14536 = x96 &  n14038 ;
  assign n14537 = ( n14535 & ~n14536 ) | ( n14535 & 1'b0 ) | ( ~n14536 & 1'b0 ) ;
  assign n14549 = ( n14319 & n14409 ) | ( n14319 & n14537 ) | ( n14409 & n14537 ) ;
  assign n14548 = n14319 | n14537 ;
  assign n14550 = ( n14547 & ~n14549 ) | ( n14547 & n14548 ) | ( ~n14549 & n14548 ) ;
  assign n14554 = n14046 &  n14408 ;
  assign n14555 = n14407 &  n14554 ;
  assign n14543 = x95 | n14046 ;
  assign n14544 = x95 &  n14046 ;
  assign n14545 = ( n14543 & ~n14544 ) | ( n14543 & 1'b0 ) | ( ~n14544 & 1'b0 ) ;
  assign n14557 = ( n14318 & n14409 ) | ( n14318 & n14545 ) | ( n14409 & n14545 ) ;
  assign n14556 = n14318 | n14545 ;
  assign n14558 = ( n14555 & ~n14557 ) | ( n14555 & n14556 ) | ( ~n14557 & n14556 ) ;
  assign n14562 = n14054 &  n14408 ;
  assign n14563 = n14407 &  n14562 ;
  assign n14551 = x94 | n14054 ;
  assign n14552 = x94 &  n14054 ;
  assign n14553 = ( n14551 & ~n14552 ) | ( n14551 & 1'b0 ) | ( ~n14552 & 1'b0 ) ;
  assign n14565 = ( n14317 & n14409 ) | ( n14317 & n14553 ) | ( n14409 & n14553 ) ;
  assign n14564 = n14317 | n14553 ;
  assign n14566 = ( n14563 & ~n14565 ) | ( n14563 & n14564 ) | ( ~n14565 & n14564 ) ;
  assign n14570 = n14062 &  n14408 ;
  assign n14571 = n14407 &  n14570 ;
  assign n14559 = x93 | n14062 ;
  assign n14560 = x93 &  n14062 ;
  assign n14561 = ( n14559 & ~n14560 ) | ( n14559 & 1'b0 ) | ( ~n14560 & 1'b0 ) ;
  assign n14573 = ( n14316 & n14409 ) | ( n14316 & n14561 ) | ( n14409 & n14561 ) ;
  assign n14572 = n14316 | n14561 ;
  assign n14574 = ( n14571 & ~n14573 ) | ( n14571 & n14572 ) | ( ~n14573 & n14572 ) ;
  assign n14578 = n14070 &  n14408 ;
  assign n14579 = n14407 &  n14578 ;
  assign n14567 = x92 | n14070 ;
  assign n14568 = x92 &  n14070 ;
  assign n14569 = ( n14567 & ~n14568 ) | ( n14567 & 1'b0 ) | ( ~n14568 & 1'b0 ) ;
  assign n14581 = ( n14315 & n14409 ) | ( n14315 & n14569 ) | ( n14409 & n14569 ) ;
  assign n14580 = n14315 | n14569 ;
  assign n14582 = ( n14579 & ~n14581 ) | ( n14579 & n14580 ) | ( ~n14581 & n14580 ) ;
  assign n14586 = n14078 &  n14408 ;
  assign n14587 = n14407 &  n14586 ;
  assign n14575 = x91 | n14078 ;
  assign n14576 = x91 &  n14078 ;
  assign n14577 = ( n14575 & ~n14576 ) | ( n14575 & 1'b0 ) | ( ~n14576 & 1'b0 ) ;
  assign n14589 = ( n14314 & n14409 ) | ( n14314 & n14577 ) | ( n14409 & n14577 ) ;
  assign n14588 = n14314 | n14577 ;
  assign n14590 = ( n14587 & ~n14589 ) | ( n14587 & n14588 ) | ( ~n14589 & n14588 ) ;
  assign n14594 = n14086 &  n14408 ;
  assign n14595 = n14407 &  n14594 ;
  assign n14583 = x90 | n14086 ;
  assign n14584 = x90 &  n14086 ;
  assign n14585 = ( n14583 & ~n14584 ) | ( n14583 & 1'b0 ) | ( ~n14584 & 1'b0 ) ;
  assign n14597 = ( n14313 & n14409 ) | ( n14313 & n14585 ) | ( n14409 & n14585 ) ;
  assign n14596 = n14313 | n14585 ;
  assign n14598 = ( n14595 & ~n14597 ) | ( n14595 & n14596 ) | ( ~n14597 & n14596 ) ;
  assign n14602 = n14094 &  n14408 ;
  assign n14603 = n14407 &  n14602 ;
  assign n14591 = x89 | n14094 ;
  assign n14592 = x89 &  n14094 ;
  assign n14593 = ( n14591 & ~n14592 ) | ( n14591 & 1'b0 ) | ( ~n14592 & 1'b0 ) ;
  assign n14605 = ( n14312 & n14409 ) | ( n14312 & n14593 ) | ( n14409 & n14593 ) ;
  assign n14604 = n14312 | n14593 ;
  assign n14606 = ( n14603 & ~n14605 ) | ( n14603 & n14604 ) | ( ~n14605 & n14604 ) ;
  assign n14610 = n14102 &  n14408 ;
  assign n14611 = n14407 &  n14610 ;
  assign n14599 = x88 | n14102 ;
  assign n14600 = x88 &  n14102 ;
  assign n14601 = ( n14599 & ~n14600 ) | ( n14599 & 1'b0 ) | ( ~n14600 & 1'b0 ) ;
  assign n14613 = ( n14311 & n14409 ) | ( n14311 & n14601 ) | ( n14409 & n14601 ) ;
  assign n14612 = n14311 | n14601 ;
  assign n14614 = ( n14611 & ~n14613 ) | ( n14611 & n14612 ) | ( ~n14613 & n14612 ) ;
  assign n14618 = n14110 &  n14408 ;
  assign n14619 = n14407 &  n14618 ;
  assign n14607 = x87 | n14110 ;
  assign n14608 = x87 &  n14110 ;
  assign n14609 = ( n14607 & ~n14608 ) | ( n14607 & 1'b0 ) | ( ~n14608 & 1'b0 ) ;
  assign n14621 = ( n14310 & n14409 ) | ( n14310 & n14609 ) | ( n14409 & n14609 ) ;
  assign n14620 = n14310 | n14609 ;
  assign n14622 = ( n14619 & ~n14621 ) | ( n14619 & n14620 ) | ( ~n14621 & n14620 ) ;
  assign n14626 = n14118 &  n14408 ;
  assign n14627 = n14407 &  n14626 ;
  assign n14615 = x86 | n14118 ;
  assign n14616 = x86 &  n14118 ;
  assign n14617 = ( n14615 & ~n14616 ) | ( n14615 & 1'b0 ) | ( ~n14616 & 1'b0 ) ;
  assign n14629 = ( n14309 & n14409 ) | ( n14309 & n14617 ) | ( n14409 & n14617 ) ;
  assign n14628 = n14309 | n14617 ;
  assign n14630 = ( n14627 & ~n14629 ) | ( n14627 & n14628 ) | ( ~n14629 & n14628 ) ;
  assign n14634 = n14126 &  n14408 ;
  assign n14635 = n14407 &  n14634 ;
  assign n14623 = x85 | n14126 ;
  assign n14624 = x85 &  n14126 ;
  assign n14625 = ( n14623 & ~n14624 ) | ( n14623 & 1'b0 ) | ( ~n14624 & 1'b0 ) ;
  assign n14637 = ( n14308 & n14409 ) | ( n14308 & n14625 ) | ( n14409 & n14625 ) ;
  assign n14636 = n14308 | n14625 ;
  assign n14638 = ( n14635 & ~n14637 ) | ( n14635 & n14636 ) | ( ~n14637 & n14636 ) ;
  assign n14642 = n14134 &  n14408 ;
  assign n14643 = n14407 &  n14642 ;
  assign n14631 = x84 | n14134 ;
  assign n14632 = x84 &  n14134 ;
  assign n14633 = ( n14631 & ~n14632 ) | ( n14631 & 1'b0 ) | ( ~n14632 & 1'b0 ) ;
  assign n14645 = ( n14307 & n14409 ) | ( n14307 & n14633 ) | ( n14409 & n14633 ) ;
  assign n14644 = n14307 | n14633 ;
  assign n14646 = ( n14643 & ~n14645 ) | ( n14643 & n14644 ) | ( ~n14645 & n14644 ) ;
  assign n14650 = n14142 &  n14408 ;
  assign n14651 = n14407 &  n14650 ;
  assign n14639 = x83 | n14142 ;
  assign n14640 = x83 &  n14142 ;
  assign n14641 = ( n14639 & ~n14640 ) | ( n14639 & 1'b0 ) | ( ~n14640 & 1'b0 ) ;
  assign n14653 = ( n14306 & n14409 ) | ( n14306 & n14641 ) | ( n14409 & n14641 ) ;
  assign n14652 = n14306 | n14641 ;
  assign n14654 = ( n14651 & ~n14653 ) | ( n14651 & n14652 ) | ( ~n14653 & n14652 ) ;
  assign n14658 = n14150 &  n14408 ;
  assign n14659 = n14407 &  n14658 ;
  assign n14647 = x82 | n14150 ;
  assign n14648 = x82 &  n14150 ;
  assign n14649 = ( n14647 & ~n14648 ) | ( n14647 & 1'b0 ) | ( ~n14648 & 1'b0 ) ;
  assign n14661 = ( n14305 & n14409 ) | ( n14305 & n14649 ) | ( n14409 & n14649 ) ;
  assign n14660 = n14305 | n14649 ;
  assign n14662 = ( n14659 & ~n14661 ) | ( n14659 & n14660 ) | ( ~n14661 & n14660 ) ;
  assign n14666 = n14158 &  n14408 ;
  assign n14667 = n14407 &  n14666 ;
  assign n14655 = x81 | n14158 ;
  assign n14656 = x81 &  n14158 ;
  assign n14657 = ( n14655 & ~n14656 ) | ( n14655 & 1'b0 ) | ( ~n14656 & 1'b0 ) ;
  assign n14669 = ( n14304 & n14409 ) | ( n14304 & n14657 ) | ( n14409 & n14657 ) ;
  assign n14668 = n14304 | n14657 ;
  assign n14670 = ( n14667 & ~n14669 ) | ( n14667 & n14668 ) | ( ~n14669 & n14668 ) ;
  assign n14674 = n14166 &  n14408 ;
  assign n14675 = n14407 &  n14674 ;
  assign n14663 = x80 | n14166 ;
  assign n14664 = x80 &  n14166 ;
  assign n14665 = ( n14663 & ~n14664 ) | ( n14663 & 1'b0 ) | ( ~n14664 & 1'b0 ) ;
  assign n14677 = ( n14303 & n14409 ) | ( n14303 & n14665 ) | ( n14409 & n14665 ) ;
  assign n14676 = n14303 | n14665 ;
  assign n14678 = ( n14675 & ~n14677 ) | ( n14675 & n14676 ) | ( ~n14677 & n14676 ) ;
  assign n14682 = n14174 &  n14408 ;
  assign n14683 = n14407 &  n14682 ;
  assign n14671 = x79 | n14174 ;
  assign n14672 = x79 &  n14174 ;
  assign n14673 = ( n14671 & ~n14672 ) | ( n14671 & 1'b0 ) | ( ~n14672 & 1'b0 ) ;
  assign n14685 = ( n14302 & n14409 ) | ( n14302 & n14673 ) | ( n14409 & n14673 ) ;
  assign n14684 = n14302 | n14673 ;
  assign n14686 = ( n14683 & ~n14685 ) | ( n14683 & n14684 ) | ( ~n14685 & n14684 ) ;
  assign n14690 = n14182 &  n14408 ;
  assign n14691 = n14407 &  n14690 ;
  assign n14679 = x78 | n14182 ;
  assign n14680 = x78 &  n14182 ;
  assign n14681 = ( n14679 & ~n14680 ) | ( n14679 & 1'b0 ) | ( ~n14680 & 1'b0 ) ;
  assign n14693 = ( n14301 & n14409 ) | ( n14301 & n14681 ) | ( n14409 & n14681 ) ;
  assign n14692 = n14301 | n14681 ;
  assign n14694 = ( n14691 & ~n14693 ) | ( n14691 & n14692 ) | ( ~n14693 & n14692 ) ;
  assign n14698 = n14190 &  n14408 ;
  assign n14699 = n14407 &  n14698 ;
  assign n14687 = x77 | n14190 ;
  assign n14688 = x77 &  n14190 ;
  assign n14689 = ( n14687 & ~n14688 ) | ( n14687 & 1'b0 ) | ( ~n14688 & 1'b0 ) ;
  assign n14701 = ( n14300 & n14409 ) | ( n14300 & n14689 ) | ( n14409 & n14689 ) ;
  assign n14700 = n14300 | n14689 ;
  assign n14702 = ( n14699 & ~n14701 ) | ( n14699 & n14700 ) | ( ~n14701 & n14700 ) ;
  assign n14706 = n14198 &  n14408 ;
  assign n14707 = n14407 &  n14706 ;
  assign n14695 = x76 | n14198 ;
  assign n14696 = x76 &  n14198 ;
  assign n14697 = ( n14695 & ~n14696 ) | ( n14695 & 1'b0 ) | ( ~n14696 & 1'b0 ) ;
  assign n14709 = ( n14299 & n14409 ) | ( n14299 & n14697 ) | ( n14409 & n14697 ) ;
  assign n14708 = n14299 | n14697 ;
  assign n14710 = ( n14707 & ~n14709 ) | ( n14707 & n14708 ) | ( ~n14709 & n14708 ) ;
  assign n14714 = n14206 &  n14408 ;
  assign n14715 = n14407 &  n14714 ;
  assign n14703 = x75 | n14206 ;
  assign n14704 = x75 &  n14206 ;
  assign n14705 = ( n14703 & ~n14704 ) | ( n14703 & 1'b0 ) | ( ~n14704 & 1'b0 ) ;
  assign n14717 = ( n14298 & n14409 ) | ( n14298 & n14705 ) | ( n14409 & n14705 ) ;
  assign n14716 = n14298 | n14705 ;
  assign n14718 = ( n14715 & ~n14717 ) | ( n14715 & n14716 ) | ( ~n14717 & n14716 ) ;
  assign n14722 = n14214 &  n14408 ;
  assign n14723 = n14407 &  n14722 ;
  assign n14711 = x74 | n14214 ;
  assign n14712 = x74 &  n14214 ;
  assign n14713 = ( n14711 & ~n14712 ) | ( n14711 & 1'b0 ) | ( ~n14712 & 1'b0 ) ;
  assign n14725 = ( n14297 & n14409 ) | ( n14297 & n14713 ) | ( n14409 & n14713 ) ;
  assign n14724 = n14297 | n14713 ;
  assign n14726 = ( n14723 & ~n14725 ) | ( n14723 & n14724 ) | ( ~n14725 & n14724 ) ;
  assign n14730 = n14222 &  n14408 ;
  assign n14731 = n14407 &  n14730 ;
  assign n14719 = x73 | n14222 ;
  assign n14720 = x73 &  n14222 ;
  assign n14721 = ( n14719 & ~n14720 ) | ( n14719 & 1'b0 ) | ( ~n14720 & 1'b0 ) ;
  assign n14733 = ( n14296 & n14409 ) | ( n14296 & n14721 ) | ( n14409 & n14721 ) ;
  assign n14732 = n14296 | n14721 ;
  assign n14734 = ( n14731 & ~n14733 ) | ( n14731 & n14732 ) | ( ~n14733 & n14732 ) ;
  assign n14738 = n14230 &  n14408 ;
  assign n14739 = n14407 &  n14738 ;
  assign n14727 = x72 | n14230 ;
  assign n14728 = x72 &  n14230 ;
  assign n14729 = ( n14727 & ~n14728 ) | ( n14727 & 1'b0 ) | ( ~n14728 & 1'b0 ) ;
  assign n14741 = ( n14295 & n14409 ) | ( n14295 & n14729 ) | ( n14409 & n14729 ) ;
  assign n14740 = n14295 | n14729 ;
  assign n14742 = ( n14739 & ~n14741 ) | ( n14739 & n14740 ) | ( ~n14741 & n14740 ) ;
  assign n14746 = n14238 &  n14408 ;
  assign n14747 = n14407 &  n14746 ;
  assign n14735 = x71 | n14238 ;
  assign n14736 = x71 &  n14238 ;
  assign n14737 = ( n14735 & ~n14736 ) | ( n14735 & 1'b0 ) | ( ~n14736 & 1'b0 ) ;
  assign n14749 = ( n14294 & n14409 ) | ( n14294 & n14737 ) | ( n14409 & n14737 ) ;
  assign n14748 = n14294 | n14737 ;
  assign n14750 = ( n14747 & ~n14749 ) | ( n14747 & n14748 ) | ( ~n14749 & n14748 ) ;
  assign n14754 = n14246 &  n14408 ;
  assign n14755 = n14407 &  n14754 ;
  assign n14743 = x70 | n14246 ;
  assign n14744 = x70 &  n14246 ;
  assign n14745 = ( n14743 & ~n14744 ) | ( n14743 & 1'b0 ) | ( ~n14744 & 1'b0 ) ;
  assign n14757 = ( n14293 & n14409 ) | ( n14293 & n14745 ) | ( n14409 & n14745 ) ;
  assign n14756 = n14293 | n14745 ;
  assign n14758 = ( n14755 & ~n14757 ) | ( n14755 & n14756 ) | ( ~n14757 & n14756 ) ;
  assign n14762 = n14254 &  n14408 ;
  assign n14763 = n14407 &  n14762 ;
  assign n14751 = x69 | n14254 ;
  assign n14752 = x69 &  n14254 ;
  assign n14753 = ( n14751 & ~n14752 ) | ( n14751 & 1'b0 ) | ( ~n14752 & 1'b0 ) ;
  assign n14765 = ( n14292 & n14409 ) | ( n14292 & n14753 ) | ( n14409 & n14753 ) ;
  assign n14764 = n14292 | n14753 ;
  assign n14766 = ( n14763 & ~n14765 ) | ( n14763 & n14764 ) | ( ~n14765 & n14764 ) ;
  assign n14770 = n14262 &  n14408 ;
  assign n14771 = n14407 &  n14770 ;
  assign n14759 = x68 | n14262 ;
  assign n14760 = x68 &  n14262 ;
  assign n14761 = ( n14759 & ~n14760 ) | ( n14759 & 1'b0 ) | ( ~n14760 & 1'b0 ) ;
  assign n14773 = ( n14291 & n14409 ) | ( n14291 & n14761 ) | ( n14409 & n14761 ) ;
  assign n14772 = n14291 | n14761 ;
  assign n14774 = ( n14771 & ~n14773 ) | ( n14771 & n14772 ) | ( ~n14773 & n14772 ) ;
  assign n14778 = n14271 &  n14408 ;
  assign n14779 = n14407 &  n14778 ;
  assign n14767 = x67 | n14271 ;
  assign n14768 = x67 &  n14271 ;
  assign n14769 = ( n14767 & ~n14768 ) | ( n14767 & 1'b0 ) | ( ~n14768 & 1'b0 ) ;
  assign n14781 = ( n14290 & n14409 ) | ( n14290 & n14769 ) | ( n14409 & n14769 ) ;
  assign n14780 = n14290 | n14769 ;
  assign n14782 = ( n14779 & ~n14781 ) | ( n14779 & n14780 ) | ( ~n14781 & n14780 ) ;
  assign n14783 = n14277 &  n14408 ;
  assign n14784 = n14407 &  n14783 ;
  assign n14775 = x66 | n14277 ;
  assign n14776 = x66 &  n14277 ;
  assign n14777 = ( n14775 & ~n14776 ) | ( n14775 & 1'b0 ) | ( ~n14776 & 1'b0 ) ;
  assign n14785 = n14289 &  n14777 ;
  assign n14786 = ( n14289 & ~n14409 ) | ( n14289 & n14777 ) | ( ~n14409 & n14777 ) ;
  assign n14787 = ( n14784 & ~n14785 ) | ( n14784 & n14786 ) | ( ~n14785 & n14786 ) ;
  assign n14788 = ( n14287 & ~x65 ) | ( n14287 & n14288 ) | ( ~x65 & n14288 ) ;
  assign n14789 = ( n14289 & ~n14288 ) | ( n14289 & n14788 ) | ( ~n14288 & n14788 ) ;
  assign n14790 = ~n14409 & n14789 ;
  assign n14791 = n14287 &  n14408 ;
  assign n14792 = n14407 &  n14791 ;
  assign n14793 = n14790 | n14792 ;
  assign n14794 = ( x64 & ~n14409 ) | ( x64 & 1'b0 ) | ( ~n14409 & 1'b0 ) ;
  assign n14795 = ( x8 & ~n14794 ) | ( x8 & 1'b0 ) | ( ~n14794 & 1'b0 ) ;
  assign n14796 = ( n14288 & ~n14409 ) | ( n14288 & 1'b0 ) | ( ~n14409 & 1'b0 ) ;
  assign n14797 = n14795 | n14796 ;
  assign n14798 = ~x7 & x64 ;
  assign n14799 = ( x65 & ~n14797 ) | ( x65 & n14798 ) | ( ~n14797 & n14798 ) ;
  assign n14800 = ( x66 & ~n14793 ) | ( x66 & n14799 ) | ( ~n14793 & n14799 ) ;
  assign n14801 = ( x67 & ~n14787 ) | ( x67 & n14800 ) | ( ~n14787 & n14800 ) ;
  assign n14802 = ( x68 & ~n14782 ) | ( x68 & n14801 ) | ( ~n14782 & n14801 ) ;
  assign n14803 = ( x69 & ~n14774 ) | ( x69 & n14802 ) | ( ~n14774 & n14802 ) ;
  assign n14804 = ( x70 & ~n14766 ) | ( x70 & n14803 ) | ( ~n14766 & n14803 ) ;
  assign n14805 = ( x71 & ~n14758 ) | ( x71 & n14804 ) | ( ~n14758 & n14804 ) ;
  assign n14806 = ( x72 & ~n14750 ) | ( x72 & n14805 ) | ( ~n14750 & n14805 ) ;
  assign n14807 = ( x73 & ~n14742 ) | ( x73 & n14806 ) | ( ~n14742 & n14806 ) ;
  assign n14808 = ( x74 & ~n14734 ) | ( x74 & n14807 ) | ( ~n14734 & n14807 ) ;
  assign n14809 = ( x75 & ~n14726 ) | ( x75 & n14808 ) | ( ~n14726 & n14808 ) ;
  assign n14810 = ( x76 & ~n14718 ) | ( x76 & n14809 ) | ( ~n14718 & n14809 ) ;
  assign n14811 = ( x77 & ~n14710 ) | ( x77 & n14810 ) | ( ~n14710 & n14810 ) ;
  assign n14812 = ( x78 & ~n14702 ) | ( x78 & n14811 ) | ( ~n14702 & n14811 ) ;
  assign n14813 = ( x79 & ~n14694 ) | ( x79 & n14812 ) | ( ~n14694 & n14812 ) ;
  assign n14814 = ( x80 & ~n14686 ) | ( x80 & n14813 ) | ( ~n14686 & n14813 ) ;
  assign n14815 = ( x81 & ~n14678 ) | ( x81 & n14814 ) | ( ~n14678 & n14814 ) ;
  assign n14816 = ( x82 & ~n14670 ) | ( x82 & n14815 ) | ( ~n14670 & n14815 ) ;
  assign n14817 = ( x83 & ~n14662 ) | ( x83 & n14816 ) | ( ~n14662 & n14816 ) ;
  assign n14818 = ( x84 & ~n14654 ) | ( x84 & n14817 ) | ( ~n14654 & n14817 ) ;
  assign n14819 = ( x85 & ~n14646 ) | ( x85 & n14818 ) | ( ~n14646 & n14818 ) ;
  assign n14820 = ( x86 & ~n14638 ) | ( x86 & n14819 ) | ( ~n14638 & n14819 ) ;
  assign n14821 = ( x87 & ~n14630 ) | ( x87 & n14820 ) | ( ~n14630 & n14820 ) ;
  assign n14822 = ( x88 & ~n14622 ) | ( x88 & n14821 ) | ( ~n14622 & n14821 ) ;
  assign n14823 = ( x89 & ~n14614 ) | ( x89 & n14822 ) | ( ~n14614 & n14822 ) ;
  assign n14824 = ( x90 & ~n14606 ) | ( x90 & n14823 ) | ( ~n14606 & n14823 ) ;
  assign n14825 = ( x91 & ~n14598 ) | ( x91 & n14824 ) | ( ~n14598 & n14824 ) ;
  assign n14826 = ( x92 & ~n14590 ) | ( x92 & n14825 ) | ( ~n14590 & n14825 ) ;
  assign n14827 = ( x93 & ~n14582 ) | ( x93 & n14826 ) | ( ~n14582 & n14826 ) ;
  assign n14828 = ( x94 & ~n14574 ) | ( x94 & n14827 ) | ( ~n14574 & n14827 ) ;
  assign n14829 = ( x95 & ~n14566 ) | ( x95 & n14828 ) | ( ~n14566 & n14828 ) ;
  assign n14830 = ( x96 & ~n14558 ) | ( x96 & n14829 ) | ( ~n14558 & n14829 ) ;
  assign n14831 = ( x97 & ~n14550 ) | ( x97 & n14830 ) | ( ~n14550 & n14830 ) ;
  assign n14832 = ( x98 & ~n14542 ) | ( x98 & n14831 ) | ( ~n14542 & n14831 ) ;
  assign n14833 = ( x99 & ~n14534 ) | ( x99 & n14832 ) | ( ~n14534 & n14832 ) ;
  assign n14834 = ( x100 & ~n14526 ) | ( x100 & n14833 ) | ( ~n14526 & n14833 ) ;
  assign n14835 = ( x101 & ~n14518 ) | ( x101 & n14834 ) | ( ~n14518 & n14834 ) ;
  assign n14836 = ( x102 & ~n14510 ) | ( x102 & n14835 ) | ( ~n14510 & n14835 ) ;
  assign n14837 = ( x103 & ~n14502 ) | ( x103 & n14836 ) | ( ~n14502 & n14836 ) ;
  assign n14838 = ( x104 & ~n14494 ) | ( x104 & n14837 ) | ( ~n14494 & n14837 ) ;
  assign n14839 = ( x105 & ~n14486 ) | ( x105 & n14838 ) | ( ~n14486 & n14838 ) ;
  assign n14840 = ( x106 & ~n14478 ) | ( x106 & n14839 ) | ( ~n14478 & n14839 ) ;
  assign n14841 = ( x107 & ~n14470 ) | ( x107 & n14840 ) | ( ~n14470 & n14840 ) ;
  assign n14842 = ( x108 & ~n14462 ) | ( x108 & n14841 ) | ( ~n14462 & n14841 ) ;
  assign n14843 = ( x109 & ~n14454 ) | ( x109 & n14842 ) | ( ~n14454 & n14842 ) ;
  assign n14844 = ( x110 & ~n14446 ) | ( x110 & n14843 ) | ( ~n14446 & n14843 ) ;
  assign n14845 = ( x111 & ~n14438 ) | ( x111 & n14844 ) | ( ~n14438 & n14844 ) ;
  assign n14846 = ( x112 & ~n14430 ) | ( x112 & n14845 ) | ( ~n14430 & n14845 ) ;
  assign n14847 = ( x113 & ~n14422 ) | ( x113 & n14846 ) | ( ~n14422 & n14846 ) ;
  assign n14851 = ( x114 & ~n14414 ) | ( x114 & n14847 ) | ( ~n14414 & n14847 ) ;
  assign n14895 = ( x115 & ~n14859 ) | ( x115 & n14851 ) | ( ~n14859 & n14851 ) ;
  assign n14896 = ( x116 & ~n14894 ) | ( x116 & n14895 ) | ( ~n14894 & n14895 ) ;
  assign n14897 = ( x117 & ~n14889 ) | ( x117 & n14896 ) | ( ~n14889 & n14896 ) ;
  assign n14898 = ( x118 & ~n14881 ) | ( x118 & n14897 ) | ( ~n14881 & n14897 ) ;
  assign n14899 = ( x119 & ~n14873 ) | ( x119 & n14898 ) | ( ~n14873 & n14898 ) ;
  assign n14900 = n14402 | n14404 ;
  assign n14901 = ( n14396 & ~n14900 ) | ( n14396 & 1'b0 ) | ( ~n14900 & 1'b0 ) ;
  assign n14902 = ~n14396 & n14900 ;
  assign n14903 = ( n14901 & ~n14409 ) | ( n14901 & n14902 ) | ( ~n14409 & n14902 ) ;
  assign n14904 = n13437 &  n13898 ;
  assign n14905 = n14407 &  n14904 ;
  assign n14906 = n14903 | n14905 ;
  assign n14907 = ~x120 & n14906 ;
  assign n14908 = ( x120 & ~n14905 ) | ( x120 & 1'b0 ) | ( ~n14905 & 1'b0 ) ;
  assign n14909 = ~n14903 & n14908 ;
  assign n14910 = n239 | n14909 ;
  assign n14911 = n14907 | n14910 ;
  assign n14912 = n14899 | n14911 ;
  assign n14913 = ~n14906 |  n269 ;
  assign n14932 = n14873 &  n14913 ;
  assign n14933 = n14912 &  n14932 ;
  assign n14920 = x119 | n14873 ;
  assign n14921 = x119 &  n14873 ;
  assign n14922 = ( n14920 & ~n14921 ) | ( n14920 & 1'b0 ) | ( ~n14921 & 1'b0 ) ;
  assign n14934 = n14898 &  n14922 ;
  assign n14914 = n14912 &  n14913 ;
  assign n14935 = ( n14898 & ~n14914 ) | ( n14898 & n14922 ) | ( ~n14914 & n14922 ) ;
  assign n14936 = ( n14933 & ~n14934 ) | ( n14933 & n14935 ) | ( ~n14934 & n14935 ) ;
  assign n14924 = n269 &  n14906 ;
  assign n14925 = n14912 &  n14924 ;
  assign n14923 = n14907 | n14909 ;
  assign n14927 = ( n14899 & n14914 ) | ( n14899 & n14923 ) | ( n14914 & n14923 ) ;
  assign n14926 = n14899 | n14923 ;
  assign n14928 = ( n14925 & ~n14927 ) | ( n14925 & n14926 ) | ( ~n14927 & n14926 ) ;
  assign n14940 = n14881 &  n14913 ;
  assign n14941 = n14912 &  n14940 ;
  assign n14929 = x118 | n14881 ;
  assign n14930 = x118 &  n14881 ;
  assign n14931 = ( n14929 & ~n14930 ) | ( n14929 & 1'b0 ) | ( ~n14930 & 1'b0 ) ;
  assign n14942 = n14897 &  n14931 ;
  assign n14943 = ( n14897 & ~n14914 ) | ( n14897 & n14931 ) | ( ~n14914 & n14931 ) ;
  assign n14944 = ( n14941 & ~n14942 ) | ( n14941 & n14943 ) | ( ~n14942 & n14943 ) ;
  assign n14948 = n14889 &  n14913 ;
  assign n14949 = n14912 &  n14948 ;
  assign n14937 = x117 | n14889 ;
  assign n14938 = x117 &  n14889 ;
  assign n14939 = ( n14937 & ~n14938 ) | ( n14937 & 1'b0 ) | ( ~n14938 & 1'b0 ) ;
  assign n14950 = n14896 &  n14939 ;
  assign n14951 = ( n14896 & ~n14914 ) | ( n14896 & n14939 ) | ( ~n14914 & n14939 ) ;
  assign n14952 = ( n14949 & ~n14950 ) | ( n14949 & n14951 ) | ( ~n14950 & n14951 ) ;
  assign n14953 = n14894 &  n14913 ;
  assign n14954 = n14912 &  n14953 ;
  assign n14945 = x116 | n14894 ;
  assign n14946 = x116 &  n14894 ;
  assign n14947 = ( n14945 & ~n14946 ) | ( n14945 & 1'b0 ) | ( ~n14946 & 1'b0 ) ;
  assign n14955 = n14895 &  n14947 ;
  assign n14956 = ( n14895 & ~n14914 ) | ( n14895 & n14947 ) | ( ~n14914 & n14947 ) ;
  assign n14957 = ( n14954 & ~n14955 ) | ( n14954 & n14956 ) | ( ~n14955 & n14956 ) ;
  assign n14915 = n14859 &  n14913 ;
  assign n14916 = n14912 &  n14915 ;
  assign n14860 = x115 | n14859 ;
  assign n14861 = x115 &  n14859 ;
  assign n14862 = ( n14860 & ~n14861 ) | ( n14860 & 1'b0 ) | ( ~n14861 & 1'b0 ) ;
  assign n14917 = n14851 &  n14862 ;
  assign n14918 = ( n14851 & ~n14914 ) | ( n14851 & n14862 ) | ( ~n14914 & n14862 ) ;
  assign n14919 = ( n14916 & ~n14917 ) | ( n14916 & n14918 ) | ( ~n14917 & n14918 ) ;
  assign n14961 = n14414 &  n14913 ;
  assign n14962 = n14912 &  n14961 ;
  assign n14848 = x114 | n14414 ;
  assign n14849 = x114 &  n14414 ;
  assign n14850 = ( n14848 & ~n14849 ) | ( n14848 & 1'b0 ) | ( ~n14849 & 1'b0 ) ;
  assign n14963 = n14847 &  n14850 ;
  assign n14964 = ( n14847 & ~n14914 ) | ( n14847 & n14850 ) | ( ~n14914 & n14850 ) ;
  assign n14965 = ( n14962 & ~n14963 ) | ( n14962 & n14964 ) | ( ~n14963 & n14964 ) ;
  assign n14969 = n14422 &  n14913 ;
  assign n14970 = n14912 &  n14969 ;
  assign n14958 = x113 | n14422 ;
  assign n14959 = x113 &  n14422 ;
  assign n14960 = ( n14958 & ~n14959 ) | ( n14958 & 1'b0 ) | ( ~n14959 & 1'b0 ) ;
  assign n14972 = ( n14846 & n14914 ) | ( n14846 & n14960 ) | ( n14914 & n14960 ) ;
  assign n14971 = n14846 | n14960 ;
  assign n14973 = ( n14970 & ~n14972 ) | ( n14970 & n14971 ) | ( ~n14972 & n14971 ) ;
  assign n14977 = n14430 &  n14913 ;
  assign n14978 = n14912 &  n14977 ;
  assign n14966 = x112 | n14430 ;
  assign n14967 = x112 &  n14430 ;
  assign n14968 = ( n14966 & ~n14967 ) | ( n14966 & 1'b0 ) | ( ~n14967 & 1'b0 ) ;
  assign n14980 = ( n14845 & n14914 ) | ( n14845 & n14968 ) | ( n14914 & n14968 ) ;
  assign n14979 = n14845 | n14968 ;
  assign n14981 = ( n14978 & ~n14980 ) | ( n14978 & n14979 ) | ( ~n14980 & n14979 ) ;
  assign n14985 = n14438 &  n14913 ;
  assign n14986 = n14912 &  n14985 ;
  assign n14974 = x111 | n14438 ;
  assign n14975 = x111 &  n14438 ;
  assign n14976 = ( n14974 & ~n14975 ) | ( n14974 & 1'b0 ) | ( ~n14975 & 1'b0 ) ;
  assign n14988 = ( n14844 & n14914 ) | ( n14844 & n14976 ) | ( n14914 & n14976 ) ;
  assign n14987 = n14844 | n14976 ;
  assign n14989 = ( n14986 & ~n14988 ) | ( n14986 & n14987 ) | ( ~n14988 & n14987 ) ;
  assign n14993 = n14446 &  n14913 ;
  assign n14994 = n14912 &  n14993 ;
  assign n14982 = x110 | n14446 ;
  assign n14983 = x110 &  n14446 ;
  assign n14984 = ( n14982 & ~n14983 ) | ( n14982 & 1'b0 ) | ( ~n14983 & 1'b0 ) ;
  assign n14996 = ( n14843 & n14914 ) | ( n14843 & n14984 ) | ( n14914 & n14984 ) ;
  assign n14995 = n14843 | n14984 ;
  assign n14997 = ( n14994 & ~n14996 ) | ( n14994 & n14995 ) | ( ~n14996 & n14995 ) ;
  assign n15001 = n14454 &  n14913 ;
  assign n15002 = n14912 &  n15001 ;
  assign n14990 = x109 | n14454 ;
  assign n14991 = x109 &  n14454 ;
  assign n14992 = ( n14990 & ~n14991 ) | ( n14990 & 1'b0 ) | ( ~n14991 & 1'b0 ) ;
  assign n15004 = ( n14842 & n14914 ) | ( n14842 & n14992 ) | ( n14914 & n14992 ) ;
  assign n15003 = n14842 | n14992 ;
  assign n15005 = ( n15002 & ~n15004 ) | ( n15002 & n15003 ) | ( ~n15004 & n15003 ) ;
  assign n15009 = n14462 &  n14913 ;
  assign n15010 = n14912 &  n15009 ;
  assign n14998 = x108 | n14462 ;
  assign n14999 = x108 &  n14462 ;
  assign n15000 = ( n14998 & ~n14999 ) | ( n14998 & 1'b0 ) | ( ~n14999 & 1'b0 ) ;
  assign n15012 = ( n14841 & n14914 ) | ( n14841 & n15000 ) | ( n14914 & n15000 ) ;
  assign n15011 = n14841 | n15000 ;
  assign n15013 = ( n15010 & ~n15012 ) | ( n15010 & n15011 ) | ( ~n15012 & n15011 ) ;
  assign n15017 = n14470 &  n14913 ;
  assign n15018 = n14912 &  n15017 ;
  assign n15006 = x107 | n14470 ;
  assign n15007 = x107 &  n14470 ;
  assign n15008 = ( n15006 & ~n15007 ) | ( n15006 & 1'b0 ) | ( ~n15007 & 1'b0 ) ;
  assign n15020 = ( n14840 & n14914 ) | ( n14840 & n15008 ) | ( n14914 & n15008 ) ;
  assign n15019 = n14840 | n15008 ;
  assign n15021 = ( n15018 & ~n15020 ) | ( n15018 & n15019 ) | ( ~n15020 & n15019 ) ;
  assign n15025 = n14478 &  n14913 ;
  assign n15026 = n14912 &  n15025 ;
  assign n15014 = x106 | n14478 ;
  assign n15015 = x106 &  n14478 ;
  assign n15016 = ( n15014 & ~n15015 ) | ( n15014 & 1'b0 ) | ( ~n15015 & 1'b0 ) ;
  assign n15028 = ( n14839 & n14914 ) | ( n14839 & n15016 ) | ( n14914 & n15016 ) ;
  assign n15027 = n14839 | n15016 ;
  assign n15029 = ( n15026 & ~n15028 ) | ( n15026 & n15027 ) | ( ~n15028 & n15027 ) ;
  assign n15033 = n14486 &  n14913 ;
  assign n15034 = n14912 &  n15033 ;
  assign n15022 = x105 | n14486 ;
  assign n15023 = x105 &  n14486 ;
  assign n15024 = ( n15022 & ~n15023 ) | ( n15022 & 1'b0 ) | ( ~n15023 & 1'b0 ) ;
  assign n15036 = ( n14838 & n14914 ) | ( n14838 & n15024 ) | ( n14914 & n15024 ) ;
  assign n15035 = n14838 | n15024 ;
  assign n15037 = ( n15034 & ~n15036 ) | ( n15034 & n15035 ) | ( ~n15036 & n15035 ) ;
  assign n15041 = n14494 &  n14913 ;
  assign n15042 = n14912 &  n15041 ;
  assign n15030 = x104 | n14494 ;
  assign n15031 = x104 &  n14494 ;
  assign n15032 = ( n15030 & ~n15031 ) | ( n15030 & 1'b0 ) | ( ~n15031 & 1'b0 ) ;
  assign n15044 = ( n14837 & n14914 ) | ( n14837 & n15032 ) | ( n14914 & n15032 ) ;
  assign n15043 = n14837 | n15032 ;
  assign n15045 = ( n15042 & ~n15044 ) | ( n15042 & n15043 ) | ( ~n15044 & n15043 ) ;
  assign n15049 = n14502 &  n14913 ;
  assign n15050 = n14912 &  n15049 ;
  assign n15038 = x103 | n14502 ;
  assign n15039 = x103 &  n14502 ;
  assign n15040 = ( n15038 & ~n15039 ) | ( n15038 & 1'b0 ) | ( ~n15039 & 1'b0 ) ;
  assign n15052 = ( n14836 & n14914 ) | ( n14836 & n15040 ) | ( n14914 & n15040 ) ;
  assign n15051 = n14836 | n15040 ;
  assign n15053 = ( n15050 & ~n15052 ) | ( n15050 & n15051 ) | ( ~n15052 & n15051 ) ;
  assign n15057 = n14510 &  n14913 ;
  assign n15058 = n14912 &  n15057 ;
  assign n15046 = x102 | n14510 ;
  assign n15047 = x102 &  n14510 ;
  assign n15048 = ( n15046 & ~n15047 ) | ( n15046 & 1'b0 ) | ( ~n15047 & 1'b0 ) ;
  assign n15060 = ( n14835 & n14914 ) | ( n14835 & n15048 ) | ( n14914 & n15048 ) ;
  assign n15059 = n14835 | n15048 ;
  assign n15061 = ( n15058 & ~n15060 ) | ( n15058 & n15059 ) | ( ~n15060 & n15059 ) ;
  assign n15065 = n14518 &  n14913 ;
  assign n15066 = n14912 &  n15065 ;
  assign n15054 = x101 | n14518 ;
  assign n15055 = x101 &  n14518 ;
  assign n15056 = ( n15054 & ~n15055 ) | ( n15054 & 1'b0 ) | ( ~n15055 & 1'b0 ) ;
  assign n15068 = ( n14834 & n14914 ) | ( n14834 & n15056 ) | ( n14914 & n15056 ) ;
  assign n15067 = n14834 | n15056 ;
  assign n15069 = ( n15066 & ~n15068 ) | ( n15066 & n15067 ) | ( ~n15068 & n15067 ) ;
  assign n15073 = n14526 &  n14913 ;
  assign n15074 = n14912 &  n15073 ;
  assign n15062 = x100 | n14526 ;
  assign n15063 = x100 &  n14526 ;
  assign n15064 = ( n15062 & ~n15063 ) | ( n15062 & 1'b0 ) | ( ~n15063 & 1'b0 ) ;
  assign n15076 = ( n14833 & n14914 ) | ( n14833 & n15064 ) | ( n14914 & n15064 ) ;
  assign n15075 = n14833 | n15064 ;
  assign n15077 = ( n15074 & ~n15076 ) | ( n15074 & n15075 ) | ( ~n15076 & n15075 ) ;
  assign n15081 = n14534 &  n14913 ;
  assign n15082 = n14912 &  n15081 ;
  assign n15070 = x99 | n14534 ;
  assign n15071 = x99 &  n14534 ;
  assign n15072 = ( n15070 & ~n15071 ) | ( n15070 & 1'b0 ) | ( ~n15071 & 1'b0 ) ;
  assign n15084 = ( n14832 & n14914 ) | ( n14832 & n15072 ) | ( n14914 & n15072 ) ;
  assign n15083 = n14832 | n15072 ;
  assign n15085 = ( n15082 & ~n15084 ) | ( n15082 & n15083 ) | ( ~n15084 & n15083 ) ;
  assign n15089 = n14542 &  n14913 ;
  assign n15090 = n14912 &  n15089 ;
  assign n15078 = x98 | n14542 ;
  assign n15079 = x98 &  n14542 ;
  assign n15080 = ( n15078 & ~n15079 ) | ( n15078 & 1'b0 ) | ( ~n15079 & 1'b0 ) ;
  assign n15092 = ( n14831 & n14914 ) | ( n14831 & n15080 ) | ( n14914 & n15080 ) ;
  assign n15091 = n14831 | n15080 ;
  assign n15093 = ( n15090 & ~n15092 ) | ( n15090 & n15091 ) | ( ~n15092 & n15091 ) ;
  assign n15097 = n14550 &  n14913 ;
  assign n15098 = n14912 &  n15097 ;
  assign n15086 = x97 | n14550 ;
  assign n15087 = x97 &  n14550 ;
  assign n15088 = ( n15086 & ~n15087 ) | ( n15086 & 1'b0 ) | ( ~n15087 & 1'b0 ) ;
  assign n15100 = ( n14830 & n14914 ) | ( n14830 & n15088 ) | ( n14914 & n15088 ) ;
  assign n15099 = n14830 | n15088 ;
  assign n15101 = ( n15098 & ~n15100 ) | ( n15098 & n15099 ) | ( ~n15100 & n15099 ) ;
  assign n15105 = n14558 &  n14913 ;
  assign n15106 = n14912 &  n15105 ;
  assign n15094 = x96 | n14558 ;
  assign n15095 = x96 &  n14558 ;
  assign n15096 = ( n15094 & ~n15095 ) | ( n15094 & 1'b0 ) | ( ~n15095 & 1'b0 ) ;
  assign n15108 = ( n14829 & n14914 ) | ( n14829 & n15096 ) | ( n14914 & n15096 ) ;
  assign n15107 = n14829 | n15096 ;
  assign n15109 = ( n15106 & ~n15108 ) | ( n15106 & n15107 ) | ( ~n15108 & n15107 ) ;
  assign n15113 = n14566 &  n14913 ;
  assign n15114 = n14912 &  n15113 ;
  assign n15102 = x95 | n14566 ;
  assign n15103 = x95 &  n14566 ;
  assign n15104 = ( n15102 & ~n15103 ) | ( n15102 & 1'b0 ) | ( ~n15103 & 1'b0 ) ;
  assign n15116 = ( n14828 & n14914 ) | ( n14828 & n15104 ) | ( n14914 & n15104 ) ;
  assign n15115 = n14828 | n15104 ;
  assign n15117 = ( n15114 & ~n15116 ) | ( n15114 & n15115 ) | ( ~n15116 & n15115 ) ;
  assign n15121 = n14574 &  n14913 ;
  assign n15122 = n14912 &  n15121 ;
  assign n15110 = x94 | n14574 ;
  assign n15111 = x94 &  n14574 ;
  assign n15112 = ( n15110 & ~n15111 ) | ( n15110 & 1'b0 ) | ( ~n15111 & 1'b0 ) ;
  assign n15124 = ( n14827 & n14914 ) | ( n14827 & n15112 ) | ( n14914 & n15112 ) ;
  assign n15123 = n14827 | n15112 ;
  assign n15125 = ( n15122 & ~n15124 ) | ( n15122 & n15123 ) | ( ~n15124 & n15123 ) ;
  assign n15129 = n14582 &  n14913 ;
  assign n15130 = n14912 &  n15129 ;
  assign n15118 = x93 | n14582 ;
  assign n15119 = x93 &  n14582 ;
  assign n15120 = ( n15118 & ~n15119 ) | ( n15118 & 1'b0 ) | ( ~n15119 & 1'b0 ) ;
  assign n15132 = ( n14826 & n14914 ) | ( n14826 & n15120 ) | ( n14914 & n15120 ) ;
  assign n15131 = n14826 | n15120 ;
  assign n15133 = ( n15130 & ~n15132 ) | ( n15130 & n15131 ) | ( ~n15132 & n15131 ) ;
  assign n15137 = n14590 &  n14913 ;
  assign n15138 = n14912 &  n15137 ;
  assign n15126 = x92 | n14590 ;
  assign n15127 = x92 &  n14590 ;
  assign n15128 = ( n15126 & ~n15127 ) | ( n15126 & 1'b0 ) | ( ~n15127 & 1'b0 ) ;
  assign n15140 = ( n14825 & n14914 ) | ( n14825 & n15128 ) | ( n14914 & n15128 ) ;
  assign n15139 = n14825 | n15128 ;
  assign n15141 = ( n15138 & ~n15140 ) | ( n15138 & n15139 ) | ( ~n15140 & n15139 ) ;
  assign n15145 = n14598 &  n14913 ;
  assign n15146 = n14912 &  n15145 ;
  assign n15134 = x91 | n14598 ;
  assign n15135 = x91 &  n14598 ;
  assign n15136 = ( n15134 & ~n15135 ) | ( n15134 & 1'b0 ) | ( ~n15135 & 1'b0 ) ;
  assign n15148 = ( n14824 & n14914 ) | ( n14824 & n15136 ) | ( n14914 & n15136 ) ;
  assign n15147 = n14824 | n15136 ;
  assign n15149 = ( n15146 & ~n15148 ) | ( n15146 & n15147 ) | ( ~n15148 & n15147 ) ;
  assign n15153 = n14606 &  n14913 ;
  assign n15154 = n14912 &  n15153 ;
  assign n15142 = x90 | n14606 ;
  assign n15143 = x90 &  n14606 ;
  assign n15144 = ( n15142 & ~n15143 ) | ( n15142 & 1'b0 ) | ( ~n15143 & 1'b0 ) ;
  assign n15156 = ( n14823 & n14914 ) | ( n14823 & n15144 ) | ( n14914 & n15144 ) ;
  assign n15155 = n14823 | n15144 ;
  assign n15157 = ( n15154 & ~n15156 ) | ( n15154 & n15155 ) | ( ~n15156 & n15155 ) ;
  assign n15161 = n14614 &  n14913 ;
  assign n15162 = n14912 &  n15161 ;
  assign n15150 = x89 | n14614 ;
  assign n15151 = x89 &  n14614 ;
  assign n15152 = ( n15150 & ~n15151 ) | ( n15150 & 1'b0 ) | ( ~n15151 & 1'b0 ) ;
  assign n15164 = ( n14822 & n14914 ) | ( n14822 & n15152 ) | ( n14914 & n15152 ) ;
  assign n15163 = n14822 | n15152 ;
  assign n15165 = ( n15162 & ~n15164 ) | ( n15162 & n15163 ) | ( ~n15164 & n15163 ) ;
  assign n15169 = n14622 &  n14913 ;
  assign n15170 = n14912 &  n15169 ;
  assign n15158 = x88 | n14622 ;
  assign n15159 = x88 &  n14622 ;
  assign n15160 = ( n15158 & ~n15159 ) | ( n15158 & 1'b0 ) | ( ~n15159 & 1'b0 ) ;
  assign n15172 = ( n14821 & n14914 ) | ( n14821 & n15160 ) | ( n14914 & n15160 ) ;
  assign n15171 = n14821 | n15160 ;
  assign n15173 = ( n15170 & ~n15172 ) | ( n15170 & n15171 ) | ( ~n15172 & n15171 ) ;
  assign n15177 = n14630 &  n14913 ;
  assign n15178 = n14912 &  n15177 ;
  assign n15166 = x87 | n14630 ;
  assign n15167 = x87 &  n14630 ;
  assign n15168 = ( n15166 & ~n15167 ) | ( n15166 & 1'b0 ) | ( ~n15167 & 1'b0 ) ;
  assign n15180 = ( n14820 & n14914 ) | ( n14820 & n15168 ) | ( n14914 & n15168 ) ;
  assign n15179 = n14820 | n15168 ;
  assign n15181 = ( n15178 & ~n15180 ) | ( n15178 & n15179 ) | ( ~n15180 & n15179 ) ;
  assign n15185 = n14638 &  n14913 ;
  assign n15186 = n14912 &  n15185 ;
  assign n15174 = x86 | n14638 ;
  assign n15175 = x86 &  n14638 ;
  assign n15176 = ( n15174 & ~n15175 ) | ( n15174 & 1'b0 ) | ( ~n15175 & 1'b0 ) ;
  assign n15188 = ( n14819 & n14914 ) | ( n14819 & n15176 ) | ( n14914 & n15176 ) ;
  assign n15187 = n14819 | n15176 ;
  assign n15189 = ( n15186 & ~n15188 ) | ( n15186 & n15187 ) | ( ~n15188 & n15187 ) ;
  assign n15193 = n14646 &  n14913 ;
  assign n15194 = n14912 &  n15193 ;
  assign n15182 = x85 | n14646 ;
  assign n15183 = x85 &  n14646 ;
  assign n15184 = ( n15182 & ~n15183 ) | ( n15182 & 1'b0 ) | ( ~n15183 & 1'b0 ) ;
  assign n15196 = ( n14818 & n14914 ) | ( n14818 & n15184 ) | ( n14914 & n15184 ) ;
  assign n15195 = n14818 | n15184 ;
  assign n15197 = ( n15194 & ~n15196 ) | ( n15194 & n15195 ) | ( ~n15196 & n15195 ) ;
  assign n15201 = n14654 &  n14913 ;
  assign n15202 = n14912 &  n15201 ;
  assign n15190 = x84 | n14654 ;
  assign n15191 = x84 &  n14654 ;
  assign n15192 = ( n15190 & ~n15191 ) | ( n15190 & 1'b0 ) | ( ~n15191 & 1'b0 ) ;
  assign n15204 = ( n14817 & n14914 ) | ( n14817 & n15192 ) | ( n14914 & n15192 ) ;
  assign n15203 = n14817 | n15192 ;
  assign n15205 = ( n15202 & ~n15204 ) | ( n15202 & n15203 ) | ( ~n15204 & n15203 ) ;
  assign n15209 = n14662 &  n14913 ;
  assign n15210 = n14912 &  n15209 ;
  assign n15198 = x83 | n14662 ;
  assign n15199 = x83 &  n14662 ;
  assign n15200 = ( n15198 & ~n15199 ) | ( n15198 & 1'b0 ) | ( ~n15199 & 1'b0 ) ;
  assign n15212 = ( n14816 & n14914 ) | ( n14816 & n15200 ) | ( n14914 & n15200 ) ;
  assign n15211 = n14816 | n15200 ;
  assign n15213 = ( n15210 & ~n15212 ) | ( n15210 & n15211 ) | ( ~n15212 & n15211 ) ;
  assign n15217 = n14670 &  n14913 ;
  assign n15218 = n14912 &  n15217 ;
  assign n15206 = x82 | n14670 ;
  assign n15207 = x82 &  n14670 ;
  assign n15208 = ( n15206 & ~n15207 ) | ( n15206 & 1'b0 ) | ( ~n15207 & 1'b0 ) ;
  assign n15220 = ( n14815 & n14914 ) | ( n14815 & n15208 ) | ( n14914 & n15208 ) ;
  assign n15219 = n14815 | n15208 ;
  assign n15221 = ( n15218 & ~n15220 ) | ( n15218 & n15219 ) | ( ~n15220 & n15219 ) ;
  assign n15225 = n14678 &  n14913 ;
  assign n15226 = n14912 &  n15225 ;
  assign n15214 = x81 | n14678 ;
  assign n15215 = x81 &  n14678 ;
  assign n15216 = ( n15214 & ~n15215 ) | ( n15214 & 1'b0 ) | ( ~n15215 & 1'b0 ) ;
  assign n15228 = ( n14814 & n14914 ) | ( n14814 & n15216 ) | ( n14914 & n15216 ) ;
  assign n15227 = n14814 | n15216 ;
  assign n15229 = ( n15226 & ~n15228 ) | ( n15226 & n15227 ) | ( ~n15228 & n15227 ) ;
  assign n15233 = n14686 &  n14913 ;
  assign n15234 = n14912 &  n15233 ;
  assign n15222 = x80 | n14686 ;
  assign n15223 = x80 &  n14686 ;
  assign n15224 = ( n15222 & ~n15223 ) | ( n15222 & 1'b0 ) | ( ~n15223 & 1'b0 ) ;
  assign n15236 = ( n14813 & n14914 ) | ( n14813 & n15224 ) | ( n14914 & n15224 ) ;
  assign n15235 = n14813 | n15224 ;
  assign n15237 = ( n15234 & ~n15236 ) | ( n15234 & n15235 ) | ( ~n15236 & n15235 ) ;
  assign n15241 = n14694 &  n14913 ;
  assign n15242 = n14912 &  n15241 ;
  assign n15230 = x79 | n14694 ;
  assign n15231 = x79 &  n14694 ;
  assign n15232 = ( n15230 & ~n15231 ) | ( n15230 & 1'b0 ) | ( ~n15231 & 1'b0 ) ;
  assign n15244 = ( n14812 & n14914 ) | ( n14812 & n15232 ) | ( n14914 & n15232 ) ;
  assign n15243 = n14812 | n15232 ;
  assign n15245 = ( n15242 & ~n15244 ) | ( n15242 & n15243 ) | ( ~n15244 & n15243 ) ;
  assign n15249 = n14702 &  n14913 ;
  assign n15250 = n14912 &  n15249 ;
  assign n15238 = x78 | n14702 ;
  assign n15239 = x78 &  n14702 ;
  assign n15240 = ( n15238 & ~n15239 ) | ( n15238 & 1'b0 ) | ( ~n15239 & 1'b0 ) ;
  assign n15252 = ( n14811 & n14914 ) | ( n14811 & n15240 ) | ( n14914 & n15240 ) ;
  assign n15251 = n14811 | n15240 ;
  assign n15253 = ( n15250 & ~n15252 ) | ( n15250 & n15251 ) | ( ~n15252 & n15251 ) ;
  assign n15257 = n14710 &  n14913 ;
  assign n15258 = n14912 &  n15257 ;
  assign n15246 = x77 | n14710 ;
  assign n15247 = x77 &  n14710 ;
  assign n15248 = ( n15246 & ~n15247 ) | ( n15246 & 1'b0 ) | ( ~n15247 & 1'b0 ) ;
  assign n15260 = ( n14810 & n14914 ) | ( n14810 & n15248 ) | ( n14914 & n15248 ) ;
  assign n15259 = n14810 | n15248 ;
  assign n15261 = ( n15258 & ~n15260 ) | ( n15258 & n15259 ) | ( ~n15260 & n15259 ) ;
  assign n15265 = n14718 &  n14913 ;
  assign n15266 = n14912 &  n15265 ;
  assign n15254 = x76 | n14718 ;
  assign n15255 = x76 &  n14718 ;
  assign n15256 = ( n15254 & ~n15255 ) | ( n15254 & 1'b0 ) | ( ~n15255 & 1'b0 ) ;
  assign n15268 = ( n14809 & n14914 ) | ( n14809 & n15256 ) | ( n14914 & n15256 ) ;
  assign n15267 = n14809 | n15256 ;
  assign n15269 = ( n15266 & ~n15268 ) | ( n15266 & n15267 ) | ( ~n15268 & n15267 ) ;
  assign n15273 = n14726 &  n14913 ;
  assign n15274 = n14912 &  n15273 ;
  assign n15262 = x75 | n14726 ;
  assign n15263 = x75 &  n14726 ;
  assign n15264 = ( n15262 & ~n15263 ) | ( n15262 & 1'b0 ) | ( ~n15263 & 1'b0 ) ;
  assign n15276 = ( n14808 & n14914 ) | ( n14808 & n15264 ) | ( n14914 & n15264 ) ;
  assign n15275 = n14808 | n15264 ;
  assign n15277 = ( n15274 & ~n15276 ) | ( n15274 & n15275 ) | ( ~n15276 & n15275 ) ;
  assign n15281 = n14734 &  n14913 ;
  assign n15282 = n14912 &  n15281 ;
  assign n15270 = x74 | n14734 ;
  assign n15271 = x74 &  n14734 ;
  assign n15272 = ( n15270 & ~n15271 ) | ( n15270 & 1'b0 ) | ( ~n15271 & 1'b0 ) ;
  assign n15284 = ( n14807 & n14914 ) | ( n14807 & n15272 ) | ( n14914 & n15272 ) ;
  assign n15283 = n14807 | n15272 ;
  assign n15285 = ( n15282 & ~n15284 ) | ( n15282 & n15283 ) | ( ~n15284 & n15283 ) ;
  assign n15289 = n14742 &  n14913 ;
  assign n15290 = n14912 &  n15289 ;
  assign n15278 = x73 | n14742 ;
  assign n15279 = x73 &  n14742 ;
  assign n15280 = ( n15278 & ~n15279 ) | ( n15278 & 1'b0 ) | ( ~n15279 & 1'b0 ) ;
  assign n15292 = ( n14806 & n14914 ) | ( n14806 & n15280 ) | ( n14914 & n15280 ) ;
  assign n15291 = n14806 | n15280 ;
  assign n15293 = ( n15290 & ~n15292 ) | ( n15290 & n15291 ) | ( ~n15292 & n15291 ) ;
  assign n15297 = n14750 &  n14913 ;
  assign n15298 = n14912 &  n15297 ;
  assign n15286 = x72 | n14750 ;
  assign n15287 = x72 &  n14750 ;
  assign n15288 = ( n15286 & ~n15287 ) | ( n15286 & 1'b0 ) | ( ~n15287 & 1'b0 ) ;
  assign n15300 = ( n14805 & n14914 ) | ( n14805 & n15288 ) | ( n14914 & n15288 ) ;
  assign n15299 = n14805 | n15288 ;
  assign n15301 = ( n15298 & ~n15300 ) | ( n15298 & n15299 ) | ( ~n15300 & n15299 ) ;
  assign n15305 = n14758 &  n14913 ;
  assign n15306 = n14912 &  n15305 ;
  assign n15294 = x71 | n14758 ;
  assign n15295 = x71 &  n14758 ;
  assign n15296 = ( n15294 & ~n15295 ) | ( n15294 & 1'b0 ) | ( ~n15295 & 1'b0 ) ;
  assign n15308 = ( n14804 & n14914 ) | ( n14804 & n15296 ) | ( n14914 & n15296 ) ;
  assign n15307 = n14804 | n15296 ;
  assign n15309 = ( n15306 & ~n15308 ) | ( n15306 & n15307 ) | ( ~n15308 & n15307 ) ;
  assign n15313 = n14766 &  n14913 ;
  assign n15314 = n14912 &  n15313 ;
  assign n15302 = x70 | n14766 ;
  assign n15303 = x70 &  n14766 ;
  assign n15304 = ( n15302 & ~n15303 ) | ( n15302 & 1'b0 ) | ( ~n15303 & 1'b0 ) ;
  assign n15316 = ( n14803 & n14914 ) | ( n14803 & n15304 ) | ( n14914 & n15304 ) ;
  assign n15315 = n14803 | n15304 ;
  assign n15317 = ( n15314 & ~n15316 ) | ( n15314 & n15315 ) | ( ~n15316 & n15315 ) ;
  assign n15321 = n14774 &  n14913 ;
  assign n15322 = n14912 &  n15321 ;
  assign n15310 = x69 | n14774 ;
  assign n15311 = x69 &  n14774 ;
  assign n15312 = ( n15310 & ~n15311 ) | ( n15310 & 1'b0 ) | ( ~n15311 & 1'b0 ) ;
  assign n15324 = ( n14802 & n14914 ) | ( n14802 & n15312 ) | ( n14914 & n15312 ) ;
  assign n15323 = n14802 | n15312 ;
  assign n15325 = ( n15322 & ~n15324 ) | ( n15322 & n15323 ) | ( ~n15324 & n15323 ) ;
  assign n15329 = n14782 &  n14913 ;
  assign n15330 = n14912 &  n15329 ;
  assign n15318 = x68 | n14782 ;
  assign n15319 = x68 &  n14782 ;
  assign n15320 = ( n15318 & ~n15319 ) | ( n15318 & 1'b0 ) | ( ~n15319 & 1'b0 ) ;
  assign n15332 = ( n14801 & n14914 ) | ( n14801 & n15320 ) | ( n14914 & n15320 ) ;
  assign n15331 = n14801 | n15320 ;
  assign n15333 = ( n15330 & ~n15332 ) | ( n15330 & n15331 ) | ( ~n15332 & n15331 ) ;
  assign n15337 = n14787 &  n14913 ;
  assign n15338 = n14912 &  n15337 ;
  assign n15326 = x67 | n14787 ;
  assign n15327 = x67 &  n14787 ;
  assign n15328 = ( n15326 & ~n15327 ) | ( n15326 & 1'b0 ) | ( ~n15327 & 1'b0 ) ;
  assign n15340 = ( n14800 & n14914 ) | ( n14800 & n15328 ) | ( n14914 & n15328 ) ;
  assign n15339 = n14800 | n15328 ;
  assign n15341 = ( n15338 & ~n15340 ) | ( n15338 & n15339 ) | ( ~n15340 & n15339 ) ;
  assign n15342 = n14793 &  n14913 ;
  assign n15343 = n14912 &  n15342 ;
  assign n15334 = x66 | n14793 ;
  assign n15335 = x66 &  n14793 ;
  assign n15336 = ( n15334 & ~n15335 ) | ( n15334 & 1'b0 ) | ( ~n15335 & 1'b0 ) ;
  assign n15344 = n14799 &  n15336 ;
  assign n15345 = ( n14799 & ~n14914 ) | ( n14799 & n15336 ) | ( ~n14914 & n15336 ) ;
  assign n15346 = ( n15343 & ~n15344 ) | ( n15343 & n15345 ) | ( ~n15344 & n15345 ) ;
  assign n15347 = ( n14797 & ~x65 ) | ( n14797 & n14798 ) | ( ~x65 & n14798 ) ;
  assign n15348 = ( n14799 & ~n14798 ) | ( n14799 & n15347 ) | ( ~n14798 & n15347 ) ;
  assign n15349 = ~n14914 & n15348 ;
  assign n15350 = n14797 &  n14913 ;
  assign n15351 = n14912 &  n15350 ;
  assign n15352 = n15349 | n15351 ;
  assign n15353 = ( x64 & ~n14914 ) | ( x64 & 1'b0 ) | ( ~n14914 & 1'b0 ) ;
  assign n15354 = ( x7 & ~n15353 ) | ( x7 & 1'b0 ) | ( ~n15353 & 1'b0 ) ;
  assign n15355 = ( n14798 & ~n14914 ) | ( n14798 & 1'b0 ) | ( ~n14914 & 1'b0 ) ;
  assign n15356 = n15354 | n15355 ;
  assign n15357 = ~x6 & x64 ;
  assign n15358 = ( x65 & ~n15356 ) | ( x65 & n15357 ) | ( ~n15356 & n15357 ) ;
  assign n15359 = ( x66 & ~n15352 ) | ( x66 & n15358 ) | ( ~n15352 & n15358 ) ;
  assign n15360 = ( x67 & ~n15346 ) | ( x67 & n15359 ) | ( ~n15346 & n15359 ) ;
  assign n15361 = ( x68 & ~n15341 ) | ( x68 & n15360 ) | ( ~n15341 & n15360 ) ;
  assign n15362 = ( x69 & ~n15333 ) | ( x69 & n15361 ) | ( ~n15333 & n15361 ) ;
  assign n15363 = ( x70 & ~n15325 ) | ( x70 & n15362 ) | ( ~n15325 & n15362 ) ;
  assign n15364 = ( x71 & ~n15317 ) | ( x71 & n15363 ) | ( ~n15317 & n15363 ) ;
  assign n15365 = ( x72 & ~n15309 ) | ( x72 & n15364 ) | ( ~n15309 & n15364 ) ;
  assign n15366 = ( x73 & ~n15301 ) | ( x73 & n15365 ) | ( ~n15301 & n15365 ) ;
  assign n15367 = ( x74 & ~n15293 ) | ( x74 & n15366 ) | ( ~n15293 & n15366 ) ;
  assign n15368 = ( x75 & ~n15285 ) | ( x75 & n15367 ) | ( ~n15285 & n15367 ) ;
  assign n15369 = ( x76 & ~n15277 ) | ( x76 & n15368 ) | ( ~n15277 & n15368 ) ;
  assign n15370 = ( x77 & ~n15269 ) | ( x77 & n15369 ) | ( ~n15269 & n15369 ) ;
  assign n15371 = ( x78 & ~n15261 ) | ( x78 & n15370 ) | ( ~n15261 & n15370 ) ;
  assign n15372 = ( x79 & ~n15253 ) | ( x79 & n15371 ) | ( ~n15253 & n15371 ) ;
  assign n15373 = ( x80 & ~n15245 ) | ( x80 & n15372 ) | ( ~n15245 & n15372 ) ;
  assign n15374 = ( x81 & ~n15237 ) | ( x81 & n15373 ) | ( ~n15237 & n15373 ) ;
  assign n15375 = ( x82 & ~n15229 ) | ( x82 & n15374 ) | ( ~n15229 & n15374 ) ;
  assign n15376 = ( x83 & ~n15221 ) | ( x83 & n15375 ) | ( ~n15221 & n15375 ) ;
  assign n15377 = ( x84 & ~n15213 ) | ( x84 & n15376 ) | ( ~n15213 & n15376 ) ;
  assign n15378 = ( x85 & ~n15205 ) | ( x85 & n15377 ) | ( ~n15205 & n15377 ) ;
  assign n15379 = ( x86 & ~n15197 ) | ( x86 & n15378 ) | ( ~n15197 & n15378 ) ;
  assign n15380 = ( x87 & ~n15189 ) | ( x87 & n15379 ) | ( ~n15189 & n15379 ) ;
  assign n15381 = ( x88 & ~n15181 ) | ( x88 & n15380 ) | ( ~n15181 & n15380 ) ;
  assign n15382 = ( x89 & ~n15173 ) | ( x89 & n15381 ) | ( ~n15173 & n15381 ) ;
  assign n15383 = ( x90 & ~n15165 ) | ( x90 & n15382 ) | ( ~n15165 & n15382 ) ;
  assign n15384 = ( x91 & ~n15157 ) | ( x91 & n15383 ) | ( ~n15157 & n15383 ) ;
  assign n15385 = ( x92 & ~n15149 ) | ( x92 & n15384 ) | ( ~n15149 & n15384 ) ;
  assign n15386 = ( x93 & ~n15141 ) | ( x93 & n15385 ) | ( ~n15141 & n15385 ) ;
  assign n15387 = ( x94 & ~n15133 ) | ( x94 & n15386 ) | ( ~n15133 & n15386 ) ;
  assign n15388 = ( x95 & ~n15125 ) | ( x95 & n15387 ) | ( ~n15125 & n15387 ) ;
  assign n15389 = ( x96 & ~n15117 ) | ( x96 & n15388 ) | ( ~n15117 & n15388 ) ;
  assign n15390 = ( x97 & ~n15109 ) | ( x97 & n15389 ) | ( ~n15109 & n15389 ) ;
  assign n15391 = ( x98 & ~n15101 ) | ( x98 & n15390 ) | ( ~n15101 & n15390 ) ;
  assign n15392 = ( x99 & ~n15093 ) | ( x99 & n15391 ) | ( ~n15093 & n15391 ) ;
  assign n15393 = ( x100 & ~n15085 ) | ( x100 & n15392 ) | ( ~n15085 & n15392 ) ;
  assign n15394 = ( x101 & ~n15077 ) | ( x101 & n15393 ) | ( ~n15077 & n15393 ) ;
  assign n15395 = ( x102 & ~n15069 ) | ( x102 & n15394 ) | ( ~n15069 & n15394 ) ;
  assign n15396 = ( x103 & ~n15061 ) | ( x103 & n15395 ) | ( ~n15061 & n15395 ) ;
  assign n15397 = ( x104 & ~n15053 ) | ( x104 & n15396 ) | ( ~n15053 & n15396 ) ;
  assign n15398 = ( x105 & ~n15045 ) | ( x105 & n15397 ) | ( ~n15045 & n15397 ) ;
  assign n15399 = ( x106 & ~n15037 ) | ( x106 & n15398 ) | ( ~n15037 & n15398 ) ;
  assign n15400 = ( x107 & ~n15029 ) | ( x107 & n15399 ) | ( ~n15029 & n15399 ) ;
  assign n15401 = ( x108 & ~n15021 ) | ( x108 & n15400 ) | ( ~n15021 & n15400 ) ;
  assign n15402 = ( x109 & ~n15013 ) | ( x109 & n15401 ) | ( ~n15013 & n15401 ) ;
  assign n15403 = ( x110 & ~n15005 ) | ( x110 & n15402 ) | ( ~n15005 & n15402 ) ;
  assign n15404 = ( x111 & ~n14997 ) | ( x111 & n15403 ) | ( ~n14997 & n15403 ) ;
  assign n15405 = ( x112 & ~n14989 ) | ( x112 & n15404 ) | ( ~n14989 & n15404 ) ;
  assign n15406 = ( x113 & ~n14981 ) | ( x113 & n15405 ) | ( ~n14981 & n15405 ) ;
  assign n15407 = ( x114 & ~n14973 ) | ( x114 & n15406 ) | ( ~n14973 & n15406 ) ;
  assign n15408 = ( x115 & ~n14965 ) | ( x115 & n15407 ) | ( ~n14965 & n15407 ) ;
  assign n15409 = ( x116 & ~n14919 ) | ( x116 & n15408 ) | ( ~n14919 & n15408 ) ;
  assign n15410 = ( x117 & ~n14957 ) | ( x117 & n15409 ) | ( ~n14957 & n15409 ) ;
  assign n15411 = ( x118 & ~n14952 ) | ( x118 & n15410 ) | ( ~n14952 & n15410 ) ;
  assign n15412 = ( x119 & ~n14944 ) | ( x119 & n15411 ) | ( ~n14944 & n15411 ) ;
  assign n15413 = ( x120 & ~n14936 ) | ( x120 & n15412 ) | ( ~n14936 & n15412 ) ;
  assign n15414 = ( x121 & ~n14928 ) | ( x121 & n15413 ) | ( ~n14928 & n15413 ) ;
  assign n15415 = n152 | n154 ;
  assign n15416 = n15414 | n15415 ;
  assign n15912 = n14936 &  n15416 ;
  assign n15916 = x120 | n14936 ;
  assign n15917 = x120 &  n14936 ;
  assign n15918 = ( n15916 & ~n15917 ) | ( n15916 & 1'b0 ) | ( ~n15917 & 1'b0 ) ;
  assign n15919 = ( n15412 & n15414 ) | ( n15412 & n15918 ) | ( n15414 & n15918 ) ;
  assign n15920 = ( n15412 & ~n15415 ) | ( n15412 & n15918 ) | ( ~n15415 & n15918 ) ;
  assign n15921 = ~n15919 & n15920 ;
  assign n15922 = n15912 | n15921 ;
  assign n15923 = n14944 &  n15416 ;
  assign n15913 = x119 | n14944 ;
  assign n15914 = x119 &  n14944 ;
  assign n15915 = ( n15913 & ~n15914 ) | ( n15913 & 1'b0 ) | ( ~n15914 & 1'b0 ) ;
  assign n15927 = ( n15411 & n15414 ) | ( n15411 & n15915 ) | ( n15414 & n15915 ) ;
  assign n15928 = ( n15411 & ~n15415 ) | ( n15411 & n15915 ) | ( ~n15415 & n15915 ) ;
  assign n15929 = ~n15927 & n15928 ;
  assign n15930 = n15923 | n15929 ;
  assign n15931 = n14952 &  n15416 ;
  assign n15924 = x118 | n14952 ;
  assign n15925 = x118 &  n14952 ;
  assign n15926 = ( n15924 & ~n15925 ) | ( n15924 & 1'b0 ) | ( ~n15925 & 1'b0 ) ;
  assign n15932 = ( n15410 & n15414 ) | ( n15410 & n15926 ) | ( n15414 & n15926 ) ;
  assign n15933 = ( n15410 & ~n15415 ) | ( n15410 & n15926 ) | ( ~n15415 & n15926 ) ;
  assign n15934 = ~n15932 & n15933 ;
  assign n15935 = n15931 | n15934 ;
  assign n15901 = n14957 &  n15416 ;
  assign n15902 = x117 | n14957 ;
  assign n15903 = x117 &  n14957 ;
  assign n15904 = ( n15902 & ~n15903 ) | ( n15902 & 1'b0 ) | ( ~n15903 & 1'b0 ) ;
  assign n15905 = ( n15409 & n15414 ) | ( n15409 & n15904 ) | ( n15414 & n15904 ) ;
  assign n15906 = ( n15409 & ~n15415 ) | ( n15409 & n15904 ) | ( ~n15415 & n15904 ) ;
  assign n15907 = ~n15905 & n15906 ;
  assign n15908 = n15901 | n15907 ;
  assign n15417 = n14919 &  n15416 ;
  assign n15421 = x116 | n14919 ;
  assign n15422 = x116 &  n14919 ;
  assign n15423 = ( n15421 & ~n15422 ) | ( n15421 & 1'b0 ) | ( ~n15422 & 1'b0 ) ;
  assign n15424 = ( n15408 & n15414 ) | ( n15408 & n15423 ) | ( n15414 & n15423 ) ;
  assign n15425 = ( n15408 & ~n15415 ) | ( n15408 & n15423 ) | ( ~n15415 & n15423 ) ;
  assign n15426 = ~n15424 & n15425 ;
  assign n15427 = n15417 | n15426 ;
  assign n15428 = n14965 &  n15416 ;
  assign n15418 = x115 | n14965 ;
  assign n15419 = x115 &  n14965 ;
  assign n15420 = ( n15418 & ~n15419 ) | ( n15418 & 1'b0 ) | ( ~n15419 & 1'b0 ) ;
  assign n15432 = ( n15407 & n15414 ) | ( n15407 & n15420 ) | ( n15414 & n15420 ) ;
  assign n15433 = ( n15407 & ~n15415 ) | ( n15407 & n15420 ) | ( ~n15415 & n15420 ) ;
  assign n15434 = ~n15432 & n15433 ;
  assign n15435 = n15428 | n15434 ;
  assign n15436 = n14973 &  n15416 ;
  assign n15429 = x114 | n14973 ;
  assign n15430 = x114 &  n14973 ;
  assign n15431 = ( n15429 & ~n15430 ) | ( n15429 & 1'b0 ) | ( ~n15430 & 1'b0 ) ;
  assign n15440 = ( n15406 & n15414 ) | ( n15406 & n15431 ) | ( n15414 & n15431 ) ;
  assign n15441 = ( n15406 & ~n15415 ) | ( n15406 & n15431 ) | ( ~n15415 & n15431 ) ;
  assign n15442 = ~n15440 & n15441 ;
  assign n15443 = n15436 | n15442 ;
  assign n15444 = n14981 &  n15416 ;
  assign n15437 = x113 | n14981 ;
  assign n15438 = x113 &  n14981 ;
  assign n15439 = ( n15437 & ~n15438 ) | ( n15437 & 1'b0 ) | ( ~n15438 & 1'b0 ) ;
  assign n15448 = ( n15405 & n15414 ) | ( n15405 & n15439 ) | ( n15414 & n15439 ) ;
  assign n15449 = ( n15405 & ~n15415 ) | ( n15405 & n15439 ) | ( ~n15415 & n15439 ) ;
  assign n15450 = ~n15448 & n15449 ;
  assign n15451 = n15444 | n15450 ;
  assign n15452 = n14989 &  n15416 ;
  assign n15445 = x112 | n14989 ;
  assign n15446 = x112 &  n14989 ;
  assign n15447 = ( n15445 & ~n15446 ) | ( n15445 & 1'b0 ) | ( ~n15446 & 1'b0 ) ;
  assign n15456 = ( n15404 & n15414 ) | ( n15404 & n15447 ) | ( n15414 & n15447 ) ;
  assign n15457 = ( n15404 & ~n15415 ) | ( n15404 & n15447 ) | ( ~n15415 & n15447 ) ;
  assign n15458 = ~n15456 & n15457 ;
  assign n15459 = n15452 | n15458 ;
  assign n15460 = n14997 &  n15416 ;
  assign n15453 = x111 | n14997 ;
  assign n15454 = x111 &  n14997 ;
  assign n15455 = ( n15453 & ~n15454 ) | ( n15453 & 1'b0 ) | ( ~n15454 & 1'b0 ) ;
  assign n15464 = ( n15403 & n15414 ) | ( n15403 & n15455 ) | ( n15414 & n15455 ) ;
  assign n15465 = ( n15403 & ~n15415 ) | ( n15403 & n15455 ) | ( ~n15415 & n15455 ) ;
  assign n15466 = ~n15464 & n15465 ;
  assign n15467 = n15460 | n15466 ;
  assign n15468 = n15005 &  n15416 ;
  assign n15461 = x110 | n15005 ;
  assign n15462 = x110 &  n15005 ;
  assign n15463 = ( n15461 & ~n15462 ) | ( n15461 & 1'b0 ) | ( ~n15462 & 1'b0 ) ;
  assign n15472 = ( n15402 & n15414 ) | ( n15402 & n15463 ) | ( n15414 & n15463 ) ;
  assign n15473 = ( n15402 & ~n15415 ) | ( n15402 & n15463 ) | ( ~n15415 & n15463 ) ;
  assign n15474 = ~n15472 & n15473 ;
  assign n15475 = n15468 | n15474 ;
  assign n15476 = n15013 &  n15416 ;
  assign n15469 = x109 | n15013 ;
  assign n15470 = x109 &  n15013 ;
  assign n15471 = ( n15469 & ~n15470 ) | ( n15469 & 1'b0 ) | ( ~n15470 & 1'b0 ) ;
  assign n15480 = ( n15401 & n15414 ) | ( n15401 & n15471 ) | ( n15414 & n15471 ) ;
  assign n15481 = ( n15401 & ~n15415 ) | ( n15401 & n15471 ) | ( ~n15415 & n15471 ) ;
  assign n15482 = ~n15480 & n15481 ;
  assign n15483 = n15476 | n15482 ;
  assign n15484 = n15021 &  n15416 ;
  assign n15477 = x108 | n15021 ;
  assign n15478 = x108 &  n15021 ;
  assign n15479 = ( n15477 & ~n15478 ) | ( n15477 & 1'b0 ) | ( ~n15478 & 1'b0 ) ;
  assign n15488 = ( n15400 & n15414 ) | ( n15400 & n15479 ) | ( n15414 & n15479 ) ;
  assign n15489 = ( n15400 & ~n15415 ) | ( n15400 & n15479 ) | ( ~n15415 & n15479 ) ;
  assign n15490 = ~n15488 & n15489 ;
  assign n15491 = n15484 | n15490 ;
  assign n15492 = n15029 &  n15416 ;
  assign n15485 = x107 | n15029 ;
  assign n15486 = x107 &  n15029 ;
  assign n15487 = ( n15485 & ~n15486 ) | ( n15485 & 1'b0 ) | ( ~n15486 & 1'b0 ) ;
  assign n15496 = ( n15399 & n15414 ) | ( n15399 & n15487 ) | ( n15414 & n15487 ) ;
  assign n15497 = ( n15399 & ~n15415 ) | ( n15399 & n15487 ) | ( ~n15415 & n15487 ) ;
  assign n15498 = ~n15496 & n15497 ;
  assign n15499 = n15492 | n15498 ;
  assign n15500 = n15037 &  n15416 ;
  assign n15493 = x106 | n15037 ;
  assign n15494 = x106 &  n15037 ;
  assign n15495 = ( n15493 & ~n15494 ) | ( n15493 & 1'b0 ) | ( ~n15494 & 1'b0 ) ;
  assign n15504 = ( n15398 & n15414 ) | ( n15398 & n15495 ) | ( n15414 & n15495 ) ;
  assign n15505 = ( n15398 & ~n15415 ) | ( n15398 & n15495 ) | ( ~n15415 & n15495 ) ;
  assign n15506 = ~n15504 & n15505 ;
  assign n15507 = n15500 | n15506 ;
  assign n15508 = n15045 &  n15416 ;
  assign n15501 = x105 | n15045 ;
  assign n15502 = x105 &  n15045 ;
  assign n15503 = ( n15501 & ~n15502 ) | ( n15501 & 1'b0 ) | ( ~n15502 & 1'b0 ) ;
  assign n15512 = ( n15397 & n15414 ) | ( n15397 & n15503 ) | ( n15414 & n15503 ) ;
  assign n15513 = ( n15397 & ~n15415 ) | ( n15397 & n15503 ) | ( ~n15415 & n15503 ) ;
  assign n15514 = ~n15512 & n15513 ;
  assign n15515 = n15508 | n15514 ;
  assign n15516 = n15053 &  n15416 ;
  assign n15509 = x104 | n15053 ;
  assign n15510 = x104 &  n15053 ;
  assign n15511 = ( n15509 & ~n15510 ) | ( n15509 & 1'b0 ) | ( ~n15510 & 1'b0 ) ;
  assign n15520 = ( n15396 & n15414 ) | ( n15396 & n15511 ) | ( n15414 & n15511 ) ;
  assign n15521 = ( n15396 & ~n15415 ) | ( n15396 & n15511 ) | ( ~n15415 & n15511 ) ;
  assign n15522 = ~n15520 & n15521 ;
  assign n15523 = n15516 | n15522 ;
  assign n15524 = n15061 &  n15416 ;
  assign n15517 = x103 | n15061 ;
  assign n15518 = x103 &  n15061 ;
  assign n15519 = ( n15517 & ~n15518 ) | ( n15517 & 1'b0 ) | ( ~n15518 & 1'b0 ) ;
  assign n15528 = ( n15395 & n15414 ) | ( n15395 & n15519 ) | ( n15414 & n15519 ) ;
  assign n15529 = ( n15395 & ~n15415 ) | ( n15395 & n15519 ) | ( ~n15415 & n15519 ) ;
  assign n15530 = ~n15528 & n15529 ;
  assign n15531 = n15524 | n15530 ;
  assign n15532 = n15069 &  n15416 ;
  assign n15525 = x102 | n15069 ;
  assign n15526 = x102 &  n15069 ;
  assign n15527 = ( n15525 & ~n15526 ) | ( n15525 & 1'b0 ) | ( ~n15526 & 1'b0 ) ;
  assign n15536 = ( n15394 & n15414 ) | ( n15394 & n15527 ) | ( n15414 & n15527 ) ;
  assign n15537 = ( n15394 & ~n15415 ) | ( n15394 & n15527 ) | ( ~n15415 & n15527 ) ;
  assign n15538 = ~n15536 & n15537 ;
  assign n15539 = n15532 | n15538 ;
  assign n15540 = n15077 &  n15416 ;
  assign n15533 = x101 | n15077 ;
  assign n15534 = x101 &  n15077 ;
  assign n15535 = ( n15533 & ~n15534 ) | ( n15533 & 1'b0 ) | ( ~n15534 & 1'b0 ) ;
  assign n15544 = ( n15393 & n15414 ) | ( n15393 & n15535 ) | ( n15414 & n15535 ) ;
  assign n15545 = ( n15393 & ~n15415 ) | ( n15393 & n15535 ) | ( ~n15415 & n15535 ) ;
  assign n15546 = ~n15544 & n15545 ;
  assign n15547 = n15540 | n15546 ;
  assign n15548 = n15085 &  n15416 ;
  assign n15541 = x100 | n15085 ;
  assign n15542 = x100 &  n15085 ;
  assign n15543 = ( n15541 & ~n15542 ) | ( n15541 & 1'b0 ) | ( ~n15542 & 1'b0 ) ;
  assign n15552 = ( n15392 & n15414 ) | ( n15392 & n15543 ) | ( n15414 & n15543 ) ;
  assign n15553 = ( n15392 & ~n15415 ) | ( n15392 & n15543 ) | ( ~n15415 & n15543 ) ;
  assign n15554 = ~n15552 & n15553 ;
  assign n15555 = n15548 | n15554 ;
  assign n15556 = n15093 &  n15416 ;
  assign n15549 = x99 | n15093 ;
  assign n15550 = x99 &  n15093 ;
  assign n15551 = ( n15549 & ~n15550 ) | ( n15549 & 1'b0 ) | ( ~n15550 & 1'b0 ) ;
  assign n15560 = ( n15391 & n15414 ) | ( n15391 & n15551 ) | ( n15414 & n15551 ) ;
  assign n15561 = ( n15391 & ~n15415 ) | ( n15391 & n15551 ) | ( ~n15415 & n15551 ) ;
  assign n15562 = ~n15560 & n15561 ;
  assign n15563 = n15556 | n15562 ;
  assign n15564 = n15101 &  n15416 ;
  assign n15557 = x98 | n15101 ;
  assign n15558 = x98 &  n15101 ;
  assign n15559 = ( n15557 & ~n15558 ) | ( n15557 & 1'b0 ) | ( ~n15558 & 1'b0 ) ;
  assign n15568 = ( n15390 & n15414 ) | ( n15390 & n15559 ) | ( n15414 & n15559 ) ;
  assign n15569 = ( n15390 & ~n15415 ) | ( n15390 & n15559 ) | ( ~n15415 & n15559 ) ;
  assign n15570 = ~n15568 & n15569 ;
  assign n15571 = n15564 | n15570 ;
  assign n15572 = n15109 &  n15416 ;
  assign n15565 = x97 | n15109 ;
  assign n15566 = x97 &  n15109 ;
  assign n15567 = ( n15565 & ~n15566 ) | ( n15565 & 1'b0 ) | ( ~n15566 & 1'b0 ) ;
  assign n15576 = ( n15389 & n15414 ) | ( n15389 & n15567 ) | ( n15414 & n15567 ) ;
  assign n15577 = ( n15389 & ~n15415 ) | ( n15389 & n15567 ) | ( ~n15415 & n15567 ) ;
  assign n15578 = ~n15576 & n15577 ;
  assign n15579 = n15572 | n15578 ;
  assign n15580 = n15117 &  n15416 ;
  assign n15573 = x96 | n15117 ;
  assign n15574 = x96 &  n15117 ;
  assign n15575 = ( n15573 & ~n15574 ) | ( n15573 & 1'b0 ) | ( ~n15574 & 1'b0 ) ;
  assign n15584 = ( n15388 & n15414 ) | ( n15388 & n15575 ) | ( n15414 & n15575 ) ;
  assign n15585 = ( n15388 & ~n15415 ) | ( n15388 & n15575 ) | ( ~n15415 & n15575 ) ;
  assign n15586 = ~n15584 & n15585 ;
  assign n15587 = n15580 | n15586 ;
  assign n15588 = n15125 &  n15416 ;
  assign n15581 = x95 | n15125 ;
  assign n15582 = x95 &  n15125 ;
  assign n15583 = ( n15581 & ~n15582 ) | ( n15581 & 1'b0 ) | ( ~n15582 & 1'b0 ) ;
  assign n15592 = ( n15387 & n15414 ) | ( n15387 & n15583 ) | ( n15414 & n15583 ) ;
  assign n15593 = ( n15387 & ~n15415 ) | ( n15387 & n15583 ) | ( ~n15415 & n15583 ) ;
  assign n15594 = ~n15592 & n15593 ;
  assign n15595 = n15588 | n15594 ;
  assign n15596 = n15133 &  n15416 ;
  assign n15589 = x94 | n15133 ;
  assign n15590 = x94 &  n15133 ;
  assign n15591 = ( n15589 & ~n15590 ) | ( n15589 & 1'b0 ) | ( ~n15590 & 1'b0 ) ;
  assign n15600 = ( n15386 & n15414 ) | ( n15386 & n15591 ) | ( n15414 & n15591 ) ;
  assign n15601 = ( n15386 & ~n15415 ) | ( n15386 & n15591 ) | ( ~n15415 & n15591 ) ;
  assign n15602 = ~n15600 & n15601 ;
  assign n15603 = n15596 | n15602 ;
  assign n15604 = n15141 &  n15416 ;
  assign n15597 = x93 | n15141 ;
  assign n15598 = x93 &  n15141 ;
  assign n15599 = ( n15597 & ~n15598 ) | ( n15597 & 1'b0 ) | ( ~n15598 & 1'b0 ) ;
  assign n15608 = ( n15385 & n15414 ) | ( n15385 & n15599 ) | ( n15414 & n15599 ) ;
  assign n15609 = ( n15385 & ~n15415 ) | ( n15385 & n15599 ) | ( ~n15415 & n15599 ) ;
  assign n15610 = ~n15608 & n15609 ;
  assign n15611 = n15604 | n15610 ;
  assign n15612 = n15149 &  n15416 ;
  assign n15605 = x92 | n15149 ;
  assign n15606 = x92 &  n15149 ;
  assign n15607 = ( n15605 & ~n15606 ) | ( n15605 & 1'b0 ) | ( ~n15606 & 1'b0 ) ;
  assign n15616 = ( n15384 & n15414 ) | ( n15384 & n15607 ) | ( n15414 & n15607 ) ;
  assign n15617 = ( n15384 & ~n15415 ) | ( n15384 & n15607 ) | ( ~n15415 & n15607 ) ;
  assign n15618 = ~n15616 & n15617 ;
  assign n15619 = n15612 | n15618 ;
  assign n15620 = n15157 &  n15416 ;
  assign n15613 = x91 | n15157 ;
  assign n15614 = x91 &  n15157 ;
  assign n15615 = ( n15613 & ~n15614 ) | ( n15613 & 1'b0 ) | ( ~n15614 & 1'b0 ) ;
  assign n15624 = ( n15383 & n15414 ) | ( n15383 & n15615 ) | ( n15414 & n15615 ) ;
  assign n15625 = ( n15383 & ~n15415 ) | ( n15383 & n15615 ) | ( ~n15415 & n15615 ) ;
  assign n15626 = ~n15624 & n15625 ;
  assign n15627 = n15620 | n15626 ;
  assign n15628 = n15165 &  n15416 ;
  assign n15621 = x90 | n15165 ;
  assign n15622 = x90 &  n15165 ;
  assign n15623 = ( n15621 & ~n15622 ) | ( n15621 & 1'b0 ) | ( ~n15622 & 1'b0 ) ;
  assign n15632 = ( n15382 & n15414 ) | ( n15382 & n15623 ) | ( n15414 & n15623 ) ;
  assign n15633 = ( n15382 & ~n15415 ) | ( n15382 & n15623 ) | ( ~n15415 & n15623 ) ;
  assign n15634 = ~n15632 & n15633 ;
  assign n15635 = n15628 | n15634 ;
  assign n15636 = n15173 &  n15416 ;
  assign n15629 = x89 | n15173 ;
  assign n15630 = x89 &  n15173 ;
  assign n15631 = ( n15629 & ~n15630 ) | ( n15629 & 1'b0 ) | ( ~n15630 & 1'b0 ) ;
  assign n15640 = ( n15381 & n15414 ) | ( n15381 & n15631 ) | ( n15414 & n15631 ) ;
  assign n15641 = ( n15381 & ~n15415 ) | ( n15381 & n15631 ) | ( ~n15415 & n15631 ) ;
  assign n15642 = ~n15640 & n15641 ;
  assign n15643 = n15636 | n15642 ;
  assign n15644 = n15181 &  n15416 ;
  assign n15637 = x88 | n15181 ;
  assign n15638 = x88 &  n15181 ;
  assign n15639 = ( n15637 & ~n15638 ) | ( n15637 & 1'b0 ) | ( ~n15638 & 1'b0 ) ;
  assign n15648 = ( n15380 & n15414 ) | ( n15380 & n15639 ) | ( n15414 & n15639 ) ;
  assign n15649 = ( n15380 & ~n15415 ) | ( n15380 & n15639 ) | ( ~n15415 & n15639 ) ;
  assign n15650 = ~n15648 & n15649 ;
  assign n15651 = n15644 | n15650 ;
  assign n15652 = n15189 &  n15416 ;
  assign n15645 = x87 | n15189 ;
  assign n15646 = x87 &  n15189 ;
  assign n15647 = ( n15645 & ~n15646 ) | ( n15645 & 1'b0 ) | ( ~n15646 & 1'b0 ) ;
  assign n15656 = ( n15379 & n15414 ) | ( n15379 & n15647 ) | ( n15414 & n15647 ) ;
  assign n15657 = ( n15379 & ~n15415 ) | ( n15379 & n15647 ) | ( ~n15415 & n15647 ) ;
  assign n15658 = ~n15656 & n15657 ;
  assign n15659 = n15652 | n15658 ;
  assign n15660 = n15197 &  n15416 ;
  assign n15653 = x86 | n15197 ;
  assign n15654 = x86 &  n15197 ;
  assign n15655 = ( n15653 & ~n15654 ) | ( n15653 & 1'b0 ) | ( ~n15654 & 1'b0 ) ;
  assign n15664 = ( n15378 & n15414 ) | ( n15378 & n15655 ) | ( n15414 & n15655 ) ;
  assign n15665 = ( n15378 & ~n15415 ) | ( n15378 & n15655 ) | ( ~n15415 & n15655 ) ;
  assign n15666 = ~n15664 & n15665 ;
  assign n15667 = n15660 | n15666 ;
  assign n15668 = n15205 &  n15416 ;
  assign n15661 = x85 | n15205 ;
  assign n15662 = x85 &  n15205 ;
  assign n15663 = ( n15661 & ~n15662 ) | ( n15661 & 1'b0 ) | ( ~n15662 & 1'b0 ) ;
  assign n15672 = ( n15377 & n15414 ) | ( n15377 & n15663 ) | ( n15414 & n15663 ) ;
  assign n15673 = ( n15377 & ~n15415 ) | ( n15377 & n15663 ) | ( ~n15415 & n15663 ) ;
  assign n15674 = ~n15672 & n15673 ;
  assign n15675 = n15668 | n15674 ;
  assign n15676 = n15213 &  n15416 ;
  assign n15669 = x84 | n15213 ;
  assign n15670 = x84 &  n15213 ;
  assign n15671 = ( n15669 & ~n15670 ) | ( n15669 & 1'b0 ) | ( ~n15670 & 1'b0 ) ;
  assign n15680 = ( n15376 & n15414 ) | ( n15376 & n15671 ) | ( n15414 & n15671 ) ;
  assign n15681 = ( n15376 & ~n15415 ) | ( n15376 & n15671 ) | ( ~n15415 & n15671 ) ;
  assign n15682 = ~n15680 & n15681 ;
  assign n15683 = n15676 | n15682 ;
  assign n15684 = n15221 &  n15416 ;
  assign n15677 = x83 | n15221 ;
  assign n15678 = x83 &  n15221 ;
  assign n15679 = ( n15677 & ~n15678 ) | ( n15677 & 1'b0 ) | ( ~n15678 & 1'b0 ) ;
  assign n15688 = ( n15375 & n15414 ) | ( n15375 & n15679 ) | ( n15414 & n15679 ) ;
  assign n15689 = ( n15375 & ~n15415 ) | ( n15375 & n15679 ) | ( ~n15415 & n15679 ) ;
  assign n15690 = ~n15688 & n15689 ;
  assign n15691 = n15684 | n15690 ;
  assign n15692 = n15229 &  n15416 ;
  assign n15685 = x82 | n15229 ;
  assign n15686 = x82 &  n15229 ;
  assign n15687 = ( n15685 & ~n15686 ) | ( n15685 & 1'b0 ) | ( ~n15686 & 1'b0 ) ;
  assign n15696 = ( n15374 & n15414 ) | ( n15374 & n15687 ) | ( n15414 & n15687 ) ;
  assign n15697 = ( n15374 & ~n15415 ) | ( n15374 & n15687 ) | ( ~n15415 & n15687 ) ;
  assign n15698 = ~n15696 & n15697 ;
  assign n15699 = n15692 | n15698 ;
  assign n15700 = n15237 &  n15416 ;
  assign n15693 = x81 | n15237 ;
  assign n15694 = x81 &  n15237 ;
  assign n15695 = ( n15693 & ~n15694 ) | ( n15693 & 1'b0 ) | ( ~n15694 & 1'b0 ) ;
  assign n15704 = ( n15373 & n15414 ) | ( n15373 & n15695 ) | ( n15414 & n15695 ) ;
  assign n15705 = ( n15373 & ~n15415 ) | ( n15373 & n15695 ) | ( ~n15415 & n15695 ) ;
  assign n15706 = ~n15704 & n15705 ;
  assign n15707 = n15700 | n15706 ;
  assign n15708 = n15245 &  n15416 ;
  assign n15701 = x80 | n15245 ;
  assign n15702 = x80 &  n15245 ;
  assign n15703 = ( n15701 & ~n15702 ) | ( n15701 & 1'b0 ) | ( ~n15702 & 1'b0 ) ;
  assign n15712 = ( n15372 & n15414 ) | ( n15372 & n15703 ) | ( n15414 & n15703 ) ;
  assign n15713 = ( n15372 & ~n15415 ) | ( n15372 & n15703 ) | ( ~n15415 & n15703 ) ;
  assign n15714 = ~n15712 & n15713 ;
  assign n15715 = n15708 | n15714 ;
  assign n15716 = n15253 &  n15416 ;
  assign n15709 = x79 | n15253 ;
  assign n15710 = x79 &  n15253 ;
  assign n15711 = ( n15709 & ~n15710 ) | ( n15709 & 1'b0 ) | ( ~n15710 & 1'b0 ) ;
  assign n15720 = ( n15371 & n15414 ) | ( n15371 & n15711 ) | ( n15414 & n15711 ) ;
  assign n15721 = ( n15371 & ~n15415 ) | ( n15371 & n15711 ) | ( ~n15415 & n15711 ) ;
  assign n15722 = ~n15720 & n15721 ;
  assign n15723 = n15716 | n15722 ;
  assign n15724 = n15261 &  n15416 ;
  assign n15717 = x78 | n15261 ;
  assign n15718 = x78 &  n15261 ;
  assign n15719 = ( n15717 & ~n15718 ) | ( n15717 & 1'b0 ) | ( ~n15718 & 1'b0 ) ;
  assign n15728 = ( n15370 & n15414 ) | ( n15370 & n15719 ) | ( n15414 & n15719 ) ;
  assign n15729 = ( n15370 & ~n15415 ) | ( n15370 & n15719 ) | ( ~n15415 & n15719 ) ;
  assign n15730 = ~n15728 & n15729 ;
  assign n15731 = n15724 | n15730 ;
  assign n15732 = n15269 &  n15416 ;
  assign n15725 = x77 | n15269 ;
  assign n15726 = x77 &  n15269 ;
  assign n15727 = ( n15725 & ~n15726 ) | ( n15725 & 1'b0 ) | ( ~n15726 & 1'b0 ) ;
  assign n15736 = ( n15369 & n15414 ) | ( n15369 & n15727 ) | ( n15414 & n15727 ) ;
  assign n15737 = ( n15369 & ~n15415 ) | ( n15369 & n15727 ) | ( ~n15415 & n15727 ) ;
  assign n15738 = ~n15736 & n15737 ;
  assign n15739 = n15732 | n15738 ;
  assign n15740 = n15277 &  n15416 ;
  assign n15733 = x76 | n15277 ;
  assign n15734 = x76 &  n15277 ;
  assign n15735 = ( n15733 & ~n15734 ) | ( n15733 & 1'b0 ) | ( ~n15734 & 1'b0 ) ;
  assign n15744 = ( n15368 & n15414 ) | ( n15368 & n15735 ) | ( n15414 & n15735 ) ;
  assign n15745 = ( n15368 & ~n15415 ) | ( n15368 & n15735 ) | ( ~n15415 & n15735 ) ;
  assign n15746 = ~n15744 & n15745 ;
  assign n15747 = n15740 | n15746 ;
  assign n15748 = n15285 &  n15416 ;
  assign n15741 = x75 | n15285 ;
  assign n15742 = x75 &  n15285 ;
  assign n15743 = ( n15741 & ~n15742 ) | ( n15741 & 1'b0 ) | ( ~n15742 & 1'b0 ) ;
  assign n15752 = ( n15367 & n15414 ) | ( n15367 & n15743 ) | ( n15414 & n15743 ) ;
  assign n15753 = ( n15367 & ~n15415 ) | ( n15367 & n15743 ) | ( ~n15415 & n15743 ) ;
  assign n15754 = ~n15752 & n15753 ;
  assign n15755 = n15748 | n15754 ;
  assign n15756 = n15293 &  n15416 ;
  assign n15749 = x74 | n15293 ;
  assign n15750 = x74 &  n15293 ;
  assign n15751 = ( n15749 & ~n15750 ) | ( n15749 & 1'b0 ) | ( ~n15750 & 1'b0 ) ;
  assign n15760 = ( n15366 & n15414 ) | ( n15366 & n15751 ) | ( n15414 & n15751 ) ;
  assign n15761 = ( n15366 & ~n15415 ) | ( n15366 & n15751 ) | ( ~n15415 & n15751 ) ;
  assign n15762 = ~n15760 & n15761 ;
  assign n15763 = n15756 | n15762 ;
  assign n15764 = n15301 &  n15416 ;
  assign n15757 = x73 | n15301 ;
  assign n15758 = x73 &  n15301 ;
  assign n15759 = ( n15757 & ~n15758 ) | ( n15757 & 1'b0 ) | ( ~n15758 & 1'b0 ) ;
  assign n15768 = ( n15365 & n15414 ) | ( n15365 & n15759 ) | ( n15414 & n15759 ) ;
  assign n15769 = ( n15365 & ~n15415 ) | ( n15365 & n15759 ) | ( ~n15415 & n15759 ) ;
  assign n15770 = ~n15768 & n15769 ;
  assign n15771 = n15764 | n15770 ;
  assign n15772 = n15309 &  n15416 ;
  assign n15765 = x72 | n15309 ;
  assign n15766 = x72 &  n15309 ;
  assign n15767 = ( n15765 & ~n15766 ) | ( n15765 & 1'b0 ) | ( ~n15766 & 1'b0 ) ;
  assign n15776 = ( n15364 & n15414 ) | ( n15364 & n15767 ) | ( n15414 & n15767 ) ;
  assign n15777 = ( n15364 & ~n15415 ) | ( n15364 & n15767 ) | ( ~n15415 & n15767 ) ;
  assign n15778 = ~n15776 & n15777 ;
  assign n15779 = n15772 | n15778 ;
  assign n15780 = n15317 &  n15416 ;
  assign n15773 = x71 | n15317 ;
  assign n15774 = x71 &  n15317 ;
  assign n15775 = ( n15773 & ~n15774 ) | ( n15773 & 1'b0 ) | ( ~n15774 & 1'b0 ) ;
  assign n15784 = ( n15363 & n15414 ) | ( n15363 & n15775 ) | ( n15414 & n15775 ) ;
  assign n15785 = ( n15363 & ~n15415 ) | ( n15363 & n15775 ) | ( ~n15415 & n15775 ) ;
  assign n15786 = ~n15784 & n15785 ;
  assign n15787 = n15780 | n15786 ;
  assign n15788 = n15325 &  n15416 ;
  assign n15781 = x70 | n15325 ;
  assign n15782 = x70 &  n15325 ;
  assign n15783 = ( n15781 & ~n15782 ) | ( n15781 & 1'b0 ) | ( ~n15782 & 1'b0 ) ;
  assign n15792 = ( n15362 & n15414 ) | ( n15362 & n15783 ) | ( n15414 & n15783 ) ;
  assign n15793 = ( n15362 & ~n15415 ) | ( n15362 & n15783 ) | ( ~n15415 & n15783 ) ;
  assign n15794 = ~n15792 & n15793 ;
  assign n15795 = n15788 | n15794 ;
  assign n15796 = n15333 &  n15416 ;
  assign n15789 = x69 | n15333 ;
  assign n15790 = x69 &  n15333 ;
  assign n15791 = ( n15789 & ~n15790 ) | ( n15789 & 1'b0 ) | ( ~n15790 & 1'b0 ) ;
  assign n15800 = ( n15361 & n15414 ) | ( n15361 & n15791 ) | ( n15414 & n15791 ) ;
  assign n15801 = ( n15361 & ~n15415 ) | ( n15361 & n15791 ) | ( ~n15415 & n15791 ) ;
  assign n15802 = ~n15800 & n15801 ;
  assign n15803 = n15796 | n15802 ;
  assign n15804 = n15341 &  n15416 ;
  assign n15797 = x68 | n15341 ;
  assign n15798 = x68 &  n15341 ;
  assign n15799 = ( n15797 & ~n15798 ) | ( n15797 & 1'b0 ) | ( ~n15798 & 1'b0 ) ;
  assign n15808 = ( n15360 & n15414 ) | ( n15360 & n15799 ) | ( n15414 & n15799 ) ;
  assign n15809 = ( n15360 & ~n15415 ) | ( n15360 & n15799 ) | ( ~n15415 & n15799 ) ;
  assign n15810 = ~n15808 & n15809 ;
  assign n15811 = n15804 | n15810 ;
  assign n15812 = n15346 &  n15416 ;
  assign n15805 = x67 | n15346 ;
  assign n15806 = x67 &  n15346 ;
  assign n15807 = ( n15805 & ~n15806 ) | ( n15805 & 1'b0 ) | ( ~n15806 & 1'b0 ) ;
  assign n15816 = ( n15359 & n15414 ) | ( n15359 & n15807 ) | ( n15414 & n15807 ) ;
  assign n15817 = ( n15359 & ~n15415 ) | ( n15359 & n15807 ) | ( ~n15415 & n15807 ) ;
  assign n15818 = ~n15816 & n15817 ;
  assign n15819 = n15812 | n15818 ;
  assign n15820 = n15352 &  n15416 ;
  assign n15813 = x66 | n15352 ;
  assign n15814 = x66 &  n15352 ;
  assign n15815 = ( n15813 & ~n15814 ) | ( n15813 & 1'b0 ) | ( ~n15814 & 1'b0 ) ;
  assign n15825 = ( n15358 & ~n15414 ) | ( n15358 & n15815 ) | ( ~n15414 & n15815 ) ;
  assign n15826 = ( n15358 & n15415 ) | ( n15358 & n15815 ) | ( n15415 & n15815 ) ;
  assign n15827 = ( n15825 & ~n15826 ) | ( n15825 & 1'b0 ) | ( ~n15826 & 1'b0 ) ;
  assign n15828 = n15820 | n15827 ;
  assign n15829 = n15356 &  n15416 ;
  assign n15821 = x65 &  n15356 ;
  assign n15822 = ( n15354 & ~x65 ) | ( n15354 & n15355 ) | ( ~x65 & n15355 ) ;
  assign n15823 = x65 | n15822 ;
  assign n15824 = ( n15357 & ~n15821 ) | ( n15357 & n15823 ) | ( ~n15821 & n15823 ) ;
  assign n15830 = ( x65 & n15356 ) | ( x65 & n15357 ) | ( n15356 & n15357 ) ;
  assign n15831 = ( n15415 & ~n15821 ) | ( n15415 & n15830 ) | ( ~n15821 & n15830 ) ;
  assign n15832 = ( n15414 & n15824 ) | ( n15414 & n15831 ) | ( n15824 & n15831 ) ;
  assign n15833 = ( n15824 & ~n15832 ) | ( n15824 & 1'b0 ) | ( ~n15832 & 1'b0 ) ;
  assign n15834 = n15829 | n15833 ;
  assign n15835 = ( x64 & ~x122 ) | ( x64 & 1'b0 ) | ( ~x122 & 1'b0 ) ;
  assign n15836 = ( n235 & ~n237 ) | ( n235 & n15835 ) | ( ~n237 & n15835 ) ;
  assign n15837 = ~n235 & n15836 ;
  assign n15838 = n15414 &  n15837 ;
  assign n15839 = ( x6 & ~n15837 ) | ( x6 & n15838 ) | ( ~n15837 & n15838 ) ;
  assign n15840 = ~n154 & n15357 ;
  assign n15841 = ~n152 & n15840 ;
  assign n15842 = ~n15414 & n15841 ;
  assign n15843 = n15839 | n15842 ;
  assign n15844 = ~x5 & x64 ;
  assign n15845 = ( x65 & ~n15843 ) | ( x65 & n15844 ) | ( ~n15843 & n15844 ) ;
  assign n15846 = ( x66 & ~n15834 ) | ( x66 & n15845 ) | ( ~n15834 & n15845 ) ;
  assign n15847 = ( x67 & ~n15828 ) | ( x67 & n15846 ) | ( ~n15828 & n15846 ) ;
  assign n15848 = ( x68 & ~n15819 ) | ( x68 & n15847 ) | ( ~n15819 & n15847 ) ;
  assign n15849 = ( x69 & ~n15811 ) | ( x69 & n15848 ) | ( ~n15811 & n15848 ) ;
  assign n15850 = ( x70 & ~n15803 ) | ( x70 & n15849 ) | ( ~n15803 & n15849 ) ;
  assign n15851 = ( x71 & ~n15795 ) | ( x71 & n15850 ) | ( ~n15795 & n15850 ) ;
  assign n15852 = ( x72 & ~n15787 ) | ( x72 & n15851 ) | ( ~n15787 & n15851 ) ;
  assign n15853 = ( x73 & ~n15779 ) | ( x73 & n15852 ) | ( ~n15779 & n15852 ) ;
  assign n15854 = ( x74 & ~n15771 ) | ( x74 & n15853 ) | ( ~n15771 & n15853 ) ;
  assign n15855 = ( x75 & ~n15763 ) | ( x75 & n15854 ) | ( ~n15763 & n15854 ) ;
  assign n15856 = ( x76 & ~n15755 ) | ( x76 & n15855 ) | ( ~n15755 & n15855 ) ;
  assign n15857 = ( x77 & ~n15747 ) | ( x77 & n15856 ) | ( ~n15747 & n15856 ) ;
  assign n15858 = ( x78 & ~n15739 ) | ( x78 & n15857 ) | ( ~n15739 & n15857 ) ;
  assign n15859 = ( x79 & ~n15731 ) | ( x79 & n15858 ) | ( ~n15731 & n15858 ) ;
  assign n15860 = ( x80 & ~n15723 ) | ( x80 & n15859 ) | ( ~n15723 & n15859 ) ;
  assign n15861 = ( x81 & ~n15715 ) | ( x81 & n15860 ) | ( ~n15715 & n15860 ) ;
  assign n15862 = ( x82 & ~n15707 ) | ( x82 & n15861 ) | ( ~n15707 & n15861 ) ;
  assign n15863 = ( x83 & ~n15699 ) | ( x83 & n15862 ) | ( ~n15699 & n15862 ) ;
  assign n15864 = ( x84 & ~n15691 ) | ( x84 & n15863 ) | ( ~n15691 & n15863 ) ;
  assign n15865 = ( x85 & ~n15683 ) | ( x85 & n15864 ) | ( ~n15683 & n15864 ) ;
  assign n15866 = ( x86 & ~n15675 ) | ( x86 & n15865 ) | ( ~n15675 & n15865 ) ;
  assign n15867 = ( x87 & ~n15667 ) | ( x87 & n15866 ) | ( ~n15667 & n15866 ) ;
  assign n15868 = ( x88 & ~n15659 ) | ( x88 & n15867 ) | ( ~n15659 & n15867 ) ;
  assign n15869 = ( x89 & ~n15651 ) | ( x89 & n15868 ) | ( ~n15651 & n15868 ) ;
  assign n15870 = ( x90 & ~n15643 ) | ( x90 & n15869 ) | ( ~n15643 & n15869 ) ;
  assign n15871 = ( x91 & ~n15635 ) | ( x91 & n15870 ) | ( ~n15635 & n15870 ) ;
  assign n15872 = ( x92 & ~n15627 ) | ( x92 & n15871 ) | ( ~n15627 & n15871 ) ;
  assign n15873 = ( x93 & ~n15619 ) | ( x93 & n15872 ) | ( ~n15619 & n15872 ) ;
  assign n15874 = ( x94 & ~n15611 ) | ( x94 & n15873 ) | ( ~n15611 & n15873 ) ;
  assign n15875 = ( x95 & ~n15603 ) | ( x95 & n15874 ) | ( ~n15603 & n15874 ) ;
  assign n15876 = ( x96 & ~n15595 ) | ( x96 & n15875 ) | ( ~n15595 & n15875 ) ;
  assign n15877 = ( x97 & ~n15587 ) | ( x97 & n15876 ) | ( ~n15587 & n15876 ) ;
  assign n15878 = ( x98 & ~n15579 ) | ( x98 & n15877 ) | ( ~n15579 & n15877 ) ;
  assign n15879 = ( x99 & ~n15571 ) | ( x99 & n15878 ) | ( ~n15571 & n15878 ) ;
  assign n15880 = ( x100 & ~n15563 ) | ( x100 & n15879 ) | ( ~n15563 & n15879 ) ;
  assign n15881 = ( x101 & ~n15555 ) | ( x101 & n15880 ) | ( ~n15555 & n15880 ) ;
  assign n15882 = ( x102 & ~n15547 ) | ( x102 & n15881 ) | ( ~n15547 & n15881 ) ;
  assign n15883 = ( x103 & ~n15539 ) | ( x103 & n15882 ) | ( ~n15539 & n15882 ) ;
  assign n15884 = ( x104 & ~n15531 ) | ( x104 & n15883 ) | ( ~n15531 & n15883 ) ;
  assign n15885 = ( x105 & ~n15523 ) | ( x105 & n15884 ) | ( ~n15523 & n15884 ) ;
  assign n15886 = ( x106 & ~n15515 ) | ( x106 & n15885 ) | ( ~n15515 & n15885 ) ;
  assign n15887 = ( x107 & ~n15507 ) | ( x107 & n15886 ) | ( ~n15507 & n15886 ) ;
  assign n15888 = ( x108 & ~n15499 ) | ( x108 & n15887 ) | ( ~n15499 & n15887 ) ;
  assign n15889 = ( x109 & ~n15491 ) | ( x109 & n15888 ) | ( ~n15491 & n15888 ) ;
  assign n15890 = ( x110 & ~n15483 ) | ( x110 & n15889 ) | ( ~n15483 & n15889 ) ;
  assign n15891 = ( x111 & ~n15475 ) | ( x111 & n15890 ) | ( ~n15475 & n15890 ) ;
  assign n15892 = ( x112 & ~n15467 ) | ( x112 & n15891 ) | ( ~n15467 & n15891 ) ;
  assign n15893 = ( x113 & ~n15459 ) | ( x113 & n15892 ) | ( ~n15459 & n15892 ) ;
  assign n15894 = ( x114 & ~n15451 ) | ( x114 & n15893 ) | ( ~n15451 & n15893 ) ;
  assign n15895 = ( x115 & ~n15443 ) | ( x115 & n15894 ) | ( ~n15443 & n15894 ) ;
  assign n15896 = ( x116 & ~n15435 ) | ( x116 & n15895 ) | ( ~n15435 & n15895 ) ;
  assign n15900 = ( x117 & ~n15427 ) | ( x117 & n15896 ) | ( ~n15427 & n15896 ) ;
  assign n15936 = ( x118 & ~n15908 ) | ( x118 & n15900 ) | ( ~n15908 & n15900 ) ;
  assign n15937 = ( x119 & ~n15935 ) | ( x119 & n15936 ) | ( ~n15935 & n15936 ) ;
  assign n15938 = ( x120 & ~n15930 ) | ( x120 & n15937 ) | ( ~n15930 & n15937 ) ;
  assign n15939 = ( x121 & ~n15922 ) | ( x121 & n15938 ) | ( ~n15922 & n15938 ) ;
  assign n15943 = n235 | n237 ;
  assign n15940 = x121 | n15413 ;
  assign n15941 = ( x121 & n15413 ) | ( x121 & n15415 ) | ( n15413 & n15415 ) ;
  assign n15942 = ( n14928 & ~n15940 ) | ( n14928 & n15941 ) | ( ~n15940 & n15941 ) ;
  assign n15945 = x122 &  n15942 ;
  assign n15944 = x122 | n15942 ;
  assign n15946 = ( n15943 & ~n15945 ) | ( n15943 & n15944 ) | ( ~n15945 & n15944 ) ;
  assign n15947 = n15939 | n15946 ;
  assign n15948 = ~n15942 |  n15415 ;
  assign n16454 = n15922 &  n15948 ;
  assign n16455 = n15947 &  n16454 ;
  assign n16451 = x121 | n15922 ;
  assign n16452 = x121 &  n15922 ;
  assign n16453 = ( n16451 & ~n16452 ) | ( n16451 & 1'b0 ) | ( ~n16452 & 1'b0 ) ;
  assign n16456 = n15938 &  n16453 ;
  assign n15949 = n15947 &  n15948 ;
  assign n16457 = ( n15938 & ~n15949 ) | ( n15938 & n16453 ) | ( ~n15949 & n16453 ) ;
  assign n16458 = ( n16455 & ~n16456 ) | ( n16455 & n16457 ) | ( ~n16456 & n16457 ) ;
  assign n16459 = n15930 &  n15948 ;
  assign n16460 = n15947 &  n16459 ;
  assign n16448 = x120 | n15930 ;
  assign n16449 = x120 &  n15930 ;
  assign n16450 = ( n16448 & ~n16449 ) | ( n16448 & 1'b0 ) | ( ~n16449 & 1'b0 ) ;
  assign n16461 = n15937 &  n16450 ;
  assign n16462 = ( n15937 & ~n15949 ) | ( n15937 & n16450 ) | ( ~n15949 & n16450 ) ;
  assign n16463 = ( n16460 & ~n16461 ) | ( n16460 & n16462 ) | ( ~n16461 & n16462 ) ;
  assign n16440 = n15935 &  n15948 ;
  assign n16441 = n15947 &  n16440 ;
  assign n16437 = x119 | n15935 ;
  assign n16438 = x119 &  n15935 ;
  assign n16439 = ( n16437 & ~n16438 ) | ( n16437 & 1'b0 ) | ( ~n16438 & 1'b0 ) ;
  assign n16442 = n15936 &  n16439 ;
  assign n16443 = ( n15936 & ~n15949 ) | ( n15936 & n16439 ) | ( ~n15949 & n16439 ) ;
  assign n16444 = ( n16441 & ~n16442 ) | ( n16441 & n16443 ) | ( ~n16442 & n16443 ) ;
  assign n15950 = n15908 &  n15948 ;
  assign n15951 = n15947 &  n15950 ;
  assign n15909 = x118 | n15908 ;
  assign n15910 = x118 &  n15908 ;
  assign n15911 = ( n15909 & ~n15910 ) | ( n15909 & 1'b0 ) | ( ~n15910 & 1'b0 ) ;
  assign n15952 = n15900 &  n15911 ;
  assign n15953 = ( n15900 & ~n15949 ) | ( n15900 & n15911 ) | ( ~n15949 & n15911 ) ;
  assign n15954 = ( n15951 & ~n15952 ) | ( n15951 & n15953 ) | ( ~n15952 & n15953 ) ;
  assign n15958 = n15427 &  n15948 ;
  assign n15959 = n15947 &  n15958 ;
  assign n15897 = x117 | n15427 ;
  assign n15898 = x117 &  n15427 ;
  assign n15899 = ( n15897 & ~n15898 ) | ( n15897 & 1'b0 ) | ( ~n15898 & 1'b0 ) ;
  assign n15961 = ( n15896 & n15899 ) | ( n15896 & n15949 ) | ( n15899 & n15949 ) ;
  assign n15960 = n15896 | n15899 ;
  assign n15962 = ( n15959 & ~n15961 ) | ( n15959 & n15960 ) | ( ~n15961 & n15960 ) ;
  assign n15966 = n15435 &  n15948 ;
  assign n15967 = n15947 &  n15966 ;
  assign n15955 = x116 | n15435 ;
  assign n15956 = x116 &  n15435 ;
  assign n15957 = ( n15955 & ~n15956 ) | ( n15955 & 1'b0 ) | ( ~n15956 & 1'b0 ) ;
  assign n15969 = ( n15895 & n15949 ) | ( n15895 & n15957 ) | ( n15949 & n15957 ) ;
  assign n15968 = n15895 | n15957 ;
  assign n15970 = ( n15967 & ~n15969 ) | ( n15967 & n15968 ) | ( ~n15969 & n15968 ) ;
  assign n15974 = n15443 &  n15948 ;
  assign n15975 = n15947 &  n15974 ;
  assign n15963 = x115 | n15443 ;
  assign n15964 = x115 &  n15443 ;
  assign n15965 = ( n15963 & ~n15964 ) | ( n15963 & 1'b0 ) | ( ~n15964 & 1'b0 ) ;
  assign n15977 = ( n15894 & n15949 ) | ( n15894 & n15965 ) | ( n15949 & n15965 ) ;
  assign n15976 = n15894 | n15965 ;
  assign n15978 = ( n15975 & ~n15977 ) | ( n15975 & n15976 ) | ( ~n15977 & n15976 ) ;
  assign n15982 = n15451 &  n15948 ;
  assign n15983 = n15947 &  n15982 ;
  assign n15971 = x114 | n15451 ;
  assign n15972 = x114 &  n15451 ;
  assign n15973 = ( n15971 & ~n15972 ) | ( n15971 & 1'b0 ) | ( ~n15972 & 1'b0 ) ;
  assign n15985 = ( n15893 & n15949 ) | ( n15893 & n15973 ) | ( n15949 & n15973 ) ;
  assign n15984 = n15893 | n15973 ;
  assign n15986 = ( n15983 & ~n15985 ) | ( n15983 & n15984 ) | ( ~n15985 & n15984 ) ;
  assign n15990 = n15459 &  n15948 ;
  assign n15991 = n15947 &  n15990 ;
  assign n15979 = x113 | n15459 ;
  assign n15980 = x113 &  n15459 ;
  assign n15981 = ( n15979 & ~n15980 ) | ( n15979 & 1'b0 ) | ( ~n15980 & 1'b0 ) ;
  assign n15993 = ( n15892 & n15949 ) | ( n15892 & n15981 ) | ( n15949 & n15981 ) ;
  assign n15992 = n15892 | n15981 ;
  assign n15994 = ( n15991 & ~n15993 ) | ( n15991 & n15992 ) | ( ~n15993 & n15992 ) ;
  assign n15998 = n15467 &  n15948 ;
  assign n15999 = n15947 &  n15998 ;
  assign n15987 = x112 | n15467 ;
  assign n15988 = x112 &  n15467 ;
  assign n15989 = ( n15987 & ~n15988 ) | ( n15987 & 1'b0 ) | ( ~n15988 & 1'b0 ) ;
  assign n16001 = ( n15891 & n15949 ) | ( n15891 & n15989 ) | ( n15949 & n15989 ) ;
  assign n16000 = n15891 | n15989 ;
  assign n16002 = ( n15999 & ~n16001 ) | ( n15999 & n16000 ) | ( ~n16001 & n16000 ) ;
  assign n16006 = n15475 &  n15948 ;
  assign n16007 = n15947 &  n16006 ;
  assign n15995 = x111 | n15475 ;
  assign n15996 = x111 &  n15475 ;
  assign n15997 = ( n15995 & ~n15996 ) | ( n15995 & 1'b0 ) | ( ~n15996 & 1'b0 ) ;
  assign n16009 = ( n15890 & n15949 ) | ( n15890 & n15997 ) | ( n15949 & n15997 ) ;
  assign n16008 = n15890 | n15997 ;
  assign n16010 = ( n16007 & ~n16009 ) | ( n16007 & n16008 ) | ( ~n16009 & n16008 ) ;
  assign n16014 = n15483 &  n15948 ;
  assign n16015 = n15947 &  n16014 ;
  assign n16003 = x110 | n15483 ;
  assign n16004 = x110 &  n15483 ;
  assign n16005 = ( n16003 & ~n16004 ) | ( n16003 & 1'b0 ) | ( ~n16004 & 1'b0 ) ;
  assign n16017 = ( n15889 & n15949 ) | ( n15889 & n16005 ) | ( n15949 & n16005 ) ;
  assign n16016 = n15889 | n16005 ;
  assign n16018 = ( n16015 & ~n16017 ) | ( n16015 & n16016 ) | ( ~n16017 & n16016 ) ;
  assign n16022 = n15491 &  n15948 ;
  assign n16023 = n15947 &  n16022 ;
  assign n16011 = x109 | n15491 ;
  assign n16012 = x109 &  n15491 ;
  assign n16013 = ( n16011 & ~n16012 ) | ( n16011 & 1'b0 ) | ( ~n16012 & 1'b0 ) ;
  assign n16025 = ( n15888 & n15949 ) | ( n15888 & n16013 ) | ( n15949 & n16013 ) ;
  assign n16024 = n15888 | n16013 ;
  assign n16026 = ( n16023 & ~n16025 ) | ( n16023 & n16024 ) | ( ~n16025 & n16024 ) ;
  assign n16030 = n15499 &  n15948 ;
  assign n16031 = n15947 &  n16030 ;
  assign n16019 = x108 | n15499 ;
  assign n16020 = x108 &  n15499 ;
  assign n16021 = ( n16019 & ~n16020 ) | ( n16019 & 1'b0 ) | ( ~n16020 & 1'b0 ) ;
  assign n16033 = ( n15887 & n15949 ) | ( n15887 & n16021 ) | ( n15949 & n16021 ) ;
  assign n16032 = n15887 | n16021 ;
  assign n16034 = ( n16031 & ~n16033 ) | ( n16031 & n16032 ) | ( ~n16033 & n16032 ) ;
  assign n16038 = n15507 &  n15948 ;
  assign n16039 = n15947 &  n16038 ;
  assign n16027 = x107 | n15507 ;
  assign n16028 = x107 &  n15507 ;
  assign n16029 = ( n16027 & ~n16028 ) | ( n16027 & 1'b0 ) | ( ~n16028 & 1'b0 ) ;
  assign n16041 = ( n15886 & n15949 ) | ( n15886 & n16029 ) | ( n15949 & n16029 ) ;
  assign n16040 = n15886 | n16029 ;
  assign n16042 = ( n16039 & ~n16041 ) | ( n16039 & n16040 ) | ( ~n16041 & n16040 ) ;
  assign n16046 = n15515 &  n15948 ;
  assign n16047 = n15947 &  n16046 ;
  assign n16035 = x106 | n15515 ;
  assign n16036 = x106 &  n15515 ;
  assign n16037 = ( n16035 & ~n16036 ) | ( n16035 & 1'b0 ) | ( ~n16036 & 1'b0 ) ;
  assign n16049 = ( n15885 & n15949 ) | ( n15885 & n16037 ) | ( n15949 & n16037 ) ;
  assign n16048 = n15885 | n16037 ;
  assign n16050 = ( n16047 & ~n16049 ) | ( n16047 & n16048 ) | ( ~n16049 & n16048 ) ;
  assign n16054 = n15523 &  n15948 ;
  assign n16055 = n15947 &  n16054 ;
  assign n16043 = x105 | n15523 ;
  assign n16044 = x105 &  n15523 ;
  assign n16045 = ( n16043 & ~n16044 ) | ( n16043 & 1'b0 ) | ( ~n16044 & 1'b0 ) ;
  assign n16057 = ( n15884 & n15949 ) | ( n15884 & n16045 ) | ( n15949 & n16045 ) ;
  assign n16056 = n15884 | n16045 ;
  assign n16058 = ( n16055 & ~n16057 ) | ( n16055 & n16056 ) | ( ~n16057 & n16056 ) ;
  assign n16062 = n15531 &  n15948 ;
  assign n16063 = n15947 &  n16062 ;
  assign n16051 = x104 | n15531 ;
  assign n16052 = x104 &  n15531 ;
  assign n16053 = ( n16051 & ~n16052 ) | ( n16051 & 1'b0 ) | ( ~n16052 & 1'b0 ) ;
  assign n16065 = ( n15883 & n15949 ) | ( n15883 & n16053 ) | ( n15949 & n16053 ) ;
  assign n16064 = n15883 | n16053 ;
  assign n16066 = ( n16063 & ~n16065 ) | ( n16063 & n16064 ) | ( ~n16065 & n16064 ) ;
  assign n16070 = n15539 &  n15948 ;
  assign n16071 = n15947 &  n16070 ;
  assign n16059 = x103 | n15539 ;
  assign n16060 = x103 &  n15539 ;
  assign n16061 = ( n16059 & ~n16060 ) | ( n16059 & 1'b0 ) | ( ~n16060 & 1'b0 ) ;
  assign n16073 = ( n15882 & n15949 ) | ( n15882 & n16061 ) | ( n15949 & n16061 ) ;
  assign n16072 = n15882 | n16061 ;
  assign n16074 = ( n16071 & ~n16073 ) | ( n16071 & n16072 ) | ( ~n16073 & n16072 ) ;
  assign n16078 = n15547 &  n15948 ;
  assign n16079 = n15947 &  n16078 ;
  assign n16067 = x102 | n15547 ;
  assign n16068 = x102 &  n15547 ;
  assign n16069 = ( n16067 & ~n16068 ) | ( n16067 & 1'b0 ) | ( ~n16068 & 1'b0 ) ;
  assign n16081 = ( n15881 & n15949 ) | ( n15881 & n16069 ) | ( n15949 & n16069 ) ;
  assign n16080 = n15881 | n16069 ;
  assign n16082 = ( n16079 & ~n16081 ) | ( n16079 & n16080 ) | ( ~n16081 & n16080 ) ;
  assign n16086 = n15555 &  n15948 ;
  assign n16087 = n15947 &  n16086 ;
  assign n16075 = x101 | n15555 ;
  assign n16076 = x101 &  n15555 ;
  assign n16077 = ( n16075 & ~n16076 ) | ( n16075 & 1'b0 ) | ( ~n16076 & 1'b0 ) ;
  assign n16089 = ( n15880 & n15949 ) | ( n15880 & n16077 ) | ( n15949 & n16077 ) ;
  assign n16088 = n15880 | n16077 ;
  assign n16090 = ( n16087 & ~n16089 ) | ( n16087 & n16088 ) | ( ~n16089 & n16088 ) ;
  assign n16094 = n15563 &  n15948 ;
  assign n16095 = n15947 &  n16094 ;
  assign n16083 = x100 | n15563 ;
  assign n16084 = x100 &  n15563 ;
  assign n16085 = ( n16083 & ~n16084 ) | ( n16083 & 1'b0 ) | ( ~n16084 & 1'b0 ) ;
  assign n16097 = ( n15879 & n15949 ) | ( n15879 & n16085 ) | ( n15949 & n16085 ) ;
  assign n16096 = n15879 | n16085 ;
  assign n16098 = ( n16095 & ~n16097 ) | ( n16095 & n16096 ) | ( ~n16097 & n16096 ) ;
  assign n16102 = n15571 &  n15948 ;
  assign n16103 = n15947 &  n16102 ;
  assign n16091 = x99 | n15571 ;
  assign n16092 = x99 &  n15571 ;
  assign n16093 = ( n16091 & ~n16092 ) | ( n16091 & 1'b0 ) | ( ~n16092 & 1'b0 ) ;
  assign n16105 = ( n15878 & n15949 ) | ( n15878 & n16093 ) | ( n15949 & n16093 ) ;
  assign n16104 = n15878 | n16093 ;
  assign n16106 = ( n16103 & ~n16105 ) | ( n16103 & n16104 ) | ( ~n16105 & n16104 ) ;
  assign n16110 = n15579 &  n15948 ;
  assign n16111 = n15947 &  n16110 ;
  assign n16099 = x98 | n15579 ;
  assign n16100 = x98 &  n15579 ;
  assign n16101 = ( n16099 & ~n16100 ) | ( n16099 & 1'b0 ) | ( ~n16100 & 1'b0 ) ;
  assign n16113 = ( n15877 & n15949 ) | ( n15877 & n16101 ) | ( n15949 & n16101 ) ;
  assign n16112 = n15877 | n16101 ;
  assign n16114 = ( n16111 & ~n16113 ) | ( n16111 & n16112 ) | ( ~n16113 & n16112 ) ;
  assign n16118 = n15587 &  n15948 ;
  assign n16119 = n15947 &  n16118 ;
  assign n16107 = x97 | n15587 ;
  assign n16108 = x97 &  n15587 ;
  assign n16109 = ( n16107 & ~n16108 ) | ( n16107 & 1'b0 ) | ( ~n16108 & 1'b0 ) ;
  assign n16121 = ( n15876 & n15949 ) | ( n15876 & n16109 ) | ( n15949 & n16109 ) ;
  assign n16120 = n15876 | n16109 ;
  assign n16122 = ( n16119 & ~n16121 ) | ( n16119 & n16120 ) | ( ~n16121 & n16120 ) ;
  assign n16126 = n15595 &  n15948 ;
  assign n16127 = n15947 &  n16126 ;
  assign n16115 = x96 | n15595 ;
  assign n16116 = x96 &  n15595 ;
  assign n16117 = ( n16115 & ~n16116 ) | ( n16115 & 1'b0 ) | ( ~n16116 & 1'b0 ) ;
  assign n16129 = ( n15875 & n15949 ) | ( n15875 & n16117 ) | ( n15949 & n16117 ) ;
  assign n16128 = n15875 | n16117 ;
  assign n16130 = ( n16127 & ~n16129 ) | ( n16127 & n16128 ) | ( ~n16129 & n16128 ) ;
  assign n16134 = n15603 &  n15948 ;
  assign n16135 = n15947 &  n16134 ;
  assign n16123 = x95 | n15603 ;
  assign n16124 = x95 &  n15603 ;
  assign n16125 = ( n16123 & ~n16124 ) | ( n16123 & 1'b0 ) | ( ~n16124 & 1'b0 ) ;
  assign n16137 = ( n15874 & n15949 ) | ( n15874 & n16125 ) | ( n15949 & n16125 ) ;
  assign n16136 = n15874 | n16125 ;
  assign n16138 = ( n16135 & ~n16137 ) | ( n16135 & n16136 ) | ( ~n16137 & n16136 ) ;
  assign n16142 = n15611 &  n15948 ;
  assign n16143 = n15947 &  n16142 ;
  assign n16131 = x94 | n15611 ;
  assign n16132 = x94 &  n15611 ;
  assign n16133 = ( n16131 & ~n16132 ) | ( n16131 & 1'b0 ) | ( ~n16132 & 1'b0 ) ;
  assign n16145 = ( n15873 & n15949 ) | ( n15873 & n16133 ) | ( n15949 & n16133 ) ;
  assign n16144 = n15873 | n16133 ;
  assign n16146 = ( n16143 & ~n16145 ) | ( n16143 & n16144 ) | ( ~n16145 & n16144 ) ;
  assign n16150 = n15619 &  n15948 ;
  assign n16151 = n15947 &  n16150 ;
  assign n16139 = x93 | n15619 ;
  assign n16140 = x93 &  n15619 ;
  assign n16141 = ( n16139 & ~n16140 ) | ( n16139 & 1'b0 ) | ( ~n16140 & 1'b0 ) ;
  assign n16153 = ( n15872 & n15949 ) | ( n15872 & n16141 ) | ( n15949 & n16141 ) ;
  assign n16152 = n15872 | n16141 ;
  assign n16154 = ( n16151 & ~n16153 ) | ( n16151 & n16152 ) | ( ~n16153 & n16152 ) ;
  assign n16158 = n15627 &  n15948 ;
  assign n16159 = n15947 &  n16158 ;
  assign n16147 = x92 | n15627 ;
  assign n16148 = x92 &  n15627 ;
  assign n16149 = ( n16147 & ~n16148 ) | ( n16147 & 1'b0 ) | ( ~n16148 & 1'b0 ) ;
  assign n16161 = ( n15871 & n15949 ) | ( n15871 & n16149 ) | ( n15949 & n16149 ) ;
  assign n16160 = n15871 | n16149 ;
  assign n16162 = ( n16159 & ~n16161 ) | ( n16159 & n16160 ) | ( ~n16161 & n16160 ) ;
  assign n16166 = n15635 &  n15948 ;
  assign n16167 = n15947 &  n16166 ;
  assign n16155 = x91 | n15635 ;
  assign n16156 = x91 &  n15635 ;
  assign n16157 = ( n16155 & ~n16156 ) | ( n16155 & 1'b0 ) | ( ~n16156 & 1'b0 ) ;
  assign n16169 = ( n15870 & n15949 ) | ( n15870 & n16157 ) | ( n15949 & n16157 ) ;
  assign n16168 = n15870 | n16157 ;
  assign n16170 = ( n16167 & ~n16169 ) | ( n16167 & n16168 ) | ( ~n16169 & n16168 ) ;
  assign n16174 = n15643 &  n15948 ;
  assign n16175 = n15947 &  n16174 ;
  assign n16163 = x90 | n15643 ;
  assign n16164 = x90 &  n15643 ;
  assign n16165 = ( n16163 & ~n16164 ) | ( n16163 & 1'b0 ) | ( ~n16164 & 1'b0 ) ;
  assign n16177 = ( n15869 & n15949 ) | ( n15869 & n16165 ) | ( n15949 & n16165 ) ;
  assign n16176 = n15869 | n16165 ;
  assign n16178 = ( n16175 & ~n16177 ) | ( n16175 & n16176 ) | ( ~n16177 & n16176 ) ;
  assign n16182 = n15651 &  n15948 ;
  assign n16183 = n15947 &  n16182 ;
  assign n16171 = x89 | n15651 ;
  assign n16172 = x89 &  n15651 ;
  assign n16173 = ( n16171 & ~n16172 ) | ( n16171 & 1'b0 ) | ( ~n16172 & 1'b0 ) ;
  assign n16185 = ( n15868 & n15949 ) | ( n15868 & n16173 ) | ( n15949 & n16173 ) ;
  assign n16184 = n15868 | n16173 ;
  assign n16186 = ( n16183 & ~n16185 ) | ( n16183 & n16184 ) | ( ~n16185 & n16184 ) ;
  assign n16190 = n15659 &  n15948 ;
  assign n16191 = n15947 &  n16190 ;
  assign n16179 = x88 | n15659 ;
  assign n16180 = x88 &  n15659 ;
  assign n16181 = ( n16179 & ~n16180 ) | ( n16179 & 1'b0 ) | ( ~n16180 & 1'b0 ) ;
  assign n16193 = ( n15867 & n15949 ) | ( n15867 & n16181 ) | ( n15949 & n16181 ) ;
  assign n16192 = n15867 | n16181 ;
  assign n16194 = ( n16191 & ~n16193 ) | ( n16191 & n16192 ) | ( ~n16193 & n16192 ) ;
  assign n16198 = n15667 &  n15948 ;
  assign n16199 = n15947 &  n16198 ;
  assign n16187 = x87 | n15667 ;
  assign n16188 = x87 &  n15667 ;
  assign n16189 = ( n16187 & ~n16188 ) | ( n16187 & 1'b0 ) | ( ~n16188 & 1'b0 ) ;
  assign n16201 = ( n15866 & n15949 ) | ( n15866 & n16189 ) | ( n15949 & n16189 ) ;
  assign n16200 = n15866 | n16189 ;
  assign n16202 = ( n16199 & ~n16201 ) | ( n16199 & n16200 ) | ( ~n16201 & n16200 ) ;
  assign n16206 = n15675 &  n15948 ;
  assign n16207 = n15947 &  n16206 ;
  assign n16195 = x86 | n15675 ;
  assign n16196 = x86 &  n15675 ;
  assign n16197 = ( n16195 & ~n16196 ) | ( n16195 & 1'b0 ) | ( ~n16196 & 1'b0 ) ;
  assign n16209 = ( n15865 & n15949 ) | ( n15865 & n16197 ) | ( n15949 & n16197 ) ;
  assign n16208 = n15865 | n16197 ;
  assign n16210 = ( n16207 & ~n16209 ) | ( n16207 & n16208 ) | ( ~n16209 & n16208 ) ;
  assign n16214 = n15683 &  n15948 ;
  assign n16215 = n15947 &  n16214 ;
  assign n16203 = x85 | n15683 ;
  assign n16204 = x85 &  n15683 ;
  assign n16205 = ( n16203 & ~n16204 ) | ( n16203 & 1'b0 ) | ( ~n16204 & 1'b0 ) ;
  assign n16217 = ( n15864 & n15949 ) | ( n15864 & n16205 ) | ( n15949 & n16205 ) ;
  assign n16216 = n15864 | n16205 ;
  assign n16218 = ( n16215 & ~n16217 ) | ( n16215 & n16216 ) | ( ~n16217 & n16216 ) ;
  assign n16222 = n15691 &  n15948 ;
  assign n16223 = n15947 &  n16222 ;
  assign n16211 = x84 | n15691 ;
  assign n16212 = x84 &  n15691 ;
  assign n16213 = ( n16211 & ~n16212 ) | ( n16211 & 1'b0 ) | ( ~n16212 & 1'b0 ) ;
  assign n16225 = ( n15863 & n15949 ) | ( n15863 & n16213 ) | ( n15949 & n16213 ) ;
  assign n16224 = n15863 | n16213 ;
  assign n16226 = ( n16223 & ~n16225 ) | ( n16223 & n16224 ) | ( ~n16225 & n16224 ) ;
  assign n16230 = n15699 &  n15948 ;
  assign n16231 = n15947 &  n16230 ;
  assign n16219 = x83 | n15699 ;
  assign n16220 = x83 &  n15699 ;
  assign n16221 = ( n16219 & ~n16220 ) | ( n16219 & 1'b0 ) | ( ~n16220 & 1'b0 ) ;
  assign n16233 = ( n15862 & n15949 ) | ( n15862 & n16221 ) | ( n15949 & n16221 ) ;
  assign n16232 = n15862 | n16221 ;
  assign n16234 = ( n16231 & ~n16233 ) | ( n16231 & n16232 ) | ( ~n16233 & n16232 ) ;
  assign n16238 = n15707 &  n15948 ;
  assign n16239 = n15947 &  n16238 ;
  assign n16227 = x82 | n15707 ;
  assign n16228 = x82 &  n15707 ;
  assign n16229 = ( n16227 & ~n16228 ) | ( n16227 & 1'b0 ) | ( ~n16228 & 1'b0 ) ;
  assign n16241 = ( n15861 & n15949 ) | ( n15861 & n16229 ) | ( n15949 & n16229 ) ;
  assign n16240 = n15861 | n16229 ;
  assign n16242 = ( n16239 & ~n16241 ) | ( n16239 & n16240 ) | ( ~n16241 & n16240 ) ;
  assign n16246 = n15715 &  n15948 ;
  assign n16247 = n15947 &  n16246 ;
  assign n16235 = x81 | n15715 ;
  assign n16236 = x81 &  n15715 ;
  assign n16237 = ( n16235 & ~n16236 ) | ( n16235 & 1'b0 ) | ( ~n16236 & 1'b0 ) ;
  assign n16249 = ( n15860 & n15949 ) | ( n15860 & n16237 ) | ( n15949 & n16237 ) ;
  assign n16248 = n15860 | n16237 ;
  assign n16250 = ( n16247 & ~n16249 ) | ( n16247 & n16248 ) | ( ~n16249 & n16248 ) ;
  assign n16254 = n15723 &  n15948 ;
  assign n16255 = n15947 &  n16254 ;
  assign n16243 = x80 | n15723 ;
  assign n16244 = x80 &  n15723 ;
  assign n16245 = ( n16243 & ~n16244 ) | ( n16243 & 1'b0 ) | ( ~n16244 & 1'b0 ) ;
  assign n16257 = ( n15859 & n15949 ) | ( n15859 & n16245 ) | ( n15949 & n16245 ) ;
  assign n16256 = n15859 | n16245 ;
  assign n16258 = ( n16255 & ~n16257 ) | ( n16255 & n16256 ) | ( ~n16257 & n16256 ) ;
  assign n16262 = n15731 &  n15948 ;
  assign n16263 = n15947 &  n16262 ;
  assign n16251 = x79 | n15731 ;
  assign n16252 = x79 &  n15731 ;
  assign n16253 = ( n16251 & ~n16252 ) | ( n16251 & 1'b0 ) | ( ~n16252 & 1'b0 ) ;
  assign n16265 = ( n15858 & n15949 ) | ( n15858 & n16253 ) | ( n15949 & n16253 ) ;
  assign n16264 = n15858 | n16253 ;
  assign n16266 = ( n16263 & ~n16265 ) | ( n16263 & n16264 ) | ( ~n16265 & n16264 ) ;
  assign n16270 = n15739 &  n15948 ;
  assign n16271 = n15947 &  n16270 ;
  assign n16259 = x78 | n15739 ;
  assign n16260 = x78 &  n15739 ;
  assign n16261 = ( n16259 & ~n16260 ) | ( n16259 & 1'b0 ) | ( ~n16260 & 1'b0 ) ;
  assign n16273 = ( n15857 & n15949 ) | ( n15857 & n16261 ) | ( n15949 & n16261 ) ;
  assign n16272 = n15857 | n16261 ;
  assign n16274 = ( n16271 & ~n16273 ) | ( n16271 & n16272 ) | ( ~n16273 & n16272 ) ;
  assign n16278 = n15747 &  n15948 ;
  assign n16279 = n15947 &  n16278 ;
  assign n16267 = x77 | n15747 ;
  assign n16268 = x77 &  n15747 ;
  assign n16269 = ( n16267 & ~n16268 ) | ( n16267 & 1'b0 ) | ( ~n16268 & 1'b0 ) ;
  assign n16281 = ( n15856 & n15949 ) | ( n15856 & n16269 ) | ( n15949 & n16269 ) ;
  assign n16280 = n15856 | n16269 ;
  assign n16282 = ( n16279 & ~n16281 ) | ( n16279 & n16280 ) | ( ~n16281 & n16280 ) ;
  assign n16286 = n15755 &  n15948 ;
  assign n16287 = n15947 &  n16286 ;
  assign n16275 = x76 | n15755 ;
  assign n16276 = x76 &  n15755 ;
  assign n16277 = ( n16275 & ~n16276 ) | ( n16275 & 1'b0 ) | ( ~n16276 & 1'b0 ) ;
  assign n16289 = ( n15855 & n15949 ) | ( n15855 & n16277 ) | ( n15949 & n16277 ) ;
  assign n16288 = n15855 | n16277 ;
  assign n16290 = ( n16287 & ~n16289 ) | ( n16287 & n16288 ) | ( ~n16289 & n16288 ) ;
  assign n16294 = n15763 &  n15948 ;
  assign n16295 = n15947 &  n16294 ;
  assign n16283 = x75 | n15763 ;
  assign n16284 = x75 &  n15763 ;
  assign n16285 = ( n16283 & ~n16284 ) | ( n16283 & 1'b0 ) | ( ~n16284 & 1'b0 ) ;
  assign n16297 = ( n15854 & n15949 ) | ( n15854 & n16285 ) | ( n15949 & n16285 ) ;
  assign n16296 = n15854 | n16285 ;
  assign n16298 = ( n16295 & ~n16297 ) | ( n16295 & n16296 ) | ( ~n16297 & n16296 ) ;
  assign n16302 = n15771 &  n15948 ;
  assign n16303 = n15947 &  n16302 ;
  assign n16291 = x74 | n15771 ;
  assign n16292 = x74 &  n15771 ;
  assign n16293 = ( n16291 & ~n16292 ) | ( n16291 & 1'b0 ) | ( ~n16292 & 1'b0 ) ;
  assign n16305 = ( n15853 & n15949 ) | ( n15853 & n16293 ) | ( n15949 & n16293 ) ;
  assign n16304 = n15853 | n16293 ;
  assign n16306 = ( n16303 & ~n16305 ) | ( n16303 & n16304 ) | ( ~n16305 & n16304 ) ;
  assign n16310 = n15779 &  n15948 ;
  assign n16311 = n15947 &  n16310 ;
  assign n16299 = x73 | n15779 ;
  assign n16300 = x73 &  n15779 ;
  assign n16301 = ( n16299 & ~n16300 ) | ( n16299 & 1'b0 ) | ( ~n16300 & 1'b0 ) ;
  assign n16313 = ( n15852 & n15949 ) | ( n15852 & n16301 ) | ( n15949 & n16301 ) ;
  assign n16312 = n15852 | n16301 ;
  assign n16314 = ( n16311 & ~n16313 ) | ( n16311 & n16312 ) | ( ~n16313 & n16312 ) ;
  assign n16318 = n15787 &  n15948 ;
  assign n16319 = n15947 &  n16318 ;
  assign n16307 = x72 | n15787 ;
  assign n16308 = x72 &  n15787 ;
  assign n16309 = ( n16307 & ~n16308 ) | ( n16307 & 1'b0 ) | ( ~n16308 & 1'b0 ) ;
  assign n16321 = ( n15851 & n15949 ) | ( n15851 & n16309 ) | ( n15949 & n16309 ) ;
  assign n16320 = n15851 | n16309 ;
  assign n16322 = ( n16319 & ~n16321 ) | ( n16319 & n16320 ) | ( ~n16321 & n16320 ) ;
  assign n16326 = n15795 &  n15948 ;
  assign n16327 = n15947 &  n16326 ;
  assign n16315 = x71 | n15795 ;
  assign n16316 = x71 &  n15795 ;
  assign n16317 = ( n16315 & ~n16316 ) | ( n16315 & 1'b0 ) | ( ~n16316 & 1'b0 ) ;
  assign n16329 = ( n15850 & n15949 ) | ( n15850 & n16317 ) | ( n15949 & n16317 ) ;
  assign n16328 = n15850 | n16317 ;
  assign n16330 = ( n16327 & ~n16329 ) | ( n16327 & n16328 ) | ( ~n16329 & n16328 ) ;
  assign n16334 = n15803 &  n15948 ;
  assign n16335 = n15947 &  n16334 ;
  assign n16323 = x70 | n15803 ;
  assign n16324 = x70 &  n15803 ;
  assign n16325 = ( n16323 & ~n16324 ) | ( n16323 & 1'b0 ) | ( ~n16324 & 1'b0 ) ;
  assign n16337 = ( n15849 & n15949 ) | ( n15849 & n16325 ) | ( n15949 & n16325 ) ;
  assign n16336 = n15849 | n16325 ;
  assign n16338 = ( n16335 & ~n16337 ) | ( n16335 & n16336 ) | ( ~n16337 & n16336 ) ;
  assign n16342 = n15811 &  n15948 ;
  assign n16343 = n15947 &  n16342 ;
  assign n16331 = x69 | n15811 ;
  assign n16332 = x69 &  n15811 ;
  assign n16333 = ( n16331 & ~n16332 ) | ( n16331 & 1'b0 ) | ( ~n16332 & 1'b0 ) ;
  assign n16345 = ( n15848 & n15949 ) | ( n15848 & n16333 ) | ( n15949 & n16333 ) ;
  assign n16344 = n15848 | n16333 ;
  assign n16346 = ( n16343 & ~n16345 ) | ( n16343 & n16344 ) | ( ~n16345 & n16344 ) ;
  assign n16350 = n15819 &  n15948 ;
  assign n16351 = n15947 &  n16350 ;
  assign n16339 = x68 | n15819 ;
  assign n16340 = x68 &  n15819 ;
  assign n16341 = ( n16339 & ~n16340 ) | ( n16339 & 1'b0 ) | ( ~n16340 & 1'b0 ) ;
  assign n16353 = ( n15847 & n15949 ) | ( n15847 & n16341 ) | ( n15949 & n16341 ) ;
  assign n16352 = n15847 | n16341 ;
  assign n16354 = ( n16351 & ~n16353 ) | ( n16351 & n16352 ) | ( ~n16353 & n16352 ) ;
  assign n16358 = n15828 &  n15948 ;
  assign n16359 = n15947 &  n16358 ;
  assign n16347 = x67 | n15828 ;
  assign n16348 = x67 &  n15828 ;
  assign n16349 = ( n16347 & ~n16348 ) | ( n16347 & 1'b0 ) | ( ~n16348 & 1'b0 ) ;
  assign n16361 = ( n15846 & n15949 ) | ( n15846 & n16349 ) | ( n15949 & n16349 ) ;
  assign n16360 = n15846 | n16349 ;
  assign n16362 = ( n16359 & ~n16361 ) | ( n16359 & n16360 ) | ( ~n16361 & n16360 ) ;
  assign n16363 = n15834 &  n15948 ;
  assign n16364 = n15947 &  n16363 ;
  assign n16355 = x66 | n15834 ;
  assign n16356 = x66 &  n15834 ;
  assign n16357 = ( n16355 & ~n16356 ) | ( n16355 & 1'b0 ) | ( ~n16356 & 1'b0 ) ;
  assign n16365 = n15845 &  n16357 ;
  assign n16366 = ( n15845 & ~n15949 ) | ( n15845 & n16357 ) | ( ~n15949 & n16357 ) ;
  assign n16367 = ( n16364 & ~n16365 ) | ( n16364 & n16366 ) | ( ~n16365 & n16366 ) ;
  assign n16368 = ( n15843 & ~x65 ) | ( n15843 & n15844 ) | ( ~x65 & n15844 ) ;
  assign n16369 = ( n15845 & ~n15844 ) | ( n15845 & n16368 ) | ( ~n15844 & n16368 ) ;
  assign n16370 = ~n15949 & n16369 ;
  assign n16371 = n15843 &  n15948 ;
  assign n16372 = n15947 &  n16371 ;
  assign n16373 = n16370 | n16372 ;
  assign n16374 = ( x64 & ~n15949 ) | ( x64 & 1'b0 ) | ( ~n15949 & 1'b0 ) ;
  assign n16375 = ( x5 & ~n16374 ) | ( x5 & 1'b0 ) | ( ~n16374 & 1'b0 ) ;
  assign n16376 = ( n15844 & ~n15949 ) | ( n15844 & 1'b0 ) | ( ~n15949 & 1'b0 ) ;
  assign n16377 = n16375 | n16376 ;
  assign n16378 = ~x4 & x64 ;
  assign n16379 = ( x65 & ~n16377 ) | ( x65 & n16378 ) | ( ~n16377 & n16378 ) ;
  assign n16380 = ( x66 & ~n16373 ) | ( x66 & n16379 ) | ( ~n16373 & n16379 ) ;
  assign n16381 = ( x67 & ~n16367 ) | ( x67 & n16380 ) | ( ~n16367 & n16380 ) ;
  assign n16382 = ( x68 & ~n16362 ) | ( x68 & n16381 ) | ( ~n16362 & n16381 ) ;
  assign n16383 = ( x69 & ~n16354 ) | ( x69 & n16382 ) | ( ~n16354 & n16382 ) ;
  assign n16384 = ( x70 & ~n16346 ) | ( x70 & n16383 ) | ( ~n16346 & n16383 ) ;
  assign n16385 = ( x71 & ~n16338 ) | ( x71 & n16384 ) | ( ~n16338 & n16384 ) ;
  assign n16386 = ( x72 & ~n16330 ) | ( x72 & n16385 ) | ( ~n16330 & n16385 ) ;
  assign n16387 = ( x73 & ~n16322 ) | ( x73 & n16386 ) | ( ~n16322 & n16386 ) ;
  assign n16388 = ( x74 & ~n16314 ) | ( x74 & n16387 ) | ( ~n16314 & n16387 ) ;
  assign n16389 = ( x75 & ~n16306 ) | ( x75 & n16388 ) | ( ~n16306 & n16388 ) ;
  assign n16390 = ( x76 & ~n16298 ) | ( x76 & n16389 ) | ( ~n16298 & n16389 ) ;
  assign n16391 = ( x77 & ~n16290 ) | ( x77 & n16390 ) | ( ~n16290 & n16390 ) ;
  assign n16392 = ( x78 & ~n16282 ) | ( x78 & n16391 ) | ( ~n16282 & n16391 ) ;
  assign n16393 = ( x79 & ~n16274 ) | ( x79 & n16392 ) | ( ~n16274 & n16392 ) ;
  assign n16394 = ( x80 & ~n16266 ) | ( x80 & n16393 ) | ( ~n16266 & n16393 ) ;
  assign n16395 = ( x81 & ~n16258 ) | ( x81 & n16394 ) | ( ~n16258 & n16394 ) ;
  assign n16396 = ( x82 & ~n16250 ) | ( x82 & n16395 ) | ( ~n16250 & n16395 ) ;
  assign n16397 = ( x83 & ~n16242 ) | ( x83 & n16396 ) | ( ~n16242 & n16396 ) ;
  assign n16398 = ( x84 & ~n16234 ) | ( x84 & n16397 ) | ( ~n16234 & n16397 ) ;
  assign n16399 = ( x85 & ~n16226 ) | ( x85 & n16398 ) | ( ~n16226 & n16398 ) ;
  assign n16400 = ( x86 & ~n16218 ) | ( x86 & n16399 ) | ( ~n16218 & n16399 ) ;
  assign n16401 = ( x87 & ~n16210 ) | ( x87 & n16400 ) | ( ~n16210 & n16400 ) ;
  assign n16402 = ( x88 & ~n16202 ) | ( x88 & n16401 ) | ( ~n16202 & n16401 ) ;
  assign n16403 = ( x89 & ~n16194 ) | ( x89 & n16402 ) | ( ~n16194 & n16402 ) ;
  assign n16404 = ( x90 & ~n16186 ) | ( x90 & n16403 ) | ( ~n16186 & n16403 ) ;
  assign n16405 = ( x91 & ~n16178 ) | ( x91 & n16404 ) | ( ~n16178 & n16404 ) ;
  assign n16406 = ( x92 & ~n16170 ) | ( x92 & n16405 ) | ( ~n16170 & n16405 ) ;
  assign n16407 = ( x93 & ~n16162 ) | ( x93 & n16406 ) | ( ~n16162 & n16406 ) ;
  assign n16408 = ( x94 & ~n16154 ) | ( x94 & n16407 ) | ( ~n16154 & n16407 ) ;
  assign n16409 = ( x95 & ~n16146 ) | ( x95 & n16408 ) | ( ~n16146 & n16408 ) ;
  assign n16410 = ( x96 & ~n16138 ) | ( x96 & n16409 ) | ( ~n16138 & n16409 ) ;
  assign n16411 = ( x97 & ~n16130 ) | ( x97 & n16410 ) | ( ~n16130 & n16410 ) ;
  assign n16412 = ( x98 & ~n16122 ) | ( x98 & n16411 ) | ( ~n16122 & n16411 ) ;
  assign n16413 = ( x99 & ~n16114 ) | ( x99 & n16412 ) | ( ~n16114 & n16412 ) ;
  assign n16414 = ( x100 & ~n16106 ) | ( x100 & n16413 ) | ( ~n16106 & n16413 ) ;
  assign n16415 = ( x101 & ~n16098 ) | ( x101 & n16414 ) | ( ~n16098 & n16414 ) ;
  assign n16416 = ( x102 & ~n16090 ) | ( x102 & n16415 ) | ( ~n16090 & n16415 ) ;
  assign n16417 = ( x103 & ~n16082 ) | ( x103 & n16416 ) | ( ~n16082 & n16416 ) ;
  assign n16418 = ( x104 & ~n16074 ) | ( x104 & n16417 ) | ( ~n16074 & n16417 ) ;
  assign n16419 = ( x105 & ~n16066 ) | ( x105 & n16418 ) | ( ~n16066 & n16418 ) ;
  assign n16420 = ( x106 & ~n16058 ) | ( x106 & n16419 ) | ( ~n16058 & n16419 ) ;
  assign n16421 = ( x107 & ~n16050 ) | ( x107 & n16420 ) | ( ~n16050 & n16420 ) ;
  assign n16422 = ( x108 & ~n16042 ) | ( x108 & n16421 ) | ( ~n16042 & n16421 ) ;
  assign n16423 = ( x109 & ~n16034 ) | ( x109 & n16422 ) | ( ~n16034 & n16422 ) ;
  assign n16424 = ( x110 & ~n16026 ) | ( x110 & n16423 ) | ( ~n16026 & n16423 ) ;
  assign n16425 = ( x111 & ~n16018 ) | ( x111 & n16424 ) | ( ~n16018 & n16424 ) ;
  assign n16426 = ( x112 & ~n16010 ) | ( x112 & n16425 ) | ( ~n16010 & n16425 ) ;
  assign n16427 = ( x113 & ~n16002 ) | ( x113 & n16426 ) | ( ~n16002 & n16426 ) ;
  assign n16428 = ( x114 & ~n15994 ) | ( x114 & n16427 ) | ( ~n15994 & n16427 ) ;
  assign n16429 = ( x115 & ~n15986 ) | ( x115 & n16428 ) | ( ~n15986 & n16428 ) ;
  assign n16430 = ( x116 & ~n15978 ) | ( x116 & n16429 ) | ( ~n15978 & n16429 ) ;
  assign n16431 = ( x117 & ~n15970 ) | ( x117 & n16430 ) | ( ~n15970 & n16430 ) ;
  assign n16432 = ( x118 & ~n15962 ) | ( x118 & n16431 ) | ( ~n15962 & n16431 ) ;
  assign n16436 = ( x119 & ~n15954 ) | ( x119 & n16432 ) | ( ~n15954 & n16432 ) ;
  assign n16464 = ( x120 & ~n16444 ) | ( x120 & n16436 ) | ( ~n16444 & n16436 ) ;
  assign n16465 = ( x121 & ~n16463 ) | ( x121 & n16464 ) | ( ~n16463 & n16464 ) ;
  assign n16466 = ( x122 & ~n16458 ) | ( x122 & n16465 ) | ( ~n16458 & n16465 ) ;
  assign n16468 = ( x122 & n15939 ) | ( x122 & n15942 ) | ( n15939 & n15942 ) ;
  assign n16467 = ( x122 & ~n15939 ) | ( x122 & n15942 ) | ( ~n15939 & n15942 ) ;
  assign n16469 = ( n15939 & ~n16468 ) | ( n15939 & n16467 ) | ( ~n16468 & n16467 ) ;
  assign n16470 = ~n15949 & n16469 ;
  assign n16471 = n14928 &  n15415 ;
  assign n16472 = n15947 &  n16471 ;
  assign n16473 = n16470 | n16472 ;
  assign n16474 = ~x123 & n16473 ;
  assign n16475 = ( x123 & ~n16472 ) | ( x123 & 1'b0 ) | ( ~n16472 & 1'b0 ) ;
  assign n16476 = ~n16470 & n16475 ;
  assign n16477 = n152 | n16476 ;
  assign n16478 = n16474 | n16477 ;
  assign n16479 = n16466 | n16478 ;
  assign n16480 = ~n16473 |  n15943 ;
  assign n17001 = n16458 &  n16480 ;
  assign n17002 = n16479 &  n17001 ;
  assign n16998 = x122 | n16458 ;
  assign n16999 = x122 &  n16458 ;
  assign n17000 = ( n16998 & ~n16999 ) | ( n16998 & 1'b0 ) | ( ~n16999 & 1'b0 ) ;
  assign n17003 = n16465 &  n17000 ;
  assign n16481 = n16479 &  n16480 ;
  assign n17004 = ( n16465 & ~n16481 ) | ( n16465 & n17000 ) | ( ~n16481 & n17000 ) ;
  assign n17005 = ( n17002 & ~n17003 ) | ( n17002 & n17004 ) | ( ~n17003 & n17004 ) ;
  assign n16990 = n16463 &  n16480 ;
  assign n16991 = n16479 &  n16990 ;
  assign n16987 = x121 | n16463 ;
  assign n16988 = x121 &  n16463 ;
  assign n16989 = ( n16987 & ~n16988 ) | ( n16987 & 1'b0 ) | ( ~n16988 & 1'b0 ) ;
  assign n16992 = n16464 &  n16989 ;
  assign n16993 = ( n16464 & ~n16481 ) | ( n16464 & n16989 ) | ( ~n16481 & n16989 ) ;
  assign n16994 = ( n16991 & ~n16992 ) | ( n16991 & n16993 ) | ( ~n16992 & n16993 ) ;
  assign n16482 = n16444 &  n16480 ;
  assign n16483 = n16479 &  n16482 ;
  assign n16445 = x120 | n16444 ;
  assign n16446 = x120 &  n16444 ;
  assign n16447 = ( n16445 & ~n16446 ) | ( n16445 & 1'b0 ) | ( ~n16446 & 1'b0 ) ;
  assign n16484 = n16436 &  n16447 ;
  assign n16485 = ( n16436 & ~n16481 ) | ( n16436 & n16447 ) | ( ~n16481 & n16447 ) ;
  assign n16486 = ( n16483 & ~n16484 ) | ( n16483 & n16485 ) | ( ~n16484 & n16485 ) ;
  assign n16490 = n15954 &  n16480 ;
  assign n16491 = n16479 &  n16490 ;
  assign n16433 = x119 | n15954 ;
  assign n16434 = x119 &  n15954 ;
  assign n16435 = ( n16433 & ~n16434 ) | ( n16433 & 1'b0 ) | ( ~n16434 & 1'b0 ) ;
  assign n16493 = ( n16432 & n16435 ) | ( n16432 & n16481 ) | ( n16435 & n16481 ) ;
  assign n16492 = n16432 | n16435 ;
  assign n16494 = ( n16491 & ~n16493 ) | ( n16491 & n16492 ) | ( ~n16493 & n16492 ) ;
  assign n16498 = n15962 &  n16480 ;
  assign n16499 = n16479 &  n16498 ;
  assign n16487 = x118 | n15962 ;
  assign n16488 = x118 &  n15962 ;
  assign n16489 = ( n16487 & ~n16488 ) | ( n16487 & 1'b0 ) | ( ~n16488 & 1'b0 ) ;
  assign n16500 = n16431 &  n16489 ;
  assign n16501 = ( n16431 & ~n16481 ) | ( n16431 & n16489 ) | ( ~n16481 & n16489 ) ;
  assign n16502 = ( n16499 & ~n16500 ) | ( n16499 & n16501 ) | ( ~n16500 & n16501 ) ;
  assign n16506 = n15970 &  n16480 ;
  assign n16507 = n16479 &  n16506 ;
  assign n16495 = x117 | n15970 ;
  assign n16496 = x117 &  n15970 ;
  assign n16497 = ( n16495 & ~n16496 ) | ( n16495 & 1'b0 ) | ( ~n16496 & 1'b0 ) ;
  assign n16509 = ( n16430 & n16481 ) | ( n16430 & n16497 ) | ( n16481 & n16497 ) ;
  assign n16508 = n16430 | n16497 ;
  assign n16510 = ( n16507 & ~n16509 ) | ( n16507 & n16508 ) | ( ~n16509 & n16508 ) ;
  assign n16514 = n15978 &  n16480 ;
  assign n16515 = n16479 &  n16514 ;
  assign n16503 = x116 | n15978 ;
  assign n16504 = x116 &  n15978 ;
  assign n16505 = ( n16503 & ~n16504 ) | ( n16503 & 1'b0 ) | ( ~n16504 & 1'b0 ) ;
  assign n16517 = ( n16429 & n16481 ) | ( n16429 & n16505 ) | ( n16481 & n16505 ) ;
  assign n16516 = n16429 | n16505 ;
  assign n16518 = ( n16515 & ~n16517 ) | ( n16515 & n16516 ) | ( ~n16517 & n16516 ) ;
  assign n16522 = n15986 &  n16480 ;
  assign n16523 = n16479 &  n16522 ;
  assign n16511 = x115 | n15986 ;
  assign n16512 = x115 &  n15986 ;
  assign n16513 = ( n16511 & ~n16512 ) | ( n16511 & 1'b0 ) | ( ~n16512 & 1'b0 ) ;
  assign n16525 = ( n16428 & n16481 ) | ( n16428 & n16513 ) | ( n16481 & n16513 ) ;
  assign n16524 = n16428 | n16513 ;
  assign n16526 = ( n16523 & ~n16525 ) | ( n16523 & n16524 ) | ( ~n16525 & n16524 ) ;
  assign n16530 = n15994 &  n16480 ;
  assign n16531 = n16479 &  n16530 ;
  assign n16519 = x114 | n15994 ;
  assign n16520 = x114 &  n15994 ;
  assign n16521 = ( n16519 & ~n16520 ) | ( n16519 & 1'b0 ) | ( ~n16520 & 1'b0 ) ;
  assign n16533 = ( n16427 & n16481 ) | ( n16427 & n16521 ) | ( n16481 & n16521 ) ;
  assign n16532 = n16427 | n16521 ;
  assign n16534 = ( n16531 & ~n16533 ) | ( n16531 & n16532 ) | ( ~n16533 & n16532 ) ;
  assign n16538 = n16002 &  n16480 ;
  assign n16539 = n16479 &  n16538 ;
  assign n16527 = x113 | n16002 ;
  assign n16528 = x113 &  n16002 ;
  assign n16529 = ( n16527 & ~n16528 ) | ( n16527 & 1'b0 ) | ( ~n16528 & 1'b0 ) ;
  assign n16541 = ( n16426 & n16481 ) | ( n16426 & n16529 ) | ( n16481 & n16529 ) ;
  assign n16540 = n16426 | n16529 ;
  assign n16542 = ( n16539 & ~n16541 ) | ( n16539 & n16540 ) | ( ~n16541 & n16540 ) ;
  assign n16546 = n16010 &  n16480 ;
  assign n16547 = n16479 &  n16546 ;
  assign n16535 = x112 | n16010 ;
  assign n16536 = x112 &  n16010 ;
  assign n16537 = ( n16535 & ~n16536 ) | ( n16535 & 1'b0 ) | ( ~n16536 & 1'b0 ) ;
  assign n16549 = ( n16425 & n16481 ) | ( n16425 & n16537 ) | ( n16481 & n16537 ) ;
  assign n16548 = n16425 | n16537 ;
  assign n16550 = ( n16547 & ~n16549 ) | ( n16547 & n16548 ) | ( ~n16549 & n16548 ) ;
  assign n16554 = n16018 &  n16480 ;
  assign n16555 = n16479 &  n16554 ;
  assign n16543 = x111 | n16018 ;
  assign n16544 = x111 &  n16018 ;
  assign n16545 = ( n16543 & ~n16544 ) | ( n16543 & 1'b0 ) | ( ~n16544 & 1'b0 ) ;
  assign n16557 = ( n16424 & n16481 ) | ( n16424 & n16545 ) | ( n16481 & n16545 ) ;
  assign n16556 = n16424 | n16545 ;
  assign n16558 = ( n16555 & ~n16557 ) | ( n16555 & n16556 ) | ( ~n16557 & n16556 ) ;
  assign n16562 = n16026 &  n16480 ;
  assign n16563 = n16479 &  n16562 ;
  assign n16551 = x110 | n16026 ;
  assign n16552 = x110 &  n16026 ;
  assign n16553 = ( n16551 & ~n16552 ) | ( n16551 & 1'b0 ) | ( ~n16552 & 1'b0 ) ;
  assign n16565 = ( n16423 & n16481 ) | ( n16423 & n16553 ) | ( n16481 & n16553 ) ;
  assign n16564 = n16423 | n16553 ;
  assign n16566 = ( n16563 & ~n16565 ) | ( n16563 & n16564 ) | ( ~n16565 & n16564 ) ;
  assign n16570 = n16034 &  n16480 ;
  assign n16571 = n16479 &  n16570 ;
  assign n16559 = x109 | n16034 ;
  assign n16560 = x109 &  n16034 ;
  assign n16561 = ( n16559 & ~n16560 ) | ( n16559 & 1'b0 ) | ( ~n16560 & 1'b0 ) ;
  assign n16573 = ( n16422 & n16481 ) | ( n16422 & n16561 ) | ( n16481 & n16561 ) ;
  assign n16572 = n16422 | n16561 ;
  assign n16574 = ( n16571 & ~n16573 ) | ( n16571 & n16572 ) | ( ~n16573 & n16572 ) ;
  assign n16578 = n16042 &  n16480 ;
  assign n16579 = n16479 &  n16578 ;
  assign n16567 = x108 | n16042 ;
  assign n16568 = x108 &  n16042 ;
  assign n16569 = ( n16567 & ~n16568 ) | ( n16567 & 1'b0 ) | ( ~n16568 & 1'b0 ) ;
  assign n16581 = ( n16421 & n16481 ) | ( n16421 & n16569 ) | ( n16481 & n16569 ) ;
  assign n16580 = n16421 | n16569 ;
  assign n16582 = ( n16579 & ~n16581 ) | ( n16579 & n16580 ) | ( ~n16581 & n16580 ) ;
  assign n16586 = n16050 &  n16480 ;
  assign n16587 = n16479 &  n16586 ;
  assign n16575 = x107 | n16050 ;
  assign n16576 = x107 &  n16050 ;
  assign n16577 = ( n16575 & ~n16576 ) | ( n16575 & 1'b0 ) | ( ~n16576 & 1'b0 ) ;
  assign n16589 = ( n16420 & n16481 ) | ( n16420 & n16577 ) | ( n16481 & n16577 ) ;
  assign n16588 = n16420 | n16577 ;
  assign n16590 = ( n16587 & ~n16589 ) | ( n16587 & n16588 ) | ( ~n16589 & n16588 ) ;
  assign n16594 = n16058 &  n16480 ;
  assign n16595 = n16479 &  n16594 ;
  assign n16583 = x106 | n16058 ;
  assign n16584 = x106 &  n16058 ;
  assign n16585 = ( n16583 & ~n16584 ) | ( n16583 & 1'b0 ) | ( ~n16584 & 1'b0 ) ;
  assign n16597 = ( n16419 & n16481 ) | ( n16419 & n16585 ) | ( n16481 & n16585 ) ;
  assign n16596 = n16419 | n16585 ;
  assign n16598 = ( n16595 & ~n16597 ) | ( n16595 & n16596 ) | ( ~n16597 & n16596 ) ;
  assign n16602 = n16066 &  n16480 ;
  assign n16603 = n16479 &  n16602 ;
  assign n16591 = x105 | n16066 ;
  assign n16592 = x105 &  n16066 ;
  assign n16593 = ( n16591 & ~n16592 ) | ( n16591 & 1'b0 ) | ( ~n16592 & 1'b0 ) ;
  assign n16605 = ( n16418 & n16481 ) | ( n16418 & n16593 ) | ( n16481 & n16593 ) ;
  assign n16604 = n16418 | n16593 ;
  assign n16606 = ( n16603 & ~n16605 ) | ( n16603 & n16604 ) | ( ~n16605 & n16604 ) ;
  assign n16610 = n16074 &  n16480 ;
  assign n16611 = n16479 &  n16610 ;
  assign n16599 = x104 | n16074 ;
  assign n16600 = x104 &  n16074 ;
  assign n16601 = ( n16599 & ~n16600 ) | ( n16599 & 1'b0 ) | ( ~n16600 & 1'b0 ) ;
  assign n16613 = ( n16417 & n16481 ) | ( n16417 & n16601 ) | ( n16481 & n16601 ) ;
  assign n16612 = n16417 | n16601 ;
  assign n16614 = ( n16611 & ~n16613 ) | ( n16611 & n16612 ) | ( ~n16613 & n16612 ) ;
  assign n16618 = n16082 &  n16480 ;
  assign n16619 = n16479 &  n16618 ;
  assign n16607 = x103 | n16082 ;
  assign n16608 = x103 &  n16082 ;
  assign n16609 = ( n16607 & ~n16608 ) | ( n16607 & 1'b0 ) | ( ~n16608 & 1'b0 ) ;
  assign n16621 = ( n16416 & n16481 ) | ( n16416 & n16609 ) | ( n16481 & n16609 ) ;
  assign n16620 = n16416 | n16609 ;
  assign n16622 = ( n16619 & ~n16621 ) | ( n16619 & n16620 ) | ( ~n16621 & n16620 ) ;
  assign n16626 = n16090 &  n16480 ;
  assign n16627 = n16479 &  n16626 ;
  assign n16615 = x102 | n16090 ;
  assign n16616 = x102 &  n16090 ;
  assign n16617 = ( n16615 & ~n16616 ) | ( n16615 & 1'b0 ) | ( ~n16616 & 1'b0 ) ;
  assign n16629 = ( n16415 & n16481 ) | ( n16415 & n16617 ) | ( n16481 & n16617 ) ;
  assign n16628 = n16415 | n16617 ;
  assign n16630 = ( n16627 & ~n16629 ) | ( n16627 & n16628 ) | ( ~n16629 & n16628 ) ;
  assign n16634 = n16098 &  n16480 ;
  assign n16635 = n16479 &  n16634 ;
  assign n16623 = x101 | n16098 ;
  assign n16624 = x101 &  n16098 ;
  assign n16625 = ( n16623 & ~n16624 ) | ( n16623 & 1'b0 ) | ( ~n16624 & 1'b0 ) ;
  assign n16637 = ( n16414 & n16481 ) | ( n16414 & n16625 ) | ( n16481 & n16625 ) ;
  assign n16636 = n16414 | n16625 ;
  assign n16638 = ( n16635 & ~n16637 ) | ( n16635 & n16636 ) | ( ~n16637 & n16636 ) ;
  assign n16642 = n16106 &  n16480 ;
  assign n16643 = n16479 &  n16642 ;
  assign n16631 = x100 | n16106 ;
  assign n16632 = x100 &  n16106 ;
  assign n16633 = ( n16631 & ~n16632 ) | ( n16631 & 1'b0 ) | ( ~n16632 & 1'b0 ) ;
  assign n16645 = ( n16413 & n16481 ) | ( n16413 & n16633 ) | ( n16481 & n16633 ) ;
  assign n16644 = n16413 | n16633 ;
  assign n16646 = ( n16643 & ~n16645 ) | ( n16643 & n16644 ) | ( ~n16645 & n16644 ) ;
  assign n16650 = n16114 &  n16480 ;
  assign n16651 = n16479 &  n16650 ;
  assign n16639 = x99 | n16114 ;
  assign n16640 = x99 &  n16114 ;
  assign n16641 = ( n16639 & ~n16640 ) | ( n16639 & 1'b0 ) | ( ~n16640 & 1'b0 ) ;
  assign n16653 = ( n16412 & n16481 ) | ( n16412 & n16641 ) | ( n16481 & n16641 ) ;
  assign n16652 = n16412 | n16641 ;
  assign n16654 = ( n16651 & ~n16653 ) | ( n16651 & n16652 ) | ( ~n16653 & n16652 ) ;
  assign n16658 = n16122 &  n16480 ;
  assign n16659 = n16479 &  n16658 ;
  assign n16647 = x98 | n16122 ;
  assign n16648 = x98 &  n16122 ;
  assign n16649 = ( n16647 & ~n16648 ) | ( n16647 & 1'b0 ) | ( ~n16648 & 1'b0 ) ;
  assign n16661 = ( n16411 & n16481 ) | ( n16411 & n16649 ) | ( n16481 & n16649 ) ;
  assign n16660 = n16411 | n16649 ;
  assign n16662 = ( n16659 & ~n16661 ) | ( n16659 & n16660 ) | ( ~n16661 & n16660 ) ;
  assign n16666 = n16130 &  n16480 ;
  assign n16667 = n16479 &  n16666 ;
  assign n16655 = x97 | n16130 ;
  assign n16656 = x97 &  n16130 ;
  assign n16657 = ( n16655 & ~n16656 ) | ( n16655 & 1'b0 ) | ( ~n16656 & 1'b0 ) ;
  assign n16669 = ( n16410 & n16481 ) | ( n16410 & n16657 ) | ( n16481 & n16657 ) ;
  assign n16668 = n16410 | n16657 ;
  assign n16670 = ( n16667 & ~n16669 ) | ( n16667 & n16668 ) | ( ~n16669 & n16668 ) ;
  assign n16674 = n16138 &  n16480 ;
  assign n16675 = n16479 &  n16674 ;
  assign n16663 = x96 | n16138 ;
  assign n16664 = x96 &  n16138 ;
  assign n16665 = ( n16663 & ~n16664 ) | ( n16663 & 1'b0 ) | ( ~n16664 & 1'b0 ) ;
  assign n16677 = ( n16409 & n16481 ) | ( n16409 & n16665 ) | ( n16481 & n16665 ) ;
  assign n16676 = n16409 | n16665 ;
  assign n16678 = ( n16675 & ~n16677 ) | ( n16675 & n16676 ) | ( ~n16677 & n16676 ) ;
  assign n16682 = n16146 &  n16480 ;
  assign n16683 = n16479 &  n16682 ;
  assign n16671 = x95 | n16146 ;
  assign n16672 = x95 &  n16146 ;
  assign n16673 = ( n16671 & ~n16672 ) | ( n16671 & 1'b0 ) | ( ~n16672 & 1'b0 ) ;
  assign n16685 = ( n16408 & n16481 ) | ( n16408 & n16673 ) | ( n16481 & n16673 ) ;
  assign n16684 = n16408 | n16673 ;
  assign n16686 = ( n16683 & ~n16685 ) | ( n16683 & n16684 ) | ( ~n16685 & n16684 ) ;
  assign n16690 = n16154 &  n16480 ;
  assign n16691 = n16479 &  n16690 ;
  assign n16679 = x94 | n16154 ;
  assign n16680 = x94 &  n16154 ;
  assign n16681 = ( n16679 & ~n16680 ) | ( n16679 & 1'b0 ) | ( ~n16680 & 1'b0 ) ;
  assign n16693 = ( n16407 & n16481 ) | ( n16407 & n16681 ) | ( n16481 & n16681 ) ;
  assign n16692 = n16407 | n16681 ;
  assign n16694 = ( n16691 & ~n16693 ) | ( n16691 & n16692 ) | ( ~n16693 & n16692 ) ;
  assign n16698 = n16162 &  n16480 ;
  assign n16699 = n16479 &  n16698 ;
  assign n16687 = x93 | n16162 ;
  assign n16688 = x93 &  n16162 ;
  assign n16689 = ( n16687 & ~n16688 ) | ( n16687 & 1'b0 ) | ( ~n16688 & 1'b0 ) ;
  assign n16701 = ( n16406 & n16481 ) | ( n16406 & n16689 ) | ( n16481 & n16689 ) ;
  assign n16700 = n16406 | n16689 ;
  assign n16702 = ( n16699 & ~n16701 ) | ( n16699 & n16700 ) | ( ~n16701 & n16700 ) ;
  assign n16706 = n16170 &  n16480 ;
  assign n16707 = n16479 &  n16706 ;
  assign n16695 = x92 | n16170 ;
  assign n16696 = x92 &  n16170 ;
  assign n16697 = ( n16695 & ~n16696 ) | ( n16695 & 1'b0 ) | ( ~n16696 & 1'b0 ) ;
  assign n16709 = ( n16405 & n16481 ) | ( n16405 & n16697 ) | ( n16481 & n16697 ) ;
  assign n16708 = n16405 | n16697 ;
  assign n16710 = ( n16707 & ~n16709 ) | ( n16707 & n16708 ) | ( ~n16709 & n16708 ) ;
  assign n16714 = n16178 &  n16480 ;
  assign n16715 = n16479 &  n16714 ;
  assign n16703 = x91 | n16178 ;
  assign n16704 = x91 &  n16178 ;
  assign n16705 = ( n16703 & ~n16704 ) | ( n16703 & 1'b0 ) | ( ~n16704 & 1'b0 ) ;
  assign n16717 = ( n16404 & n16481 ) | ( n16404 & n16705 ) | ( n16481 & n16705 ) ;
  assign n16716 = n16404 | n16705 ;
  assign n16718 = ( n16715 & ~n16717 ) | ( n16715 & n16716 ) | ( ~n16717 & n16716 ) ;
  assign n16722 = n16186 &  n16480 ;
  assign n16723 = n16479 &  n16722 ;
  assign n16711 = x90 | n16186 ;
  assign n16712 = x90 &  n16186 ;
  assign n16713 = ( n16711 & ~n16712 ) | ( n16711 & 1'b0 ) | ( ~n16712 & 1'b0 ) ;
  assign n16725 = ( n16403 & n16481 ) | ( n16403 & n16713 ) | ( n16481 & n16713 ) ;
  assign n16724 = n16403 | n16713 ;
  assign n16726 = ( n16723 & ~n16725 ) | ( n16723 & n16724 ) | ( ~n16725 & n16724 ) ;
  assign n16730 = n16194 &  n16480 ;
  assign n16731 = n16479 &  n16730 ;
  assign n16719 = x89 | n16194 ;
  assign n16720 = x89 &  n16194 ;
  assign n16721 = ( n16719 & ~n16720 ) | ( n16719 & 1'b0 ) | ( ~n16720 & 1'b0 ) ;
  assign n16733 = ( n16402 & n16481 ) | ( n16402 & n16721 ) | ( n16481 & n16721 ) ;
  assign n16732 = n16402 | n16721 ;
  assign n16734 = ( n16731 & ~n16733 ) | ( n16731 & n16732 ) | ( ~n16733 & n16732 ) ;
  assign n16738 = n16202 &  n16480 ;
  assign n16739 = n16479 &  n16738 ;
  assign n16727 = x88 | n16202 ;
  assign n16728 = x88 &  n16202 ;
  assign n16729 = ( n16727 & ~n16728 ) | ( n16727 & 1'b0 ) | ( ~n16728 & 1'b0 ) ;
  assign n16741 = ( n16401 & n16481 ) | ( n16401 & n16729 ) | ( n16481 & n16729 ) ;
  assign n16740 = n16401 | n16729 ;
  assign n16742 = ( n16739 & ~n16741 ) | ( n16739 & n16740 ) | ( ~n16741 & n16740 ) ;
  assign n16746 = n16210 &  n16480 ;
  assign n16747 = n16479 &  n16746 ;
  assign n16735 = x87 | n16210 ;
  assign n16736 = x87 &  n16210 ;
  assign n16737 = ( n16735 & ~n16736 ) | ( n16735 & 1'b0 ) | ( ~n16736 & 1'b0 ) ;
  assign n16749 = ( n16400 & n16481 ) | ( n16400 & n16737 ) | ( n16481 & n16737 ) ;
  assign n16748 = n16400 | n16737 ;
  assign n16750 = ( n16747 & ~n16749 ) | ( n16747 & n16748 ) | ( ~n16749 & n16748 ) ;
  assign n16754 = n16218 &  n16480 ;
  assign n16755 = n16479 &  n16754 ;
  assign n16743 = x86 | n16218 ;
  assign n16744 = x86 &  n16218 ;
  assign n16745 = ( n16743 & ~n16744 ) | ( n16743 & 1'b0 ) | ( ~n16744 & 1'b0 ) ;
  assign n16757 = ( n16399 & n16481 ) | ( n16399 & n16745 ) | ( n16481 & n16745 ) ;
  assign n16756 = n16399 | n16745 ;
  assign n16758 = ( n16755 & ~n16757 ) | ( n16755 & n16756 ) | ( ~n16757 & n16756 ) ;
  assign n16762 = n16226 &  n16480 ;
  assign n16763 = n16479 &  n16762 ;
  assign n16751 = x85 | n16226 ;
  assign n16752 = x85 &  n16226 ;
  assign n16753 = ( n16751 & ~n16752 ) | ( n16751 & 1'b0 ) | ( ~n16752 & 1'b0 ) ;
  assign n16765 = ( n16398 & n16481 ) | ( n16398 & n16753 ) | ( n16481 & n16753 ) ;
  assign n16764 = n16398 | n16753 ;
  assign n16766 = ( n16763 & ~n16765 ) | ( n16763 & n16764 ) | ( ~n16765 & n16764 ) ;
  assign n16770 = n16234 &  n16480 ;
  assign n16771 = n16479 &  n16770 ;
  assign n16759 = x84 | n16234 ;
  assign n16760 = x84 &  n16234 ;
  assign n16761 = ( n16759 & ~n16760 ) | ( n16759 & 1'b0 ) | ( ~n16760 & 1'b0 ) ;
  assign n16773 = ( n16397 & n16481 ) | ( n16397 & n16761 ) | ( n16481 & n16761 ) ;
  assign n16772 = n16397 | n16761 ;
  assign n16774 = ( n16771 & ~n16773 ) | ( n16771 & n16772 ) | ( ~n16773 & n16772 ) ;
  assign n16778 = n16242 &  n16480 ;
  assign n16779 = n16479 &  n16778 ;
  assign n16767 = x83 | n16242 ;
  assign n16768 = x83 &  n16242 ;
  assign n16769 = ( n16767 & ~n16768 ) | ( n16767 & 1'b0 ) | ( ~n16768 & 1'b0 ) ;
  assign n16781 = ( n16396 & n16481 ) | ( n16396 & n16769 ) | ( n16481 & n16769 ) ;
  assign n16780 = n16396 | n16769 ;
  assign n16782 = ( n16779 & ~n16781 ) | ( n16779 & n16780 ) | ( ~n16781 & n16780 ) ;
  assign n16786 = n16250 &  n16480 ;
  assign n16787 = n16479 &  n16786 ;
  assign n16775 = x82 | n16250 ;
  assign n16776 = x82 &  n16250 ;
  assign n16777 = ( n16775 & ~n16776 ) | ( n16775 & 1'b0 ) | ( ~n16776 & 1'b0 ) ;
  assign n16789 = ( n16395 & n16481 ) | ( n16395 & n16777 ) | ( n16481 & n16777 ) ;
  assign n16788 = n16395 | n16777 ;
  assign n16790 = ( n16787 & ~n16789 ) | ( n16787 & n16788 ) | ( ~n16789 & n16788 ) ;
  assign n16794 = n16258 &  n16480 ;
  assign n16795 = n16479 &  n16794 ;
  assign n16783 = x81 | n16258 ;
  assign n16784 = x81 &  n16258 ;
  assign n16785 = ( n16783 & ~n16784 ) | ( n16783 & 1'b0 ) | ( ~n16784 & 1'b0 ) ;
  assign n16797 = ( n16394 & n16481 ) | ( n16394 & n16785 ) | ( n16481 & n16785 ) ;
  assign n16796 = n16394 | n16785 ;
  assign n16798 = ( n16795 & ~n16797 ) | ( n16795 & n16796 ) | ( ~n16797 & n16796 ) ;
  assign n16802 = n16266 &  n16480 ;
  assign n16803 = n16479 &  n16802 ;
  assign n16791 = x80 | n16266 ;
  assign n16792 = x80 &  n16266 ;
  assign n16793 = ( n16791 & ~n16792 ) | ( n16791 & 1'b0 ) | ( ~n16792 & 1'b0 ) ;
  assign n16805 = ( n16393 & n16481 ) | ( n16393 & n16793 ) | ( n16481 & n16793 ) ;
  assign n16804 = n16393 | n16793 ;
  assign n16806 = ( n16803 & ~n16805 ) | ( n16803 & n16804 ) | ( ~n16805 & n16804 ) ;
  assign n16810 = n16274 &  n16480 ;
  assign n16811 = n16479 &  n16810 ;
  assign n16799 = x79 | n16274 ;
  assign n16800 = x79 &  n16274 ;
  assign n16801 = ( n16799 & ~n16800 ) | ( n16799 & 1'b0 ) | ( ~n16800 & 1'b0 ) ;
  assign n16813 = ( n16392 & n16481 ) | ( n16392 & n16801 ) | ( n16481 & n16801 ) ;
  assign n16812 = n16392 | n16801 ;
  assign n16814 = ( n16811 & ~n16813 ) | ( n16811 & n16812 ) | ( ~n16813 & n16812 ) ;
  assign n16818 = n16282 &  n16480 ;
  assign n16819 = n16479 &  n16818 ;
  assign n16807 = x78 | n16282 ;
  assign n16808 = x78 &  n16282 ;
  assign n16809 = ( n16807 & ~n16808 ) | ( n16807 & 1'b0 ) | ( ~n16808 & 1'b0 ) ;
  assign n16821 = ( n16391 & n16481 ) | ( n16391 & n16809 ) | ( n16481 & n16809 ) ;
  assign n16820 = n16391 | n16809 ;
  assign n16822 = ( n16819 & ~n16821 ) | ( n16819 & n16820 ) | ( ~n16821 & n16820 ) ;
  assign n16826 = n16290 &  n16480 ;
  assign n16827 = n16479 &  n16826 ;
  assign n16815 = x77 | n16290 ;
  assign n16816 = x77 &  n16290 ;
  assign n16817 = ( n16815 & ~n16816 ) | ( n16815 & 1'b0 ) | ( ~n16816 & 1'b0 ) ;
  assign n16829 = ( n16390 & n16481 ) | ( n16390 & n16817 ) | ( n16481 & n16817 ) ;
  assign n16828 = n16390 | n16817 ;
  assign n16830 = ( n16827 & ~n16829 ) | ( n16827 & n16828 ) | ( ~n16829 & n16828 ) ;
  assign n16834 = n16298 &  n16480 ;
  assign n16835 = n16479 &  n16834 ;
  assign n16823 = x76 | n16298 ;
  assign n16824 = x76 &  n16298 ;
  assign n16825 = ( n16823 & ~n16824 ) | ( n16823 & 1'b0 ) | ( ~n16824 & 1'b0 ) ;
  assign n16837 = ( n16389 & n16481 ) | ( n16389 & n16825 ) | ( n16481 & n16825 ) ;
  assign n16836 = n16389 | n16825 ;
  assign n16838 = ( n16835 & ~n16837 ) | ( n16835 & n16836 ) | ( ~n16837 & n16836 ) ;
  assign n16842 = n16306 &  n16480 ;
  assign n16843 = n16479 &  n16842 ;
  assign n16831 = x75 | n16306 ;
  assign n16832 = x75 &  n16306 ;
  assign n16833 = ( n16831 & ~n16832 ) | ( n16831 & 1'b0 ) | ( ~n16832 & 1'b0 ) ;
  assign n16845 = ( n16388 & n16481 ) | ( n16388 & n16833 ) | ( n16481 & n16833 ) ;
  assign n16844 = n16388 | n16833 ;
  assign n16846 = ( n16843 & ~n16845 ) | ( n16843 & n16844 ) | ( ~n16845 & n16844 ) ;
  assign n16850 = n16314 &  n16480 ;
  assign n16851 = n16479 &  n16850 ;
  assign n16839 = x74 | n16314 ;
  assign n16840 = x74 &  n16314 ;
  assign n16841 = ( n16839 & ~n16840 ) | ( n16839 & 1'b0 ) | ( ~n16840 & 1'b0 ) ;
  assign n16853 = ( n16387 & n16481 ) | ( n16387 & n16841 ) | ( n16481 & n16841 ) ;
  assign n16852 = n16387 | n16841 ;
  assign n16854 = ( n16851 & ~n16853 ) | ( n16851 & n16852 ) | ( ~n16853 & n16852 ) ;
  assign n16858 = n16322 &  n16480 ;
  assign n16859 = n16479 &  n16858 ;
  assign n16847 = x73 | n16322 ;
  assign n16848 = x73 &  n16322 ;
  assign n16849 = ( n16847 & ~n16848 ) | ( n16847 & 1'b0 ) | ( ~n16848 & 1'b0 ) ;
  assign n16861 = ( n16386 & n16481 ) | ( n16386 & n16849 ) | ( n16481 & n16849 ) ;
  assign n16860 = n16386 | n16849 ;
  assign n16862 = ( n16859 & ~n16861 ) | ( n16859 & n16860 ) | ( ~n16861 & n16860 ) ;
  assign n16866 = n16330 &  n16480 ;
  assign n16867 = n16479 &  n16866 ;
  assign n16855 = x72 | n16330 ;
  assign n16856 = x72 &  n16330 ;
  assign n16857 = ( n16855 & ~n16856 ) | ( n16855 & 1'b0 ) | ( ~n16856 & 1'b0 ) ;
  assign n16869 = ( n16385 & n16481 ) | ( n16385 & n16857 ) | ( n16481 & n16857 ) ;
  assign n16868 = n16385 | n16857 ;
  assign n16870 = ( n16867 & ~n16869 ) | ( n16867 & n16868 ) | ( ~n16869 & n16868 ) ;
  assign n16874 = n16338 &  n16480 ;
  assign n16875 = n16479 &  n16874 ;
  assign n16863 = x71 | n16338 ;
  assign n16864 = x71 &  n16338 ;
  assign n16865 = ( n16863 & ~n16864 ) | ( n16863 & 1'b0 ) | ( ~n16864 & 1'b0 ) ;
  assign n16877 = ( n16384 & n16481 ) | ( n16384 & n16865 ) | ( n16481 & n16865 ) ;
  assign n16876 = n16384 | n16865 ;
  assign n16878 = ( n16875 & ~n16877 ) | ( n16875 & n16876 ) | ( ~n16877 & n16876 ) ;
  assign n16882 = n16346 &  n16480 ;
  assign n16883 = n16479 &  n16882 ;
  assign n16871 = x70 | n16346 ;
  assign n16872 = x70 &  n16346 ;
  assign n16873 = ( n16871 & ~n16872 ) | ( n16871 & 1'b0 ) | ( ~n16872 & 1'b0 ) ;
  assign n16885 = ( n16383 & n16481 ) | ( n16383 & n16873 ) | ( n16481 & n16873 ) ;
  assign n16884 = n16383 | n16873 ;
  assign n16886 = ( n16883 & ~n16885 ) | ( n16883 & n16884 ) | ( ~n16885 & n16884 ) ;
  assign n16890 = n16354 &  n16480 ;
  assign n16891 = n16479 &  n16890 ;
  assign n16879 = x69 | n16354 ;
  assign n16880 = x69 &  n16354 ;
  assign n16881 = ( n16879 & ~n16880 ) | ( n16879 & 1'b0 ) | ( ~n16880 & 1'b0 ) ;
  assign n16893 = ( n16382 & n16481 ) | ( n16382 & n16881 ) | ( n16481 & n16881 ) ;
  assign n16892 = n16382 | n16881 ;
  assign n16894 = ( n16891 & ~n16893 ) | ( n16891 & n16892 ) | ( ~n16893 & n16892 ) ;
  assign n16898 = n16362 &  n16480 ;
  assign n16899 = n16479 &  n16898 ;
  assign n16887 = x68 | n16362 ;
  assign n16888 = x68 &  n16362 ;
  assign n16889 = ( n16887 & ~n16888 ) | ( n16887 & 1'b0 ) | ( ~n16888 & 1'b0 ) ;
  assign n16901 = ( n16381 & n16481 ) | ( n16381 & n16889 ) | ( n16481 & n16889 ) ;
  assign n16900 = n16381 | n16889 ;
  assign n16902 = ( n16899 & ~n16901 ) | ( n16899 & n16900 ) | ( ~n16901 & n16900 ) ;
  assign n16906 = n16367 &  n16480 ;
  assign n16907 = n16479 &  n16906 ;
  assign n16895 = x67 | n16367 ;
  assign n16896 = x67 &  n16367 ;
  assign n16897 = ( n16895 & ~n16896 ) | ( n16895 & 1'b0 ) | ( ~n16896 & 1'b0 ) ;
  assign n16909 = ( n16380 & n16481 ) | ( n16380 & n16897 ) | ( n16481 & n16897 ) ;
  assign n16908 = n16380 | n16897 ;
  assign n16910 = ( n16907 & ~n16909 ) | ( n16907 & n16908 ) | ( ~n16909 & n16908 ) ;
  assign n16911 = n16373 &  n16480 ;
  assign n16912 = n16479 &  n16911 ;
  assign n16903 = x66 | n16373 ;
  assign n16904 = x66 &  n16373 ;
  assign n16905 = ( n16903 & ~n16904 ) | ( n16903 & 1'b0 ) | ( ~n16904 & 1'b0 ) ;
  assign n16913 = n16379 &  n16905 ;
  assign n16914 = ( n16379 & ~n16481 ) | ( n16379 & n16905 ) | ( ~n16481 & n16905 ) ;
  assign n16915 = ( n16912 & ~n16913 ) | ( n16912 & n16914 ) | ( ~n16913 & n16914 ) ;
  assign n16916 = ( n16377 & ~x65 ) | ( n16377 & n16378 ) | ( ~x65 & n16378 ) ;
  assign n16917 = ( n16379 & ~n16378 ) | ( n16379 & n16916 ) | ( ~n16378 & n16916 ) ;
  assign n16918 = ~n16481 & n16917 ;
  assign n16919 = n16377 &  n16480 ;
  assign n16920 = n16479 &  n16919 ;
  assign n16921 = n16918 | n16920 ;
  assign n16922 = ( x64 & ~n16481 ) | ( x64 & 1'b0 ) | ( ~n16481 & 1'b0 ) ;
  assign n16923 = ( x4 & ~n16922 ) | ( x4 & 1'b0 ) | ( ~n16922 & 1'b0 ) ;
  assign n16924 = ( n16378 & ~n16481 ) | ( n16378 & 1'b0 ) | ( ~n16481 & 1'b0 ) ;
  assign n16925 = n16923 | n16924 ;
  assign n16926 = ~x3 & x64 ;
  assign n16927 = ( x65 & ~n16925 ) | ( x65 & n16926 ) | ( ~n16925 & n16926 ) ;
  assign n16928 = ( x66 & ~n16921 ) | ( x66 & n16927 ) | ( ~n16921 & n16927 ) ;
  assign n16929 = ( x67 & ~n16915 ) | ( x67 & n16928 ) | ( ~n16915 & n16928 ) ;
  assign n16930 = ( x68 & ~n16910 ) | ( x68 & n16929 ) | ( ~n16910 & n16929 ) ;
  assign n16931 = ( x69 & ~n16902 ) | ( x69 & n16930 ) | ( ~n16902 & n16930 ) ;
  assign n16932 = ( x70 & ~n16894 ) | ( x70 & n16931 ) | ( ~n16894 & n16931 ) ;
  assign n16933 = ( x71 & ~n16886 ) | ( x71 & n16932 ) | ( ~n16886 & n16932 ) ;
  assign n16934 = ( x72 & ~n16878 ) | ( x72 & n16933 ) | ( ~n16878 & n16933 ) ;
  assign n16935 = ( x73 & ~n16870 ) | ( x73 & n16934 ) | ( ~n16870 & n16934 ) ;
  assign n16936 = ( x74 & ~n16862 ) | ( x74 & n16935 ) | ( ~n16862 & n16935 ) ;
  assign n16937 = ( x75 & ~n16854 ) | ( x75 & n16936 ) | ( ~n16854 & n16936 ) ;
  assign n16938 = ( x76 & ~n16846 ) | ( x76 & n16937 ) | ( ~n16846 & n16937 ) ;
  assign n16939 = ( x77 & ~n16838 ) | ( x77 & n16938 ) | ( ~n16838 & n16938 ) ;
  assign n16940 = ( x78 & ~n16830 ) | ( x78 & n16939 ) | ( ~n16830 & n16939 ) ;
  assign n16941 = ( x79 & ~n16822 ) | ( x79 & n16940 ) | ( ~n16822 & n16940 ) ;
  assign n16942 = ( x80 & ~n16814 ) | ( x80 & n16941 ) | ( ~n16814 & n16941 ) ;
  assign n16943 = ( x81 & ~n16806 ) | ( x81 & n16942 ) | ( ~n16806 & n16942 ) ;
  assign n16944 = ( x82 & ~n16798 ) | ( x82 & n16943 ) | ( ~n16798 & n16943 ) ;
  assign n16945 = ( x83 & ~n16790 ) | ( x83 & n16944 ) | ( ~n16790 & n16944 ) ;
  assign n16946 = ( x84 & ~n16782 ) | ( x84 & n16945 ) | ( ~n16782 & n16945 ) ;
  assign n16947 = ( x85 & ~n16774 ) | ( x85 & n16946 ) | ( ~n16774 & n16946 ) ;
  assign n16948 = ( x86 & ~n16766 ) | ( x86 & n16947 ) | ( ~n16766 & n16947 ) ;
  assign n16949 = ( x87 & ~n16758 ) | ( x87 & n16948 ) | ( ~n16758 & n16948 ) ;
  assign n16950 = ( x88 & ~n16750 ) | ( x88 & n16949 ) | ( ~n16750 & n16949 ) ;
  assign n16951 = ( x89 & ~n16742 ) | ( x89 & n16950 ) | ( ~n16742 & n16950 ) ;
  assign n16952 = ( x90 & ~n16734 ) | ( x90 & n16951 ) | ( ~n16734 & n16951 ) ;
  assign n16953 = ( x91 & ~n16726 ) | ( x91 & n16952 ) | ( ~n16726 & n16952 ) ;
  assign n16954 = ( x92 & ~n16718 ) | ( x92 & n16953 ) | ( ~n16718 & n16953 ) ;
  assign n16955 = ( x93 & ~n16710 ) | ( x93 & n16954 ) | ( ~n16710 & n16954 ) ;
  assign n16956 = ( x94 & ~n16702 ) | ( x94 & n16955 ) | ( ~n16702 & n16955 ) ;
  assign n16957 = ( x95 & ~n16694 ) | ( x95 & n16956 ) | ( ~n16694 & n16956 ) ;
  assign n16958 = ( x96 & ~n16686 ) | ( x96 & n16957 ) | ( ~n16686 & n16957 ) ;
  assign n16959 = ( x97 & ~n16678 ) | ( x97 & n16958 ) | ( ~n16678 & n16958 ) ;
  assign n16960 = ( x98 & ~n16670 ) | ( x98 & n16959 ) | ( ~n16670 & n16959 ) ;
  assign n16961 = ( x99 & ~n16662 ) | ( x99 & n16960 ) | ( ~n16662 & n16960 ) ;
  assign n16962 = ( x100 & ~n16654 ) | ( x100 & n16961 ) | ( ~n16654 & n16961 ) ;
  assign n16963 = ( x101 & ~n16646 ) | ( x101 & n16962 ) | ( ~n16646 & n16962 ) ;
  assign n16964 = ( x102 & ~n16638 ) | ( x102 & n16963 ) | ( ~n16638 & n16963 ) ;
  assign n16965 = ( x103 & ~n16630 ) | ( x103 & n16964 ) | ( ~n16630 & n16964 ) ;
  assign n16966 = ( x104 & ~n16622 ) | ( x104 & n16965 ) | ( ~n16622 & n16965 ) ;
  assign n16967 = ( x105 & ~n16614 ) | ( x105 & n16966 ) | ( ~n16614 & n16966 ) ;
  assign n16968 = ( x106 & ~n16606 ) | ( x106 & n16967 ) | ( ~n16606 & n16967 ) ;
  assign n16969 = ( x107 & ~n16598 ) | ( x107 & n16968 ) | ( ~n16598 & n16968 ) ;
  assign n16970 = ( x108 & ~n16590 ) | ( x108 & n16969 ) | ( ~n16590 & n16969 ) ;
  assign n16971 = ( x109 & ~n16582 ) | ( x109 & n16970 ) | ( ~n16582 & n16970 ) ;
  assign n16972 = ( x110 & ~n16574 ) | ( x110 & n16971 ) | ( ~n16574 & n16971 ) ;
  assign n16973 = ( x111 & ~n16566 ) | ( x111 & n16972 ) | ( ~n16566 & n16972 ) ;
  assign n16974 = ( x112 & ~n16558 ) | ( x112 & n16973 ) | ( ~n16558 & n16973 ) ;
  assign n16975 = ( x113 & ~n16550 ) | ( x113 & n16974 ) | ( ~n16550 & n16974 ) ;
  assign n16976 = ( x114 & ~n16542 ) | ( x114 & n16975 ) | ( ~n16542 & n16975 ) ;
  assign n16977 = ( x115 & ~n16534 ) | ( x115 & n16976 ) | ( ~n16534 & n16976 ) ;
  assign n16978 = ( x116 & ~n16526 ) | ( x116 & n16977 ) | ( ~n16526 & n16977 ) ;
  assign n16979 = ( x117 & ~n16518 ) | ( x117 & n16978 ) | ( ~n16518 & n16978 ) ;
  assign n16980 = ( x118 & ~n16510 ) | ( x118 & n16979 ) | ( ~n16510 & n16979 ) ;
  assign n16981 = ( x119 & ~n16502 ) | ( x119 & n16980 ) | ( ~n16502 & n16980 ) ;
  assign n16982 = ( x120 & ~n16494 ) | ( x120 & n16981 ) | ( ~n16494 & n16981 ) ;
  assign n16986 = ( x121 & ~n16486 ) | ( x121 & n16982 ) | ( ~n16486 & n16982 ) ;
  assign n17006 = ( x122 & ~n16994 ) | ( x122 & n16986 ) | ( ~n16994 & n16986 ) ;
  assign n17007 = ( x123 & ~n17005 ) | ( x123 & n17006 ) | ( ~n17005 & n17006 ) ;
  assign n17008 = n16474 | n16476 ;
  assign n17009 = ( n16466 & ~n17008 ) | ( n16466 & 1'b0 ) | ( ~n17008 & 1'b0 ) ;
  assign n17010 = ~n16466 & n17008 ;
  assign n17011 = ( n17009 & ~n16481 ) | ( n17009 & n17010 ) | ( ~n16481 & n17010 ) ;
  assign n17012 = n15943 &  n16473 ;
  assign n17013 = n16479 &  n17012 ;
  assign n17014 = n17011 | n17013 ;
  assign n17015 = ~x124 & n17014 ;
  assign n17016 = ( x124 & ~n17013 ) | ( x124 & 1'b0 ) | ( ~n17013 & 1'b0 ) ;
  assign n17017 = ~n17011 & n17016 ;
  assign n17018 = n235 | n17017 ;
  assign n17019 = n17015 | n17018 ;
  assign n17020 = n17007 | n17019 ;
  assign n17021 = ~n17014 |  n152 ;
  assign n17549 = n17005 &  n17021 ;
  assign n17550 = n17020 &  n17549 ;
  assign n17546 = x123 | n17005 ;
  assign n17547 = x123 &  n17005 ;
  assign n17548 = ( n17546 & ~n17547 ) | ( n17546 & 1'b0 ) | ( ~n17547 & 1'b0 ) ;
  assign n17551 = n17006 &  n17548 ;
  assign n17022 = n17020 &  n17021 ;
  assign n17552 = ( n17006 & ~n17022 ) | ( n17006 & n17548 ) | ( ~n17022 & n17548 ) ;
  assign n17553 = ( n17550 & ~n17551 ) | ( n17550 & n17552 ) | ( ~n17551 & n17552 ) ;
  assign n17023 = n16994 &  n17021 ;
  assign n17024 = n17020 &  n17023 ;
  assign n16995 = x122 | n16994 ;
  assign n16996 = x122 &  n16994 ;
  assign n16997 = ( n16995 & ~n16996 ) | ( n16995 & 1'b0 ) | ( ~n16996 & 1'b0 ) ;
  assign n17025 = n16986 &  n16997 ;
  assign n17026 = ( n16986 & ~n17022 ) | ( n16986 & n16997 ) | ( ~n17022 & n16997 ) ;
  assign n17027 = ( n17024 & ~n17025 ) | ( n17024 & n17026 ) | ( ~n17025 & n17026 ) ;
  assign n17031 = n16486 &  n17021 ;
  assign n17032 = n17020 &  n17031 ;
  assign n16983 = x121 | n16486 ;
  assign n16984 = x121 &  n16486 ;
  assign n16985 = ( n16983 & ~n16984 ) | ( n16983 & 1'b0 ) | ( ~n16984 & 1'b0 ) ;
  assign n17034 = ( n16982 & n16985 ) | ( n16982 & n17022 ) | ( n16985 & n17022 ) ;
  assign n17033 = n16982 | n16985 ;
  assign n17035 = ( n17032 & ~n17034 ) | ( n17032 & n17033 ) | ( ~n17034 & n17033 ) ;
  assign n17039 = n16494 &  n17021 ;
  assign n17040 = n17020 &  n17039 ;
  assign n17028 = x120 | n16494 ;
  assign n17029 = x120 &  n16494 ;
  assign n17030 = ( n17028 & ~n17029 ) | ( n17028 & 1'b0 ) | ( ~n17029 & 1'b0 ) ;
  assign n17041 = n16981 &  n17030 ;
  assign n17042 = ( n16981 & ~n17022 ) | ( n16981 & n17030 ) | ( ~n17022 & n17030 ) ;
  assign n17043 = ( n17040 & ~n17041 ) | ( n17040 & n17042 ) | ( ~n17041 & n17042 ) ;
  assign n17047 = n16502 &  n17021 ;
  assign n17048 = n17020 &  n17047 ;
  assign n17036 = x119 | n16502 ;
  assign n17037 = x119 &  n16502 ;
  assign n17038 = ( n17036 & ~n17037 ) | ( n17036 & 1'b0 ) | ( ~n17037 & 1'b0 ) ;
  assign n17049 = n16980 &  n17038 ;
  assign n17050 = ( n16980 & ~n17022 ) | ( n16980 & n17038 ) | ( ~n17022 & n17038 ) ;
  assign n17051 = ( n17048 & ~n17049 ) | ( n17048 & n17050 ) | ( ~n17049 & n17050 ) ;
  assign n17055 = n16510 &  n17021 ;
  assign n17056 = n17020 &  n17055 ;
  assign n17044 = x118 | n16510 ;
  assign n17045 = x118 &  n16510 ;
  assign n17046 = ( n17044 & ~n17045 ) | ( n17044 & 1'b0 ) | ( ~n17045 & 1'b0 ) ;
  assign n17058 = ( n16979 & n17022 ) | ( n16979 & n17046 ) | ( n17022 & n17046 ) ;
  assign n17057 = n16979 | n17046 ;
  assign n17059 = ( n17056 & ~n17058 ) | ( n17056 & n17057 ) | ( ~n17058 & n17057 ) ;
  assign n17063 = n16518 &  n17021 ;
  assign n17064 = n17020 &  n17063 ;
  assign n17052 = x117 | n16518 ;
  assign n17053 = x117 &  n16518 ;
  assign n17054 = ( n17052 & ~n17053 ) | ( n17052 & 1'b0 ) | ( ~n17053 & 1'b0 ) ;
  assign n17066 = ( n16978 & n17022 ) | ( n16978 & n17054 ) | ( n17022 & n17054 ) ;
  assign n17065 = n16978 | n17054 ;
  assign n17067 = ( n17064 & ~n17066 ) | ( n17064 & n17065 ) | ( ~n17066 & n17065 ) ;
  assign n17071 = n16526 &  n17021 ;
  assign n17072 = n17020 &  n17071 ;
  assign n17060 = x116 | n16526 ;
  assign n17061 = x116 &  n16526 ;
  assign n17062 = ( n17060 & ~n17061 ) | ( n17060 & 1'b0 ) | ( ~n17061 & 1'b0 ) ;
  assign n17074 = ( n16977 & n17022 ) | ( n16977 & n17062 ) | ( n17022 & n17062 ) ;
  assign n17073 = n16977 | n17062 ;
  assign n17075 = ( n17072 & ~n17074 ) | ( n17072 & n17073 ) | ( ~n17074 & n17073 ) ;
  assign n17079 = n16534 &  n17021 ;
  assign n17080 = n17020 &  n17079 ;
  assign n17068 = x115 | n16534 ;
  assign n17069 = x115 &  n16534 ;
  assign n17070 = ( n17068 & ~n17069 ) | ( n17068 & 1'b0 ) | ( ~n17069 & 1'b0 ) ;
  assign n17082 = ( n16976 & n17022 ) | ( n16976 & n17070 ) | ( n17022 & n17070 ) ;
  assign n17081 = n16976 | n17070 ;
  assign n17083 = ( n17080 & ~n17082 ) | ( n17080 & n17081 ) | ( ~n17082 & n17081 ) ;
  assign n17087 = n16542 &  n17021 ;
  assign n17088 = n17020 &  n17087 ;
  assign n17076 = x114 | n16542 ;
  assign n17077 = x114 &  n16542 ;
  assign n17078 = ( n17076 & ~n17077 ) | ( n17076 & 1'b0 ) | ( ~n17077 & 1'b0 ) ;
  assign n17090 = ( n16975 & n17022 ) | ( n16975 & n17078 ) | ( n17022 & n17078 ) ;
  assign n17089 = n16975 | n17078 ;
  assign n17091 = ( n17088 & ~n17090 ) | ( n17088 & n17089 ) | ( ~n17090 & n17089 ) ;
  assign n17095 = n16550 &  n17021 ;
  assign n17096 = n17020 &  n17095 ;
  assign n17084 = x113 | n16550 ;
  assign n17085 = x113 &  n16550 ;
  assign n17086 = ( n17084 & ~n17085 ) | ( n17084 & 1'b0 ) | ( ~n17085 & 1'b0 ) ;
  assign n17098 = ( n16974 & n17022 ) | ( n16974 & n17086 ) | ( n17022 & n17086 ) ;
  assign n17097 = n16974 | n17086 ;
  assign n17099 = ( n17096 & ~n17098 ) | ( n17096 & n17097 ) | ( ~n17098 & n17097 ) ;
  assign n17103 = n16558 &  n17021 ;
  assign n17104 = n17020 &  n17103 ;
  assign n17092 = x112 | n16558 ;
  assign n17093 = x112 &  n16558 ;
  assign n17094 = ( n17092 & ~n17093 ) | ( n17092 & 1'b0 ) | ( ~n17093 & 1'b0 ) ;
  assign n17106 = ( n16973 & n17022 ) | ( n16973 & n17094 ) | ( n17022 & n17094 ) ;
  assign n17105 = n16973 | n17094 ;
  assign n17107 = ( n17104 & ~n17106 ) | ( n17104 & n17105 ) | ( ~n17106 & n17105 ) ;
  assign n17111 = n16566 &  n17021 ;
  assign n17112 = n17020 &  n17111 ;
  assign n17100 = x111 | n16566 ;
  assign n17101 = x111 &  n16566 ;
  assign n17102 = ( n17100 & ~n17101 ) | ( n17100 & 1'b0 ) | ( ~n17101 & 1'b0 ) ;
  assign n17114 = ( n16972 & n17022 ) | ( n16972 & n17102 ) | ( n17022 & n17102 ) ;
  assign n17113 = n16972 | n17102 ;
  assign n17115 = ( n17112 & ~n17114 ) | ( n17112 & n17113 ) | ( ~n17114 & n17113 ) ;
  assign n17119 = n16574 &  n17021 ;
  assign n17120 = n17020 &  n17119 ;
  assign n17108 = x110 | n16574 ;
  assign n17109 = x110 &  n16574 ;
  assign n17110 = ( n17108 & ~n17109 ) | ( n17108 & 1'b0 ) | ( ~n17109 & 1'b0 ) ;
  assign n17122 = ( n16971 & n17022 ) | ( n16971 & n17110 ) | ( n17022 & n17110 ) ;
  assign n17121 = n16971 | n17110 ;
  assign n17123 = ( n17120 & ~n17122 ) | ( n17120 & n17121 ) | ( ~n17122 & n17121 ) ;
  assign n17127 = n16582 &  n17021 ;
  assign n17128 = n17020 &  n17127 ;
  assign n17116 = x109 | n16582 ;
  assign n17117 = x109 &  n16582 ;
  assign n17118 = ( n17116 & ~n17117 ) | ( n17116 & 1'b0 ) | ( ~n17117 & 1'b0 ) ;
  assign n17130 = ( n16970 & n17022 ) | ( n16970 & n17118 ) | ( n17022 & n17118 ) ;
  assign n17129 = n16970 | n17118 ;
  assign n17131 = ( n17128 & ~n17130 ) | ( n17128 & n17129 ) | ( ~n17130 & n17129 ) ;
  assign n17135 = n16590 &  n17021 ;
  assign n17136 = n17020 &  n17135 ;
  assign n17124 = x108 | n16590 ;
  assign n17125 = x108 &  n16590 ;
  assign n17126 = ( n17124 & ~n17125 ) | ( n17124 & 1'b0 ) | ( ~n17125 & 1'b0 ) ;
  assign n17138 = ( n16969 & n17022 ) | ( n16969 & n17126 ) | ( n17022 & n17126 ) ;
  assign n17137 = n16969 | n17126 ;
  assign n17139 = ( n17136 & ~n17138 ) | ( n17136 & n17137 ) | ( ~n17138 & n17137 ) ;
  assign n17143 = n16598 &  n17021 ;
  assign n17144 = n17020 &  n17143 ;
  assign n17132 = x107 | n16598 ;
  assign n17133 = x107 &  n16598 ;
  assign n17134 = ( n17132 & ~n17133 ) | ( n17132 & 1'b0 ) | ( ~n17133 & 1'b0 ) ;
  assign n17146 = ( n16968 & n17022 ) | ( n16968 & n17134 ) | ( n17022 & n17134 ) ;
  assign n17145 = n16968 | n17134 ;
  assign n17147 = ( n17144 & ~n17146 ) | ( n17144 & n17145 ) | ( ~n17146 & n17145 ) ;
  assign n17151 = n16606 &  n17021 ;
  assign n17152 = n17020 &  n17151 ;
  assign n17140 = x106 | n16606 ;
  assign n17141 = x106 &  n16606 ;
  assign n17142 = ( n17140 & ~n17141 ) | ( n17140 & 1'b0 ) | ( ~n17141 & 1'b0 ) ;
  assign n17154 = ( n16967 & n17022 ) | ( n16967 & n17142 ) | ( n17022 & n17142 ) ;
  assign n17153 = n16967 | n17142 ;
  assign n17155 = ( n17152 & ~n17154 ) | ( n17152 & n17153 ) | ( ~n17154 & n17153 ) ;
  assign n17159 = n16614 &  n17021 ;
  assign n17160 = n17020 &  n17159 ;
  assign n17148 = x105 | n16614 ;
  assign n17149 = x105 &  n16614 ;
  assign n17150 = ( n17148 & ~n17149 ) | ( n17148 & 1'b0 ) | ( ~n17149 & 1'b0 ) ;
  assign n17162 = ( n16966 & n17022 ) | ( n16966 & n17150 ) | ( n17022 & n17150 ) ;
  assign n17161 = n16966 | n17150 ;
  assign n17163 = ( n17160 & ~n17162 ) | ( n17160 & n17161 ) | ( ~n17162 & n17161 ) ;
  assign n17167 = n16622 &  n17021 ;
  assign n17168 = n17020 &  n17167 ;
  assign n17156 = x104 | n16622 ;
  assign n17157 = x104 &  n16622 ;
  assign n17158 = ( n17156 & ~n17157 ) | ( n17156 & 1'b0 ) | ( ~n17157 & 1'b0 ) ;
  assign n17170 = ( n16965 & n17022 ) | ( n16965 & n17158 ) | ( n17022 & n17158 ) ;
  assign n17169 = n16965 | n17158 ;
  assign n17171 = ( n17168 & ~n17170 ) | ( n17168 & n17169 ) | ( ~n17170 & n17169 ) ;
  assign n17175 = n16630 &  n17021 ;
  assign n17176 = n17020 &  n17175 ;
  assign n17164 = x103 | n16630 ;
  assign n17165 = x103 &  n16630 ;
  assign n17166 = ( n17164 & ~n17165 ) | ( n17164 & 1'b0 ) | ( ~n17165 & 1'b0 ) ;
  assign n17178 = ( n16964 & n17022 ) | ( n16964 & n17166 ) | ( n17022 & n17166 ) ;
  assign n17177 = n16964 | n17166 ;
  assign n17179 = ( n17176 & ~n17178 ) | ( n17176 & n17177 ) | ( ~n17178 & n17177 ) ;
  assign n17183 = n16638 &  n17021 ;
  assign n17184 = n17020 &  n17183 ;
  assign n17172 = x102 | n16638 ;
  assign n17173 = x102 &  n16638 ;
  assign n17174 = ( n17172 & ~n17173 ) | ( n17172 & 1'b0 ) | ( ~n17173 & 1'b0 ) ;
  assign n17186 = ( n16963 & n17022 ) | ( n16963 & n17174 ) | ( n17022 & n17174 ) ;
  assign n17185 = n16963 | n17174 ;
  assign n17187 = ( n17184 & ~n17186 ) | ( n17184 & n17185 ) | ( ~n17186 & n17185 ) ;
  assign n17191 = n16646 &  n17021 ;
  assign n17192 = n17020 &  n17191 ;
  assign n17180 = x101 | n16646 ;
  assign n17181 = x101 &  n16646 ;
  assign n17182 = ( n17180 & ~n17181 ) | ( n17180 & 1'b0 ) | ( ~n17181 & 1'b0 ) ;
  assign n17194 = ( n16962 & n17022 ) | ( n16962 & n17182 ) | ( n17022 & n17182 ) ;
  assign n17193 = n16962 | n17182 ;
  assign n17195 = ( n17192 & ~n17194 ) | ( n17192 & n17193 ) | ( ~n17194 & n17193 ) ;
  assign n17199 = n16654 &  n17021 ;
  assign n17200 = n17020 &  n17199 ;
  assign n17188 = x100 | n16654 ;
  assign n17189 = x100 &  n16654 ;
  assign n17190 = ( n17188 & ~n17189 ) | ( n17188 & 1'b0 ) | ( ~n17189 & 1'b0 ) ;
  assign n17202 = ( n16961 & n17022 ) | ( n16961 & n17190 ) | ( n17022 & n17190 ) ;
  assign n17201 = n16961 | n17190 ;
  assign n17203 = ( n17200 & ~n17202 ) | ( n17200 & n17201 ) | ( ~n17202 & n17201 ) ;
  assign n17207 = n16662 &  n17021 ;
  assign n17208 = n17020 &  n17207 ;
  assign n17196 = x99 | n16662 ;
  assign n17197 = x99 &  n16662 ;
  assign n17198 = ( n17196 & ~n17197 ) | ( n17196 & 1'b0 ) | ( ~n17197 & 1'b0 ) ;
  assign n17210 = ( n16960 & n17022 ) | ( n16960 & n17198 ) | ( n17022 & n17198 ) ;
  assign n17209 = n16960 | n17198 ;
  assign n17211 = ( n17208 & ~n17210 ) | ( n17208 & n17209 ) | ( ~n17210 & n17209 ) ;
  assign n17215 = n16670 &  n17021 ;
  assign n17216 = n17020 &  n17215 ;
  assign n17204 = x98 | n16670 ;
  assign n17205 = x98 &  n16670 ;
  assign n17206 = ( n17204 & ~n17205 ) | ( n17204 & 1'b0 ) | ( ~n17205 & 1'b0 ) ;
  assign n17218 = ( n16959 & n17022 ) | ( n16959 & n17206 ) | ( n17022 & n17206 ) ;
  assign n17217 = n16959 | n17206 ;
  assign n17219 = ( n17216 & ~n17218 ) | ( n17216 & n17217 ) | ( ~n17218 & n17217 ) ;
  assign n17223 = n16678 &  n17021 ;
  assign n17224 = n17020 &  n17223 ;
  assign n17212 = x97 | n16678 ;
  assign n17213 = x97 &  n16678 ;
  assign n17214 = ( n17212 & ~n17213 ) | ( n17212 & 1'b0 ) | ( ~n17213 & 1'b0 ) ;
  assign n17226 = ( n16958 & n17022 ) | ( n16958 & n17214 ) | ( n17022 & n17214 ) ;
  assign n17225 = n16958 | n17214 ;
  assign n17227 = ( n17224 & ~n17226 ) | ( n17224 & n17225 ) | ( ~n17226 & n17225 ) ;
  assign n17231 = n16686 &  n17021 ;
  assign n17232 = n17020 &  n17231 ;
  assign n17220 = x96 | n16686 ;
  assign n17221 = x96 &  n16686 ;
  assign n17222 = ( n17220 & ~n17221 ) | ( n17220 & 1'b0 ) | ( ~n17221 & 1'b0 ) ;
  assign n17234 = ( n16957 & n17022 ) | ( n16957 & n17222 ) | ( n17022 & n17222 ) ;
  assign n17233 = n16957 | n17222 ;
  assign n17235 = ( n17232 & ~n17234 ) | ( n17232 & n17233 ) | ( ~n17234 & n17233 ) ;
  assign n17239 = n16694 &  n17021 ;
  assign n17240 = n17020 &  n17239 ;
  assign n17228 = x95 | n16694 ;
  assign n17229 = x95 &  n16694 ;
  assign n17230 = ( n17228 & ~n17229 ) | ( n17228 & 1'b0 ) | ( ~n17229 & 1'b0 ) ;
  assign n17242 = ( n16956 & n17022 ) | ( n16956 & n17230 ) | ( n17022 & n17230 ) ;
  assign n17241 = n16956 | n17230 ;
  assign n17243 = ( n17240 & ~n17242 ) | ( n17240 & n17241 ) | ( ~n17242 & n17241 ) ;
  assign n17247 = n16702 &  n17021 ;
  assign n17248 = n17020 &  n17247 ;
  assign n17236 = x94 | n16702 ;
  assign n17237 = x94 &  n16702 ;
  assign n17238 = ( n17236 & ~n17237 ) | ( n17236 & 1'b0 ) | ( ~n17237 & 1'b0 ) ;
  assign n17250 = ( n16955 & n17022 ) | ( n16955 & n17238 ) | ( n17022 & n17238 ) ;
  assign n17249 = n16955 | n17238 ;
  assign n17251 = ( n17248 & ~n17250 ) | ( n17248 & n17249 ) | ( ~n17250 & n17249 ) ;
  assign n17255 = n16710 &  n17021 ;
  assign n17256 = n17020 &  n17255 ;
  assign n17244 = x93 | n16710 ;
  assign n17245 = x93 &  n16710 ;
  assign n17246 = ( n17244 & ~n17245 ) | ( n17244 & 1'b0 ) | ( ~n17245 & 1'b0 ) ;
  assign n17258 = ( n16954 & n17022 ) | ( n16954 & n17246 ) | ( n17022 & n17246 ) ;
  assign n17257 = n16954 | n17246 ;
  assign n17259 = ( n17256 & ~n17258 ) | ( n17256 & n17257 ) | ( ~n17258 & n17257 ) ;
  assign n17263 = n16718 &  n17021 ;
  assign n17264 = n17020 &  n17263 ;
  assign n17252 = x92 | n16718 ;
  assign n17253 = x92 &  n16718 ;
  assign n17254 = ( n17252 & ~n17253 ) | ( n17252 & 1'b0 ) | ( ~n17253 & 1'b0 ) ;
  assign n17266 = ( n16953 & n17022 ) | ( n16953 & n17254 ) | ( n17022 & n17254 ) ;
  assign n17265 = n16953 | n17254 ;
  assign n17267 = ( n17264 & ~n17266 ) | ( n17264 & n17265 ) | ( ~n17266 & n17265 ) ;
  assign n17271 = n16726 &  n17021 ;
  assign n17272 = n17020 &  n17271 ;
  assign n17260 = x91 | n16726 ;
  assign n17261 = x91 &  n16726 ;
  assign n17262 = ( n17260 & ~n17261 ) | ( n17260 & 1'b0 ) | ( ~n17261 & 1'b0 ) ;
  assign n17274 = ( n16952 & n17022 ) | ( n16952 & n17262 ) | ( n17022 & n17262 ) ;
  assign n17273 = n16952 | n17262 ;
  assign n17275 = ( n17272 & ~n17274 ) | ( n17272 & n17273 ) | ( ~n17274 & n17273 ) ;
  assign n17279 = n16734 &  n17021 ;
  assign n17280 = n17020 &  n17279 ;
  assign n17268 = x90 | n16734 ;
  assign n17269 = x90 &  n16734 ;
  assign n17270 = ( n17268 & ~n17269 ) | ( n17268 & 1'b0 ) | ( ~n17269 & 1'b0 ) ;
  assign n17282 = ( n16951 & n17022 ) | ( n16951 & n17270 ) | ( n17022 & n17270 ) ;
  assign n17281 = n16951 | n17270 ;
  assign n17283 = ( n17280 & ~n17282 ) | ( n17280 & n17281 ) | ( ~n17282 & n17281 ) ;
  assign n17287 = n16742 &  n17021 ;
  assign n17288 = n17020 &  n17287 ;
  assign n17276 = x89 | n16742 ;
  assign n17277 = x89 &  n16742 ;
  assign n17278 = ( n17276 & ~n17277 ) | ( n17276 & 1'b0 ) | ( ~n17277 & 1'b0 ) ;
  assign n17290 = ( n16950 & n17022 ) | ( n16950 & n17278 ) | ( n17022 & n17278 ) ;
  assign n17289 = n16950 | n17278 ;
  assign n17291 = ( n17288 & ~n17290 ) | ( n17288 & n17289 ) | ( ~n17290 & n17289 ) ;
  assign n17295 = n16750 &  n17021 ;
  assign n17296 = n17020 &  n17295 ;
  assign n17284 = x88 | n16750 ;
  assign n17285 = x88 &  n16750 ;
  assign n17286 = ( n17284 & ~n17285 ) | ( n17284 & 1'b0 ) | ( ~n17285 & 1'b0 ) ;
  assign n17298 = ( n16949 & n17022 ) | ( n16949 & n17286 ) | ( n17022 & n17286 ) ;
  assign n17297 = n16949 | n17286 ;
  assign n17299 = ( n17296 & ~n17298 ) | ( n17296 & n17297 ) | ( ~n17298 & n17297 ) ;
  assign n17303 = n16758 &  n17021 ;
  assign n17304 = n17020 &  n17303 ;
  assign n17292 = x87 | n16758 ;
  assign n17293 = x87 &  n16758 ;
  assign n17294 = ( n17292 & ~n17293 ) | ( n17292 & 1'b0 ) | ( ~n17293 & 1'b0 ) ;
  assign n17306 = ( n16948 & n17022 ) | ( n16948 & n17294 ) | ( n17022 & n17294 ) ;
  assign n17305 = n16948 | n17294 ;
  assign n17307 = ( n17304 & ~n17306 ) | ( n17304 & n17305 ) | ( ~n17306 & n17305 ) ;
  assign n17311 = n16766 &  n17021 ;
  assign n17312 = n17020 &  n17311 ;
  assign n17300 = x86 | n16766 ;
  assign n17301 = x86 &  n16766 ;
  assign n17302 = ( n17300 & ~n17301 ) | ( n17300 & 1'b0 ) | ( ~n17301 & 1'b0 ) ;
  assign n17314 = ( n16947 & n17022 ) | ( n16947 & n17302 ) | ( n17022 & n17302 ) ;
  assign n17313 = n16947 | n17302 ;
  assign n17315 = ( n17312 & ~n17314 ) | ( n17312 & n17313 ) | ( ~n17314 & n17313 ) ;
  assign n17319 = n16774 &  n17021 ;
  assign n17320 = n17020 &  n17319 ;
  assign n17308 = x85 | n16774 ;
  assign n17309 = x85 &  n16774 ;
  assign n17310 = ( n17308 & ~n17309 ) | ( n17308 & 1'b0 ) | ( ~n17309 & 1'b0 ) ;
  assign n17322 = ( n16946 & n17022 ) | ( n16946 & n17310 ) | ( n17022 & n17310 ) ;
  assign n17321 = n16946 | n17310 ;
  assign n17323 = ( n17320 & ~n17322 ) | ( n17320 & n17321 ) | ( ~n17322 & n17321 ) ;
  assign n17327 = n16782 &  n17021 ;
  assign n17328 = n17020 &  n17327 ;
  assign n17316 = x84 | n16782 ;
  assign n17317 = x84 &  n16782 ;
  assign n17318 = ( n17316 & ~n17317 ) | ( n17316 & 1'b0 ) | ( ~n17317 & 1'b0 ) ;
  assign n17330 = ( n16945 & n17022 ) | ( n16945 & n17318 ) | ( n17022 & n17318 ) ;
  assign n17329 = n16945 | n17318 ;
  assign n17331 = ( n17328 & ~n17330 ) | ( n17328 & n17329 ) | ( ~n17330 & n17329 ) ;
  assign n17335 = n16790 &  n17021 ;
  assign n17336 = n17020 &  n17335 ;
  assign n17324 = x83 | n16790 ;
  assign n17325 = x83 &  n16790 ;
  assign n17326 = ( n17324 & ~n17325 ) | ( n17324 & 1'b0 ) | ( ~n17325 & 1'b0 ) ;
  assign n17338 = ( n16944 & n17022 ) | ( n16944 & n17326 ) | ( n17022 & n17326 ) ;
  assign n17337 = n16944 | n17326 ;
  assign n17339 = ( n17336 & ~n17338 ) | ( n17336 & n17337 ) | ( ~n17338 & n17337 ) ;
  assign n17343 = n16798 &  n17021 ;
  assign n17344 = n17020 &  n17343 ;
  assign n17332 = x82 | n16798 ;
  assign n17333 = x82 &  n16798 ;
  assign n17334 = ( n17332 & ~n17333 ) | ( n17332 & 1'b0 ) | ( ~n17333 & 1'b0 ) ;
  assign n17346 = ( n16943 & n17022 ) | ( n16943 & n17334 ) | ( n17022 & n17334 ) ;
  assign n17345 = n16943 | n17334 ;
  assign n17347 = ( n17344 & ~n17346 ) | ( n17344 & n17345 ) | ( ~n17346 & n17345 ) ;
  assign n17351 = n16806 &  n17021 ;
  assign n17352 = n17020 &  n17351 ;
  assign n17340 = x81 | n16806 ;
  assign n17341 = x81 &  n16806 ;
  assign n17342 = ( n17340 & ~n17341 ) | ( n17340 & 1'b0 ) | ( ~n17341 & 1'b0 ) ;
  assign n17354 = ( n16942 & n17022 ) | ( n16942 & n17342 ) | ( n17022 & n17342 ) ;
  assign n17353 = n16942 | n17342 ;
  assign n17355 = ( n17352 & ~n17354 ) | ( n17352 & n17353 ) | ( ~n17354 & n17353 ) ;
  assign n17359 = n16814 &  n17021 ;
  assign n17360 = n17020 &  n17359 ;
  assign n17348 = x80 | n16814 ;
  assign n17349 = x80 &  n16814 ;
  assign n17350 = ( n17348 & ~n17349 ) | ( n17348 & 1'b0 ) | ( ~n17349 & 1'b0 ) ;
  assign n17362 = ( n16941 & n17022 ) | ( n16941 & n17350 ) | ( n17022 & n17350 ) ;
  assign n17361 = n16941 | n17350 ;
  assign n17363 = ( n17360 & ~n17362 ) | ( n17360 & n17361 ) | ( ~n17362 & n17361 ) ;
  assign n17367 = n16822 &  n17021 ;
  assign n17368 = n17020 &  n17367 ;
  assign n17356 = x79 | n16822 ;
  assign n17357 = x79 &  n16822 ;
  assign n17358 = ( n17356 & ~n17357 ) | ( n17356 & 1'b0 ) | ( ~n17357 & 1'b0 ) ;
  assign n17370 = ( n16940 & n17022 ) | ( n16940 & n17358 ) | ( n17022 & n17358 ) ;
  assign n17369 = n16940 | n17358 ;
  assign n17371 = ( n17368 & ~n17370 ) | ( n17368 & n17369 ) | ( ~n17370 & n17369 ) ;
  assign n17375 = n16830 &  n17021 ;
  assign n17376 = n17020 &  n17375 ;
  assign n17364 = x78 | n16830 ;
  assign n17365 = x78 &  n16830 ;
  assign n17366 = ( n17364 & ~n17365 ) | ( n17364 & 1'b0 ) | ( ~n17365 & 1'b0 ) ;
  assign n17378 = ( n16939 & n17022 ) | ( n16939 & n17366 ) | ( n17022 & n17366 ) ;
  assign n17377 = n16939 | n17366 ;
  assign n17379 = ( n17376 & ~n17378 ) | ( n17376 & n17377 ) | ( ~n17378 & n17377 ) ;
  assign n17383 = n16838 &  n17021 ;
  assign n17384 = n17020 &  n17383 ;
  assign n17372 = x77 | n16838 ;
  assign n17373 = x77 &  n16838 ;
  assign n17374 = ( n17372 & ~n17373 ) | ( n17372 & 1'b0 ) | ( ~n17373 & 1'b0 ) ;
  assign n17386 = ( n16938 & n17022 ) | ( n16938 & n17374 ) | ( n17022 & n17374 ) ;
  assign n17385 = n16938 | n17374 ;
  assign n17387 = ( n17384 & ~n17386 ) | ( n17384 & n17385 ) | ( ~n17386 & n17385 ) ;
  assign n17391 = n16846 &  n17021 ;
  assign n17392 = n17020 &  n17391 ;
  assign n17380 = x76 | n16846 ;
  assign n17381 = x76 &  n16846 ;
  assign n17382 = ( n17380 & ~n17381 ) | ( n17380 & 1'b0 ) | ( ~n17381 & 1'b0 ) ;
  assign n17394 = ( n16937 & n17022 ) | ( n16937 & n17382 ) | ( n17022 & n17382 ) ;
  assign n17393 = n16937 | n17382 ;
  assign n17395 = ( n17392 & ~n17394 ) | ( n17392 & n17393 ) | ( ~n17394 & n17393 ) ;
  assign n17399 = n16854 &  n17021 ;
  assign n17400 = n17020 &  n17399 ;
  assign n17388 = x75 | n16854 ;
  assign n17389 = x75 &  n16854 ;
  assign n17390 = ( n17388 & ~n17389 ) | ( n17388 & 1'b0 ) | ( ~n17389 & 1'b0 ) ;
  assign n17402 = ( n16936 & n17022 ) | ( n16936 & n17390 ) | ( n17022 & n17390 ) ;
  assign n17401 = n16936 | n17390 ;
  assign n17403 = ( n17400 & ~n17402 ) | ( n17400 & n17401 ) | ( ~n17402 & n17401 ) ;
  assign n17407 = n16862 &  n17021 ;
  assign n17408 = n17020 &  n17407 ;
  assign n17396 = x74 | n16862 ;
  assign n17397 = x74 &  n16862 ;
  assign n17398 = ( n17396 & ~n17397 ) | ( n17396 & 1'b0 ) | ( ~n17397 & 1'b0 ) ;
  assign n17410 = ( n16935 & n17022 ) | ( n16935 & n17398 ) | ( n17022 & n17398 ) ;
  assign n17409 = n16935 | n17398 ;
  assign n17411 = ( n17408 & ~n17410 ) | ( n17408 & n17409 ) | ( ~n17410 & n17409 ) ;
  assign n17415 = n16870 &  n17021 ;
  assign n17416 = n17020 &  n17415 ;
  assign n17404 = x73 | n16870 ;
  assign n17405 = x73 &  n16870 ;
  assign n17406 = ( n17404 & ~n17405 ) | ( n17404 & 1'b0 ) | ( ~n17405 & 1'b0 ) ;
  assign n17418 = ( n16934 & n17022 ) | ( n16934 & n17406 ) | ( n17022 & n17406 ) ;
  assign n17417 = n16934 | n17406 ;
  assign n17419 = ( n17416 & ~n17418 ) | ( n17416 & n17417 ) | ( ~n17418 & n17417 ) ;
  assign n17423 = n16878 &  n17021 ;
  assign n17424 = n17020 &  n17423 ;
  assign n17412 = x72 | n16878 ;
  assign n17413 = x72 &  n16878 ;
  assign n17414 = ( n17412 & ~n17413 ) | ( n17412 & 1'b0 ) | ( ~n17413 & 1'b0 ) ;
  assign n17426 = ( n16933 & n17022 ) | ( n16933 & n17414 ) | ( n17022 & n17414 ) ;
  assign n17425 = n16933 | n17414 ;
  assign n17427 = ( n17424 & ~n17426 ) | ( n17424 & n17425 ) | ( ~n17426 & n17425 ) ;
  assign n17431 = n16886 &  n17021 ;
  assign n17432 = n17020 &  n17431 ;
  assign n17420 = x71 | n16886 ;
  assign n17421 = x71 &  n16886 ;
  assign n17422 = ( n17420 & ~n17421 ) | ( n17420 & 1'b0 ) | ( ~n17421 & 1'b0 ) ;
  assign n17434 = ( n16932 & n17022 ) | ( n16932 & n17422 ) | ( n17022 & n17422 ) ;
  assign n17433 = n16932 | n17422 ;
  assign n17435 = ( n17432 & ~n17434 ) | ( n17432 & n17433 ) | ( ~n17434 & n17433 ) ;
  assign n17439 = n16894 &  n17021 ;
  assign n17440 = n17020 &  n17439 ;
  assign n17428 = x70 | n16894 ;
  assign n17429 = x70 &  n16894 ;
  assign n17430 = ( n17428 & ~n17429 ) | ( n17428 & 1'b0 ) | ( ~n17429 & 1'b0 ) ;
  assign n17442 = ( n16931 & n17022 ) | ( n16931 & n17430 ) | ( n17022 & n17430 ) ;
  assign n17441 = n16931 | n17430 ;
  assign n17443 = ( n17440 & ~n17442 ) | ( n17440 & n17441 ) | ( ~n17442 & n17441 ) ;
  assign n17447 = n16902 &  n17021 ;
  assign n17448 = n17020 &  n17447 ;
  assign n17436 = x69 | n16902 ;
  assign n17437 = x69 &  n16902 ;
  assign n17438 = ( n17436 & ~n17437 ) | ( n17436 & 1'b0 ) | ( ~n17437 & 1'b0 ) ;
  assign n17450 = ( n16930 & n17022 ) | ( n16930 & n17438 ) | ( n17022 & n17438 ) ;
  assign n17449 = n16930 | n17438 ;
  assign n17451 = ( n17448 & ~n17450 ) | ( n17448 & n17449 ) | ( ~n17450 & n17449 ) ;
  assign n17455 = n16910 &  n17021 ;
  assign n17456 = n17020 &  n17455 ;
  assign n17444 = x68 | n16910 ;
  assign n17445 = x68 &  n16910 ;
  assign n17446 = ( n17444 & ~n17445 ) | ( n17444 & 1'b0 ) | ( ~n17445 & 1'b0 ) ;
  assign n17458 = ( n16929 & n17022 ) | ( n16929 & n17446 ) | ( n17022 & n17446 ) ;
  assign n17457 = n16929 | n17446 ;
  assign n17459 = ( n17456 & ~n17458 ) | ( n17456 & n17457 ) | ( ~n17458 & n17457 ) ;
  assign n17463 = n16915 &  n17021 ;
  assign n17464 = n17020 &  n17463 ;
  assign n17452 = x67 | n16915 ;
  assign n17453 = x67 &  n16915 ;
  assign n17454 = ( n17452 & ~n17453 ) | ( n17452 & 1'b0 ) | ( ~n17453 & 1'b0 ) ;
  assign n17466 = ( n16928 & n17022 ) | ( n16928 & n17454 ) | ( n17022 & n17454 ) ;
  assign n17465 = n16928 | n17454 ;
  assign n17467 = ( n17464 & ~n17466 ) | ( n17464 & n17465 ) | ( ~n17466 & n17465 ) ;
  assign n17468 = n16921 &  n17021 ;
  assign n17469 = n17020 &  n17468 ;
  assign n17460 = x66 | n16921 ;
  assign n17461 = x66 &  n16921 ;
  assign n17462 = ( n17460 & ~n17461 ) | ( n17460 & 1'b0 ) | ( ~n17461 & 1'b0 ) ;
  assign n17470 = n16927 &  n17462 ;
  assign n17471 = ( n16927 & ~n17022 ) | ( n16927 & n17462 ) | ( ~n17022 & n17462 ) ;
  assign n17472 = ( n17469 & ~n17470 ) | ( n17469 & n17471 ) | ( ~n17470 & n17471 ) ;
  assign n17473 = ( n16925 & ~x65 ) | ( n16925 & n16926 ) | ( ~x65 & n16926 ) ;
  assign n17474 = ( n16927 & ~n16926 ) | ( n16927 & n17473 ) | ( ~n16926 & n17473 ) ;
  assign n17475 = ~n17022 & n17474 ;
  assign n17476 = n16925 &  n17021 ;
  assign n17477 = n17020 &  n17476 ;
  assign n17478 = n17475 | n17477 ;
  assign n17479 = ( x64 & ~n17022 ) | ( x64 & 1'b0 ) | ( ~n17022 & 1'b0 ) ;
  assign n17480 = ( x3 & ~n17479 ) | ( x3 & 1'b0 ) | ( ~n17479 & 1'b0 ) ;
  assign n17481 = ( n16926 & ~n17022 ) | ( n16926 & 1'b0 ) | ( ~n17022 & 1'b0 ) ;
  assign n17482 = n17480 | n17481 ;
  assign n17483 = ~x2 & x64 ;
  assign n17484 = ( x65 & ~n17482 ) | ( x65 & n17483 ) | ( ~n17482 & n17483 ) ;
  assign n17485 = ( x66 & ~n17478 ) | ( x66 & n17484 ) | ( ~n17478 & n17484 ) ;
  assign n17486 = ( x67 & ~n17472 ) | ( x67 & n17485 ) | ( ~n17472 & n17485 ) ;
  assign n17487 = ( x68 & ~n17467 ) | ( x68 & n17486 ) | ( ~n17467 & n17486 ) ;
  assign n17488 = ( x69 & ~n17459 ) | ( x69 & n17487 ) | ( ~n17459 & n17487 ) ;
  assign n17489 = ( x70 & ~n17451 ) | ( x70 & n17488 ) | ( ~n17451 & n17488 ) ;
  assign n17490 = ( x71 & ~n17443 ) | ( x71 & n17489 ) | ( ~n17443 & n17489 ) ;
  assign n17491 = ( x72 & ~n17435 ) | ( x72 & n17490 ) | ( ~n17435 & n17490 ) ;
  assign n17492 = ( x73 & ~n17427 ) | ( x73 & n17491 ) | ( ~n17427 & n17491 ) ;
  assign n17493 = ( x74 & ~n17419 ) | ( x74 & n17492 ) | ( ~n17419 & n17492 ) ;
  assign n17494 = ( x75 & ~n17411 ) | ( x75 & n17493 ) | ( ~n17411 & n17493 ) ;
  assign n17495 = ( x76 & ~n17403 ) | ( x76 & n17494 ) | ( ~n17403 & n17494 ) ;
  assign n17496 = ( x77 & ~n17395 ) | ( x77 & n17495 ) | ( ~n17395 & n17495 ) ;
  assign n17497 = ( x78 & ~n17387 ) | ( x78 & n17496 ) | ( ~n17387 & n17496 ) ;
  assign n17498 = ( x79 & ~n17379 ) | ( x79 & n17497 ) | ( ~n17379 & n17497 ) ;
  assign n17499 = ( x80 & ~n17371 ) | ( x80 & n17498 ) | ( ~n17371 & n17498 ) ;
  assign n17500 = ( x81 & ~n17363 ) | ( x81 & n17499 ) | ( ~n17363 & n17499 ) ;
  assign n17501 = ( x82 & ~n17355 ) | ( x82 & n17500 ) | ( ~n17355 & n17500 ) ;
  assign n17502 = ( x83 & ~n17347 ) | ( x83 & n17501 ) | ( ~n17347 & n17501 ) ;
  assign n17503 = ( x84 & ~n17339 ) | ( x84 & n17502 ) | ( ~n17339 & n17502 ) ;
  assign n17504 = ( x85 & ~n17331 ) | ( x85 & n17503 ) | ( ~n17331 & n17503 ) ;
  assign n17505 = ( x86 & ~n17323 ) | ( x86 & n17504 ) | ( ~n17323 & n17504 ) ;
  assign n17506 = ( x87 & ~n17315 ) | ( x87 & n17505 ) | ( ~n17315 & n17505 ) ;
  assign n17507 = ( x88 & ~n17307 ) | ( x88 & n17506 ) | ( ~n17307 & n17506 ) ;
  assign n17508 = ( x89 & ~n17299 ) | ( x89 & n17507 ) | ( ~n17299 & n17507 ) ;
  assign n17509 = ( x90 & ~n17291 ) | ( x90 & n17508 ) | ( ~n17291 & n17508 ) ;
  assign n17510 = ( x91 & ~n17283 ) | ( x91 & n17509 ) | ( ~n17283 & n17509 ) ;
  assign n17511 = ( x92 & ~n17275 ) | ( x92 & n17510 ) | ( ~n17275 & n17510 ) ;
  assign n17512 = ( x93 & ~n17267 ) | ( x93 & n17511 ) | ( ~n17267 & n17511 ) ;
  assign n17513 = ( x94 & ~n17259 ) | ( x94 & n17512 ) | ( ~n17259 & n17512 ) ;
  assign n17514 = ( x95 & ~n17251 ) | ( x95 & n17513 ) | ( ~n17251 & n17513 ) ;
  assign n17515 = ( x96 & ~n17243 ) | ( x96 & n17514 ) | ( ~n17243 & n17514 ) ;
  assign n17516 = ( x97 & ~n17235 ) | ( x97 & n17515 ) | ( ~n17235 & n17515 ) ;
  assign n17517 = ( x98 & ~n17227 ) | ( x98 & n17516 ) | ( ~n17227 & n17516 ) ;
  assign n17518 = ( x99 & ~n17219 ) | ( x99 & n17517 ) | ( ~n17219 & n17517 ) ;
  assign n17519 = ( x100 & ~n17211 ) | ( x100 & n17518 ) | ( ~n17211 & n17518 ) ;
  assign n17520 = ( x101 & ~n17203 ) | ( x101 & n17519 ) | ( ~n17203 & n17519 ) ;
  assign n17521 = ( x102 & ~n17195 ) | ( x102 & n17520 ) | ( ~n17195 & n17520 ) ;
  assign n17522 = ( x103 & ~n17187 ) | ( x103 & n17521 ) | ( ~n17187 & n17521 ) ;
  assign n17523 = ( x104 & ~n17179 ) | ( x104 & n17522 ) | ( ~n17179 & n17522 ) ;
  assign n17524 = ( x105 & ~n17171 ) | ( x105 & n17523 ) | ( ~n17171 & n17523 ) ;
  assign n17525 = ( x106 & ~n17163 ) | ( x106 & n17524 ) | ( ~n17163 & n17524 ) ;
  assign n17526 = ( x107 & ~n17155 ) | ( x107 & n17525 ) | ( ~n17155 & n17525 ) ;
  assign n17527 = ( x108 & ~n17147 ) | ( x108 & n17526 ) | ( ~n17147 & n17526 ) ;
  assign n17528 = ( x109 & ~n17139 ) | ( x109 & n17527 ) | ( ~n17139 & n17527 ) ;
  assign n17529 = ( x110 & ~n17131 ) | ( x110 & n17528 ) | ( ~n17131 & n17528 ) ;
  assign n17530 = ( x111 & ~n17123 ) | ( x111 & n17529 ) | ( ~n17123 & n17529 ) ;
  assign n17531 = ( x112 & ~n17115 ) | ( x112 & n17530 ) | ( ~n17115 & n17530 ) ;
  assign n17532 = ( x113 & ~n17107 ) | ( x113 & n17531 ) | ( ~n17107 & n17531 ) ;
  assign n17533 = ( x114 & ~n17099 ) | ( x114 & n17532 ) | ( ~n17099 & n17532 ) ;
  assign n17534 = ( x115 & ~n17091 ) | ( x115 & n17533 ) | ( ~n17091 & n17533 ) ;
  assign n17535 = ( x116 & ~n17083 ) | ( x116 & n17534 ) | ( ~n17083 & n17534 ) ;
  assign n17536 = ( x117 & ~n17075 ) | ( x117 & n17535 ) | ( ~n17075 & n17535 ) ;
  assign n17537 = ( x118 & ~n17067 ) | ( x118 & n17536 ) | ( ~n17067 & n17536 ) ;
  assign n17538 = ( x119 & ~n17059 ) | ( x119 & n17537 ) | ( ~n17059 & n17537 ) ;
  assign n17539 = ( x120 & ~n17051 ) | ( x120 & n17538 ) | ( ~n17051 & n17538 ) ;
  assign n17540 = ( x121 & ~n17043 ) | ( x121 & n17539 ) | ( ~n17043 & n17539 ) ;
  assign n17541 = ( x122 & ~n17035 ) | ( x122 & n17540 ) | ( ~n17035 & n17540 ) ;
  assign n17545 = ( x123 & ~n17027 ) | ( x123 & n17541 ) | ( ~n17027 & n17541 ) ;
  assign n17557 = ( x124 & ~n17553 ) | ( x124 & n17545 ) | ( ~n17553 & n17545 ) ;
  assign n17558 = n17015 | n17017 ;
  assign n17559 = ( n17007 & ~n17558 ) | ( n17007 & 1'b0 ) | ( ~n17558 & 1'b0 ) ;
  assign n17560 = ~n17007 & n17558 ;
  assign n17561 = ( n17559 & ~n17022 ) | ( n17559 & n17560 ) | ( ~n17022 & n17560 ) ;
  assign n17562 = n152 &  n17014 ;
  assign n17563 = n17020 &  n17562 ;
  assign n17564 = n17561 | n17563 ;
  assign n17565 = ~x125 & n17564 ;
  assign n17566 = ( x125 & ~n17563 ) | ( x125 & 1'b0 ) | ( ~n17563 & 1'b0 ) ;
  assign n17567 = ~n17561 & n17566 ;
  assign n17568 = n151 | n17567 ;
  assign n17569 = n17565 | n17568 ;
  assign n17570 = n17557 | n17569 ;
  assign n17571 = ~n17564 |  n235 ;
  assign n17573 = n17553 &  n17571 ;
  assign n17574 = n17570 &  n17573 ;
  assign n17554 = x124 | n17553 ;
  assign n17555 = x124 &  n17553 ;
  assign n17556 = ( n17554 & ~n17555 ) | ( n17554 & 1'b0 ) | ( ~n17555 & 1'b0 ) ;
  assign n17575 = n17545 &  n17556 ;
  assign n17572 = n17570 &  n17571 ;
  assign n17576 = ( n17545 & ~n17572 ) | ( n17545 & n17556 ) | ( ~n17572 & n17556 ) ;
  assign n17577 = ( n17574 & ~n17575 ) | ( n17574 & n17576 ) | ( ~n17575 & n17576 ) ;
  assign n17581 = n17027 &  n17571 ;
  assign n17582 = n17570 &  n17581 ;
  assign n17542 = x123 | n17027 ;
  assign n17543 = x123 &  n17027 ;
  assign n17544 = ( n17542 & ~n17543 ) | ( n17542 & 1'b0 ) | ( ~n17543 & 1'b0 ) ;
  assign n17584 = ( n17541 & n17544 ) | ( n17541 & n17572 ) | ( n17544 & n17572 ) ;
  assign n17583 = n17541 | n17544 ;
  assign n17585 = ( n17582 & ~n17584 ) | ( n17582 & n17583 ) | ( ~n17584 & n17583 ) ;
  assign n17589 = n17035 &  n17571 ;
  assign n17590 = n17570 &  n17589 ;
  assign n17578 = x122 | n17035 ;
  assign n17579 = x122 &  n17035 ;
  assign n17580 = ( n17578 & ~n17579 ) | ( n17578 & 1'b0 ) | ( ~n17579 & 1'b0 ) ;
  assign n17591 = n17540 &  n17580 ;
  assign n17592 = ( n17540 & ~n17572 ) | ( n17540 & n17580 ) | ( ~n17572 & n17580 ) ;
  assign n17593 = ( n17590 & ~n17591 ) | ( n17590 & n17592 ) | ( ~n17591 & n17592 ) ;
  assign n17597 = n17043 &  n17571 ;
  assign n17598 = n17570 &  n17597 ;
  assign n17586 = x121 | n17043 ;
  assign n17587 = x121 &  n17043 ;
  assign n17588 = ( n17586 & ~n17587 ) | ( n17586 & 1'b0 ) | ( ~n17587 & 1'b0 ) ;
  assign n17599 = n17539 &  n17588 ;
  assign n17600 = ( n17539 & ~n17572 ) | ( n17539 & n17588 ) | ( ~n17572 & n17588 ) ;
  assign n17601 = ( n17598 & ~n17599 ) | ( n17598 & n17600 ) | ( ~n17599 & n17600 ) ;
  assign n17605 = n17051 &  n17571 ;
  assign n17606 = n17570 &  n17605 ;
  assign n17594 = x120 | n17051 ;
  assign n17595 = x120 &  n17051 ;
  assign n17596 = ( n17594 & ~n17595 ) | ( n17594 & 1'b0 ) | ( ~n17595 & 1'b0 ) ;
  assign n17607 = n17538 &  n17596 ;
  assign n17608 = ( n17538 & ~n17572 ) | ( n17538 & n17596 ) | ( ~n17572 & n17596 ) ;
  assign n17609 = ( n17606 & ~n17607 ) | ( n17606 & n17608 ) | ( ~n17607 & n17608 ) ;
  assign n17613 = n17059 &  n17571 ;
  assign n17614 = n17570 &  n17613 ;
  assign n17602 = x119 | n17059 ;
  assign n17603 = x119 &  n17059 ;
  assign n17604 = ( n17602 & ~n17603 ) | ( n17602 & 1'b0 ) | ( ~n17603 & 1'b0 ) ;
  assign n17616 = ( n17537 & n17572 ) | ( n17537 & n17604 ) | ( n17572 & n17604 ) ;
  assign n17615 = n17537 | n17604 ;
  assign n17617 = ( n17614 & ~n17616 ) | ( n17614 & n17615 ) | ( ~n17616 & n17615 ) ;
  assign n17621 = n17067 &  n17571 ;
  assign n17622 = n17570 &  n17621 ;
  assign n17610 = x118 | n17067 ;
  assign n17611 = x118 &  n17067 ;
  assign n17612 = ( n17610 & ~n17611 ) | ( n17610 & 1'b0 ) | ( ~n17611 & 1'b0 ) ;
  assign n17624 = ( n17536 & n17572 ) | ( n17536 & n17612 ) | ( n17572 & n17612 ) ;
  assign n17623 = n17536 | n17612 ;
  assign n17625 = ( n17622 & ~n17624 ) | ( n17622 & n17623 ) | ( ~n17624 & n17623 ) ;
  assign n17629 = n17075 &  n17571 ;
  assign n17630 = n17570 &  n17629 ;
  assign n17618 = x117 | n17075 ;
  assign n17619 = x117 &  n17075 ;
  assign n17620 = ( n17618 & ~n17619 ) | ( n17618 & 1'b0 ) | ( ~n17619 & 1'b0 ) ;
  assign n17632 = ( n17535 & n17572 ) | ( n17535 & n17620 ) | ( n17572 & n17620 ) ;
  assign n17631 = n17535 | n17620 ;
  assign n17633 = ( n17630 & ~n17632 ) | ( n17630 & n17631 ) | ( ~n17632 & n17631 ) ;
  assign n17637 = n17083 &  n17571 ;
  assign n17638 = n17570 &  n17637 ;
  assign n17626 = x116 | n17083 ;
  assign n17627 = x116 &  n17083 ;
  assign n17628 = ( n17626 & ~n17627 ) | ( n17626 & 1'b0 ) | ( ~n17627 & 1'b0 ) ;
  assign n17640 = ( n17534 & n17572 ) | ( n17534 & n17628 ) | ( n17572 & n17628 ) ;
  assign n17639 = n17534 | n17628 ;
  assign n17641 = ( n17638 & ~n17640 ) | ( n17638 & n17639 ) | ( ~n17640 & n17639 ) ;
  assign n17645 = n17091 &  n17571 ;
  assign n17646 = n17570 &  n17645 ;
  assign n17634 = x115 | n17091 ;
  assign n17635 = x115 &  n17091 ;
  assign n17636 = ( n17634 & ~n17635 ) | ( n17634 & 1'b0 ) | ( ~n17635 & 1'b0 ) ;
  assign n17648 = ( n17533 & n17572 ) | ( n17533 & n17636 ) | ( n17572 & n17636 ) ;
  assign n17647 = n17533 | n17636 ;
  assign n17649 = ( n17646 & ~n17648 ) | ( n17646 & n17647 ) | ( ~n17648 & n17647 ) ;
  assign n17653 = n17099 &  n17571 ;
  assign n17654 = n17570 &  n17653 ;
  assign n17642 = x114 | n17099 ;
  assign n17643 = x114 &  n17099 ;
  assign n17644 = ( n17642 & ~n17643 ) | ( n17642 & 1'b0 ) | ( ~n17643 & 1'b0 ) ;
  assign n17656 = ( n17532 & n17572 ) | ( n17532 & n17644 ) | ( n17572 & n17644 ) ;
  assign n17655 = n17532 | n17644 ;
  assign n17657 = ( n17654 & ~n17656 ) | ( n17654 & n17655 ) | ( ~n17656 & n17655 ) ;
  assign n17661 = n17107 &  n17571 ;
  assign n17662 = n17570 &  n17661 ;
  assign n17650 = x113 | n17107 ;
  assign n17651 = x113 &  n17107 ;
  assign n17652 = ( n17650 & ~n17651 ) | ( n17650 & 1'b0 ) | ( ~n17651 & 1'b0 ) ;
  assign n17664 = ( n17531 & n17572 ) | ( n17531 & n17652 ) | ( n17572 & n17652 ) ;
  assign n17663 = n17531 | n17652 ;
  assign n17665 = ( n17662 & ~n17664 ) | ( n17662 & n17663 ) | ( ~n17664 & n17663 ) ;
  assign n17669 = n17115 &  n17571 ;
  assign n17670 = n17570 &  n17669 ;
  assign n17658 = x112 | n17115 ;
  assign n17659 = x112 &  n17115 ;
  assign n17660 = ( n17658 & ~n17659 ) | ( n17658 & 1'b0 ) | ( ~n17659 & 1'b0 ) ;
  assign n17672 = ( n17530 & n17572 ) | ( n17530 & n17660 ) | ( n17572 & n17660 ) ;
  assign n17671 = n17530 | n17660 ;
  assign n17673 = ( n17670 & ~n17672 ) | ( n17670 & n17671 ) | ( ~n17672 & n17671 ) ;
  assign n17677 = n17123 &  n17571 ;
  assign n17678 = n17570 &  n17677 ;
  assign n17666 = x111 | n17123 ;
  assign n17667 = x111 &  n17123 ;
  assign n17668 = ( n17666 & ~n17667 ) | ( n17666 & 1'b0 ) | ( ~n17667 & 1'b0 ) ;
  assign n17680 = ( n17529 & n17572 ) | ( n17529 & n17668 ) | ( n17572 & n17668 ) ;
  assign n17679 = n17529 | n17668 ;
  assign n17681 = ( n17678 & ~n17680 ) | ( n17678 & n17679 ) | ( ~n17680 & n17679 ) ;
  assign n17685 = n17131 &  n17571 ;
  assign n17686 = n17570 &  n17685 ;
  assign n17674 = x110 | n17131 ;
  assign n17675 = x110 &  n17131 ;
  assign n17676 = ( n17674 & ~n17675 ) | ( n17674 & 1'b0 ) | ( ~n17675 & 1'b0 ) ;
  assign n17688 = ( n17528 & n17572 ) | ( n17528 & n17676 ) | ( n17572 & n17676 ) ;
  assign n17687 = n17528 | n17676 ;
  assign n17689 = ( n17686 & ~n17688 ) | ( n17686 & n17687 ) | ( ~n17688 & n17687 ) ;
  assign n17693 = n17139 &  n17571 ;
  assign n17694 = n17570 &  n17693 ;
  assign n17682 = x109 | n17139 ;
  assign n17683 = x109 &  n17139 ;
  assign n17684 = ( n17682 & ~n17683 ) | ( n17682 & 1'b0 ) | ( ~n17683 & 1'b0 ) ;
  assign n17696 = ( n17527 & n17572 ) | ( n17527 & n17684 ) | ( n17572 & n17684 ) ;
  assign n17695 = n17527 | n17684 ;
  assign n17697 = ( n17694 & ~n17696 ) | ( n17694 & n17695 ) | ( ~n17696 & n17695 ) ;
  assign n17701 = n17147 &  n17571 ;
  assign n17702 = n17570 &  n17701 ;
  assign n17690 = x108 | n17147 ;
  assign n17691 = x108 &  n17147 ;
  assign n17692 = ( n17690 & ~n17691 ) | ( n17690 & 1'b0 ) | ( ~n17691 & 1'b0 ) ;
  assign n17704 = ( n17526 & n17572 ) | ( n17526 & n17692 ) | ( n17572 & n17692 ) ;
  assign n17703 = n17526 | n17692 ;
  assign n17705 = ( n17702 & ~n17704 ) | ( n17702 & n17703 ) | ( ~n17704 & n17703 ) ;
  assign n17709 = n17155 &  n17571 ;
  assign n17710 = n17570 &  n17709 ;
  assign n17698 = x107 | n17155 ;
  assign n17699 = x107 &  n17155 ;
  assign n17700 = ( n17698 & ~n17699 ) | ( n17698 & 1'b0 ) | ( ~n17699 & 1'b0 ) ;
  assign n17712 = ( n17525 & n17572 ) | ( n17525 & n17700 ) | ( n17572 & n17700 ) ;
  assign n17711 = n17525 | n17700 ;
  assign n17713 = ( n17710 & ~n17712 ) | ( n17710 & n17711 ) | ( ~n17712 & n17711 ) ;
  assign n17717 = n17163 &  n17571 ;
  assign n17718 = n17570 &  n17717 ;
  assign n17706 = x106 | n17163 ;
  assign n17707 = x106 &  n17163 ;
  assign n17708 = ( n17706 & ~n17707 ) | ( n17706 & 1'b0 ) | ( ~n17707 & 1'b0 ) ;
  assign n17720 = ( n17524 & n17572 ) | ( n17524 & n17708 ) | ( n17572 & n17708 ) ;
  assign n17719 = n17524 | n17708 ;
  assign n17721 = ( n17718 & ~n17720 ) | ( n17718 & n17719 ) | ( ~n17720 & n17719 ) ;
  assign n17725 = n17171 &  n17571 ;
  assign n17726 = n17570 &  n17725 ;
  assign n17714 = x105 | n17171 ;
  assign n17715 = x105 &  n17171 ;
  assign n17716 = ( n17714 & ~n17715 ) | ( n17714 & 1'b0 ) | ( ~n17715 & 1'b0 ) ;
  assign n17728 = ( n17523 & n17572 ) | ( n17523 & n17716 ) | ( n17572 & n17716 ) ;
  assign n17727 = n17523 | n17716 ;
  assign n17729 = ( n17726 & ~n17728 ) | ( n17726 & n17727 ) | ( ~n17728 & n17727 ) ;
  assign n17733 = n17179 &  n17571 ;
  assign n17734 = n17570 &  n17733 ;
  assign n17722 = x104 | n17179 ;
  assign n17723 = x104 &  n17179 ;
  assign n17724 = ( n17722 & ~n17723 ) | ( n17722 & 1'b0 ) | ( ~n17723 & 1'b0 ) ;
  assign n17736 = ( n17522 & n17572 ) | ( n17522 & n17724 ) | ( n17572 & n17724 ) ;
  assign n17735 = n17522 | n17724 ;
  assign n17737 = ( n17734 & ~n17736 ) | ( n17734 & n17735 ) | ( ~n17736 & n17735 ) ;
  assign n17741 = n17187 &  n17571 ;
  assign n17742 = n17570 &  n17741 ;
  assign n17730 = x103 | n17187 ;
  assign n17731 = x103 &  n17187 ;
  assign n17732 = ( n17730 & ~n17731 ) | ( n17730 & 1'b0 ) | ( ~n17731 & 1'b0 ) ;
  assign n17744 = ( n17521 & n17572 ) | ( n17521 & n17732 ) | ( n17572 & n17732 ) ;
  assign n17743 = n17521 | n17732 ;
  assign n17745 = ( n17742 & ~n17744 ) | ( n17742 & n17743 ) | ( ~n17744 & n17743 ) ;
  assign n17749 = n17195 &  n17571 ;
  assign n17750 = n17570 &  n17749 ;
  assign n17738 = x102 | n17195 ;
  assign n17739 = x102 &  n17195 ;
  assign n17740 = ( n17738 & ~n17739 ) | ( n17738 & 1'b0 ) | ( ~n17739 & 1'b0 ) ;
  assign n17752 = ( n17520 & n17572 ) | ( n17520 & n17740 ) | ( n17572 & n17740 ) ;
  assign n17751 = n17520 | n17740 ;
  assign n17753 = ( n17750 & ~n17752 ) | ( n17750 & n17751 ) | ( ~n17752 & n17751 ) ;
  assign n17757 = n17203 &  n17571 ;
  assign n17758 = n17570 &  n17757 ;
  assign n17746 = x101 | n17203 ;
  assign n17747 = x101 &  n17203 ;
  assign n17748 = ( n17746 & ~n17747 ) | ( n17746 & 1'b0 ) | ( ~n17747 & 1'b0 ) ;
  assign n17760 = ( n17519 & n17572 ) | ( n17519 & n17748 ) | ( n17572 & n17748 ) ;
  assign n17759 = n17519 | n17748 ;
  assign n17761 = ( n17758 & ~n17760 ) | ( n17758 & n17759 ) | ( ~n17760 & n17759 ) ;
  assign n17765 = n17211 &  n17571 ;
  assign n17766 = n17570 &  n17765 ;
  assign n17754 = x100 | n17211 ;
  assign n17755 = x100 &  n17211 ;
  assign n17756 = ( n17754 & ~n17755 ) | ( n17754 & 1'b0 ) | ( ~n17755 & 1'b0 ) ;
  assign n17768 = ( n17518 & n17572 ) | ( n17518 & n17756 ) | ( n17572 & n17756 ) ;
  assign n17767 = n17518 | n17756 ;
  assign n17769 = ( n17766 & ~n17768 ) | ( n17766 & n17767 ) | ( ~n17768 & n17767 ) ;
  assign n17773 = n17219 &  n17571 ;
  assign n17774 = n17570 &  n17773 ;
  assign n17762 = x99 | n17219 ;
  assign n17763 = x99 &  n17219 ;
  assign n17764 = ( n17762 & ~n17763 ) | ( n17762 & 1'b0 ) | ( ~n17763 & 1'b0 ) ;
  assign n17776 = ( n17517 & n17572 ) | ( n17517 & n17764 ) | ( n17572 & n17764 ) ;
  assign n17775 = n17517 | n17764 ;
  assign n17777 = ( n17774 & ~n17776 ) | ( n17774 & n17775 ) | ( ~n17776 & n17775 ) ;
  assign n17781 = n17227 &  n17571 ;
  assign n17782 = n17570 &  n17781 ;
  assign n17770 = x98 | n17227 ;
  assign n17771 = x98 &  n17227 ;
  assign n17772 = ( n17770 & ~n17771 ) | ( n17770 & 1'b0 ) | ( ~n17771 & 1'b0 ) ;
  assign n17784 = ( n17516 & n17572 ) | ( n17516 & n17772 ) | ( n17572 & n17772 ) ;
  assign n17783 = n17516 | n17772 ;
  assign n17785 = ( n17782 & ~n17784 ) | ( n17782 & n17783 ) | ( ~n17784 & n17783 ) ;
  assign n17789 = n17235 &  n17571 ;
  assign n17790 = n17570 &  n17789 ;
  assign n17778 = x97 | n17235 ;
  assign n17779 = x97 &  n17235 ;
  assign n17780 = ( n17778 & ~n17779 ) | ( n17778 & 1'b0 ) | ( ~n17779 & 1'b0 ) ;
  assign n17792 = ( n17515 & n17572 ) | ( n17515 & n17780 ) | ( n17572 & n17780 ) ;
  assign n17791 = n17515 | n17780 ;
  assign n17793 = ( n17790 & ~n17792 ) | ( n17790 & n17791 ) | ( ~n17792 & n17791 ) ;
  assign n17797 = n17243 &  n17571 ;
  assign n17798 = n17570 &  n17797 ;
  assign n17786 = x96 | n17243 ;
  assign n17787 = x96 &  n17243 ;
  assign n17788 = ( n17786 & ~n17787 ) | ( n17786 & 1'b0 ) | ( ~n17787 & 1'b0 ) ;
  assign n17800 = ( n17514 & n17572 ) | ( n17514 & n17788 ) | ( n17572 & n17788 ) ;
  assign n17799 = n17514 | n17788 ;
  assign n17801 = ( n17798 & ~n17800 ) | ( n17798 & n17799 ) | ( ~n17800 & n17799 ) ;
  assign n17805 = n17251 &  n17571 ;
  assign n17806 = n17570 &  n17805 ;
  assign n17794 = x95 | n17251 ;
  assign n17795 = x95 &  n17251 ;
  assign n17796 = ( n17794 & ~n17795 ) | ( n17794 & 1'b0 ) | ( ~n17795 & 1'b0 ) ;
  assign n17808 = ( n17513 & n17572 ) | ( n17513 & n17796 ) | ( n17572 & n17796 ) ;
  assign n17807 = n17513 | n17796 ;
  assign n17809 = ( n17806 & ~n17808 ) | ( n17806 & n17807 ) | ( ~n17808 & n17807 ) ;
  assign n17813 = n17259 &  n17571 ;
  assign n17814 = n17570 &  n17813 ;
  assign n17802 = x94 | n17259 ;
  assign n17803 = x94 &  n17259 ;
  assign n17804 = ( n17802 & ~n17803 ) | ( n17802 & 1'b0 ) | ( ~n17803 & 1'b0 ) ;
  assign n17816 = ( n17512 & n17572 ) | ( n17512 & n17804 ) | ( n17572 & n17804 ) ;
  assign n17815 = n17512 | n17804 ;
  assign n17817 = ( n17814 & ~n17816 ) | ( n17814 & n17815 ) | ( ~n17816 & n17815 ) ;
  assign n17821 = n17267 &  n17571 ;
  assign n17822 = n17570 &  n17821 ;
  assign n17810 = x93 | n17267 ;
  assign n17811 = x93 &  n17267 ;
  assign n17812 = ( n17810 & ~n17811 ) | ( n17810 & 1'b0 ) | ( ~n17811 & 1'b0 ) ;
  assign n17824 = ( n17511 & n17572 ) | ( n17511 & n17812 ) | ( n17572 & n17812 ) ;
  assign n17823 = n17511 | n17812 ;
  assign n17825 = ( n17822 & ~n17824 ) | ( n17822 & n17823 ) | ( ~n17824 & n17823 ) ;
  assign n17829 = n17275 &  n17571 ;
  assign n17830 = n17570 &  n17829 ;
  assign n17818 = x92 | n17275 ;
  assign n17819 = x92 &  n17275 ;
  assign n17820 = ( n17818 & ~n17819 ) | ( n17818 & 1'b0 ) | ( ~n17819 & 1'b0 ) ;
  assign n17832 = ( n17510 & n17572 ) | ( n17510 & n17820 ) | ( n17572 & n17820 ) ;
  assign n17831 = n17510 | n17820 ;
  assign n17833 = ( n17830 & ~n17832 ) | ( n17830 & n17831 ) | ( ~n17832 & n17831 ) ;
  assign n17837 = n17283 &  n17571 ;
  assign n17838 = n17570 &  n17837 ;
  assign n17826 = x91 | n17283 ;
  assign n17827 = x91 &  n17283 ;
  assign n17828 = ( n17826 & ~n17827 ) | ( n17826 & 1'b0 ) | ( ~n17827 & 1'b0 ) ;
  assign n17840 = ( n17509 & n17572 ) | ( n17509 & n17828 ) | ( n17572 & n17828 ) ;
  assign n17839 = n17509 | n17828 ;
  assign n17841 = ( n17838 & ~n17840 ) | ( n17838 & n17839 ) | ( ~n17840 & n17839 ) ;
  assign n17845 = n17291 &  n17571 ;
  assign n17846 = n17570 &  n17845 ;
  assign n17834 = x90 | n17291 ;
  assign n17835 = x90 &  n17291 ;
  assign n17836 = ( n17834 & ~n17835 ) | ( n17834 & 1'b0 ) | ( ~n17835 & 1'b0 ) ;
  assign n17848 = ( n17508 & n17572 ) | ( n17508 & n17836 ) | ( n17572 & n17836 ) ;
  assign n17847 = n17508 | n17836 ;
  assign n17849 = ( n17846 & ~n17848 ) | ( n17846 & n17847 ) | ( ~n17848 & n17847 ) ;
  assign n17853 = n17299 &  n17571 ;
  assign n17854 = n17570 &  n17853 ;
  assign n17842 = x89 | n17299 ;
  assign n17843 = x89 &  n17299 ;
  assign n17844 = ( n17842 & ~n17843 ) | ( n17842 & 1'b0 ) | ( ~n17843 & 1'b0 ) ;
  assign n17856 = ( n17507 & n17572 ) | ( n17507 & n17844 ) | ( n17572 & n17844 ) ;
  assign n17855 = n17507 | n17844 ;
  assign n17857 = ( n17854 & ~n17856 ) | ( n17854 & n17855 ) | ( ~n17856 & n17855 ) ;
  assign n17861 = n17307 &  n17571 ;
  assign n17862 = n17570 &  n17861 ;
  assign n17850 = x88 | n17307 ;
  assign n17851 = x88 &  n17307 ;
  assign n17852 = ( n17850 & ~n17851 ) | ( n17850 & 1'b0 ) | ( ~n17851 & 1'b0 ) ;
  assign n17864 = ( n17506 & n17572 ) | ( n17506 & n17852 ) | ( n17572 & n17852 ) ;
  assign n17863 = n17506 | n17852 ;
  assign n17865 = ( n17862 & ~n17864 ) | ( n17862 & n17863 ) | ( ~n17864 & n17863 ) ;
  assign n17869 = n17315 &  n17571 ;
  assign n17870 = n17570 &  n17869 ;
  assign n17858 = x87 | n17315 ;
  assign n17859 = x87 &  n17315 ;
  assign n17860 = ( n17858 & ~n17859 ) | ( n17858 & 1'b0 ) | ( ~n17859 & 1'b0 ) ;
  assign n17872 = ( n17505 & n17572 ) | ( n17505 & n17860 ) | ( n17572 & n17860 ) ;
  assign n17871 = n17505 | n17860 ;
  assign n17873 = ( n17870 & ~n17872 ) | ( n17870 & n17871 ) | ( ~n17872 & n17871 ) ;
  assign n17877 = n17323 &  n17571 ;
  assign n17878 = n17570 &  n17877 ;
  assign n17866 = x86 | n17323 ;
  assign n17867 = x86 &  n17323 ;
  assign n17868 = ( n17866 & ~n17867 ) | ( n17866 & 1'b0 ) | ( ~n17867 & 1'b0 ) ;
  assign n17880 = ( n17504 & n17572 ) | ( n17504 & n17868 ) | ( n17572 & n17868 ) ;
  assign n17879 = n17504 | n17868 ;
  assign n17881 = ( n17878 & ~n17880 ) | ( n17878 & n17879 ) | ( ~n17880 & n17879 ) ;
  assign n17885 = n17331 &  n17571 ;
  assign n17886 = n17570 &  n17885 ;
  assign n17874 = x85 | n17331 ;
  assign n17875 = x85 &  n17331 ;
  assign n17876 = ( n17874 & ~n17875 ) | ( n17874 & 1'b0 ) | ( ~n17875 & 1'b0 ) ;
  assign n17888 = ( n17503 & n17572 ) | ( n17503 & n17876 ) | ( n17572 & n17876 ) ;
  assign n17887 = n17503 | n17876 ;
  assign n17889 = ( n17886 & ~n17888 ) | ( n17886 & n17887 ) | ( ~n17888 & n17887 ) ;
  assign n17893 = n17339 &  n17571 ;
  assign n17894 = n17570 &  n17893 ;
  assign n17882 = x84 | n17339 ;
  assign n17883 = x84 &  n17339 ;
  assign n17884 = ( n17882 & ~n17883 ) | ( n17882 & 1'b0 ) | ( ~n17883 & 1'b0 ) ;
  assign n17896 = ( n17502 & n17572 ) | ( n17502 & n17884 ) | ( n17572 & n17884 ) ;
  assign n17895 = n17502 | n17884 ;
  assign n17897 = ( n17894 & ~n17896 ) | ( n17894 & n17895 ) | ( ~n17896 & n17895 ) ;
  assign n17901 = n17347 &  n17571 ;
  assign n17902 = n17570 &  n17901 ;
  assign n17890 = x83 | n17347 ;
  assign n17891 = x83 &  n17347 ;
  assign n17892 = ( n17890 & ~n17891 ) | ( n17890 & 1'b0 ) | ( ~n17891 & 1'b0 ) ;
  assign n17904 = ( n17501 & n17572 ) | ( n17501 & n17892 ) | ( n17572 & n17892 ) ;
  assign n17903 = n17501 | n17892 ;
  assign n17905 = ( n17902 & ~n17904 ) | ( n17902 & n17903 ) | ( ~n17904 & n17903 ) ;
  assign n17909 = n17355 &  n17571 ;
  assign n17910 = n17570 &  n17909 ;
  assign n17898 = x82 | n17355 ;
  assign n17899 = x82 &  n17355 ;
  assign n17900 = ( n17898 & ~n17899 ) | ( n17898 & 1'b0 ) | ( ~n17899 & 1'b0 ) ;
  assign n17912 = ( n17500 & n17572 ) | ( n17500 & n17900 ) | ( n17572 & n17900 ) ;
  assign n17911 = n17500 | n17900 ;
  assign n17913 = ( n17910 & ~n17912 ) | ( n17910 & n17911 ) | ( ~n17912 & n17911 ) ;
  assign n17917 = n17363 &  n17571 ;
  assign n17918 = n17570 &  n17917 ;
  assign n17906 = x81 | n17363 ;
  assign n17907 = x81 &  n17363 ;
  assign n17908 = ( n17906 & ~n17907 ) | ( n17906 & 1'b0 ) | ( ~n17907 & 1'b0 ) ;
  assign n17920 = ( n17499 & n17572 ) | ( n17499 & n17908 ) | ( n17572 & n17908 ) ;
  assign n17919 = n17499 | n17908 ;
  assign n17921 = ( n17918 & ~n17920 ) | ( n17918 & n17919 ) | ( ~n17920 & n17919 ) ;
  assign n17925 = n17371 &  n17571 ;
  assign n17926 = n17570 &  n17925 ;
  assign n17914 = x80 | n17371 ;
  assign n17915 = x80 &  n17371 ;
  assign n17916 = ( n17914 & ~n17915 ) | ( n17914 & 1'b0 ) | ( ~n17915 & 1'b0 ) ;
  assign n17928 = ( n17498 & n17572 ) | ( n17498 & n17916 ) | ( n17572 & n17916 ) ;
  assign n17927 = n17498 | n17916 ;
  assign n17929 = ( n17926 & ~n17928 ) | ( n17926 & n17927 ) | ( ~n17928 & n17927 ) ;
  assign n17933 = n17379 &  n17571 ;
  assign n17934 = n17570 &  n17933 ;
  assign n17922 = x79 | n17379 ;
  assign n17923 = x79 &  n17379 ;
  assign n17924 = ( n17922 & ~n17923 ) | ( n17922 & 1'b0 ) | ( ~n17923 & 1'b0 ) ;
  assign n17936 = ( n17497 & n17572 ) | ( n17497 & n17924 ) | ( n17572 & n17924 ) ;
  assign n17935 = n17497 | n17924 ;
  assign n17937 = ( n17934 & ~n17936 ) | ( n17934 & n17935 ) | ( ~n17936 & n17935 ) ;
  assign n17941 = n17387 &  n17571 ;
  assign n17942 = n17570 &  n17941 ;
  assign n17930 = x78 | n17387 ;
  assign n17931 = x78 &  n17387 ;
  assign n17932 = ( n17930 & ~n17931 ) | ( n17930 & 1'b0 ) | ( ~n17931 & 1'b0 ) ;
  assign n17944 = ( n17496 & n17572 ) | ( n17496 & n17932 ) | ( n17572 & n17932 ) ;
  assign n17943 = n17496 | n17932 ;
  assign n17945 = ( n17942 & ~n17944 ) | ( n17942 & n17943 ) | ( ~n17944 & n17943 ) ;
  assign n17949 = n17395 &  n17571 ;
  assign n17950 = n17570 &  n17949 ;
  assign n17938 = x77 | n17395 ;
  assign n17939 = x77 &  n17395 ;
  assign n17940 = ( n17938 & ~n17939 ) | ( n17938 & 1'b0 ) | ( ~n17939 & 1'b0 ) ;
  assign n17952 = ( n17495 & n17572 ) | ( n17495 & n17940 ) | ( n17572 & n17940 ) ;
  assign n17951 = n17495 | n17940 ;
  assign n17953 = ( n17950 & ~n17952 ) | ( n17950 & n17951 ) | ( ~n17952 & n17951 ) ;
  assign n17957 = n17403 &  n17571 ;
  assign n17958 = n17570 &  n17957 ;
  assign n17946 = x76 | n17403 ;
  assign n17947 = x76 &  n17403 ;
  assign n17948 = ( n17946 & ~n17947 ) | ( n17946 & 1'b0 ) | ( ~n17947 & 1'b0 ) ;
  assign n17960 = ( n17494 & n17572 ) | ( n17494 & n17948 ) | ( n17572 & n17948 ) ;
  assign n17959 = n17494 | n17948 ;
  assign n17961 = ( n17958 & ~n17960 ) | ( n17958 & n17959 ) | ( ~n17960 & n17959 ) ;
  assign n17965 = n17411 &  n17571 ;
  assign n17966 = n17570 &  n17965 ;
  assign n17954 = x75 | n17411 ;
  assign n17955 = x75 &  n17411 ;
  assign n17956 = ( n17954 & ~n17955 ) | ( n17954 & 1'b0 ) | ( ~n17955 & 1'b0 ) ;
  assign n17968 = ( n17493 & n17572 ) | ( n17493 & n17956 ) | ( n17572 & n17956 ) ;
  assign n17967 = n17493 | n17956 ;
  assign n17969 = ( n17966 & ~n17968 ) | ( n17966 & n17967 ) | ( ~n17968 & n17967 ) ;
  assign n17973 = n17419 &  n17571 ;
  assign n17974 = n17570 &  n17973 ;
  assign n17962 = x74 | n17419 ;
  assign n17963 = x74 &  n17419 ;
  assign n17964 = ( n17962 & ~n17963 ) | ( n17962 & 1'b0 ) | ( ~n17963 & 1'b0 ) ;
  assign n17976 = ( n17492 & n17572 ) | ( n17492 & n17964 ) | ( n17572 & n17964 ) ;
  assign n17975 = n17492 | n17964 ;
  assign n17977 = ( n17974 & ~n17976 ) | ( n17974 & n17975 ) | ( ~n17976 & n17975 ) ;
  assign n17981 = n17427 &  n17571 ;
  assign n17982 = n17570 &  n17981 ;
  assign n17970 = x73 | n17427 ;
  assign n17971 = x73 &  n17427 ;
  assign n17972 = ( n17970 & ~n17971 ) | ( n17970 & 1'b0 ) | ( ~n17971 & 1'b0 ) ;
  assign n17984 = ( n17491 & n17572 ) | ( n17491 & n17972 ) | ( n17572 & n17972 ) ;
  assign n17983 = n17491 | n17972 ;
  assign n17985 = ( n17982 & ~n17984 ) | ( n17982 & n17983 ) | ( ~n17984 & n17983 ) ;
  assign n17989 = n17435 &  n17571 ;
  assign n17990 = n17570 &  n17989 ;
  assign n17978 = x72 | n17435 ;
  assign n17979 = x72 &  n17435 ;
  assign n17980 = ( n17978 & ~n17979 ) | ( n17978 & 1'b0 ) | ( ~n17979 & 1'b0 ) ;
  assign n17992 = ( n17490 & n17572 ) | ( n17490 & n17980 ) | ( n17572 & n17980 ) ;
  assign n17991 = n17490 | n17980 ;
  assign n17993 = ( n17990 & ~n17992 ) | ( n17990 & n17991 ) | ( ~n17992 & n17991 ) ;
  assign n17997 = n17443 &  n17571 ;
  assign n17998 = n17570 &  n17997 ;
  assign n17986 = x71 | n17443 ;
  assign n17987 = x71 &  n17443 ;
  assign n17988 = ( n17986 & ~n17987 ) | ( n17986 & 1'b0 ) | ( ~n17987 & 1'b0 ) ;
  assign n18000 = ( n17489 & n17572 ) | ( n17489 & n17988 ) | ( n17572 & n17988 ) ;
  assign n17999 = n17489 | n17988 ;
  assign n18001 = ( n17998 & ~n18000 ) | ( n17998 & n17999 ) | ( ~n18000 & n17999 ) ;
  assign n18005 = n17451 &  n17571 ;
  assign n18006 = n17570 &  n18005 ;
  assign n17994 = x70 | n17451 ;
  assign n17995 = x70 &  n17451 ;
  assign n17996 = ( n17994 & ~n17995 ) | ( n17994 & 1'b0 ) | ( ~n17995 & 1'b0 ) ;
  assign n18008 = ( n17488 & n17572 ) | ( n17488 & n17996 ) | ( n17572 & n17996 ) ;
  assign n18007 = n17488 | n17996 ;
  assign n18009 = ( n18006 & ~n18008 ) | ( n18006 & n18007 ) | ( ~n18008 & n18007 ) ;
  assign n18013 = n17459 &  n17571 ;
  assign n18014 = n17570 &  n18013 ;
  assign n18002 = x69 | n17459 ;
  assign n18003 = x69 &  n17459 ;
  assign n18004 = ( n18002 & ~n18003 ) | ( n18002 & 1'b0 ) | ( ~n18003 & 1'b0 ) ;
  assign n18016 = ( n17487 & n17572 ) | ( n17487 & n18004 ) | ( n17572 & n18004 ) ;
  assign n18015 = n17487 | n18004 ;
  assign n18017 = ( n18014 & ~n18016 ) | ( n18014 & n18015 ) | ( ~n18016 & n18015 ) ;
  assign n18021 = n17467 &  n17571 ;
  assign n18022 = n17570 &  n18021 ;
  assign n18010 = x68 | n17467 ;
  assign n18011 = x68 &  n17467 ;
  assign n18012 = ( n18010 & ~n18011 ) | ( n18010 & 1'b0 ) | ( ~n18011 & 1'b0 ) ;
  assign n18024 = ( n17486 & n17572 ) | ( n17486 & n18012 ) | ( n17572 & n18012 ) ;
  assign n18023 = n17486 | n18012 ;
  assign n18025 = ( n18022 & ~n18024 ) | ( n18022 & n18023 ) | ( ~n18024 & n18023 ) ;
  assign n18029 = n17472 &  n17571 ;
  assign n18030 = n17570 &  n18029 ;
  assign n18018 = x67 | n17472 ;
  assign n18019 = x67 &  n17472 ;
  assign n18020 = ( n18018 & ~n18019 ) | ( n18018 & 1'b0 ) | ( ~n18019 & 1'b0 ) ;
  assign n18032 = ( n17485 & n17572 ) | ( n17485 & n18020 ) | ( n17572 & n18020 ) ;
  assign n18031 = n17485 | n18020 ;
  assign n18033 = ( n18030 & ~n18032 ) | ( n18030 & n18031 ) | ( ~n18032 & n18031 ) ;
  assign n18034 = n17478 &  n17571 ;
  assign n18035 = n17570 &  n18034 ;
  assign n18026 = x66 | n17478 ;
  assign n18027 = x66 &  n17478 ;
  assign n18028 = ( n18026 & ~n18027 ) | ( n18026 & 1'b0 ) | ( ~n18027 & 1'b0 ) ;
  assign n18036 = n17484 &  n18028 ;
  assign n18037 = ( n17484 & ~n17572 ) | ( n17484 & n18028 ) | ( ~n17572 & n18028 ) ;
  assign n18038 = ( n18035 & ~n18036 ) | ( n18035 & n18037 ) | ( ~n18036 & n18037 ) ;
  assign n18039 = ( n17482 & ~x65 ) | ( n17482 & n17483 ) | ( ~x65 & n17483 ) ;
  assign n18040 = ( n17484 & ~n17483 ) | ( n17484 & n18039 ) | ( ~n17483 & n18039 ) ;
  assign n18041 = ~n17572 & n18040 ;
  assign n18042 = n17482 &  n17571 ;
  assign n18043 = n17570 &  n18042 ;
  assign n18044 = n18041 | n18043 ;
  assign n18045 = ( x64 & ~n17572 ) | ( x64 & 1'b0 ) | ( ~n17572 & 1'b0 ) ;
  assign n18046 = ( x2 & ~n18045 ) | ( x2 & 1'b0 ) | ( ~n18045 & 1'b0 ) ;
  assign n18047 = ( n17483 & ~n17572 ) | ( n17483 & 1'b0 ) | ( ~n17572 & 1'b0 ) ;
  assign n18048 = n18046 | n18047 ;
  assign n18049 = ~x1 & x64 ;
  assign n18050 = ( x65 & ~n18048 ) | ( x65 & n18049 ) | ( ~n18048 & n18049 ) ;
  assign n18051 = ( x66 & ~n18044 ) | ( x66 & n18050 ) | ( ~n18044 & n18050 ) ;
  assign n18052 = ( x67 & ~n18038 ) | ( x67 & n18051 ) | ( ~n18038 & n18051 ) ;
  assign n18053 = ( x68 & ~n18033 ) | ( x68 & n18052 ) | ( ~n18033 & n18052 ) ;
  assign n18054 = ( x69 & ~n18025 ) | ( x69 & n18053 ) | ( ~n18025 & n18053 ) ;
  assign n18055 = ( x70 & ~n18017 ) | ( x70 & n18054 ) | ( ~n18017 & n18054 ) ;
  assign n18056 = ( x71 & ~n18009 ) | ( x71 & n18055 ) | ( ~n18009 & n18055 ) ;
  assign n18057 = ( x72 & ~n18001 ) | ( x72 & n18056 ) | ( ~n18001 & n18056 ) ;
  assign n18058 = ( x73 & ~n17993 ) | ( x73 & n18057 ) | ( ~n17993 & n18057 ) ;
  assign n18059 = ( x74 & ~n17985 ) | ( x74 & n18058 ) | ( ~n17985 & n18058 ) ;
  assign n18060 = ( x75 & ~n17977 ) | ( x75 & n18059 ) | ( ~n17977 & n18059 ) ;
  assign n18061 = ( x76 & ~n17969 ) | ( x76 & n18060 ) | ( ~n17969 & n18060 ) ;
  assign n18062 = ( x77 & ~n17961 ) | ( x77 & n18061 ) | ( ~n17961 & n18061 ) ;
  assign n18063 = ( x78 & ~n17953 ) | ( x78 & n18062 ) | ( ~n17953 & n18062 ) ;
  assign n18064 = ( x79 & ~n17945 ) | ( x79 & n18063 ) | ( ~n17945 & n18063 ) ;
  assign n18065 = ( x80 & ~n17937 ) | ( x80 & n18064 ) | ( ~n17937 & n18064 ) ;
  assign n18066 = ( x81 & ~n17929 ) | ( x81 & n18065 ) | ( ~n17929 & n18065 ) ;
  assign n18067 = ( x82 & ~n17921 ) | ( x82 & n18066 ) | ( ~n17921 & n18066 ) ;
  assign n18068 = ( x83 & ~n17913 ) | ( x83 & n18067 ) | ( ~n17913 & n18067 ) ;
  assign n18069 = ( x84 & ~n17905 ) | ( x84 & n18068 ) | ( ~n17905 & n18068 ) ;
  assign n18070 = ( x85 & ~n17897 ) | ( x85 & n18069 ) | ( ~n17897 & n18069 ) ;
  assign n18071 = ( x86 & ~n17889 ) | ( x86 & n18070 ) | ( ~n17889 & n18070 ) ;
  assign n18072 = ( x87 & ~n17881 ) | ( x87 & n18071 ) | ( ~n17881 & n18071 ) ;
  assign n18073 = ( x88 & ~n17873 ) | ( x88 & n18072 ) | ( ~n17873 & n18072 ) ;
  assign n18074 = ( x89 & ~n17865 ) | ( x89 & n18073 ) | ( ~n17865 & n18073 ) ;
  assign n18075 = ( x90 & ~n17857 ) | ( x90 & n18074 ) | ( ~n17857 & n18074 ) ;
  assign n18076 = ( x91 & ~n17849 ) | ( x91 & n18075 ) | ( ~n17849 & n18075 ) ;
  assign n18077 = ( x92 & ~n17841 ) | ( x92 & n18076 ) | ( ~n17841 & n18076 ) ;
  assign n18078 = ( x93 & ~n17833 ) | ( x93 & n18077 ) | ( ~n17833 & n18077 ) ;
  assign n18079 = ( x94 & ~n17825 ) | ( x94 & n18078 ) | ( ~n17825 & n18078 ) ;
  assign n18080 = ( x95 & ~n17817 ) | ( x95 & n18079 ) | ( ~n17817 & n18079 ) ;
  assign n18081 = ( x96 & ~n17809 ) | ( x96 & n18080 ) | ( ~n17809 & n18080 ) ;
  assign n18082 = ( x97 & ~n17801 ) | ( x97 & n18081 ) | ( ~n17801 & n18081 ) ;
  assign n18083 = ( x98 & ~n17793 ) | ( x98 & n18082 ) | ( ~n17793 & n18082 ) ;
  assign n18084 = ( x99 & ~n17785 ) | ( x99 & n18083 ) | ( ~n17785 & n18083 ) ;
  assign n18085 = ( x100 & ~n17777 ) | ( x100 & n18084 ) | ( ~n17777 & n18084 ) ;
  assign n18086 = ( x101 & ~n17769 ) | ( x101 & n18085 ) | ( ~n17769 & n18085 ) ;
  assign n18087 = ( x102 & ~n17761 ) | ( x102 & n18086 ) | ( ~n17761 & n18086 ) ;
  assign n18088 = ( x103 & ~n17753 ) | ( x103 & n18087 ) | ( ~n17753 & n18087 ) ;
  assign n18089 = ( x104 & ~n17745 ) | ( x104 & n18088 ) | ( ~n17745 & n18088 ) ;
  assign n18090 = ( x105 & ~n17737 ) | ( x105 & n18089 ) | ( ~n17737 & n18089 ) ;
  assign n18091 = ( x106 & ~n17729 ) | ( x106 & n18090 ) | ( ~n17729 & n18090 ) ;
  assign n18092 = ( x107 & ~n17721 ) | ( x107 & n18091 ) | ( ~n17721 & n18091 ) ;
  assign n18093 = ( x108 & ~n17713 ) | ( x108 & n18092 ) | ( ~n17713 & n18092 ) ;
  assign n18094 = ( x109 & ~n17705 ) | ( x109 & n18093 ) | ( ~n17705 & n18093 ) ;
  assign n18095 = ( x110 & ~n17697 ) | ( x110 & n18094 ) | ( ~n17697 & n18094 ) ;
  assign n18096 = ( x111 & ~n17689 ) | ( x111 & n18095 ) | ( ~n17689 & n18095 ) ;
  assign n18097 = ( x112 & ~n17681 ) | ( x112 & n18096 ) | ( ~n17681 & n18096 ) ;
  assign n18098 = ( x113 & ~n17673 ) | ( x113 & n18097 ) | ( ~n17673 & n18097 ) ;
  assign n18099 = ( x114 & ~n17665 ) | ( x114 & n18098 ) | ( ~n17665 & n18098 ) ;
  assign n18100 = ( x115 & ~n17657 ) | ( x115 & n18099 ) | ( ~n17657 & n18099 ) ;
  assign n18101 = ( x116 & ~n17649 ) | ( x116 & n18100 ) | ( ~n17649 & n18100 ) ;
  assign n18102 = ( x117 & ~n17641 ) | ( x117 & n18101 ) | ( ~n17641 & n18101 ) ;
  assign n18103 = ( x118 & ~n17633 ) | ( x118 & n18102 ) | ( ~n17633 & n18102 ) ;
  assign n18104 = ( x119 & ~n17625 ) | ( x119 & n18103 ) | ( ~n17625 & n18103 ) ;
  assign n18105 = ( x120 & ~n17617 ) | ( x120 & n18104 ) | ( ~n17617 & n18104 ) ;
  assign n18106 = ( x121 & ~n17609 ) | ( x121 & n18105 ) | ( ~n17609 & n18105 ) ;
  assign n18107 = ( x122 & ~n17601 ) | ( x122 & n18106 ) | ( ~n17601 & n18106 ) ;
  assign n18108 = ( x123 & ~n17593 ) | ( x123 & n18107 ) | ( ~n17593 & n18107 ) ;
  assign n18109 = ( x124 & ~n17585 ) | ( x124 & n18108 ) | ( ~n17585 & n18108 ) ;
  assign n18110 = ( x125 & ~n17577 ) | ( x125 & n18109 ) | ( ~n17577 & n18109 ) ;
  assign n18111 = n17565 | n17567 ;
  assign n18112 = ( n17557 & ~n18111 ) | ( n17557 & 1'b0 ) | ( ~n18111 & 1'b0 ) ;
  assign n18113 = ~n17557 & n18111 ;
  assign n18114 = ( n18112 & ~n17572 ) | ( n18112 & n18113 ) | ( ~n17572 & n18113 ) ;
  assign n18115 = n235 &  n17564 ;
  assign n18116 = n17570 &  n18115 ;
  assign n18117 = n18114 | n18116 ;
  assign n18118 = ~x126 & n18117 ;
  assign n18119 = ( x126 & ~n18116 ) | ( x126 & 1'b0 ) | ( ~n18116 & 1'b0 ) ;
  assign n18120 = ~n18114 & n18119 ;
  assign n18121 = x127 | n18120 ;
  assign n18122 = n18118 | n18121 ;
  assign n18123 = n18110 | n18122 ;
  assign n18130 = n151 &  n18117 ;
  assign n18131 = n18123 &  n18130 ;
  assign n18124 = ~n18117 |  n151 ;
  assign n18125 = n18123 &  n18124 ;
  assign n18129 = n18118 | n18120 ;
  assign n18133 = ( n18110 & n18125 ) | ( n18110 & n18129 ) | ( n18125 & n18129 ) ;
  assign n18132 = n18110 | n18129 ;
  assign n18134 = ( n18131 & ~n18133 ) | ( n18131 & n18132 ) | ( ~n18133 & n18132 ) ;
  assign n18997 = n17585 &  n18124 ;
  assign n18998 = n18123 &  n18997 ;
  assign n18994 = x124 | n17585 ;
  assign n18995 = x124 &  n17585 ;
  assign n18996 = ( n18994 & ~n18995 ) | ( n18994 & 1'b0 ) | ( ~n18995 & 1'b0 ) ;
  assign n18999 = n18108 &  n18996 ;
  assign n19000 = ( n18108 & ~n18125 ) | ( n18108 & n18996 ) | ( ~n18125 & n18996 ) ;
  assign n19001 = ( n18998 & ~n18999 ) | ( n18998 & n19000 ) | ( ~n18999 & n19000 ) ;
  assign n18985 = n17593 &  n18124 ;
  assign n18986 = n18123 &  n18985 ;
  assign n18982 = x123 | n17593 ;
  assign n18983 = x123 &  n17593 ;
  assign n18984 = ( n18982 & ~n18983 ) | ( n18982 & 1'b0 ) | ( ~n18983 & 1'b0 ) ;
  assign n18987 = n18107 &  n18984 ;
  assign n18988 = ( n18107 & ~n18125 ) | ( n18107 & n18984 ) | ( ~n18125 & n18984 ) ;
  assign n18989 = ( n18986 & ~n18987 ) | ( n18986 & n18988 ) | ( ~n18987 & n18988 ) ;
  assign n18968 = n17601 &  n18124 ;
  assign n18969 = n18123 &  n18968 ;
  assign n18965 = x122 | n17601 ;
  assign n18966 = x122 &  n17601 ;
  assign n18967 = ( n18965 & ~n18966 ) | ( n18965 & 1'b0 ) | ( ~n18966 & 1'b0 ) ;
  assign n18970 = n18106 &  n18967 ;
  assign n18971 = ( n18106 & ~n18125 ) | ( n18106 & n18967 ) | ( ~n18125 & n18967 ) ;
  assign n18972 = ( n18969 & ~n18970 ) | ( n18969 & n18971 ) | ( ~n18970 & n18971 ) ;
  assign n18956 = n17609 &  n18124 ;
  assign n18957 = n18123 &  n18956 ;
  assign n18953 = x121 | n17609 ;
  assign n18954 = x121 &  n17609 ;
  assign n18955 = ( n18953 & ~n18954 ) | ( n18953 & 1'b0 ) | ( ~n18954 & 1'b0 ) ;
  assign n18958 = n18105 &  n18955 ;
  assign n18959 = ( n18105 & ~n18125 ) | ( n18105 & n18955 ) | ( ~n18125 & n18955 ) ;
  assign n18960 = ( n18957 & ~n18958 ) | ( n18957 & n18959 ) | ( ~n18958 & n18959 ) ;
  assign n18939 = n17617 &  n18124 ;
  assign n18940 = n18123 &  n18939 ;
  assign n18936 = x120 | n17617 ;
  assign n18937 = x120 &  n17617 ;
  assign n18938 = ( n18936 & ~n18937 ) | ( n18936 & 1'b0 ) | ( ~n18937 & 1'b0 ) ;
  assign n18942 = ( n18104 & n18125 ) | ( n18104 & n18938 ) | ( n18125 & n18938 ) ;
  assign n18941 = n18104 | n18938 ;
  assign n18943 = ( n18940 & ~n18942 ) | ( n18940 & n18941 ) | ( ~n18942 & n18941 ) ;
  assign n18927 = n17625 &  n18124 ;
  assign n18928 = n18123 &  n18927 ;
  assign n18924 = x119 | n17625 ;
  assign n18925 = x119 &  n17625 ;
  assign n18926 = ( n18924 & ~n18925 ) | ( n18924 & 1'b0 ) | ( ~n18925 & 1'b0 ) ;
  assign n18930 = ( n18103 & n18125 ) | ( n18103 & n18926 ) | ( n18125 & n18926 ) ;
  assign n18929 = n18103 | n18926 ;
  assign n18931 = ( n18928 & ~n18930 ) | ( n18928 & n18929 ) | ( ~n18930 & n18929 ) ;
  assign n18910 = n17633 &  n18124 ;
  assign n18911 = n18123 &  n18910 ;
  assign n18907 = x118 | n17633 ;
  assign n18908 = x118 &  n17633 ;
  assign n18909 = ( n18907 & ~n18908 ) | ( n18907 & 1'b0 ) | ( ~n18908 & 1'b0 ) ;
  assign n18913 = ( n18102 & n18125 ) | ( n18102 & n18909 ) | ( n18125 & n18909 ) ;
  assign n18912 = n18102 | n18909 ;
  assign n18914 = ( n18911 & ~n18913 ) | ( n18911 & n18912 ) | ( ~n18913 & n18912 ) ;
  assign n18898 = n17641 &  n18124 ;
  assign n18899 = n18123 &  n18898 ;
  assign n18895 = x117 | n17641 ;
  assign n18896 = x117 &  n17641 ;
  assign n18897 = ( n18895 & ~n18896 ) | ( n18895 & 1'b0 ) | ( ~n18896 & 1'b0 ) ;
  assign n18901 = ( n18101 & n18125 ) | ( n18101 & n18897 ) | ( n18125 & n18897 ) ;
  assign n18900 = n18101 | n18897 ;
  assign n18902 = ( n18899 & ~n18901 ) | ( n18899 & n18900 ) | ( ~n18901 & n18900 ) ;
  assign n18881 = n17649 &  n18124 ;
  assign n18882 = n18123 &  n18881 ;
  assign n18878 = x116 | n17649 ;
  assign n18879 = x116 &  n17649 ;
  assign n18880 = ( n18878 & ~n18879 ) | ( n18878 & 1'b0 ) | ( ~n18879 & 1'b0 ) ;
  assign n18884 = ( n18100 & n18125 ) | ( n18100 & n18880 ) | ( n18125 & n18880 ) ;
  assign n18883 = n18100 | n18880 ;
  assign n18885 = ( n18882 & ~n18884 ) | ( n18882 & n18883 ) | ( ~n18884 & n18883 ) ;
  assign n18869 = n17657 &  n18124 ;
  assign n18870 = n18123 &  n18869 ;
  assign n18866 = x115 | n17657 ;
  assign n18867 = x115 &  n17657 ;
  assign n18868 = ( n18866 & ~n18867 ) | ( n18866 & 1'b0 ) | ( ~n18867 & 1'b0 ) ;
  assign n18872 = ( n18099 & n18125 ) | ( n18099 & n18868 ) | ( n18125 & n18868 ) ;
  assign n18871 = n18099 | n18868 ;
  assign n18873 = ( n18870 & ~n18872 ) | ( n18870 & n18871 ) | ( ~n18872 & n18871 ) ;
  assign n18852 = n17665 &  n18124 ;
  assign n18853 = n18123 &  n18852 ;
  assign n18849 = x114 | n17665 ;
  assign n18850 = x114 &  n17665 ;
  assign n18851 = ( n18849 & ~n18850 ) | ( n18849 & 1'b0 ) | ( ~n18850 & 1'b0 ) ;
  assign n18855 = ( n18098 & n18125 ) | ( n18098 & n18851 ) | ( n18125 & n18851 ) ;
  assign n18854 = n18098 | n18851 ;
  assign n18856 = ( n18853 & ~n18855 ) | ( n18853 & n18854 ) | ( ~n18855 & n18854 ) ;
  assign n18840 = n17673 &  n18124 ;
  assign n18841 = n18123 &  n18840 ;
  assign n18837 = x113 | n17673 ;
  assign n18838 = x113 &  n17673 ;
  assign n18839 = ( n18837 & ~n18838 ) | ( n18837 & 1'b0 ) | ( ~n18838 & 1'b0 ) ;
  assign n18843 = ( n18097 & n18125 ) | ( n18097 & n18839 ) | ( n18125 & n18839 ) ;
  assign n18842 = n18097 | n18839 ;
  assign n18844 = ( n18841 & ~n18843 ) | ( n18841 & n18842 ) | ( ~n18843 & n18842 ) ;
  assign n18823 = n17681 &  n18124 ;
  assign n18824 = n18123 &  n18823 ;
  assign n18820 = x112 | n17681 ;
  assign n18821 = x112 &  n17681 ;
  assign n18822 = ( n18820 & ~n18821 ) | ( n18820 & 1'b0 ) | ( ~n18821 & 1'b0 ) ;
  assign n18826 = ( n18096 & n18125 ) | ( n18096 & n18822 ) | ( n18125 & n18822 ) ;
  assign n18825 = n18096 | n18822 ;
  assign n18827 = ( n18824 & ~n18826 ) | ( n18824 & n18825 ) | ( ~n18826 & n18825 ) ;
  assign n18811 = n17689 &  n18124 ;
  assign n18812 = n18123 &  n18811 ;
  assign n18808 = x111 | n17689 ;
  assign n18809 = x111 &  n17689 ;
  assign n18810 = ( n18808 & ~n18809 ) | ( n18808 & 1'b0 ) | ( ~n18809 & 1'b0 ) ;
  assign n18814 = ( n18095 & n18125 ) | ( n18095 & n18810 ) | ( n18125 & n18810 ) ;
  assign n18813 = n18095 | n18810 ;
  assign n18815 = ( n18812 & ~n18814 ) | ( n18812 & n18813 ) | ( ~n18814 & n18813 ) ;
  assign n18794 = n17697 &  n18124 ;
  assign n18795 = n18123 &  n18794 ;
  assign n18791 = x110 | n17697 ;
  assign n18792 = x110 &  n17697 ;
  assign n18793 = ( n18791 & ~n18792 ) | ( n18791 & 1'b0 ) | ( ~n18792 & 1'b0 ) ;
  assign n18797 = ( n18094 & n18125 ) | ( n18094 & n18793 ) | ( n18125 & n18793 ) ;
  assign n18796 = n18094 | n18793 ;
  assign n18798 = ( n18795 & ~n18797 ) | ( n18795 & n18796 ) | ( ~n18797 & n18796 ) ;
  assign n18782 = n17705 &  n18124 ;
  assign n18783 = n18123 &  n18782 ;
  assign n18779 = x109 | n17705 ;
  assign n18780 = x109 &  n17705 ;
  assign n18781 = ( n18779 & ~n18780 ) | ( n18779 & 1'b0 ) | ( ~n18780 & 1'b0 ) ;
  assign n18785 = ( n18093 & n18125 ) | ( n18093 & n18781 ) | ( n18125 & n18781 ) ;
  assign n18784 = n18093 | n18781 ;
  assign n18786 = ( n18783 & ~n18785 ) | ( n18783 & n18784 ) | ( ~n18785 & n18784 ) ;
  assign n18765 = n17713 &  n18124 ;
  assign n18766 = n18123 &  n18765 ;
  assign n18762 = x108 | n17713 ;
  assign n18763 = x108 &  n17713 ;
  assign n18764 = ( n18762 & ~n18763 ) | ( n18762 & 1'b0 ) | ( ~n18763 & 1'b0 ) ;
  assign n18768 = ( n18092 & n18125 ) | ( n18092 & n18764 ) | ( n18125 & n18764 ) ;
  assign n18767 = n18092 | n18764 ;
  assign n18769 = ( n18766 & ~n18768 ) | ( n18766 & n18767 ) | ( ~n18768 & n18767 ) ;
  assign n18753 = n17721 &  n18124 ;
  assign n18754 = n18123 &  n18753 ;
  assign n18750 = x107 | n17721 ;
  assign n18751 = x107 &  n17721 ;
  assign n18752 = ( n18750 & ~n18751 ) | ( n18750 & 1'b0 ) | ( ~n18751 & 1'b0 ) ;
  assign n18756 = ( n18091 & n18125 ) | ( n18091 & n18752 ) | ( n18125 & n18752 ) ;
  assign n18755 = n18091 | n18752 ;
  assign n18757 = ( n18754 & ~n18756 ) | ( n18754 & n18755 ) | ( ~n18756 & n18755 ) ;
  assign n18736 = n17729 &  n18124 ;
  assign n18737 = n18123 &  n18736 ;
  assign n18733 = x106 | n17729 ;
  assign n18734 = x106 &  n17729 ;
  assign n18735 = ( n18733 & ~n18734 ) | ( n18733 & 1'b0 ) | ( ~n18734 & 1'b0 ) ;
  assign n18739 = ( n18090 & n18125 ) | ( n18090 & n18735 ) | ( n18125 & n18735 ) ;
  assign n18738 = n18090 | n18735 ;
  assign n18740 = ( n18737 & ~n18739 ) | ( n18737 & n18738 ) | ( ~n18739 & n18738 ) ;
  assign n18724 = n17737 &  n18124 ;
  assign n18725 = n18123 &  n18724 ;
  assign n18721 = x105 | n17737 ;
  assign n18722 = x105 &  n17737 ;
  assign n18723 = ( n18721 & ~n18722 ) | ( n18721 & 1'b0 ) | ( ~n18722 & 1'b0 ) ;
  assign n18727 = ( n18089 & n18125 ) | ( n18089 & n18723 ) | ( n18125 & n18723 ) ;
  assign n18726 = n18089 | n18723 ;
  assign n18728 = ( n18725 & ~n18727 ) | ( n18725 & n18726 ) | ( ~n18727 & n18726 ) ;
  assign n18707 = n17745 &  n18124 ;
  assign n18708 = n18123 &  n18707 ;
  assign n18704 = x104 | n17745 ;
  assign n18705 = x104 &  n17745 ;
  assign n18706 = ( n18704 & ~n18705 ) | ( n18704 & 1'b0 ) | ( ~n18705 & 1'b0 ) ;
  assign n18710 = ( n18088 & n18125 ) | ( n18088 & n18706 ) | ( n18125 & n18706 ) ;
  assign n18709 = n18088 | n18706 ;
  assign n18711 = ( n18708 & ~n18710 ) | ( n18708 & n18709 ) | ( ~n18710 & n18709 ) ;
  assign n18695 = n17753 &  n18124 ;
  assign n18696 = n18123 &  n18695 ;
  assign n18692 = x103 | n17753 ;
  assign n18693 = x103 &  n17753 ;
  assign n18694 = ( n18692 & ~n18693 ) | ( n18692 & 1'b0 ) | ( ~n18693 & 1'b0 ) ;
  assign n18698 = ( n18087 & n18125 ) | ( n18087 & n18694 ) | ( n18125 & n18694 ) ;
  assign n18697 = n18087 | n18694 ;
  assign n18699 = ( n18696 & ~n18698 ) | ( n18696 & n18697 ) | ( ~n18698 & n18697 ) ;
  assign n18678 = n17761 &  n18124 ;
  assign n18679 = n18123 &  n18678 ;
  assign n18675 = x102 | n17761 ;
  assign n18676 = x102 &  n17761 ;
  assign n18677 = ( n18675 & ~n18676 ) | ( n18675 & 1'b0 ) | ( ~n18676 & 1'b0 ) ;
  assign n18681 = ( n18086 & n18125 ) | ( n18086 & n18677 ) | ( n18125 & n18677 ) ;
  assign n18680 = n18086 | n18677 ;
  assign n18682 = ( n18679 & ~n18681 ) | ( n18679 & n18680 ) | ( ~n18681 & n18680 ) ;
  assign n18666 = n17769 &  n18124 ;
  assign n18667 = n18123 &  n18666 ;
  assign n18663 = x101 | n17769 ;
  assign n18664 = x101 &  n17769 ;
  assign n18665 = ( n18663 & ~n18664 ) | ( n18663 & 1'b0 ) | ( ~n18664 & 1'b0 ) ;
  assign n18669 = ( n18085 & n18125 ) | ( n18085 & n18665 ) | ( n18125 & n18665 ) ;
  assign n18668 = n18085 | n18665 ;
  assign n18670 = ( n18667 & ~n18669 ) | ( n18667 & n18668 ) | ( ~n18669 & n18668 ) ;
  assign n18649 = n17777 &  n18124 ;
  assign n18650 = n18123 &  n18649 ;
  assign n18646 = x100 | n17777 ;
  assign n18647 = x100 &  n17777 ;
  assign n18648 = ( n18646 & ~n18647 ) | ( n18646 & 1'b0 ) | ( ~n18647 & 1'b0 ) ;
  assign n18652 = ( n18084 & n18125 ) | ( n18084 & n18648 ) | ( n18125 & n18648 ) ;
  assign n18651 = n18084 | n18648 ;
  assign n18653 = ( n18650 & ~n18652 ) | ( n18650 & n18651 ) | ( ~n18652 & n18651 ) ;
  assign n18637 = n17785 &  n18124 ;
  assign n18638 = n18123 &  n18637 ;
  assign n18634 = x99 | n17785 ;
  assign n18635 = x99 &  n17785 ;
  assign n18636 = ( n18634 & ~n18635 ) | ( n18634 & 1'b0 ) | ( ~n18635 & 1'b0 ) ;
  assign n18640 = ( n18083 & n18125 ) | ( n18083 & n18636 ) | ( n18125 & n18636 ) ;
  assign n18639 = n18083 | n18636 ;
  assign n18641 = ( n18638 & ~n18640 ) | ( n18638 & n18639 ) | ( ~n18640 & n18639 ) ;
  assign n18620 = n17793 &  n18124 ;
  assign n18621 = n18123 &  n18620 ;
  assign n18617 = x98 | n17793 ;
  assign n18618 = x98 &  n17793 ;
  assign n18619 = ( n18617 & ~n18618 ) | ( n18617 & 1'b0 ) | ( ~n18618 & 1'b0 ) ;
  assign n18623 = ( n18082 & n18125 ) | ( n18082 & n18619 ) | ( n18125 & n18619 ) ;
  assign n18622 = n18082 | n18619 ;
  assign n18624 = ( n18621 & ~n18623 ) | ( n18621 & n18622 ) | ( ~n18623 & n18622 ) ;
  assign n18608 = n17801 &  n18124 ;
  assign n18609 = n18123 &  n18608 ;
  assign n18605 = x97 | n17801 ;
  assign n18606 = x97 &  n17801 ;
  assign n18607 = ( n18605 & ~n18606 ) | ( n18605 & 1'b0 ) | ( ~n18606 & 1'b0 ) ;
  assign n18611 = ( n18081 & n18125 ) | ( n18081 & n18607 ) | ( n18125 & n18607 ) ;
  assign n18610 = n18081 | n18607 ;
  assign n18612 = ( n18609 & ~n18611 ) | ( n18609 & n18610 ) | ( ~n18611 & n18610 ) ;
  assign n18591 = n17809 &  n18124 ;
  assign n18592 = n18123 &  n18591 ;
  assign n18588 = x96 | n17809 ;
  assign n18589 = x96 &  n17809 ;
  assign n18590 = ( n18588 & ~n18589 ) | ( n18588 & 1'b0 ) | ( ~n18589 & 1'b0 ) ;
  assign n18594 = ( n18080 & n18125 ) | ( n18080 & n18590 ) | ( n18125 & n18590 ) ;
  assign n18593 = n18080 | n18590 ;
  assign n18595 = ( n18592 & ~n18594 ) | ( n18592 & n18593 ) | ( ~n18594 & n18593 ) ;
  assign n18579 = n17817 &  n18124 ;
  assign n18580 = n18123 &  n18579 ;
  assign n18576 = x95 | n17817 ;
  assign n18577 = x95 &  n17817 ;
  assign n18578 = ( n18576 & ~n18577 ) | ( n18576 & 1'b0 ) | ( ~n18577 & 1'b0 ) ;
  assign n18582 = ( n18079 & n18125 ) | ( n18079 & n18578 ) | ( n18125 & n18578 ) ;
  assign n18581 = n18079 | n18578 ;
  assign n18583 = ( n18580 & ~n18582 ) | ( n18580 & n18581 ) | ( ~n18582 & n18581 ) ;
  assign n18562 = n17825 &  n18124 ;
  assign n18563 = n18123 &  n18562 ;
  assign n18559 = x94 | n17825 ;
  assign n18560 = x94 &  n17825 ;
  assign n18561 = ( n18559 & ~n18560 ) | ( n18559 & 1'b0 ) | ( ~n18560 & 1'b0 ) ;
  assign n18565 = ( n18078 & n18125 ) | ( n18078 & n18561 ) | ( n18125 & n18561 ) ;
  assign n18564 = n18078 | n18561 ;
  assign n18566 = ( n18563 & ~n18565 ) | ( n18563 & n18564 ) | ( ~n18565 & n18564 ) ;
  assign n18550 = n17833 &  n18124 ;
  assign n18551 = n18123 &  n18550 ;
  assign n18547 = x93 | n17833 ;
  assign n18548 = x93 &  n17833 ;
  assign n18549 = ( n18547 & ~n18548 ) | ( n18547 & 1'b0 ) | ( ~n18548 & 1'b0 ) ;
  assign n18553 = ( n18077 & n18125 ) | ( n18077 & n18549 ) | ( n18125 & n18549 ) ;
  assign n18552 = n18077 | n18549 ;
  assign n18554 = ( n18551 & ~n18553 ) | ( n18551 & n18552 ) | ( ~n18553 & n18552 ) ;
  assign n18533 = n17841 &  n18124 ;
  assign n18534 = n18123 &  n18533 ;
  assign n18530 = x92 | n17841 ;
  assign n18531 = x92 &  n17841 ;
  assign n18532 = ( n18530 & ~n18531 ) | ( n18530 & 1'b0 ) | ( ~n18531 & 1'b0 ) ;
  assign n18536 = ( n18076 & n18125 ) | ( n18076 & n18532 ) | ( n18125 & n18532 ) ;
  assign n18535 = n18076 | n18532 ;
  assign n18537 = ( n18534 & ~n18536 ) | ( n18534 & n18535 ) | ( ~n18536 & n18535 ) ;
  assign n18521 = n17849 &  n18124 ;
  assign n18522 = n18123 &  n18521 ;
  assign n18518 = x91 | n17849 ;
  assign n18519 = x91 &  n17849 ;
  assign n18520 = ( n18518 & ~n18519 ) | ( n18518 & 1'b0 ) | ( ~n18519 & 1'b0 ) ;
  assign n18524 = ( n18075 & n18125 ) | ( n18075 & n18520 ) | ( n18125 & n18520 ) ;
  assign n18523 = n18075 | n18520 ;
  assign n18525 = ( n18522 & ~n18524 ) | ( n18522 & n18523 ) | ( ~n18524 & n18523 ) ;
  assign n18504 = n17857 &  n18124 ;
  assign n18505 = n18123 &  n18504 ;
  assign n18501 = x90 | n17857 ;
  assign n18502 = x90 &  n17857 ;
  assign n18503 = ( n18501 & ~n18502 ) | ( n18501 & 1'b0 ) | ( ~n18502 & 1'b0 ) ;
  assign n18507 = ( n18074 & n18125 ) | ( n18074 & n18503 ) | ( n18125 & n18503 ) ;
  assign n18506 = n18074 | n18503 ;
  assign n18508 = ( n18505 & ~n18507 ) | ( n18505 & n18506 ) | ( ~n18507 & n18506 ) ;
  assign n18492 = n17865 &  n18124 ;
  assign n18493 = n18123 &  n18492 ;
  assign n18489 = x89 | n17865 ;
  assign n18490 = x89 &  n17865 ;
  assign n18491 = ( n18489 & ~n18490 ) | ( n18489 & 1'b0 ) | ( ~n18490 & 1'b0 ) ;
  assign n18495 = ( n18073 & n18125 ) | ( n18073 & n18491 ) | ( n18125 & n18491 ) ;
  assign n18494 = n18073 | n18491 ;
  assign n18496 = ( n18493 & ~n18495 ) | ( n18493 & n18494 ) | ( ~n18495 & n18494 ) ;
  assign n18475 = n17873 &  n18124 ;
  assign n18476 = n18123 &  n18475 ;
  assign n18472 = x88 | n17873 ;
  assign n18473 = x88 &  n17873 ;
  assign n18474 = ( n18472 & ~n18473 ) | ( n18472 & 1'b0 ) | ( ~n18473 & 1'b0 ) ;
  assign n18478 = ( n18072 & n18125 ) | ( n18072 & n18474 ) | ( n18125 & n18474 ) ;
  assign n18477 = n18072 | n18474 ;
  assign n18479 = ( n18476 & ~n18478 ) | ( n18476 & n18477 ) | ( ~n18478 & n18477 ) ;
  assign n18463 = n17881 &  n18124 ;
  assign n18464 = n18123 &  n18463 ;
  assign n18460 = x87 | n17881 ;
  assign n18461 = x87 &  n17881 ;
  assign n18462 = ( n18460 & ~n18461 ) | ( n18460 & 1'b0 ) | ( ~n18461 & 1'b0 ) ;
  assign n18466 = ( n18071 & n18125 ) | ( n18071 & n18462 ) | ( n18125 & n18462 ) ;
  assign n18465 = n18071 | n18462 ;
  assign n18467 = ( n18464 & ~n18466 ) | ( n18464 & n18465 ) | ( ~n18466 & n18465 ) ;
  assign n18446 = n17889 &  n18124 ;
  assign n18447 = n18123 &  n18446 ;
  assign n18443 = x86 | n17889 ;
  assign n18444 = x86 &  n17889 ;
  assign n18445 = ( n18443 & ~n18444 ) | ( n18443 & 1'b0 ) | ( ~n18444 & 1'b0 ) ;
  assign n18449 = ( n18070 & n18125 ) | ( n18070 & n18445 ) | ( n18125 & n18445 ) ;
  assign n18448 = n18070 | n18445 ;
  assign n18450 = ( n18447 & ~n18449 ) | ( n18447 & n18448 ) | ( ~n18449 & n18448 ) ;
  assign n18434 = n17897 &  n18124 ;
  assign n18435 = n18123 &  n18434 ;
  assign n18431 = x85 | n17897 ;
  assign n18432 = x85 &  n17897 ;
  assign n18433 = ( n18431 & ~n18432 ) | ( n18431 & 1'b0 ) | ( ~n18432 & 1'b0 ) ;
  assign n18437 = ( n18069 & n18125 ) | ( n18069 & n18433 ) | ( n18125 & n18433 ) ;
  assign n18436 = n18069 | n18433 ;
  assign n18438 = ( n18435 & ~n18437 ) | ( n18435 & n18436 ) | ( ~n18437 & n18436 ) ;
  assign n18417 = n17905 &  n18124 ;
  assign n18418 = n18123 &  n18417 ;
  assign n18414 = x84 | n17905 ;
  assign n18415 = x84 &  n17905 ;
  assign n18416 = ( n18414 & ~n18415 ) | ( n18414 & 1'b0 ) | ( ~n18415 & 1'b0 ) ;
  assign n18420 = ( n18068 & n18125 ) | ( n18068 & n18416 ) | ( n18125 & n18416 ) ;
  assign n18419 = n18068 | n18416 ;
  assign n18421 = ( n18418 & ~n18420 ) | ( n18418 & n18419 ) | ( ~n18420 & n18419 ) ;
  assign n18405 = n17913 &  n18124 ;
  assign n18406 = n18123 &  n18405 ;
  assign n18402 = x83 | n17913 ;
  assign n18403 = x83 &  n17913 ;
  assign n18404 = ( n18402 & ~n18403 ) | ( n18402 & 1'b0 ) | ( ~n18403 & 1'b0 ) ;
  assign n18408 = ( n18067 & n18125 ) | ( n18067 & n18404 ) | ( n18125 & n18404 ) ;
  assign n18407 = n18067 | n18404 ;
  assign n18409 = ( n18406 & ~n18408 ) | ( n18406 & n18407 ) | ( ~n18408 & n18407 ) ;
  assign n18388 = n17921 &  n18124 ;
  assign n18389 = n18123 &  n18388 ;
  assign n18385 = x82 | n17921 ;
  assign n18386 = x82 &  n17921 ;
  assign n18387 = ( n18385 & ~n18386 ) | ( n18385 & 1'b0 ) | ( ~n18386 & 1'b0 ) ;
  assign n18391 = ( n18066 & n18125 ) | ( n18066 & n18387 ) | ( n18125 & n18387 ) ;
  assign n18390 = n18066 | n18387 ;
  assign n18392 = ( n18389 & ~n18391 ) | ( n18389 & n18390 ) | ( ~n18391 & n18390 ) ;
  assign n18376 = n17929 &  n18124 ;
  assign n18377 = n18123 &  n18376 ;
  assign n18373 = x81 | n17929 ;
  assign n18374 = x81 &  n17929 ;
  assign n18375 = ( n18373 & ~n18374 ) | ( n18373 & 1'b0 ) | ( ~n18374 & 1'b0 ) ;
  assign n18379 = ( n18065 & n18125 ) | ( n18065 & n18375 ) | ( n18125 & n18375 ) ;
  assign n18378 = n18065 | n18375 ;
  assign n18380 = ( n18377 & ~n18379 ) | ( n18377 & n18378 ) | ( ~n18379 & n18378 ) ;
  assign n18359 = n17937 &  n18124 ;
  assign n18360 = n18123 &  n18359 ;
  assign n18356 = x80 | n17937 ;
  assign n18357 = x80 &  n17937 ;
  assign n18358 = ( n18356 & ~n18357 ) | ( n18356 & 1'b0 ) | ( ~n18357 & 1'b0 ) ;
  assign n18362 = ( n18064 & n18125 ) | ( n18064 & n18358 ) | ( n18125 & n18358 ) ;
  assign n18361 = n18064 | n18358 ;
  assign n18363 = ( n18360 & ~n18362 ) | ( n18360 & n18361 ) | ( ~n18362 & n18361 ) ;
  assign n18347 = n17945 &  n18124 ;
  assign n18348 = n18123 &  n18347 ;
  assign n18344 = x79 | n17945 ;
  assign n18345 = x79 &  n17945 ;
  assign n18346 = ( n18344 & ~n18345 ) | ( n18344 & 1'b0 ) | ( ~n18345 & 1'b0 ) ;
  assign n18350 = ( n18063 & n18125 ) | ( n18063 & n18346 ) | ( n18125 & n18346 ) ;
  assign n18349 = n18063 | n18346 ;
  assign n18351 = ( n18348 & ~n18350 ) | ( n18348 & n18349 ) | ( ~n18350 & n18349 ) ;
  assign n18330 = n17953 &  n18124 ;
  assign n18331 = n18123 &  n18330 ;
  assign n18327 = x78 | n17953 ;
  assign n18328 = x78 &  n17953 ;
  assign n18329 = ( n18327 & ~n18328 ) | ( n18327 & 1'b0 ) | ( ~n18328 & 1'b0 ) ;
  assign n18333 = ( n18062 & n18125 ) | ( n18062 & n18329 ) | ( n18125 & n18329 ) ;
  assign n18332 = n18062 | n18329 ;
  assign n18334 = ( n18331 & ~n18333 ) | ( n18331 & n18332 ) | ( ~n18333 & n18332 ) ;
  assign n18318 = n17961 &  n18124 ;
  assign n18319 = n18123 &  n18318 ;
  assign n18315 = x77 | n17961 ;
  assign n18316 = x77 &  n17961 ;
  assign n18317 = ( n18315 & ~n18316 ) | ( n18315 & 1'b0 ) | ( ~n18316 & 1'b0 ) ;
  assign n18321 = ( n18061 & n18125 ) | ( n18061 & n18317 ) | ( n18125 & n18317 ) ;
  assign n18320 = n18061 | n18317 ;
  assign n18322 = ( n18319 & ~n18321 ) | ( n18319 & n18320 ) | ( ~n18321 & n18320 ) ;
  assign n18301 = n17969 &  n18124 ;
  assign n18302 = n18123 &  n18301 ;
  assign n18298 = x76 | n17969 ;
  assign n18299 = x76 &  n17969 ;
  assign n18300 = ( n18298 & ~n18299 ) | ( n18298 & 1'b0 ) | ( ~n18299 & 1'b0 ) ;
  assign n18304 = ( n18060 & n18125 ) | ( n18060 & n18300 ) | ( n18125 & n18300 ) ;
  assign n18303 = n18060 | n18300 ;
  assign n18305 = ( n18302 & ~n18304 ) | ( n18302 & n18303 ) | ( ~n18304 & n18303 ) ;
  assign n18289 = n17977 &  n18124 ;
  assign n18290 = n18123 &  n18289 ;
  assign n18286 = x75 | n17977 ;
  assign n18287 = x75 &  n17977 ;
  assign n18288 = ( n18286 & ~n18287 ) | ( n18286 & 1'b0 ) | ( ~n18287 & 1'b0 ) ;
  assign n18292 = ( n18059 & n18125 ) | ( n18059 & n18288 ) | ( n18125 & n18288 ) ;
  assign n18291 = n18059 | n18288 ;
  assign n18293 = ( n18290 & ~n18292 ) | ( n18290 & n18291 ) | ( ~n18292 & n18291 ) ;
  assign n18272 = n17985 &  n18124 ;
  assign n18273 = n18123 &  n18272 ;
  assign n18269 = x74 | n17985 ;
  assign n18270 = x74 &  n17985 ;
  assign n18271 = ( n18269 & ~n18270 ) | ( n18269 & 1'b0 ) | ( ~n18270 & 1'b0 ) ;
  assign n18275 = ( n18058 & n18125 ) | ( n18058 & n18271 ) | ( n18125 & n18271 ) ;
  assign n18274 = n18058 | n18271 ;
  assign n18276 = ( n18273 & ~n18275 ) | ( n18273 & n18274 ) | ( ~n18275 & n18274 ) ;
  assign n18260 = n17993 &  n18124 ;
  assign n18261 = n18123 &  n18260 ;
  assign n18257 = x73 | n17993 ;
  assign n18258 = x73 &  n17993 ;
  assign n18259 = ( n18257 & ~n18258 ) | ( n18257 & 1'b0 ) | ( ~n18258 & 1'b0 ) ;
  assign n18263 = ( n18057 & n18125 ) | ( n18057 & n18259 ) | ( n18125 & n18259 ) ;
  assign n18262 = n18057 | n18259 ;
  assign n18264 = ( n18261 & ~n18263 ) | ( n18261 & n18262 ) | ( ~n18263 & n18262 ) ;
  assign n18243 = n18001 &  n18124 ;
  assign n18244 = n18123 &  n18243 ;
  assign n18240 = x72 | n18001 ;
  assign n18241 = x72 &  n18001 ;
  assign n18242 = ( n18240 & ~n18241 ) | ( n18240 & 1'b0 ) | ( ~n18241 & 1'b0 ) ;
  assign n18246 = ( n18056 & n18125 ) | ( n18056 & n18242 ) | ( n18125 & n18242 ) ;
  assign n18245 = n18056 | n18242 ;
  assign n18247 = ( n18244 & ~n18246 ) | ( n18244 & n18245 ) | ( ~n18246 & n18245 ) ;
  assign n18231 = n18009 &  n18124 ;
  assign n18232 = n18123 &  n18231 ;
  assign n18228 = x71 | n18009 ;
  assign n18229 = x71 &  n18009 ;
  assign n18230 = ( n18228 & ~n18229 ) | ( n18228 & 1'b0 ) | ( ~n18229 & 1'b0 ) ;
  assign n18234 = ( n18055 & n18125 ) | ( n18055 & n18230 ) | ( n18125 & n18230 ) ;
  assign n18233 = n18055 | n18230 ;
  assign n18235 = ( n18232 & ~n18234 ) | ( n18232 & n18233 ) | ( ~n18234 & n18233 ) ;
  assign n18214 = n18017 &  n18124 ;
  assign n18215 = n18123 &  n18214 ;
  assign n18211 = x70 | n18017 ;
  assign n18212 = x70 &  n18017 ;
  assign n18213 = ( n18211 & ~n18212 ) | ( n18211 & 1'b0 ) | ( ~n18212 & 1'b0 ) ;
  assign n18217 = ( n18054 & n18125 ) | ( n18054 & n18213 ) | ( n18125 & n18213 ) ;
  assign n18216 = n18054 | n18213 ;
  assign n18218 = ( n18215 & ~n18217 ) | ( n18215 & n18216 ) | ( ~n18217 & n18216 ) ;
  assign n18202 = n18025 &  n18124 ;
  assign n18203 = n18123 &  n18202 ;
  assign n18199 = x69 | n18025 ;
  assign n18200 = x69 &  n18025 ;
  assign n18201 = ( n18199 & ~n18200 ) | ( n18199 & 1'b0 ) | ( ~n18200 & 1'b0 ) ;
  assign n18205 = ( n18053 & n18125 ) | ( n18053 & n18201 ) | ( n18125 & n18201 ) ;
  assign n18204 = n18053 | n18201 ;
  assign n18206 = ( n18203 & ~n18205 ) | ( n18203 & n18204 ) | ( ~n18205 & n18204 ) ;
  assign n18185 = n18033 &  n18124 ;
  assign n18186 = n18123 &  n18185 ;
  assign n18182 = x68 | n18033 ;
  assign n18183 = x68 &  n18033 ;
  assign n18184 = ( n18182 & ~n18183 ) | ( n18182 & 1'b0 ) | ( ~n18183 & 1'b0 ) ;
  assign n18188 = ( n18052 & n18125 ) | ( n18052 & n18184 ) | ( n18125 & n18184 ) ;
  assign n18187 = n18052 | n18184 ;
  assign n18189 = ( n18186 & ~n18188 ) | ( n18186 & n18187 ) | ( ~n18188 & n18187 ) ;
  assign n18173 = n18038 &  n18124 ;
  assign n18174 = n18123 &  n18173 ;
  assign n18170 = x67 | n18038 ;
  assign n18171 = x67 &  n18038 ;
  assign n18172 = ( n18170 & ~n18171 ) | ( n18170 & 1'b0 ) | ( ~n18171 & 1'b0 ) ;
  assign n18176 = ( n18051 & n18125 ) | ( n18051 & n18172 ) | ( n18125 & n18172 ) ;
  assign n18175 = n18051 | n18172 ;
  assign n18177 = ( n18174 & ~n18176 ) | ( n18174 & n18175 ) | ( ~n18176 & n18175 ) ;
  assign n18157 = n18044 &  n18124 ;
  assign n18158 = n18123 &  n18157 ;
  assign n18154 = x66 | n18044 ;
  assign n18155 = x66 &  n18044 ;
  assign n18156 = ( n18154 & ~n18155 ) | ( n18154 & 1'b0 ) | ( ~n18155 & 1'b0 ) ;
  assign n18160 = ( n18050 & n18125 ) | ( n18050 & n18156 ) | ( n18125 & n18156 ) ;
  assign n18159 = n18050 | n18156 ;
  assign n18161 = ( n18158 & ~n18160 ) | ( n18158 & n18159 ) | ( ~n18160 & n18159 ) ;
  assign n18145 = ( n18048 & ~x65 ) | ( n18048 & n18049 ) | ( ~x65 & n18049 ) ;
  assign n18146 = ( n18050 & ~n18049 ) | ( n18050 & n18145 ) | ( ~n18049 & n18145 ) ;
  assign n18147 = ~n18125 & n18146 ;
  assign n18148 = n18048 &  n18124 ;
  assign n18149 = n18123 &  n18148 ;
  assign n18150 = n18147 | n18149 ;
  assign n18138 = ( n18049 & ~n18125 ) | ( n18049 & 1'b0 ) | ( ~n18125 & 1'b0 ) ;
  assign n18136 = ( x64 & ~n18125 ) | ( x64 & 1'b0 ) | ( ~n18125 & 1'b0 ) ;
  assign n18137 = ( x1 & ~n18136 ) | ( x1 & 1'b0 ) | ( ~n18136 & 1'b0 ) ;
  assign n18139 = ~n18138 & n18137 ;
  assign n18135 = ~x0 & x64 ;
  assign n18140 = ( n18139 & ~n18135 ) | ( n18139 & n18138 ) | ( ~n18135 & n18138 ) ;
  assign n18141 = ( x1 & ~x64 ) | ( x1 & n18125 ) | ( ~x64 & n18125 ) ;
  assign n18142 = ( x1 & ~x0 ) | ( x1 & n18125 ) | ( ~x0 & n18125 ) ;
  assign n18143 = ~n18141 & n18142 ;
  assign n18144 = x65 | n18143 ;
  assign n18167 = ~n18140 & n18144 ;
  assign n18168 = ( x66 & ~n18150 ) | ( x66 & n18167 ) | ( ~n18150 & n18167 ) ;
  assign n18169 = ( n18161 & ~n18168 ) | ( n18161 & 1'b0 ) | ( ~n18168 & 1'b0 ) ;
  assign n18151 = ( n18144 & ~n18150 ) | ( n18144 & 1'b0 ) | ( ~n18150 & 1'b0 ) ;
  assign n18152 = n18140 &  n18151 ;
  assign n18153 = ( x66 & ~n18152 ) | ( x66 & n18151 ) | ( ~n18152 & n18151 ) ;
  assign n18162 = n18137 | n18138 ;
  assign n18163 = ( x65 & ~n18162 ) | ( x65 & n18135 ) | ( ~n18162 & n18135 ) ;
  assign n18164 = ( n18150 & ~n18163 ) | ( n18150 & 1'b0 ) | ( ~n18163 & 1'b0 ) ;
  assign n18165 = n18161 | n18164 ;
  assign n18166 = ( n18153 & ~n18165 ) | ( n18153 & 1'b0 ) | ( ~n18165 & 1'b0 ) ;
  assign n18195 = x67 | n18166 ;
  assign n18196 = ~n18169 & n18195 ;
  assign n18197 = ( x68 & ~n18177 ) | ( x68 & n18196 ) | ( ~n18177 & n18196 ) ;
  assign n18198 = ( n18189 & ~n18197 ) | ( n18189 & 1'b0 ) | ( ~n18197 & 1'b0 ) ;
  assign n18178 = n18169 | n18177 ;
  assign n18179 = ~x67 & n18166 ;
  assign n18180 = ( x67 & ~n18178 ) | ( x67 & n18179 ) | ( ~n18178 & n18179 ) ;
  assign n18181 = x68 | n18180 ;
  assign n18190 = ( n18153 & ~n18164 ) | ( n18153 & 1'b0 ) | ( ~n18164 & 1'b0 ) ;
  assign n18191 = ( x67 & ~n18161 ) | ( x67 & n18190 ) | ( ~n18161 & n18190 ) ;
  assign n18192 = ( n18177 & ~n18191 ) | ( n18177 & 1'b0 ) | ( ~n18191 & 1'b0 ) ;
  assign n18193 = n18189 | n18192 ;
  assign n18194 = ( n18181 & ~n18193 ) | ( n18181 & 1'b0 ) | ( ~n18193 & 1'b0 ) ;
  assign n18224 = x69 | n18194 ;
  assign n18225 = ~n18198 & n18224 ;
  assign n18226 = ( x70 & ~n18206 ) | ( x70 & n18225 ) | ( ~n18206 & n18225 ) ;
  assign n18227 = ( n18218 & ~n18226 ) | ( n18218 & 1'b0 ) | ( ~n18226 & 1'b0 ) ;
  assign n18207 = n18198 | n18206 ;
  assign n18208 = ~x69 & n18194 ;
  assign n18209 = ( x69 & ~n18207 ) | ( x69 & n18208 ) | ( ~n18207 & n18208 ) ;
  assign n18210 = x70 | n18209 ;
  assign n18219 = ( n18181 & ~n18192 ) | ( n18181 & 1'b0 ) | ( ~n18192 & 1'b0 ) ;
  assign n18220 = ( x69 & ~n18189 ) | ( x69 & n18219 ) | ( ~n18189 & n18219 ) ;
  assign n18221 = ( n18206 & ~n18220 ) | ( n18206 & 1'b0 ) | ( ~n18220 & 1'b0 ) ;
  assign n18222 = n18218 | n18221 ;
  assign n18223 = ( n18210 & ~n18222 ) | ( n18210 & 1'b0 ) | ( ~n18222 & 1'b0 ) ;
  assign n18253 = x71 | n18223 ;
  assign n18254 = ~n18227 & n18253 ;
  assign n18255 = ( x72 & ~n18235 ) | ( x72 & n18254 ) | ( ~n18235 & n18254 ) ;
  assign n18256 = ( n18247 & ~n18255 ) | ( n18247 & 1'b0 ) | ( ~n18255 & 1'b0 ) ;
  assign n18236 = n18227 | n18235 ;
  assign n18237 = ~x71 & n18223 ;
  assign n18238 = ( x71 & ~n18236 ) | ( x71 & n18237 ) | ( ~n18236 & n18237 ) ;
  assign n18239 = x72 | n18238 ;
  assign n18248 = ( n18210 & ~n18221 ) | ( n18210 & 1'b0 ) | ( ~n18221 & 1'b0 ) ;
  assign n18249 = ( x71 & ~n18218 ) | ( x71 & n18248 ) | ( ~n18218 & n18248 ) ;
  assign n18250 = ( n18235 & ~n18249 ) | ( n18235 & 1'b0 ) | ( ~n18249 & 1'b0 ) ;
  assign n18251 = n18247 | n18250 ;
  assign n18252 = ( n18239 & ~n18251 ) | ( n18239 & 1'b0 ) | ( ~n18251 & 1'b0 ) ;
  assign n18282 = x73 | n18252 ;
  assign n18283 = ~n18256 & n18282 ;
  assign n18284 = ( x74 & ~n18264 ) | ( x74 & n18283 ) | ( ~n18264 & n18283 ) ;
  assign n18285 = ( n18276 & ~n18284 ) | ( n18276 & 1'b0 ) | ( ~n18284 & 1'b0 ) ;
  assign n18265 = n18256 | n18264 ;
  assign n18266 = ~x73 & n18252 ;
  assign n18267 = ( x73 & ~n18265 ) | ( x73 & n18266 ) | ( ~n18265 & n18266 ) ;
  assign n18268 = x74 | n18267 ;
  assign n18277 = ( n18239 & ~n18250 ) | ( n18239 & 1'b0 ) | ( ~n18250 & 1'b0 ) ;
  assign n18278 = ( x73 & ~n18247 ) | ( x73 & n18277 ) | ( ~n18247 & n18277 ) ;
  assign n18279 = ( n18264 & ~n18278 ) | ( n18264 & 1'b0 ) | ( ~n18278 & 1'b0 ) ;
  assign n18280 = n18276 | n18279 ;
  assign n18281 = ( n18268 & ~n18280 ) | ( n18268 & 1'b0 ) | ( ~n18280 & 1'b0 ) ;
  assign n18311 = x75 | n18281 ;
  assign n18312 = ~n18285 & n18311 ;
  assign n18313 = ( x76 & ~n18293 ) | ( x76 & n18312 ) | ( ~n18293 & n18312 ) ;
  assign n18314 = ( n18305 & ~n18313 ) | ( n18305 & 1'b0 ) | ( ~n18313 & 1'b0 ) ;
  assign n18294 = n18285 | n18293 ;
  assign n18295 = ~x75 & n18281 ;
  assign n18296 = ( x75 & ~n18294 ) | ( x75 & n18295 ) | ( ~n18294 & n18295 ) ;
  assign n18297 = x76 | n18296 ;
  assign n18306 = ( n18268 & ~n18279 ) | ( n18268 & 1'b0 ) | ( ~n18279 & 1'b0 ) ;
  assign n18307 = ( x75 & ~n18276 ) | ( x75 & n18306 ) | ( ~n18276 & n18306 ) ;
  assign n18308 = ( n18293 & ~n18307 ) | ( n18293 & 1'b0 ) | ( ~n18307 & 1'b0 ) ;
  assign n18309 = n18305 | n18308 ;
  assign n18310 = ( n18297 & ~n18309 ) | ( n18297 & 1'b0 ) | ( ~n18309 & 1'b0 ) ;
  assign n18340 = x77 | n18310 ;
  assign n18341 = ~n18314 & n18340 ;
  assign n18342 = ( x78 & ~n18322 ) | ( x78 & n18341 ) | ( ~n18322 & n18341 ) ;
  assign n18343 = ( n18334 & ~n18342 ) | ( n18334 & 1'b0 ) | ( ~n18342 & 1'b0 ) ;
  assign n18323 = n18314 | n18322 ;
  assign n18324 = ~x77 & n18310 ;
  assign n18325 = ( x77 & ~n18323 ) | ( x77 & n18324 ) | ( ~n18323 & n18324 ) ;
  assign n18326 = x78 | n18325 ;
  assign n18335 = ( n18297 & ~n18308 ) | ( n18297 & 1'b0 ) | ( ~n18308 & 1'b0 ) ;
  assign n18336 = ( x77 & ~n18305 ) | ( x77 & n18335 ) | ( ~n18305 & n18335 ) ;
  assign n18337 = ( n18322 & ~n18336 ) | ( n18322 & 1'b0 ) | ( ~n18336 & 1'b0 ) ;
  assign n18338 = n18334 | n18337 ;
  assign n18339 = ( n18326 & ~n18338 ) | ( n18326 & 1'b0 ) | ( ~n18338 & 1'b0 ) ;
  assign n18369 = x79 | n18339 ;
  assign n18370 = ~n18343 & n18369 ;
  assign n18371 = ( x80 & ~n18351 ) | ( x80 & n18370 ) | ( ~n18351 & n18370 ) ;
  assign n18372 = ( n18363 & ~n18371 ) | ( n18363 & 1'b0 ) | ( ~n18371 & 1'b0 ) ;
  assign n18352 = n18343 | n18351 ;
  assign n18353 = ~x79 & n18339 ;
  assign n18354 = ( x79 & ~n18352 ) | ( x79 & n18353 ) | ( ~n18352 & n18353 ) ;
  assign n18355 = x80 | n18354 ;
  assign n18364 = ( n18326 & ~n18337 ) | ( n18326 & 1'b0 ) | ( ~n18337 & 1'b0 ) ;
  assign n18365 = ( x79 & ~n18334 ) | ( x79 & n18364 ) | ( ~n18334 & n18364 ) ;
  assign n18366 = ( n18351 & ~n18365 ) | ( n18351 & 1'b0 ) | ( ~n18365 & 1'b0 ) ;
  assign n18367 = n18363 | n18366 ;
  assign n18368 = ( n18355 & ~n18367 ) | ( n18355 & 1'b0 ) | ( ~n18367 & 1'b0 ) ;
  assign n18398 = x81 | n18368 ;
  assign n18399 = ~n18372 & n18398 ;
  assign n18400 = ( x82 & ~n18380 ) | ( x82 & n18399 ) | ( ~n18380 & n18399 ) ;
  assign n18401 = ( n18392 & ~n18400 ) | ( n18392 & 1'b0 ) | ( ~n18400 & 1'b0 ) ;
  assign n18381 = n18372 | n18380 ;
  assign n18382 = ~x81 & n18368 ;
  assign n18383 = ( x81 & ~n18381 ) | ( x81 & n18382 ) | ( ~n18381 & n18382 ) ;
  assign n18384 = x82 | n18383 ;
  assign n18393 = ( n18355 & ~n18366 ) | ( n18355 & 1'b0 ) | ( ~n18366 & 1'b0 ) ;
  assign n18394 = ( x81 & ~n18363 ) | ( x81 & n18393 ) | ( ~n18363 & n18393 ) ;
  assign n18395 = ( n18380 & ~n18394 ) | ( n18380 & 1'b0 ) | ( ~n18394 & 1'b0 ) ;
  assign n18396 = n18392 | n18395 ;
  assign n18397 = ( n18384 & ~n18396 ) | ( n18384 & 1'b0 ) | ( ~n18396 & 1'b0 ) ;
  assign n18427 = x83 | n18397 ;
  assign n18428 = ~n18401 & n18427 ;
  assign n18429 = ( x84 & ~n18409 ) | ( x84 & n18428 ) | ( ~n18409 & n18428 ) ;
  assign n18430 = ( n18421 & ~n18429 ) | ( n18421 & 1'b0 ) | ( ~n18429 & 1'b0 ) ;
  assign n18410 = n18401 | n18409 ;
  assign n18411 = ~x83 & n18397 ;
  assign n18412 = ( x83 & ~n18410 ) | ( x83 & n18411 ) | ( ~n18410 & n18411 ) ;
  assign n18413 = x84 | n18412 ;
  assign n18422 = ( n18384 & ~n18395 ) | ( n18384 & 1'b0 ) | ( ~n18395 & 1'b0 ) ;
  assign n18423 = ( x83 & ~n18392 ) | ( x83 & n18422 ) | ( ~n18392 & n18422 ) ;
  assign n18424 = ( n18409 & ~n18423 ) | ( n18409 & 1'b0 ) | ( ~n18423 & 1'b0 ) ;
  assign n18425 = n18421 | n18424 ;
  assign n18426 = ( n18413 & ~n18425 ) | ( n18413 & 1'b0 ) | ( ~n18425 & 1'b0 ) ;
  assign n18456 = x85 | n18426 ;
  assign n18457 = ~n18430 & n18456 ;
  assign n18458 = ( x86 & ~n18438 ) | ( x86 & n18457 ) | ( ~n18438 & n18457 ) ;
  assign n18459 = ( n18450 & ~n18458 ) | ( n18450 & 1'b0 ) | ( ~n18458 & 1'b0 ) ;
  assign n18439 = n18430 | n18438 ;
  assign n18440 = ~x85 & n18426 ;
  assign n18441 = ( x85 & ~n18439 ) | ( x85 & n18440 ) | ( ~n18439 & n18440 ) ;
  assign n18442 = x86 | n18441 ;
  assign n18451 = ( n18413 & ~n18424 ) | ( n18413 & 1'b0 ) | ( ~n18424 & 1'b0 ) ;
  assign n18452 = ( x85 & ~n18421 ) | ( x85 & n18451 ) | ( ~n18421 & n18451 ) ;
  assign n18453 = ( n18438 & ~n18452 ) | ( n18438 & 1'b0 ) | ( ~n18452 & 1'b0 ) ;
  assign n18454 = n18450 | n18453 ;
  assign n18455 = ( n18442 & ~n18454 ) | ( n18442 & 1'b0 ) | ( ~n18454 & 1'b0 ) ;
  assign n18485 = x87 | n18455 ;
  assign n18486 = ~n18459 & n18485 ;
  assign n18487 = ( x88 & ~n18467 ) | ( x88 & n18486 ) | ( ~n18467 & n18486 ) ;
  assign n18488 = ( n18479 & ~n18487 ) | ( n18479 & 1'b0 ) | ( ~n18487 & 1'b0 ) ;
  assign n18468 = n18459 | n18467 ;
  assign n18469 = ~x87 & n18455 ;
  assign n18470 = ( x87 & ~n18468 ) | ( x87 & n18469 ) | ( ~n18468 & n18469 ) ;
  assign n18471 = x88 | n18470 ;
  assign n18480 = ( n18442 & ~n18453 ) | ( n18442 & 1'b0 ) | ( ~n18453 & 1'b0 ) ;
  assign n18481 = ( x87 & ~n18450 ) | ( x87 & n18480 ) | ( ~n18450 & n18480 ) ;
  assign n18482 = ( n18467 & ~n18481 ) | ( n18467 & 1'b0 ) | ( ~n18481 & 1'b0 ) ;
  assign n18483 = n18479 | n18482 ;
  assign n18484 = ( n18471 & ~n18483 ) | ( n18471 & 1'b0 ) | ( ~n18483 & 1'b0 ) ;
  assign n18514 = x89 | n18484 ;
  assign n18515 = ~n18488 & n18514 ;
  assign n18516 = ( x90 & ~n18496 ) | ( x90 & n18515 ) | ( ~n18496 & n18515 ) ;
  assign n18517 = ( n18508 & ~n18516 ) | ( n18508 & 1'b0 ) | ( ~n18516 & 1'b0 ) ;
  assign n18497 = n18488 | n18496 ;
  assign n18498 = ~x89 & n18484 ;
  assign n18499 = ( x89 & ~n18497 ) | ( x89 & n18498 ) | ( ~n18497 & n18498 ) ;
  assign n18500 = x90 | n18499 ;
  assign n18509 = ( n18471 & ~n18482 ) | ( n18471 & 1'b0 ) | ( ~n18482 & 1'b0 ) ;
  assign n18510 = ( x89 & ~n18479 ) | ( x89 & n18509 ) | ( ~n18479 & n18509 ) ;
  assign n18511 = ( n18496 & ~n18510 ) | ( n18496 & 1'b0 ) | ( ~n18510 & 1'b0 ) ;
  assign n18512 = n18508 | n18511 ;
  assign n18513 = ( n18500 & ~n18512 ) | ( n18500 & 1'b0 ) | ( ~n18512 & 1'b0 ) ;
  assign n18543 = x91 | n18513 ;
  assign n18544 = ~n18517 & n18543 ;
  assign n18545 = ( x92 & ~n18525 ) | ( x92 & n18544 ) | ( ~n18525 & n18544 ) ;
  assign n18546 = ( n18537 & ~n18545 ) | ( n18537 & 1'b0 ) | ( ~n18545 & 1'b0 ) ;
  assign n18526 = n18517 | n18525 ;
  assign n18527 = ~x91 & n18513 ;
  assign n18528 = ( x91 & ~n18526 ) | ( x91 & n18527 ) | ( ~n18526 & n18527 ) ;
  assign n18529 = x92 | n18528 ;
  assign n18538 = ( n18500 & ~n18511 ) | ( n18500 & 1'b0 ) | ( ~n18511 & 1'b0 ) ;
  assign n18539 = ( x91 & ~n18508 ) | ( x91 & n18538 ) | ( ~n18508 & n18538 ) ;
  assign n18540 = ( n18525 & ~n18539 ) | ( n18525 & 1'b0 ) | ( ~n18539 & 1'b0 ) ;
  assign n18541 = n18537 | n18540 ;
  assign n18542 = ( n18529 & ~n18541 ) | ( n18529 & 1'b0 ) | ( ~n18541 & 1'b0 ) ;
  assign n18572 = x93 | n18542 ;
  assign n18573 = ~n18546 & n18572 ;
  assign n18574 = ( x94 & ~n18554 ) | ( x94 & n18573 ) | ( ~n18554 & n18573 ) ;
  assign n18575 = ( n18566 & ~n18574 ) | ( n18566 & 1'b0 ) | ( ~n18574 & 1'b0 ) ;
  assign n18555 = n18546 | n18554 ;
  assign n18556 = ~x93 & n18542 ;
  assign n18557 = ( x93 & ~n18555 ) | ( x93 & n18556 ) | ( ~n18555 & n18556 ) ;
  assign n18558 = x94 | n18557 ;
  assign n18567 = ( n18529 & ~n18540 ) | ( n18529 & 1'b0 ) | ( ~n18540 & 1'b0 ) ;
  assign n18568 = ( x93 & ~n18537 ) | ( x93 & n18567 ) | ( ~n18537 & n18567 ) ;
  assign n18569 = ( n18554 & ~n18568 ) | ( n18554 & 1'b0 ) | ( ~n18568 & 1'b0 ) ;
  assign n18570 = n18566 | n18569 ;
  assign n18571 = ( n18558 & ~n18570 ) | ( n18558 & 1'b0 ) | ( ~n18570 & 1'b0 ) ;
  assign n18601 = x95 | n18571 ;
  assign n18602 = ~n18575 & n18601 ;
  assign n18603 = ( x96 & ~n18583 ) | ( x96 & n18602 ) | ( ~n18583 & n18602 ) ;
  assign n18604 = ( n18595 & ~n18603 ) | ( n18595 & 1'b0 ) | ( ~n18603 & 1'b0 ) ;
  assign n18584 = n18575 | n18583 ;
  assign n18585 = ~x95 & n18571 ;
  assign n18586 = ( x95 & ~n18584 ) | ( x95 & n18585 ) | ( ~n18584 & n18585 ) ;
  assign n18587 = x96 | n18586 ;
  assign n18596 = ( n18558 & ~n18569 ) | ( n18558 & 1'b0 ) | ( ~n18569 & 1'b0 ) ;
  assign n18597 = ( x95 & ~n18566 ) | ( x95 & n18596 ) | ( ~n18566 & n18596 ) ;
  assign n18598 = ( n18583 & ~n18597 ) | ( n18583 & 1'b0 ) | ( ~n18597 & 1'b0 ) ;
  assign n18599 = n18595 | n18598 ;
  assign n18600 = ( n18587 & ~n18599 ) | ( n18587 & 1'b0 ) | ( ~n18599 & 1'b0 ) ;
  assign n18630 = x97 | n18600 ;
  assign n18631 = ~n18604 & n18630 ;
  assign n18632 = ( x98 & ~n18612 ) | ( x98 & n18631 ) | ( ~n18612 & n18631 ) ;
  assign n18633 = ( n18624 & ~n18632 ) | ( n18624 & 1'b0 ) | ( ~n18632 & 1'b0 ) ;
  assign n18613 = n18604 | n18612 ;
  assign n18614 = ~x97 & n18600 ;
  assign n18615 = ( x97 & ~n18613 ) | ( x97 & n18614 ) | ( ~n18613 & n18614 ) ;
  assign n18616 = x98 | n18615 ;
  assign n18625 = ( n18587 & ~n18598 ) | ( n18587 & 1'b0 ) | ( ~n18598 & 1'b0 ) ;
  assign n18626 = ( x97 & ~n18595 ) | ( x97 & n18625 ) | ( ~n18595 & n18625 ) ;
  assign n18627 = ( n18612 & ~n18626 ) | ( n18612 & 1'b0 ) | ( ~n18626 & 1'b0 ) ;
  assign n18628 = n18624 | n18627 ;
  assign n18629 = ( n18616 & ~n18628 ) | ( n18616 & 1'b0 ) | ( ~n18628 & 1'b0 ) ;
  assign n18659 = x99 | n18629 ;
  assign n18660 = ~n18633 & n18659 ;
  assign n18661 = ( x100 & ~n18641 ) | ( x100 & n18660 ) | ( ~n18641 & n18660 ) ;
  assign n18662 = ( n18653 & ~n18661 ) | ( n18653 & 1'b0 ) | ( ~n18661 & 1'b0 ) ;
  assign n18642 = n18633 | n18641 ;
  assign n18643 = ~x99 & n18629 ;
  assign n18644 = ( x99 & ~n18642 ) | ( x99 & n18643 ) | ( ~n18642 & n18643 ) ;
  assign n18645 = x100 | n18644 ;
  assign n18654 = ( n18616 & ~n18627 ) | ( n18616 & 1'b0 ) | ( ~n18627 & 1'b0 ) ;
  assign n18655 = ( x99 & ~n18624 ) | ( x99 & n18654 ) | ( ~n18624 & n18654 ) ;
  assign n18656 = ( n18641 & ~n18655 ) | ( n18641 & 1'b0 ) | ( ~n18655 & 1'b0 ) ;
  assign n18657 = n18653 | n18656 ;
  assign n18658 = ( n18645 & ~n18657 ) | ( n18645 & 1'b0 ) | ( ~n18657 & 1'b0 ) ;
  assign n18688 = x101 | n18658 ;
  assign n18689 = ~n18662 & n18688 ;
  assign n18690 = ( x102 & ~n18670 ) | ( x102 & n18689 ) | ( ~n18670 & n18689 ) ;
  assign n18691 = ( n18682 & ~n18690 ) | ( n18682 & 1'b0 ) | ( ~n18690 & 1'b0 ) ;
  assign n18671 = n18662 | n18670 ;
  assign n18672 = ~x101 & n18658 ;
  assign n18673 = ( x101 & ~n18671 ) | ( x101 & n18672 ) | ( ~n18671 & n18672 ) ;
  assign n18674 = x102 | n18673 ;
  assign n18683 = ( n18645 & ~n18656 ) | ( n18645 & 1'b0 ) | ( ~n18656 & 1'b0 ) ;
  assign n18684 = ( x101 & ~n18653 ) | ( x101 & n18683 ) | ( ~n18653 & n18683 ) ;
  assign n18685 = ( n18670 & ~n18684 ) | ( n18670 & 1'b0 ) | ( ~n18684 & 1'b0 ) ;
  assign n18686 = n18682 | n18685 ;
  assign n18687 = ( n18674 & ~n18686 ) | ( n18674 & 1'b0 ) | ( ~n18686 & 1'b0 ) ;
  assign n18717 = x103 | n18687 ;
  assign n18718 = ~n18691 & n18717 ;
  assign n18719 = ( x104 & ~n18699 ) | ( x104 & n18718 ) | ( ~n18699 & n18718 ) ;
  assign n18720 = ( n18711 & ~n18719 ) | ( n18711 & 1'b0 ) | ( ~n18719 & 1'b0 ) ;
  assign n18700 = n18691 | n18699 ;
  assign n18701 = ~x103 & n18687 ;
  assign n18702 = ( x103 & ~n18700 ) | ( x103 & n18701 ) | ( ~n18700 & n18701 ) ;
  assign n18703 = x104 | n18702 ;
  assign n18712 = ( n18674 & ~n18685 ) | ( n18674 & 1'b0 ) | ( ~n18685 & 1'b0 ) ;
  assign n18713 = ( x103 & ~n18682 ) | ( x103 & n18712 ) | ( ~n18682 & n18712 ) ;
  assign n18714 = ( n18699 & ~n18713 ) | ( n18699 & 1'b0 ) | ( ~n18713 & 1'b0 ) ;
  assign n18715 = n18711 | n18714 ;
  assign n18716 = ( n18703 & ~n18715 ) | ( n18703 & 1'b0 ) | ( ~n18715 & 1'b0 ) ;
  assign n18746 = x105 | n18716 ;
  assign n18747 = ~n18720 & n18746 ;
  assign n18748 = ( x106 & ~n18728 ) | ( x106 & n18747 ) | ( ~n18728 & n18747 ) ;
  assign n18749 = ( n18740 & ~n18748 ) | ( n18740 & 1'b0 ) | ( ~n18748 & 1'b0 ) ;
  assign n18729 = n18720 | n18728 ;
  assign n18730 = ~x105 & n18716 ;
  assign n18731 = ( x105 & ~n18729 ) | ( x105 & n18730 ) | ( ~n18729 & n18730 ) ;
  assign n18732 = x106 | n18731 ;
  assign n18741 = ( n18703 & ~n18714 ) | ( n18703 & 1'b0 ) | ( ~n18714 & 1'b0 ) ;
  assign n18742 = ( x105 & ~n18711 ) | ( x105 & n18741 ) | ( ~n18711 & n18741 ) ;
  assign n18743 = ( n18728 & ~n18742 ) | ( n18728 & 1'b0 ) | ( ~n18742 & 1'b0 ) ;
  assign n18744 = n18740 | n18743 ;
  assign n18745 = ( n18732 & ~n18744 ) | ( n18732 & 1'b0 ) | ( ~n18744 & 1'b0 ) ;
  assign n18775 = x107 | n18745 ;
  assign n18776 = ~n18749 & n18775 ;
  assign n18777 = ( x108 & ~n18757 ) | ( x108 & n18776 ) | ( ~n18757 & n18776 ) ;
  assign n18778 = ( n18769 & ~n18777 ) | ( n18769 & 1'b0 ) | ( ~n18777 & 1'b0 ) ;
  assign n18758 = n18749 | n18757 ;
  assign n18759 = ~x107 & n18745 ;
  assign n18760 = ( x107 & ~n18758 ) | ( x107 & n18759 ) | ( ~n18758 & n18759 ) ;
  assign n18761 = x108 | n18760 ;
  assign n18770 = ( n18732 & ~n18743 ) | ( n18732 & 1'b0 ) | ( ~n18743 & 1'b0 ) ;
  assign n18771 = ( x107 & ~n18740 ) | ( x107 & n18770 ) | ( ~n18740 & n18770 ) ;
  assign n18772 = ( n18757 & ~n18771 ) | ( n18757 & 1'b0 ) | ( ~n18771 & 1'b0 ) ;
  assign n18773 = n18769 | n18772 ;
  assign n18774 = ( n18761 & ~n18773 ) | ( n18761 & 1'b0 ) | ( ~n18773 & 1'b0 ) ;
  assign n18804 = x109 | n18774 ;
  assign n18805 = ~n18778 & n18804 ;
  assign n18806 = ( x110 & ~n18786 ) | ( x110 & n18805 ) | ( ~n18786 & n18805 ) ;
  assign n18807 = ( n18798 & ~n18806 ) | ( n18798 & 1'b0 ) | ( ~n18806 & 1'b0 ) ;
  assign n18787 = n18778 | n18786 ;
  assign n18788 = ~x109 & n18774 ;
  assign n18789 = ( x109 & ~n18787 ) | ( x109 & n18788 ) | ( ~n18787 & n18788 ) ;
  assign n18790 = x110 | n18789 ;
  assign n18799 = ( n18761 & ~n18772 ) | ( n18761 & 1'b0 ) | ( ~n18772 & 1'b0 ) ;
  assign n18800 = ( x109 & ~n18769 ) | ( x109 & n18799 ) | ( ~n18769 & n18799 ) ;
  assign n18801 = ( n18786 & ~n18800 ) | ( n18786 & 1'b0 ) | ( ~n18800 & 1'b0 ) ;
  assign n18802 = n18798 | n18801 ;
  assign n18803 = ( n18790 & ~n18802 ) | ( n18790 & 1'b0 ) | ( ~n18802 & 1'b0 ) ;
  assign n18833 = x111 | n18803 ;
  assign n18834 = ~n18807 & n18833 ;
  assign n18835 = ( x112 & ~n18815 ) | ( x112 & n18834 ) | ( ~n18815 & n18834 ) ;
  assign n18836 = ( n18827 & ~n18835 ) | ( n18827 & 1'b0 ) | ( ~n18835 & 1'b0 ) ;
  assign n18816 = n18807 | n18815 ;
  assign n18817 = ~x111 & n18803 ;
  assign n18818 = ( x111 & ~n18816 ) | ( x111 & n18817 ) | ( ~n18816 & n18817 ) ;
  assign n18819 = x112 | n18818 ;
  assign n18828 = ( n18790 & ~n18801 ) | ( n18790 & 1'b0 ) | ( ~n18801 & 1'b0 ) ;
  assign n18829 = ( x111 & ~n18798 ) | ( x111 & n18828 ) | ( ~n18798 & n18828 ) ;
  assign n18830 = ( n18815 & ~n18829 ) | ( n18815 & 1'b0 ) | ( ~n18829 & 1'b0 ) ;
  assign n18831 = n18827 | n18830 ;
  assign n18832 = ( n18819 & ~n18831 ) | ( n18819 & 1'b0 ) | ( ~n18831 & 1'b0 ) ;
  assign n18862 = x113 | n18832 ;
  assign n18863 = ~n18836 & n18862 ;
  assign n18864 = ( x114 & ~n18844 ) | ( x114 & n18863 ) | ( ~n18844 & n18863 ) ;
  assign n18865 = ( n18856 & ~n18864 ) | ( n18856 & 1'b0 ) | ( ~n18864 & 1'b0 ) ;
  assign n18845 = n18836 | n18844 ;
  assign n18846 = ~x113 & n18832 ;
  assign n18847 = ( x113 & ~n18845 ) | ( x113 & n18846 ) | ( ~n18845 & n18846 ) ;
  assign n18848 = x114 | n18847 ;
  assign n18857 = ( n18819 & ~n18830 ) | ( n18819 & 1'b0 ) | ( ~n18830 & 1'b0 ) ;
  assign n18858 = ( x113 & ~n18827 ) | ( x113 & n18857 ) | ( ~n18827 & n18857 ) ;
  assign n18859 = ( n18844 & ~n18858 ) | ( n18844 & 1'b0 ) | ( ~n18858 & 1'b0 ) ;
  assign n18860 = n18856 | n18859 ;
  assign n18861 = ( n18848 & ~n18860 ) | ( n18848 & 1'b0 ) | ( ~n18860 & 1'b0 ) ;
  assign n18891 = x115 | n18861 ;
  assign n18892 = ~n18865 & n18891 ;
  assign n18893 = ( x116 & ~n18873 ) | ( x116 & n18892 ) | ( ~n18873 & n18892 ) ;
  assign n18894 = ( n18885 & ~n18893 ) | ( n18885 & 1'b0 ) | ( ~n18893 & 1'b0 ) ;
  assign n18874 = n18865 | n18873 ;
  assign n18875 = ~x115 & n18861 ;
  assign n18876 = ( x115 & ~n18874 ) | ( x115 & n18875 ) | ( ~n18874 & n18875 ) ;
  assign n18877 = x116 | n18876 ;
  assign n18886 = ( n18848 & ~n18859 ) | ( n18848 & 1'b0 ) | ( ~n18859 & 1'b0 ) ;
  assign n18887 = ( x115 & ~n18856 ) | ( x115 & n18886 ) | ( ~n18856 & n18886 ) ;
  assign n18888 = ( n18873 & ~n18887 ) | ( n18873 & 1'b0 ) | ( ~n18887 & 1'b0 ) ;
  assign n18889 = n18885 | n18888 ;
  assign n18890 = ( n18877 & ~n18889 ) | ( n18877 & 1'b0 ) | ( ~n18889 & 1'b0 ) ;
  assign n18920 = x117 | n18890 ;
  assign n18921 = ~n18894 & n18920 ;
  assign n18922 = ( x118 & ~n18902 ) | ( x118 & n18921 ) | ( ~n18902 & n18921 ) ;
  assign n18923 = ( n18914 & ~n18922 ) | ( n18914 & 1'b0 ) | ( ~n18922 & 1'b0 ) ;
  assign n18903 = n18894 | n18902 ;
  assign n18904 = ~x117 & n18890 ;
  assign n18905 = ( x117 & ~n18903 ) | ( x117 & n18904 ) | ( ~n18903 & n18904 ) ;
  assign n18906 = x118 | n18905 ;
  assign n18915 = ( n18877 & ~n18888 ) | ( n18877 & 1'b0 ) | ( ~n18888 & 1'b0 ) ;
  assign n18916 = ( x117 & ~n18885 ) | ( x117 & n18915 ) | ( ~n18885 & n18915 ) ;
  assign n18917 = ( n18902 & ~n18916 ) | ( n18902 & 1'b0 ) | ( ~n18916 & 1'b0 ) ;
  assign n18918 = n18914 | n18917 ;
  assign n18919 = ( n18906 & ~n18918 ) | ( n18906 & 1'b0 ) | ( ~n18918 & 1'b0 ) ;
  assign n18949 = x119 | n18919 ;
  assign n18950 = ~n18923 & n18949 ;
  assign n18951 = ( x120 & ~n18931 ) | ( x120 & n18950 ) | ( ~n18931 & n18950 ) ;
  assign n18952 = ( n18943 & ~n18951 ) | ( n18943 & 1'b0 ) | ( ~n18951 & 1'b0 ) ;
  assign n18932 = n18923 | n18931 ;
  assign n18933 = ~x119 & n18919 ;
  assign n18934 = ( x119 & ~n18932 ) | ( x119 & n18933 ) | ( ~n18932 & n18933 ) ;
  assign n18935 = x120 | n18934 ;
  assign n18944 = ( n18906 & ~n18917 ) | ( n18906 & 1'b0 ) | ( ~n18917 & 1'b0 ) ;
  assign n18945 = ( x119 & ~n18914 ) | ( x119 & n18944 ) | ( ~n18914 & n18944 ) ;
  assign n18946 = ( n18931 & ~n18945 ) | ( n18931 & 1'b0 ) | ( ~n18945 & 1'b0 ) ;
  assign n18947 = n18943 | n18946 ;
  assign n18948 = ( n18935 & ~n18947 ) | ( n18935 & 1'b0 ) | ( ~n18947 & 1'b0 ) ;
  assign n18978 = x121 | n18948 ;
  assign n18979 = ~n18952 & n18978 ;
  assign n18980 = ( x122 & ~n18960 ) | ( x122 & n18979 ) | ( ~n18960 & n18979 ) ;
  assign n18981 = ( n18972 & ~n18980 ) | ( n18972 & 1'b0 ) | ( ~n18980 & 1'b0 ) ;
  assign n18961 = n18952 | n18960 ;
  assign n18962 = ~x121 & n18948 ;
  assign n18963 = ( x121 & ~n18961 ) | ( x121 & n18962 ) | ( ~n18961 & n18962 ) ;
  assign n18964 = x122 | n18963 ;
  assign n18973 = ( n18935 & ~n18946 ) | ( n18935 & 1'b0 ) | ( ~n18946 & 1'b0 ) ;
  assign n18974 = ( x121 & ~n18943 ) | ( x121 & n18973 ) | ( ~n18943 & n18973 ) ;
  assign n18975 = ( n18960 & ~n18974 ) | ( n18960 & 1'b0 ) | ( ~n18974 & 1'b0 ) ;
  assign n18976 = n18972 | n18975 ;
  assign n18977 = ( n18964 & ~n18976 ) | ( n18964 & 1'b0 ) | ( ~n18976 & 1'b0 ) ;
  assign n19007 = x123 | n18977 ;
  assign n19008 = ~n18981 & n19007 ;
  assign n19009 = ( x124 & ~n18989 ) | ( x124 & n19008 ) | ( ~n18989 & n19008 ) ;
  assign n19010 = ( n19001 & ~n19009 ) | ( n19001 & 1'b0 ) | ( ~n19009 & 1'b0 ) ;
  assign n19011 = n17577 &  n18124 ;
  assign n19012 = n18123 &  n19011 ;
  assign n18126 = x125 | n17577 ;
  assign n18127 = x125 &  n17577 ;
  assign n18128 = ( n18126 & ~n18127 ) | ( n18126 & 1'b0 ) | ( ~n18127 & 1'b0 ) ;
  assign n19013 = n18109 &  n18128 ;
  assign n19014 = ( n18109 & ~n18125 ) | ( n18109 & n18128 ) | ( ~n18125 & n18128 ) ;
  assign n19015 = ( n19012 & ~n19013 ) | ( n19012 & n19014 ) | ( ~n19013 & n19014 ) ;
  assign n19016 = n19010 | n19015 ;
  assign n18990 = n18981 | n18989 ;
  assign n18991 = ~x123 & n18977 ;
  assign n18992 = ( x123 & ~n18990 ) | ( x123 & n18991 ) | ( ~n18990 & n18991 ) ;
  assign n18993 = x124 | n18992 ;
  assign n19002 = ( n18964 & ~n18975 ) | ( n18964 & 1'b0 ) | ( ~n18975 & 1'b0 ) ;
  assign n19003 = ( x123 & ~n18972 ) | ( x123 & n19002 ) | ( ~n18972 & n19002 ) ;
  assign n19004 = ( n18989 & ~n19003 ) | ( n18989 & 1'b0 ) | ( ~n19003 & 1'b0 ) ;
  assign n19005 = n19001 | n19004 ;
  assign n19006 = ( n18993 & ~n19005 ) | ( n18993 & 1'b0 ) | ( ~n19005 & 1'b0 ) ;
  assign n19017 = ~x125 & n19006 ;
  assign n19018 = ( x125 & ~n19016 ) | ( x125 & n19017 ) | ( ~n19016 & n19017 ) ;
  assign n19019 = x126 | n19018 ;
  assign n19020 = ( n18993 & ~n19004 ) | ( n18993 & 1'b0 ) | ( ~n19004 & 1'b0 ) ;
  assign n19021 = ( x125 & ~n19001 ) | ( x125 & n19020 ) | ( ~n19001 & n19020 ) ;
  assign n19022 = ( n19015 & ~n19021 ) | ( n19015 & 1'b0 ) | ( ~n19021 & 1'b0 ) ;
  assign n19023 = ( n19019 & ~n19022 ) | ( n19019 & 1'b0 ) | ( ~n19022 & 1'b0 ) ;
  assign n19024 = ( x127 & ~n18134 ) | ( x127 & n19023 ) | ( ~n18134 & n19023 ) ;
  assign n19025 = n262 | n279 ;
  assign n19026 = ( n274 & ~n195 ) | ( n274 & n19025 ) | ( ~n195 & n19025 ) ;
  assign n19027 = n195 | n19026 ;
  assign n19028 = x65 | x66 ;
  assign n19029 = ( n215 & ~n130 ) | ( n215 & n19028 ) | ( ~n130 & n19028 ) ;
  assign n19030 = n130 | n19029 ;
  assign n19031 = ( n462 & ~n423 ) | ( n462 & n19030 ) | ( ~n423 & n19030 ) ;
  assign n19032 = n423 | n19031 ;
  assign n19033 = ( n133 & ~n139 ) | ( n133 & 1'b0 ) | ( ~n139 & 1'b0 ) ;
  assign n19034 = ~n263 & n19033 ;
  assign n19035 = ~n262 & n19034 ;
  assign n19036 = ~n274 & n19035 ;
  assign n19037 = ( x63 & ~n19036 ) | ( x63 & 1'b0 ) | ( ~n19036 & 1'b0 ) ;
  assign n19038 = ( x65 & ~n19037 ) | ( x65 & n129 ) | ( ~n19037 & n129 ) ;
  assign n19039 = ( n257 & ~n19038 ) | ( n257 & 1'b0 ) | ( ~n19038 & 1'b0 ) ;
  assign n19040 = ( x62 & ~n19039 ) | ( x62 & 1'b0 ) | ( ~n19039 & 1'b0 ) ;
  assign n19041 = ( n275 & ~n19038 ) | ( n275 & 1'b0 ) | ( ~n19038 & 1'b0 ) ;
  assign n19042 = n19040 | n19041 ;
  assign n19043 = ( n284 & ~n19037 ) | ( n284 & 1'b0 ) | ( ~n19037 & 1'b0 ) ;
  assign n19044 = ~n19038 & n19043 ;
  assign n19045 = ( n295 & ~n19038 ) | ( n295 & 1'b0 ) | ( ~n19038 & 1'b0 ) ;
  assign n19046 = ( n19037 & ~n19045 ) | ( n19037 & 1'b0 ) | ( ~n19045 & 1'b0 ) ;
  assign n19047 = n19044 | n19046 ;
  assign n19048 = ( x65 & ~n19042 ) | ( x65 & n299 ) | ( ~n19042 & n299 ) ;
  assign n19049 = ( x66 & ~n19047 ) | ( x66 & n19048 ) | ( ~n19047 & n19048 ) ;
  assign n19050 = ( n311 & ~n19049 ) | ( n311 & 1'b0 ) | ( ~n19049 & 1'b0 ) ;
  assign n19051 = ( n19042 & ~n19050 ) | ( n19042 & 1'b0 ) | ( ~n19050 & 1'b0 ) ;
  assign n19052 = ( n319 & ~n19041 ) | ( n319 & 1'b0 ) | ( ~n19041 & 1'b0 ) ;
  assign n19053 = ( n19040 & ~n19049 ) | ( n19040 & n19052 ) | ( ~n19049 & n19052 ) ;
  assign n19054 = ~n19040 & n19053 ;
  assign n19055 = n19051 | n19054 ;
  assign n19056 = ( n328 & ~n19049 ) | ( n328 & 1'b0 ) | ( ~n19049 & 1'b0 ) ;
  assign n19057 = ( x61 & ~n19056 ) | ( x61 & 1'b0 ) | ( ~n19056 & 1'b0 ) ;
  assign n19058 = ( n335 & ~n19049 ) | ( n335 & 1'b0 ) | ( ~n19049 & 1'b0 ) ;
  assign n19059 = n19057 | n19058 ;
  assign n19060 = ( x65 & ~n19059 ) | ( x65 & n338 ) | ( ~n19059 & n338 ) ;
  assign n19061 = ( x66 & ~n19055 ) | ( x66 & n19060 ) | ( ~n19055 & n19060 ) ;
  assign n19062 = ( n19046 & ~n19044 ) | ( n19046 & n19048 ) | ( ~n19044 & n19048 ) ;
  assign n19063 = ~n19046 & n19062 ;
  assign n19064 = ( x66 & ~n19063 ) | ( x66 & n19048 ) | ( ~n19063 & n19048 ) ;
  assign n19065 = ( n345 & n19049 ) | ( n345 & n19064 ) | ( n19049 & n19064 ) ;
  assign n19066 = n19064 | n19065 ;
  assign n19067 = ( n19047 & ~n19066 ) | ( n19047 & n19065 ) | ( ~n19066 & n19065 ) ;
  assign n19070 = ~x66 & n19047 ;
  assign n19068 = ( x66 & ~n19044 ) | ( x66 & 1'b0 ) | ( ~n19044 & 1'b0 ) ;
  assign n19069 = ~n19046 & n19068 ;
  assign n19071 = ( n19048 & ~n19070 ) | ( n19048 & n19069 ) | ( ~n19070 & n19069 ) ;
  assign n19072 = ( n345 & ~n19071 ) | ( n345 & n19069 ) | ( ~n19071 & n19069 ) ;
  assign n19073 = ~n345 & n19072 ;
  assign n19074 = n19067 | n19073 ;
  assign n19103 = ~x67 & n19074 ;
  assign n19104 = ( n357 & ~n19061 ) | ( n357 & n19103 ) | ( ~n19061 & n19103 ) ;
  assign n19105 = ~n357 & n19104 ;
  assign n19075 = ( x67 & ~n19074 ) | ( x67 & n19061 ) | ( ~n19074 & n19061 ) ;
  assign n19106 = ~n357 & n19075 ;
  assign n19107 = ( n357 & n19106 ) | ( n357 & n19074 ) | ( n19106 & n19074 ) ;
  assign n19108 = n19105 | n19107 ;
  assign n19076 = ( x66 & ~n19054 ) | ( x66 & 1'b0 ) | ( ~n19054 & 1'b0 ) ;
  assign n19077 = ~n19051 & n19076 ;
  assign n19078 = ~n19060 & n19077 ;
  assign n19079 = n19055 | x66 ;
  assign n19080 = ( n19079 & ~x66 ) | ( n19079 & n19077 ) | ( ~x66 & n19077 ) ;
  assign n19081 = ( n19060 & ~n19080 ) | ( n19060 & 1'b0 ) | ( ~n19080 & 1'b0 ) ;
  assign n19082 = ( n19078 & ~n357 ) | ( n19078 & n19081 ) | ( ~n357 & n19081 ) ;
  assign n19083 = ~n19075 & n19082 ;
  assign n19084 = ~n19060 & n19080 ;
  assign n19085 = ( x66 & ~n19084 ) | ( x66 & n19080 ) | ( ~n19084 & n19080 ) ;
  assign n19086 = ( n357 & ~n19075 ) | ( n357 & n19085 ) | ( ~n19075 & n19085 ) ;
  assign n19087 = ~n357 & n19086 ;
  assign n19088 = ( n19055 & ~n19087 ) | ( n19055 & 1'b0 ) | ( ~n19087 & 1'b0 ) ;
  assign n19089 = n19083 | n19088 ;
  assign n19090 = ( n375 & ~n19075 ) | ( n375 & 1'b0 ) | ( ~n19075 & 1'b0 ) ;
  assign n19091 = ( n19059 & ~n19090 ) | ( n19059 & 1'b0 ) | ( ~n19090 & 1'b0 ) ;
  assign n19092 = ( n380 & ~n19058 ) | ( n380 & 1'b0 ) | ( ~n19058 & 1'b0 ) ;
  assign n19093 = ( n19057 & ~n19075 ) | ( n19057 & n19092 ) | ( ~n19075 & n19092 ) ;
  assign n19094 = ~n19057 & n19093 ;
  assign n19095 = n19091 | n19094 ;
  assign n19096 = ( n390 & ~n19075 ) | ( n390 & 1'b0 ) | ( ~n19075 & 1'b0 ) ;
  assign n19097 = ( x60 & ~n19096 ) | ( x60 & 1'b0 ) | ( ~n19096 & 1'b0 ) ;
  assign n19098 = ( n396 & ~n19075 ) | ( n396 & 1'b0 ) | ( ~n19075 & 1'b0 ) ;
  assign n19099 = n19097 | n19098 ;
  assign n19100 = ( x65 & ~n19099 ) | ( x65 & n385 ) | ( ~n19099 & n385 ) ;
  assign n19101 = ( x66 & ~n19095 ) | ( x66 & n19100 ) | ( ~n19095 & n19100 ) ;
  assign n19102 = ( x67 & ~n19089 ) | ( x67 & n19101 ) | ( ~n19089 & n19101 ) ;
  assign n19109 = ( x68 & ~n19108 ) | ( x68 & n19102 ) | ( ~n19108 & n19102 ) ;
  assign n19110 = ( x67 & ~n19083 ) | ( x67 & 1'b0 ) | ( ~n19083 & 1'b0 ) ;
  assign n19111 = ~n19088 & n19110 ;
  assign n19113 = ~x67 & n19089 ;
  assign n19114 = ~x66 & n19095 ;
  assign n19115 = ( x66 & ~n19094 ) | ( x66 & 1'b0 ) | ( ~n19094 & 1'b0 ) ;
  assign n19116 = ~n19091 & n19115 ;
  assign n19117 = n19100 | n19116 ;
  assign n19118 = ~n19114 & n19117 ;
  assign n19119 = ( n19111 & n19113 ) | ( n19111 & n19118 ) | ( n19113 & n19118 ) ;
  assign n19112 = n19101 | n19111 ;
  assign n19120 = ( n19109 & ~n19119 ) | ( n19109 & n19112 ) | ( ~n19119 & n19112 ) ;
  assign n19121 = ( n431 & ~n19109 ) | ( n431 & n19120 ) | ( ~n19109 & n19120 ) ;
  assign n19122 = ~n431 & n19121 ;
  assign n19123 = n431 | n19109 ;
  assign n19124 = ~x67 & n19119 ;
  assign n19125 = ( x67 & ~n19123 ) | ( x67 & n19124 ) | ( ~n19123 & n19124 ) ;
  assign n19126 = ( n19089 & ~n19125 ) | ( n19089 & 1'b0 ) | ( ~n19125 & 1'b0 ) ;
  assign n19127 = n19122 | n19126 ;
  assign n19131 = n19114 | n19116 ;
  assign n19132 = n19100 &  n19131 ;
  assign n19133 = ~n431 & n19117 ;
  assign n19134 = ( n19109 & ~n19132 ) | ( n19109 & n19133 ) | ( ~n19132 & n19133 ) ;
  assign n19135 = ~n19109 & n19134 ;
  assign n19136 = ~x66 & n19132 ;
  assign n19137 = ( x66 & ~n19123 ) | ( x66 & n19136 ) | ( ~n19123 & n19136 ) ;
  assign n19138 = ( n19095 & ~n19137 ) | ( n19095 & 1'b0 ) | ( ~n19137 & 1'b0 ) ;
  assign n19139 = n19135 | n19138 ;
  assign n19140 = ( n457 & ~n19109 ) | ( n457 & 1'b0 ) | ( ~n19109 & 1'b0 ) ;
  assign n19141 = ( n19099 & ~n19140 ) | ( n19099 & 1'b0 ) | ( ~n19140 & 1'b0 ) ;
  assign n19142 = ( n464 & ~n19098 ) | ( n464 & 1'b0 ) | ( ~n19098 & 1'b0 ) ;
  assign n19143 = ( n19097 & ~n19109 ) | ( n19097 & n19142 ) | ( ~n19109 & n19142 ) ;
  assign n19144 = ~n19097 & n19143 ;
  assign n19145 = n19141 | n19144 ;
  assign n19146 = ( n474 & ~n19109 ) | ( n474 & 1'b0 ) | ( ~n19109 & 1'b0 ) ;
  assign n19147 = ( x59 & ~n19146 ) | ( x59 & 1'b0 ) | ( ~n19146 & 1'b0 ) ;
  assign n19148 = ( n480 & ~n19109 ) | ( n480 & 1'b0 ) | ( ~n19109 & 1'b0 ) ;
  assign n19149 = n19147 | n19148 ;
  assign n19150 = ( x65 & ~n19149 ) | ( x65 & n483 ) | ( ~n19149 & n483 ) ;
  assign n19151 = ( x66 & ~n19145 ) | ( x66 & n19150 ) | ( ~n19145 & n19150 ) ;
  assign n19152 = ( x67 & ~n19139 ) | ( x67 & n19151 ) | ( ~n19139 & n19151 ) ;
  assign n19153 = ( x68 & ~n19127 ) | ( x68 & n19152 ) | ( ~n19127 & n19152 ) ;
  assign n19156 = n19108 | x68 ;
  assign n19154 = ( x68 & ~n19107 ) | ( x68 & 1'b0 ) | ( ~n19107 & 1'b0 ) ;
  assign n19155 = ~n19105 & n19154 ;
  assign n19157 = ( n19156 & ~x68 ) | ( n19156 & n19155 ) | ( ~x68 & n19155 ) ;
  assign n19158 = ( n19112 & n19113 ) | ( n19112 & n19157 ) | ( n19113 & n19157 ) ;
  assign n19159 = ~n19113 & n19158 ;
  assign n19160 = n431 | n19159 ;
  assign n19161 = ~n19102 & n19155 ;
  assign n19162 = ( n19102 & ~n19160 ) | ( n19102 & n19161 ) | ( ~n19160 & n19161 ) ;
  assign n19163 = ~n19109 & n19162 ;
  assign n19164 = ~x68 & n19159 ;
  assign n19165 = ( x68 & ~n19123 ) | ( x68 & n19164 ) | ( ~n19123 & n19164 ) ;
  assign n19166 = ( n19108 & ~n19165 ) | ( n19108 & 1'b0 ) | ( ~n19165 & 1'b0 ) ;
  assign n19167 = n19163 | n19166 ;
  assign n19168 = x69 | n19167 ;
  assign n19169 = x69 &  n19167 ;
  assign n19170 = ( n19168 & ~n19169 ) | ( n19168 & 1'b0 ) | ( ~n19169 & 1'b0 ) ;
  assign n19171 = n509 | n19170 ;
  assign n19172 = n19153 | n19171 ;
  assign n19175 = n431 &  n19167 ;
  assign n19176 = n19172 &  n19175 ;
  assign n19177 = n19153 &  n19170 ;
  assign n19173 = ~n431 & n19167 ;
  assign n19178 = ( n19153 & n19170 ) | ( n19153 & n19173 ) | ( n19170 & n19173 ) ;
  assign n19179 = ( n19176 & ~n19177 ) | ( n19176 & n19178 ) | ( ~n19177 & n19178 ) ;
  assign n19183 = ( n19127 & ~n19173 ) | ( n19127 & 1'b0 ) | ( ~n19173 & 1'b0 ) ;
  assign n19184 = n19172 &  n19183 ;
  assign n19128 = x68 | n19127 ;
  assign n19129 = x68 &  n19127 ;
  assign n19130 = ( n19128 & ~n19129 ) | ( n19128 & 1'b0 ) | ( ~n19129 & 1'b0 ) ;
  assign n19185 = n19130 &  n19152 ;
  assign n19174 = ( n19172 & ~n19173 ) | ( n19172 & 1'b0 ) | ( ~n19173 & 1'b0 ) ;
  assign n19186 = ( n19130 & ~n19174 ) | ( n19130 & n19152 ) | ( ~n19174 & n19152 ) ;
  assign n19187 = ( n19184 & ~n19185 ) | ( n19184 & n19186 ) | ( ~n19185 & n19186 ) ;
  assign n19191 = ( n19139 & ~n19173 ) | ( n19139 & 1'b0 ) | ( ~n19173 & 1'b0 ) ;
  assign n19192 = n19172 &  n19191 ;
  assign n19180 = x67 | n19139 ;
  assign n19181 = x67 &  n19139 ;
  assign n19182 = ( n19180 & ~n19181 ) | ( n19180 & 1'b0 ) | ( ~n19181 & 1'b0 ) ;
  assign n19194 = ( n19151 & n19174 ) | ( n19151 & n19182 ) | ( n19174 & n19182 ) ;
  assign n19193 = n19151 | n19182 ;
  assign n19195 = ( n19192 & ~n19194 ) | ( n19192 & n19193 ) | ( ~n19194 & n19193 ) ;
  assign n19196 = ( n19145 & ~n19173 ) | ( n19145 & 1'b0 ) | ( ~n19173 & 1'b0 ) ;
  assign n19197 = n19172 &  n19196 ;
  assign n19188 = x66 | n19145 ;
  assign n19189 = x66 &  n19145 ;
  assign n19190 = ( n19188 & ~n19189 ) | ( n19188 & 1'b0 ) | ( ~n19189 & 1'b0 ) ;
  assign n19199 = ( n19150 & n19174 ) | ( n19150 & n19190 ) | ( n19174 & n19190 ) ;
  assign n19198 = n19150 | n19190 ;
  assign n19200 = ( n19197 & ~n19199 ) | ( n19197 & n19198 ) | ( ~n19199 & n19198 ) ;
  assign n19201 = ( x65 & ~n483 ) | ( x65 & n19149 ) | ( ~n483 & n19149 ) ;
  assign n19202 = ( n19150 & ~x65 ) | ( n19150 & n19201 ) | ( ~x65 & n19201 ) ;
  assign n19203 = ~n19174 & n19202 ;
  assign n19204 = ( n19149 & ~n19173 ) | ( n19149 & 1'b0 ) | ( ~n19173 & 1'b0 ) ;
  assign n19205 = n19172 &  n19204 ;
  assign n19206 = n19203 | n19205 ;
  assign n19207 = ( x64 & ~n19174 ) | ( x64 & 1'b0 ) | ( ~n19174 & 1'b0 ) ;
  assign n19208 = ( x58 & ~n19207 ) | ( x58 & 1'b0 ) | ( ~n19207 & 1'b0 ) ;
  assign n19209 = ( n483 & ~n19174 ) | ( n483 & 1'b0 ) | ( ~n19174 & 1'b0 ) ;
  assign n19210 = n19208 | n19209 ;
  assign n19211 = ( x65 & ~n19210 ) | ( x65 & n553 ) | ( ~n19210 & n553 ) ;
  assign n19212 = ( x66 & ~n19206 ) | ( x66 & n19211 ) | ( ~n19206 & n19211 ) ;
  assign n19213 = ( x67 & ~n19200 ) | ( x67 & n19212 ) | ( ~n19200 & n19212 ) ;
  assign n19214 = ( x68 & ~n19195 ) | ( x68 & n19213 ) | ( ~n19195 & n19213 ) ;
  assign n19215 = ( x69 & ~n19187 ) | ( x69 & n19214 ) | ( ~n19187 & n19214 ) ;
  assign n19222 = ( x70 & ~n563 ) | ( x70 & n19215 ) | ( ~n563 & n19215 ) ;
  assign n19221 = x70 &  n19215 ;
  assign n19223 = ( n19179 & ~n19222 ) | ( n19179 & n19221 ) | ( ~n19222 & n19221 ) ;
  assign n19216 = ( x70 & ~n19179 ) | ( x70 & n19215 ) | ( ~n19179 & n19215 ) ;
  assign n19217 = n563 | n19216 ;
  assign n19224 = n19187 &  n19217 ;
  assign n19218 = x69 | n19187 ;
  assign n19219 = x69 &  n19187 ;
  assign n19220 = ( n19218 & ~n19219 ) | ( n19218 & 1'b0 ) | ( ~n19219 & 1'b0 ) ;
  assign n19228 = ( n563 & n19214 ) | ( n563 & n19220 ) | ( n19214 & n19220 ) ;
  assign n19229 = ( n19214 & ~n19216 ) | ( n19214 & n19220 ) | ( ~n19216 & n19220 ) ;
  assign n19230 = ~n19228 & n19229 ;
  assign n19231 = n19224 | n19230 ;
  assign n19232 = n19195 &  n19217 ;
  assign n19225 = x68 | n19195 ;
  assign n19226 = x68 &  n19195 ;
  assign n19227 = ( n19225 & ~n19226 ) | ( n19225 & 1'b0 ) | ( ~n19226 & 1'b0 ) ;
  assign n19236 = ( n563 & n19213 ) | ( n563 & n19227 ) | ( n19213 & n19227 ) ;
  assign n19237 = ( n19213 & ~n19216 ) | ( n19213 & n19227 ) | ( ~n19216 & n19227 ) ;
  assign n19238 = ~n19236 & n19237 ;
  assign n19239 = n19232 | n19238 ;
  assign n19240 = n19200 &  n19217 ;
  assign n19233 = x67 | n19200 ;
  assign n19234 = x67 &  n19200 ;
  assign n19235 = ( n19233 & ~n19234 ) | ( n19233 & 1'b0 ) | ( ~n19234 & 1'b0 ) ;
  assign n19244 = ( n563 & n19212 ) | ( n563 & n19235 ) | ( n19212 & n19235 ) ;
  assign n19245 = ( n19212 & ~n19216 ) | ( n19212 & n19235 ) | ( ~n19216 & n19235 ) ;
  assign n19246 = ~n19244 & n19245 ;
  assign n19247 = n19240 | n19246 ;
  assign n19248 = n19206 &  n19217 ;
  assign n19241 = x66 | n19206 ;
  assign n19242 = x66 &  n19206 ;
  assign n19243 = ( n19241 & ~n19242 ) | ( n19241 & 1'b0 ) | ( ~n19242 & 1'b0 ) ;
  assign n19249 = ( n563 & n19211 ) | ( n563 & n19243 ) | ( n19211 & n19243 ) ;
  assign n19250 = ( n19211 & ~n19216 ) | ( n19211 & n19243 ) | ( ~n19216 & n19243 ) ;
  assign n19251 = ~n19249 & n19250 ;
  assign n19252 = n19248 | n19251 ;
  assign n19253 = n19210 &  n19217 ;
  assign n19254 = ( x65 & ~x58 ) | ( x65 & n19207 ) | ( ~x58 & n19207 ) ;
  assign n19255 = ( x58 & ~n19207 ) | ( x58 & x65 ) | ( ~n19207 & x65 ) ;
  assign n19256 = ( n19254 & ~x65 ) | ( n19254 & n19255 ) | ( ~x65 & n19255 ) ;
  assign n19257 = ( n553 & ~n563 ) | ( n553 & n19256 ) | ( ~n563 & n19256 ) ;
  assign n19258 = ( n553 & n19216 ) | ( n553 & n19256 ) | ( n19216 & n19256 ) ;
  assign n19259 = ( n19257 & ~n19258 ) | ( n19257 & 1'b0 ) | ( ~n19258 & 1'b0 ) ;
  assign n19260 = n19253 | n19259 ;
  assign n19261 = ( n614 & ~n19216 ) | ( n614 & 1'b0 ) | ( ~n19216 & 1'b0 ) ;
  assign n19262 = ( x57 & ~n19261 ) | ( x57 & 1'b0 ) | ( ~n19261 & 1'b0 ) ;
  assign n19263 = ( n621 & ~n19216 ) | ( n621 & 1'b0 ) | ( ~n19216 & 1'b0 ) ;
  assign n19264 = n19262 | n19263 ;
  assign n19265 = ( x65 & ~n19264 ) | ( x65 & n624 ) | ( ~n19264 & n624 ) ;
  assign n19266 = ( x66 & ~n19260 ) | ( x66 & n19265 ) | ( ~n19260 & n19265 ) ;
  assign n19267 = ( x67 & ~n19252 ) | ( x67 & n19266 ) | ( ~n19252 & n19266 ) ;
  assign n19268 = ( x68 & ~n19247 ) | ( x68 & n19267 ) | ( ~n19247 & n19267 ) ;
  assign n19269 = ( x69 & ~n19239 ) | ( x69 & n19268 ) | ( ~n19239 & n19268 ) ;
  assign n19270 = ( x70 & ~n19231 ) | ( x70 & n19269 ) | ( ~n19231 & n19269 ) ;
  assign n19271 = ( x71 & ~n19223 ) | ( x71 & n19270 ) | ( ~n19223 & n19270 ) ;
  assign n19272 = n633 | n19271 ;
  assign n19273 = n19223 &  n19272 ;
  assign n19277 = ( n633 & n19223 ) | ( n633 & n19270 ) | ( n19223 & n19270 ) ;
  assign n19278 = ( x71 & ~n19277 ) | ( x71 & n19223 ) | ( ~n19277 & n19223 ) ;
  assign n19279 = ~x71 & n19278 ;
  assign n19280 = n19273 | n19279 ;
  assign n19281 = ~x72 & n19280 ;
  assign n19282 = n19231 &  n19272 ;
  assign n19274 = x70 | n19231 ;
  assign n19275 = x70 &  n19231 ;
  assign n19276 = ( n19274 & ~n19275 ) | ( n19274 & 1'b0 ) | ( ~n19275 & 1'b0 ) ;
  assign n19286 = ( n633 & n19269 ) | ( n633 & n19276 ) | ( n19269 & n19276 ) ;
  assign n19287 = ( n19269 & ~n19271 ) | ( n19269 & n19276 ) | ( ~n19271 & n19276 ) ;
  assign n19288 = ~n19286 & n19287 ;
  assign n19289 = n19282 | n19288 ;
  assign n19290 = n19239 &  n19272 ;
  assign n19283 = x69 | n19239 ;
  assign n19284 = x69 &  n19239 ;
  assign n19285 = ( n19283 & ~n19284 ) | ( n19283 & 1'b0 ) | ( ~n19284 & 1'b0 ) ;
  assign n19294 = ( n633 & n19268 ) | ( n633 & n19285 ) | ( n19268 & n19285 ) ;
  assign n19295 = ( n19268 & ~n19271 ) | ( n19268 & n19285 ) | ( ~n19271 & n19285 ) ;
  assign n19296 = ~n19294 & n19295 ;
  assign n19297 = n19290 | n19296 ;
  assign n19298 = n19247 &  n19272 ;
  assign n19291 = x68 | n19247 ;
  assign n19292 = x68 &  n19247 ;
  assign n19293 = ( n19291 & ~n19292 ) | ( n19291 & 1'b0 ) | ( ~n19292 & 1'b0 ) ;
  assign n19302 = ( n633 & n19267 ) | ( n633 & n19293 ) | ( n19267 & n19293 ) ;
  assign n19303 = ( n19267 & ~n19271 ) | ( n19267 & n19293 ) | ( ~n19271 & n19293 ) ;
  assign n19304 = ~n19302 & n19303 ;
  assign n19305 = n19298 | n19304 ;
  assign n19306 = n19252 &  n19272 ;
  assign n19299 = x67 | n19252 ;
  assign n19300 = x67 &  n19252 ;
  assign n19301 = ( n19299 & ~n19300 ) | ( n19299 & 1'b0 ) | ( ~n19300 & 1'b0 ) ;
  assign n19310 = ( n633 & n19266 ) | ( n633 & n19301 ) | ( n19266 & n19301 ) ;
  assign n19311 = ( n19266 & ~n19271 ) | ( n19266 & n19301 ) | ( ~n19271 & n19301 ) ;
  assign n19312 = ~n19310 & n19311 ;
  assign n19313 = n19306 | n19312 ;
  assign n19314 = n19260 &  n19272 ;
  assign n19307 = x66 | n19260 ;
  assign n19308 = x66 &  n19260 ;
  assign n19309 = ( n19307 & ~n19308 ) | ( n19307 & 1'b0 ) | ( ~n19308 & 1'b0 ) ;
  assign n19318 = ( n633 & n19265 ) | ( n633 & n19309 ) | ( n19265 & n19309 ) ;
  assign n19319 = ( n19265 & ~n19271 ) | ( n19265 & n19309 ) | ( ~n19271 & n19309 ) ;
  assign n19320 = ~n19318 & n19319 ;
  assign n19321 = n19314 | n19320 ;
  assign n19322 = n19264 &  n19272 ;
  assign n19315 = x65 &  n19264 ;
  assign n19316 = x65 | n19263 ;
  assign n19317 = n19262 | n19316 ;
  assign n19323 = ~n19315 & n19317 ;
  assign n19324 = ( n624 & ~n633 ) | ( n624 & n19323 ) | ( ~n633 & n19323 ) ;
  assign n19325 = ( n624 & n19271 ) | ( n624 & n19323 ) | ( n19271 & n19323 ) ;
  assign n19326 = ( n19324 & ~n19325 ) | ( n19324 & 1'b0 ) | ( ~n19325 & 1'b0 ) ;
  assign n19327 = n19322 | n19326 ;
  assign n19328 = ( n657 & ~n19271 ) | ( n657 & 1'b0 ) | ( ~n19271 & 1'b0 ) ;
  assign n19329 = ( x56 & ~n19328 ) | ( x56 & 1'b0 ) | ( ~n19328 & 1'b0 ) ;
  assign n19330 = ( n663 & ~n19271 ) | ( n663 & 1'b0 ) | ( ~n19271 & 1'b0 ) ;
  assign n19331 = n19329 | n19330 ;
  assign n19332 = ( x65 & ~n19331 ) | ( x65 & n666 ) | ( ~n19331 & n666 ) ;
  assign n19333 = ( x66 & ~n19327 ) | ( x66 & n19332 ) | ( ~n19327 & n19332 ) ;
  assign n19334 = ( x67 & ~n19321 ) | ( x67 & n19333 ) | ( ~n19321 & n19333 ) ;
  assign n19335 = ( x68 & ~n19313 ) | ( x68 & n19334 ) | ( ~n19313 & n19334 ) ;
  assign n19336 = ( x69 & ~n19305 ) | ( x69 & n19335 ) | ( ~n19305 & n19335 ) ;
  assign n19337 = ( x70 & ~n19297 ) | ( x70 & n19336 ) | ( ~n19297 & n19336 ) ;
  assign n19338 = ( x71 & ~n19289 ) | ( x71 & n19337 ) | ( ~n19289 & n19337 ) ;
  assign n19339 = ( x72 & ~n19273 ) | ( x72 & 1'b0 ) | ( ~n19273 & 1'b0 ) ;
  assign n19340 = ~n19279 & n19339 ;
  assign n19341 = ( n19338 & ~n19281 ) | ( n19338 & n19340 ) | ( ~n19281 & n19340 ) ;
  assign n19342 = ( n19281 & ~n716 ) | ( n19281 & n19341 ) | ( ~n716 & n19341 ) ;
  assign n19343 = n716 | n19342 ;
  assign n19350 = n633 &  n19223 ;
  assign n19351 = n19343 &  n19350 ;
  assign n19344 = ~n633 & n19280 ;
  assign n19345 = ( n19343 & ~n19344 ) | ( n19343 & 1'b0 ) | ( ~n19344 & 1'b0 ) ;
  assign n19349 = n19281 | n19340 ;
  assign n19353 = ( n19338 & n19345 ) | ( n19338 & n19349 ) | ( n19345 & n19349 ) ;
  assign n19352 = n19338 | n19349 ;
  assign n19354 = ( n19351 & ~n19353 ) | ( n19351 & n19352 ) | ( ~n19353 & n19352 ) ;
  assign n19358 = ( n19289 & ~n19344 ) | ( n19289 & 1'b0 ) | ( ~n19344 & 1'b0 ) ;
  assign n19359 = n19343 &  n19358 ;
  assign n19346 = x71 | n19289 ;
  assign n19347 = x71 &  n19289 ;
  assign n19348 = ( n19346 & ~n19347 ) | ( n19346 & 1'b0 ) | ( ~n19347 & 1'b0 ) ;
  assign n19361 = ( n19337 & n19345 ) | ( n19337 & n19348 ) | ( n19345 & n19348 ) ;
  assign n19360 = n19337 | n19348 ;
  assign n19362 = ( n19359 & ~n19361 ) | ( n19359 & n19360 ) | ( ~n19361 & n19360 ) ;
  assign n19366 = ( n19297 & ~n19344 ) | ( n19297 & 1'b0 ) | ( ~n19344 & 1'b0 ) ;
  assign n19367 = n19343 &  n19366 ;
  assign n19355 = x70 | n19297 ;
  assign n19356 = x70 &  n19297 ;
  assign n19357 = ( n19355 & ~n19356 ) | ( n19355 & 1'b0 ) | ( ~n19356 & 1'b0 ) ;
  assign n19369 = ( n19336 & n19345 ) | ( n19336 & n19357 ) | ( n19345 & n19357 ) ;
  assign n19368 = n19336 | n19357 ;
  assign n19370 = ( n19367 & ~n19369 ) | ( n19367 & n19368 ) | ( ~n19369 & n19368 ) ;
  assign n19374 = ( n19305 & ~n19344 ) | ( n19305 & 1'b0 ) | ( ~n19344 & 1'b0 ) ;
  assign n19375 = n19343 &  n19374 ;
  assign n19363 = x69 | n19305 ;
  assign n19364 = x69 &  n19305 ;
  assign n19365 = ( n19363 & ~n19364 ) | ( n19363 & 1'b0 ) | ( ~n19364 & 1'b0 ) ;
  assign n19377 = ( n19335 & n19345 ) | ( n19335 & n19365 ) | ( n19345 & n19365 ) ;
  assign n19376 = n19335 | n19365 ;
  assign n19378 = ( n19375 & ~n19377 ) | ( n19375 & n19376 ) | ( ~n19377 & n19376 ) ;
  assign n19382 = ( n19313 & ~n19344 ) | ( n19313 & 1'b0 ) | ( ~n19344 & 1'b0 ) ;
  assign n19383 = n19343 &  n19382 ;
  assign n19371 = x68 | n19313 ;
  assign n19372 = x68 &  n19313 ;
  assign n19373 = ( n19371 & ~n19372 ) | ( n19371 & 1'b0 ) | ( ~n19372 & 1'b0 ) ;
  assign n19385 = ( n19334 & n19345 ) | ( n19334 & n19373 ) | ( n19345 & n19373 ) ;
  assign n19384 = n19334 | n19373 ;
  assign n19386 = ( n19383 & ~n19385 ) | ( n19383 & n19384 ) | ( ~n19385 & n19384 ) ;
  assign n19390 = ( n19321 & ~n19344 ) | ( n19321 & 1'b0 ) | ( ~n19344 & 1'b0 ) ;
  assign n19391 = n19343 &  n19390 ;
  assign n19379 = x67 | n19321 ;
  assign n19380 = x67 &  n19321 ;
  assign n19381 = ( n19379 & ~n19380 ) | ( n19379 & 1'b0 ) | ( ~n19380 & 1'b0 ) ;
  assign n19393 = ( n19333 & n19345 ) | ( n19333 & n19381 ) | ( n19345 & n19381 ) ;
  assign n19392 = n19333 | n19381 ;
  assign n19394 = ( n19391 & ~n19393 ) | ( n19391 & n19392 ) | ( ~n19393 & n19392 ) ;
  assign n19395 = ( n19327 & ~n19344 ) | ( n19327 & 1'b0 ) | ( ~n19344 & 1'b0 ) ;
  assign n19396 = n19343 &  n19395 ;
  assign n19387 = x66 | n19327 ;
  assign n19388 = x66 &  n19327 ;
  assign n19389 = ( n19387 & ~n19388 ) | ( n19387 & 1'b0 ) | ( ~n19388 & 1'b0 ) ;
  assign n19398 = ( n19332 & n19345 ) | ( n19332 & n19389 ) | ( n19345 & n19389 ) ;
  assign n19397 = n19332 | n19389 ;
  assign n19399 = ( n19396 & ~n19398 ) | ( n19396 & n19397 ) | ( ~n19398 & n19397 ) ;
  assign n19400 = ( x65 & ~n666 ) | ( x65 & n19331 ) | ( ~n666 & n19331 ) ;
  assign n19401 = ( n19332 & ~x65 ) | ( n19332 & n19400 ) | ( ~x65 & n19400 ) ;
  assign n19402 = ~n19345 & n19401 ;
  assign n19403 = ( n19331 & ~n19344 ) | ( n19331 & 1'b0 ) | ( ~n19344 & 1'b0 ) ;
  assign n19404 = n19343 &  n19403 ;
  assign n19405 = n19402 | n19404 ;
  assign n19406 = ( x64 & ~n19345 ) | ( x64 & 1'b0 ) | ( ~n19345 & 1'b0 ) ;
  assign n19407 = ( x55 & ~n19406 ) | ( x55 & 1'b0 ) | ( ~n19406 & 1'b0 ) ;
  assign n19408 = ( n666 & ~n19345 ) | ( n666 & 1'b0 ) | ( ~n19345 & 1'b0 ) ;
  assign n19409 = n19407 | n19408 ;
  assign n19410 = ( x65 & ~n19409 ) | ( x65 & n782 ) | ( ~n19409 & n782 ) ;
  assign n19411 = ( x66 & ~n19405 ) | ( x66 & n19410 ) | ( ~n19405 & n19410 ) ;
  assign n19412 = ( x67 & ~n19399 ) | ( x67 & n19411 ) | ( ~n19399 & n19411 ) ;
  assign n19413 = ( x68 & ~n19394 ) | ( x68 & n19412 ) | ( ~n19394 & n19412 ) ;
  assign n19414 = ( x69 & ~n19386 ) | ( x69 & n19413 ) | ( ~n19386 & n19413 ) ;
  assign n19415 = ( x70 & ~n19378 ) | ( x70 & n19414 ) | ( ~n19378 & n19414 ) ;
  assign n19416 = ( x71 & ~n19370 ) | ( x71 & n19415 ) | ( ~n19370 & n19415 ) ;
  assign n19417 = ( x72 & ~n19362 ) | ( x72 & n19416 ) | ( ~n19362 & n19416 ) ;
  assign n19424 = ( x73 & ~n794 ) | ( x73 & n19417 ) | ( ~n794 & n19417 ) ;
  assign n19423 = x73 &  n19417 ;
  assign n19425 = ( n19354 & ~n19424 ) | ( n19354 & n19423 ) | ( ~n19424 & n19423 ) ;
  assign n19418 = ( x73 & ~n19354 ) | ( x73 & n19417 ) | ( ~n19354 & n19417 ) ;
  assign n19419 = n794 | n19418 ;
  assign n19426 = n19362 &  n19419 ;
  assign n19420 = x72 | n19362 ;
  assign n19421 = x72 &  n19362 ;
  assign n19422 = ( n19420 & ~n19421 ) | ( n19420 & 1'b0 ) | ( ~n19421 & 1'b0 ) ;
  assign n19430 = ( n794 & n19416 ) | ( n794 & n19422 ) | ( n19416 & n19422 ) ;
  assign n19431 = ( n19416 & ~n19418 ) | ( n19416 & n19422 ) | ( ~n19418 & n19422 ) ;
  assign n19432 = ~n19430 & n19431 ;
  assign n19433 = n19426 | n19432 ;
  assign n19434 = n19370 &  n19419 ;
  assign n19427 = x71 | n19370 ;
  assign n19428 = x71 &  n19370 ;
  assign n19429 = ( n19427 & ~n19428 ) | ( n19427 & 1'b0 ) | ( ~n19428 & 1'b0 ) ;
  assign n19438 = ( n794 & n19415 ) | ( n794 & n19429 ) | ( n19415 & n19429 ) ;
  assign n19439 = ( n19415 & ~n19418 ) | ( n19415 & n19429 ) | ( ~n19418 & n19429 ) ;
  assign n19440 = ~n19438 & n19439 ;
  assign n19441 = n19434 | n19440 ;
  assign n19442 = n19378 &  n19419 ;
  assign n19435 = x70 | n19378 ;
  assign n19436 = x70 &  n19378 ;
  assign n19437 = ( n19435 & ~n19436 ) | ( n19435 & 1'b0 ) | ( ~n19436 & 1'b0 ) ;
  assign n19446 = ( n794 & n19414 ) | ( n794 & n19437 ) | ( n19414 & n19437 ) ;
  assign n19447 = ( n19414 & ~n19418 ) | ( n19414 & n19437 ) | ( ~n19418 & n19437 ) ;
  assign n19448 = ~n19446 & n19447 ;
  assign n19449 = n19442 | n19448 ;
  assign n19450 = n19386 &  n19419 ;
  assign n19443 = x69 | n19386 ;
  assign n19444 = x69 &  n19386 ;
  assign n19445 = ( n19443 & ~n19444 ) | ( n19443 & 1'b0 ) | ( ~n19444 & 1'b0 ) ;
  assign n19454 = ( n794 & n19413 ) | ( n794 & n19445 ) | ( n19413 & n19445 ) ;
  assign n19455 = ( n19413 & ~n19418 ) | ( n19413 & n19445 ) | ( ~n19418 & n19445 ) ;
  assign n19456 = ~n19454 & n19455 ;
  assign n19457 = n19450 | n19456 ;
  assign n19458 = n19394 &  n19419 ;
  assign n19451 = x68 | n19394 ;
  assign n19452 = x68 &  n19394 ;
  assign n19453 = ( n19451 & ~n19452 ) | ( n19451 & 1'b0 ) | ( ~n19452 & 1'b0 ) ;
  assign n19462 = ( n794 & n19412 ) | ( n794 & n19453 ) | ( n19412 & n19453 ) ;
  assign n19463 = ( n19412 & ~n19418 ) | ( n19412 & n19453 ) | ( ~n19418 & n19453 ) ;
  assign n19464 = ~n19462 & n19463 ;
  assign n19465 = n19458 | n19464 ;
  assign n19466 = n19399 &  n19419 ;
  assign n19459 = x67 | n19399 ;
  assign n19460 = x67 &  n19399 ;
  assign n19461 = ( n19459 & ~n19460 ) | ( n19459 & 1'b0 ) | ( ~n19460 & 1'b0 ) ;
  assign n19470 = ( n794 & n19411 ) | ( n794 & n19461 ) | ( n19411 & n19461 ) ;
  assign n19471 = ( n19411 & ~n19418 ) | ( n19411 & n19461 ) | ( ~n19418 & n19461 ) ;
  assign n19472 = ~n19470 & n19471 ;
  assign n19473 = n19466 | n19472 ;
  assign n19474 = n19405 &  n19419 ;
  assign n19467 = x66 | n19405 ;
  assign n19468 = x66 &  n19405 ;
  assign n19469 = ( n19467 & ~n19468 ) | ( n19467 & 1'b0 ) | ( ~n19468 & 1'b0 ) ;
  assign n19475 = ( n794 & n19410 ) | ( n794 & n19469 ) | ( n19410 & n19469 ) ;
  assign n19476 = ( n19410 & ~n19418 ) | ( n19410 & n19469 ) | ( ~n19418 & n19469 ) ;
  assign n19477 = ~n19475 & n19476 ;
  assign n19478 = n19474 | n19477 ;
  assign n19479 = n19409 &  n19419 ;
  assign n19480 = ( x65 & ~x55 ) | ( x65 & n19406 ) | ( ~x55 & n19406 ) ;
  assign n19481 = ( x55 & ~n19406 ) | ( x55 & x65 ) | ( ~n19406 & x65 ) ;
  assign n19482 = ( n19480 & ~x65 ) | ( n19480 & n19481 ) | ( ~x65 & n19481 ) ;
  assign n19483 = ( n782 & ~n794 ) | ( n782 & n19482 ) | ( ~n794 & n19482 ) ;
  assign n19484 = ( n782 & n19418 ) | ( n782 & n19482 ) | ( n19418 & n19482 ) ;
  assign n19485 = ( n19483 & ~n19484 ) | ( n19483 & 1'b0 ) | ( ~n19484 & 1'b0 ) ;
  assign n19486 = n19479 | n19485 ;
  assign n19487 = ( n869 & ~n19418 ) | ( n869 & 1'b0 ) | ( ~n19418 & 1'b0 ) ;
  assign n19488 = ( x54 & ~n19487 ) | ( x54 & 1'b0 ) | ( ~n19487 & 1'b0 ) ;
  assign n19489 = ( n875 & ~n19418 ) | ( n875 & 1'b0 ) | ( ~n19418 & 1'b0 ) ;
  assign n19490 = n19488 | n19489 ;
  assign n19491 = ( x65 & ~n19490 ) | ( x65 & n878 ) | ( ~n19490 & n878 ) ;
  assign n19492 = ( x66 & ~n19486 ) | ( x66 & n19491 ) | ( ~n19486 & n19491 ) ;
  assign n19493 = ( x67 & ~n19478 ) | ( x67 & n19492 ) | ( ~n19478 & n19492 ) ;
  assign n19494 = ( x68 & ~n19473 ) | ( x68 & n19493 ) | ( ~n19473 & n19493 ) ;
  assign n19495 = ( x69 & ~n19465 ) | ( x69 & n19494 ) | ( ~n19465 & n19494 ) ;
  assign n19496 = ( x70 & ~n19457 ) | ( x70 & n19495 ) | ( ~n19457 & n19495 ) ;
  assign n19497 = ( x71 & ~n19449 ) | ( x71 & n19496 ) | ( ~n19449 & n19496 ) ;
  assign n19498 = ( x72 & ~n19441 ) | ( x72 & n19497 ) | ( ~n19441 & n19497 ) ;
  assign n19499 = ( x73 & ~n19433 ) | ( x73 & n19498 ) | ( ~n19433 & n19498 ) ;
  assign n19500 = ( x74 & ~n19425 ) | ( x74 & n19499 ) | ( ~n19425 & n19499 ) ;
  assign n19501 = n891 | n19500 ;
  assign n19502 = n19425 &  n19501 ;
  assign n19506 = ( n891 & n19425 ) | ( n891 & n19499 ) | ( n19425 & n19499 ) ;
  assign n19507 = ( x74 & ~n19506 ) | ( x74 & n19425 ) | ( ~n19506 & n19425 ) ;
  assign n19508 = ~x74 & n19507 ;
  assign n19509 = n19502 | n19508 ;
  assign n19510 = ~x75 & n19509 ;
  assign n19511 = n19433 &  n19501 ;
  assign n19503 = x73 | n19433 ;
  assign n19504 = x73 &  n19433 ;
  assign n19505 = ( n19503 & ~n19504 ) | ( n19503 & 1'b0 ) | ( ~n19504 & 1'b0 ) ;
  assign n19515 = ( n891 & n19498 ) | ( n891 & n19505 ) | ( n19498 & n19505 ) ;
  assign n19516 = ( n19498 & ~n19500 ) | ( n19498 & n19505 ) | ( ~n19500 & n19505 ) ;
  assign n19517 = ~n19515 & n19516 ;
  assign n19518 = n19511 | n19517 ;
  assign n19519 = n19441 &  n19501 ;
  assign n19512 = x72 | n19441 ;
  assign n19513 = x72 &  n19441 ;
  assign n19514 = ( n19512 & ~n19513 ) | ( n19512 & 1'b0 ) | ( ~n19513 & 1'b0 ) ;
  assign n19523 = ( n891 & n19497 ) | ( n891 & n19514 ) | ( n19497 & n19514 ) ;
  assign n19524 = ( n19497 & ~n19500 ) | ( n19497 & n19514 ) | ( ~n19500 & n19514 ) ;
  assign n19525 = ~n19523 & n19524 ;
  assign n19526 = n19519 | n19525 ;
  assign n19527 = n19449 &  n19501 ;
  assign n19520 = x71 | n19449 ;
  assign n19521 = x71 &  n19449 ;
  assign n19522 = ( n19520 & ~n19521 ) | ( n19520 & 1'b0 ) | ( ~n19521 & 1'b0 ) ;
  assign n19531 = ( n891 & n19496 ) | ( n891 & n19522 ) | ( n19496 & n19522 ) ;
  assign n19532 = ( n19496 & ~n19500 ) | ( n19496 & n19522 ) | ( ~n19500 & n19522 ) ;
  assign n19533 = ~n19531 & n19532 ;
  assign n19534 = n19527 | n19533 ;
  assign n19535 = n19457 &  n19501 ;
  assign n19528 = x70 | n19457 ;
  assign n19529 = x70 &  n19457 ;
  assign n19530 = ( n19528 & ~n19529 ) | ( n19528 & 1'b0 ) | ( ~n19529 & 1'b0 ) ;
  assign n19539 = ( n891 & n19495 ) | ( n891 & n19530 ) | ( n19495 & n19530 ) ;
  assign n19540 = ( n19495 & ~n19500 ) | ( n19495 & n19530 ) | ( ~n19500 & n19530 ) ;
  assign n19541 = ~n19539 & n19540 ;
  assign n19542 = n19535 | n19541 ;
  assign n19543 = n19465 &  n19501 ;
  assign n19536 = x69 | n19465 ;
  assign n19537 = x69 &  n19465 ;
  assign n19538 = ( n19536 & ~n19537 ) | ( n19536 & 1'b0 ) | ( ~n19537 & 1'b0 ) ;
  assign n19547 = ( n891 & n19494 ) | ( n891 & n19538 ) | ( n19494 & n19538 ) ;
  assign n19548 = ( n19494 & ~n19500 ) | ( n19494 & n19538 ) | ( ~n19500 & n19538 ) ;
  assign n19549 = ~n19547 & n19548 ;
  assign n19550 = n19543 | n19549 ;
  assign n19551 = n19473 &  n19501 ;
  assign n19544 = x68 | n19473 ;
  assign n19545 = x68 &  n19473 ;
  assign n19546 = ( n19544 & ~n19545 ) | ( n19544 & 1'b0 ) | ( ~n19545 & 1'b0 ) ;
  assign n19555 = ( n891 & n19493 ) | ( n891 & n19546 ) | ( n19493 & n19546 ) ;
  assign n19556 = ( n19493 & ~n19500 ) | ( n19493 & n19546 ) | ( ~n19500 & n19546 ) ;
  assign n19557 = ~n19555 & n19556 ;
  assign n19558 = n19551 | n19557 ;
  assign n19559 = n19478 &  n19501 ;
  assign n19552 = x67 | n19478 ;
  assign n19553 = x67 &  n19478 ;
  assign n19554 = ( n19552 & ~n19553 ) | ( n19552 & 1'b0 ) | ( ~n19553 & 1'b0 ) ;
  assign n19563 = ( n891 & n19492 ) | ( n891 & n19554 ) | ( n19492 & n19554 ) ;
  assign n19564 = ( n19492 & ~n19500 ) | ( n19492 & n19554 ) | ( ~n19500 & n19554 ) ;
  assign n19565 = ~n19563 & n19564 ;
  assign n19566 = n19559 | n19565 ;
  assign n19567 = n19486 &  n19501 ;
  assign n19560 = x66 | n19486 ;
  assign n19561 = x66 &  n19486 ;
  assign n19562 = ( n19560 & ~n19561 ) | ( n19560 & 1'b0 ) | ( ~n19561 & 1'b0 ) ;
  assign n19571 = ( n891 & n19491 ) | ( n891 & n19562 ) | ( n19491 & n19562 ) ;
  assign n19572 = ( n19491 & ~n19500 ) | ( n19491 & n19562 ) | ( ~n19500 & n19562 ) ;
  assign n19573 = ~n19571 & n19572 ;
  assign n19574 = n19567 | n19573 ;
  assign n19575 = n19490 &  n19501 ;
  assign n19568 = x65 &  n19490 ;
  assign n19569 = x65 | n19489 ;
  assign n19570 = n19488 | n19569 ;
  assign n19576 = ~n19568 & n19570 ;
  assign n19577 = ( n878 & ~n891 ) | ( n878 & n19576 ) | ( ~n891 & n19576 ) ;
  assign n19578 = ( n878 & n19500 ) | ( n878 & n19576 ) | ( n19500 & n19576 ) ;
  assign n19579 = ( n19577 & ~n19578 ) | ( n19577 & 1'b0 ) | ( ~n19578 & 1'b0 ) ;
  assign n19580 = n19575 | n19579 ;
  assign n19581 = ( n946 & ~n19500 ) | ( n946 & 1'b0 ) | ( ~n19500 & 1'b0 ) ;
  assign n19582 = ( x53 & ~n19581 ) | ( x53 & 1'b0 ) | ( ~n19581 & 1'b0 ) ;
  assign n19583 = ( n952 & ~n19500 ) | ( n952 & 1'b0 ) | ( ~n19500 & 1'b0 ) ;
  assign n19584 = n19582 | n19583 ;
  assign n19585 = ( x65 & ~n19584 ) | ( x65 & n955 ) | ( ~n19584 & n955 ) ;
  assign n19586 = ( x66 & ~n19580 ) | ( x66 & n19585 ) | ( ~n19580 & n19585 ) ;
  assign n19587 = ( x67 & ~n19574 ) | ( x67 & n19586 ) | ( ~n19574 & n19586 ) ;
  assign n19588 = ( x68 & ~n19566 ) | ( x68 & n19587 ) | ( ~n19566 & n19587 ) ;
  assign n19589 = ( x69 & ~n19558 ) | ( x69 & n19588 ) | ( ~n19558 & n19588 ) ;
  assign n19590 = ( x70 & ~n19550 ) | ( x70 & n19589 ) | ( ~n19550 & n19589 ) ;
  assign n19591 = ( x71 & ~n19542 ) | ( x71 & n19590 ) | ( ~n19542 & n19590 ) ;
  assign n19592 = ( x72 & ~n19534 ) | ( x72 & n19591 ) | ( ~n19534 & n19591 ) ;
  assign n19593 = ( x73 & ~n19526 ) | ( x73 & n19592 ) | ( ~n19526 & n19592 ) ;
  assign n19594 = ( x74 & ~n19518 ) | ( x74 & n19593 ) | ( ~n19518 & n19593 ) ;
  assign n19595 = ( x75 & ~n19502 ) | ( x75 & 1'b0 ) | ( ~n19502 & 1'b0 ) ;
  assign n19596 = ~n19508 & n19595 ;
  assign n19597 = ( n19594 & ~n19510 ) | ( n19594 & n19596 ) | ( ~n19510 & n19596 ) ;
  assign n19598 = ( n19510 & ~n1000 ) | ( n19510 & n19597 ) | ( ~n1000 & n19597 ) ;
  assign n19599 = n1000 | n19598 ;
  assign n19606 = n891 &  n19425 ;
  assign n19607 = n19599 &  n19606 ;
  assign n19600 = ~n891 & n19509 ;
  assign n19601 = ( n19599 & ~n19600 ) | ( n19599 & 1'b0 ) | ( ~n19600 & 1'b0 ) ;
  assign n19605 = n19510 | n19596 ;
  assign n19609 = ( n19594 & n19601 ) | ( n19594 & n19605 ) | ( n19601 & n19605 ) ;
  assign n19608 = n19594 | n19605 ;
  assign n19610 = ( n19607 & ~n19609 ) | ( n19607 & n19608 ) | ( ~n19609 & n19608 ) ;
  assign n19614 = ( n19518 & ~n19600 ) | ( n19518 & 1'b0 ) | ( ~n19600 & 1'b0 ) ;
  assign n19615 = n19599 &  n19614 ;
  assign n19602 = x74 | n19518 ;
  assign n19603 = x74 &  n19518 ;
  assign n19604 = ( n19602 & ~n19603 ) | ( n19602 & 1'b0 ) | ( ~n19603 & 1'b0 ) ;
  assign n19617 = ( n19593 & n19601 ) | ( n19593 & n19604 ) | ( n19601 & n19604 ) ;
  assign n19616 = n19593 | n19604 ;
  assign n19618 = ( n19615 & ~n19617 ) | ( n19615 & n19616 ) | ( ~n19617 & n19616 ) ;
  assign n19622 = ( n19526 & ~n19600 ) | ( n19526 & 1'b0 ) | ( ~n19600 & 1'b0 ) ;
  assign n19623 = n19599 &  n19622 ;
  assign n19611 = x73 | n19526 ;
  assign n19612 = x73 &  n19526 ;
  assign n19613 = ( n19611 & ~n19612 ) | ( n19611 & 1'b0 ) | ( ~n19612 & 1'b0 ) ;
  assign n19625 = ( n19592 & n19601 ) | ( n19592 & n19613 ) | ( n19601 & n19613 ) ;
  assign n19624 = n19592 | n19613 ;
  assign n19626 = ( n19623 & ~n19625 ) | ( n19623 & n19624 ) | ( ~n19625 & n19624 ) ;
  assign n19630 = ( n19534 & ~n19600 ) | ( n19534 & 1'b0 ) | ( ~n19600 & 1'b0 ) ;
  assign n19631 = n19599 &  n19630 ;
  assign n19619 = x72 | n19534 ;
  assign n19620 = x72 &  n19534 ;
  assign n19621 = ( n19619 & ~n19620 ) | ( n19619 & 1'b0 ) | ( ~n19620 & 1'b0 ) ;
  assign n19633 = ( n19591 & n19601 ) | ( n19591 & n19621 ) | ( n19601 & n19621 ) ;
  assign n19632 = n19591 | n19621 ;
  assign n19634 = ( n19631 & ~n19633 ) | ( n19631 & n19632 ) | ( ~n19633 & n19632 ) ;
  assign n19638 = ( n19542 & ~n19600 ) | ( n19542 & 1'b0 ) | ( ~n19600 & 1'b0 ) ;
  assign n19639 = n19599 &  n19638 ;
  assign n19627 = x71 | n19542 ;
  assign n19628 = x71 &  n19542 ;
  assign n19629 = ( n19627 & ~n19628 ) | ( n19627 & 1'b0 ) | ( ~n19628 & 1'b0 ) ;
  assign n19641 = ( n19590 & n19601 ) | ( n19590 & n19629 ) | ( n19601 & n19629 ) ;
  assign n19640 = n19590 | n19629 ;
  assign n19642 = ( n19639 & ~n19641 ) | ( n19639 & n19640 ) | ( ~n19641 & n19640 ) ;
  assign n19646 = ( n19550 & ~n19600 ) | ( n19550 & 1'b0 ) | ( ~n19600 & 1'b0 ) ;
  assign n19647 = n19599 &  n19646 ;
  assign n19635 = x70 | n19550 ;
  assign n19636 = x70 &  n19550 ;
  assign n19637 = ( n19635 & ~n19636 ) | ( n19635 & 1'b0 ) | ( ~n19636 & 1'b0 ) ;
  assign n19649 = ( n19589 & n19601 ) | ( n19589 & n19637 ) | ( n19601 & n19637 ) ;
  assign n19648 = n19589 | n19637 ;
  assign n19650 = ( n19647 & ~n19649 ) | ( n19647 & n19648 ) | ( ~n19649 & n19648 ) ;
  assign n19654 = ( n19558 & ~n19600 ) | ( n19558 & 1'b0 ) | ( ~n19600 & 1'b0 ) ;
  assign n19655 = n19599 &  n19654 ;
  assign n19643 = x69 | n19558 ;
  assign n19644 = x69 &  n19558 ;
  assign n19645 = ( n19643 & ~n19644 ) | ( n19643 & 1'b0 ) | ( ~n19644 & 1'b0 ) ;
  assign n19657 = ( n19588 & n19601 ) | ( n19588 & n19645 ) | ( n19601 & n19645 ) ;
  assign n19656 = n19588 | n19645 ;
  assign n19658 = ( n19655 & ~n19657 ) | ( n19655 & n19656 ) | ( ~n19657 & n19656 ) ;
  assign n19662 = ( n19566 & ~n19600 ) | ( n19566 & 1'b0 ) | ( ~n19600 & 1'b0 ) ;
  assign n19663 = n19599 &  n19662 ;
  assign n19651 = x68 | n19566 ;
  assign n19652 = x68 &  n19566 ;
  assign n19653 = ( n19651 & ~n19652 ) | ( n19651 & 1'b0 ) | ( ~n19652 & 1'b0 ) ;
  assign n19665 = ( n19587 & n19601 ) | ( n19587 & n19653 ) | ( n19601 & n19653 ) ;
  assign n19664 = n19587 | n19653 ;
  assign n19666 = ( n19663 & ~n19665 ) | ( n19663 & n19664 ) | ( ~n19665 & n19664 ) ;
  assign n19670 = ( n19574 & ~n19600 ) | ( n19574 & 1'b0 ) | ( ~n19600 & 1'b0 ) ;
  assign n19671 = n19599 &  n19670 ;
  assign n19659 = x67 | n19574 ;
  assign n19660 = x67 &  n19574 ;
  assign n19661 = ( n19659 & ~n19660 ) | ( n19659 & 1'b0 ) | ( ~n19660 & 1'b0 ) ;
  assign n19673 = ( n19586 & n19601 ) | ( n19586 & n19661 ) | ( n19601 & n19661 ) ;
  assign n19672 = n19586 | n19661 ;
  assign n19674 = ( n19671 & ~n19673 ) | ( n19671 & n19672 ) | ( ~n19673 & n19672 ) ;
  assign n19675 = ( n19580 & ~n19600 ) | ( n19580 & 1'b0 ) | ( ~n19600 & 1'b0 ) ;
  assign n19676 = n19599 &  n19675 ;
  assign n19667 = x66 | n19580 ;
  assign n19668 = x66 &  n19580 ;
  assign n19669 = ( n19667 & ~n19668 ) | ( n19667 & 1'b0 ) | ( ~n19668 & 1'b0 ) ;
  assign n19678 = ( n19585 & n19601 ) | ( n19585 & n19669 ) | ( n19601 & n19669 ) ;
  assign n19677 = n19585 | n19669 ;
  assign n19679 = ( n19676 & ~n19678 ) | ( n19676 & n19677 ) | ( ~n19678 & n19677 ) ;
  assign n19680 = ( x65 & ~n955 ) | ( x65 & n19584 ) | ( ~n955 & n19584 ) ;
  assign n19681 = ( n19585 & ~x65 ) | ( n19585 & n19680 ) | ( ~x65 & n19680 ) ;
  assign n19682 = ~n19601 & n19681 ;
  assign n19683 = ( n19584 & ~n19600 ) | ( n19584 & 1'b0 ) | ( ~n19600 & 1'b0 ) ;
  assign n19684 = n19599 &  n19683 ;
  assign n19685 = n19682 | n19684 ;
  assign n19686 = ( x64 & ~n19601 ) | ( x64 & 1'b0 ) | ( ~n19601 & 1'b0 ) ;
  assign n19687 = ( x52 & ~n19686 ) | ( x52 & 1'b0 ) | ( ~n19686 & 1'b0 ) ;
  assign n19688 = ( n955 & ~n19601 ) | ( n955 & 1'b0 ) | ( ~n19601 & 1'b0 ) ;
  assign n19689 = n19687 | n19688 ;
  assign n19690 = ( x65 & ~n19689 ) | ( x65 & n1090 ) | ( ~n19689 & n1090 ) ;
  assign n19691 = ( x66 & ~n19685 ) | ( x66 & n19690 ) | ( ~n19685 & n19690 ) ;
  assign n19692 = ( x67 & ~n19679 ) | ( x67 & n19691 ) | ( ~n19679 & n19691 ) ;
  assign n19693 = ( x68 & ~n19674 ) | ( x68 & n19692 ) | ( ~n19674 & n19692 ) ;
  assign n19694 = ( x69 & ~n19666 ) | ( x69 & n19693 ) | ( ~n19666 & n19693 ) ;
  assign n19695 = ( x70 & ~n19658 ) | ( x70 & n19694 ) | ( ~n19658 & n19694 ) ;
  assign n19696 = ( x71 & ~n19650 ) | ( x71 & n19695 ) | ( ~n19650 & n19695 ) ;
  assign n19697 = ( x72 & ~n19642 ) | ( x72 & n19696 ) | ( ~n19642 & n19696 ) ;
  assign n19698 = ( x73 & ~n19634 ) | ( x73 & n19697 ) | ( ~n19634 & n19697 ) ;
  assign n19699 = ( x74 & ~n19626 ) | ( x74 & n19698 ) | ( ~n19626 & n19698 ) ;
  assign n19700 = ( x75 & ~n19618 ) | ( x75 & n19699 ) | ( ~n19618 & n19699 ) ;
  assign n19707 = ( x76 & ~n1104 ) | ( x76 & n19700 ) | ( ~n1104 & n19700 ) ;
  assign n19706 = x76 &  n19700 ;
  assign n19708 = ( n19610 & ~n19707 ) | ( n19610 & n19706 ) | ( ~n19707 & n19706 ) ;
  assign n19701 = ( x76 & ~n19610 ) | ( x76 & n19700 ) | ( ~n19610 & n19700 ) ;
  assign n19702 = n1104 | n19701 ;
  assign n19709 = n19618 &  n19702 ;
  assign n19703 = x75 | n19618 ;
  assign n19704 = x75 &  n19618 ;
  assign n19705 = ( n19703 & ~n19704 ) | ( n19703 & 1'b0 ) | ( ~n19704 & 1'b0 ) ;
  assign n19713 = ( n1104 & n19699 ) | ( n1104 & n19705 ) | ( n19699 & n19705 ) ;
  assign n19714 = ( n19699 & ~n19701 ) | ( n19699 & n19705 ) | ( ~n19701 & n19705 ) ;
  assign n19715 = ~n19713 & n19714 ;
  assign n19716 = n19709 | n19715 ;
  assign n19717 = n19626 &  n19702 ;
  assign n19710 = x74 | n19626 ;
  assign n19711 = x74 &  n19626 ;
  assign n19712 = ( n19710 & ~n19711 ) | ( n19710 & 1'b0 ) | ( ~n19711 & 1'b0 ) ;
  assign n19721 = ( n1104 & n19698 ) | ( n1104 & n19712 ) | ( n19698 & n19712 ) ;
  assign n19722 = ( n19698 & ~n19701 ) | ( n19698 & n19712 ) | ( ~n19701 & n19712 ) ;
  assign n19723 = ~n19721 & n19722 ;
  assign n19724 = n19717 | n19723 ;
  assign n19725 = n19634 &  n19702 ;
  assign n19718 = x73 | n19634 ;
  assign n19719 = x73 &  n19634 ;
  assign n19720 = ( n19718 & ~n19719 ) | ( n19718 & 1'b0 ) | ( ~n19719 & 1'b0 ) ;
  assign n19729 = ( n1104 & n19697 ) | ( n1104 & n19720 ) | ( n19697 & n19720 ) ;
  assign n19730 = ( n19697 & ~n19701 ) | ( n19697 & n19720 ) | ( ~n19701 & n19720 ) ;
  assign n19731 = ~n19729 & n19730 ;
  assign n19732 = n19725 | n19731 ;
  assign n19733 = n19642 &  n19702 ;
  assign n19726 = x72 | n19642 ;
  assign n19727 = x72 &  n19642 ;
  assign n19728 = ( n19726 & ~n19727 ) | ( n19726 & 1'b0 ) | ( ~n19727 & 1'b0 ) ;
  assign n19737 = ( n1104 & n19696 ) | ( n1104 & n19728 ) | ( n19696 & n19728 ) ;
  assign n19738 = ( n19696 & ~n19701 ) | ( n19696 & n19728 ) | ( ~n19701 & n19728 ) ;
  assign n19739 = ~n19737 & n19738 ;
  assign n19740 = n19733 | n19739 ;
  assign n19741 = n19650 &  n19702 ;
  assign n19734 = x71 | n19650 ;
  assign n19735 = x71 &  n19650 ;
  assign n19736 = ( n19734 & ~n19735 ) | ( n19734 & 1'b0 ) | ( ~n19735 & 1'b0 ) ;
  assign n19745 = ( n1104 & n19695 ) | ( n1104 & n19736 ) | ( n19695 & n19736 ) ;
  assign n19746 = ( n19695 & ~n19701 ) | ( n19695 & n19736 ) | ( ~n19701 & n19736 ) ;
  assign n19747 = ~n19745 & n19746 ;
  assign n19748 = n19741 | n19747 ;
  assign n19749 = n19658 &  n19702 ;
  assign n19742 = x70 | n19658 ;
  assign n19743 = x70 &  n19658 ;
  assign n19744 = ( n19742 & ~n19743 ) | ( n19742 & 1'b0 ) | ( ~n19743 & 1'b0 ) ;
  assign n19753 = ( n1104 & n19694 ) | ( n1104 & n19744 ) | ( n19694 & n19744 ) ;
  assign n19754 = ( n19694 & ~n19701 ) | ( n19694 & n19744 ) | ( ~n19701 & n19744 ) ;
  assign n19755 = ~n19753 & n19754 ;
  assign n19756 = n19749 | n19755 ;
  assign n19757 = n19666 &  n19702 ;
  assign n19750 = x69 | n19666 ;
  assign n19751 = x69 &  n19666 ;
  assign n19752 = ( n19750 & ~n19751 ) | ( n19750 & 1'b0 ) | ( ~n19751 & 1'b0 ) ;
  assign n19761 = ( n1104 & n19693 ) | ( n1104 & n19752 ) | ( n19693 & n19752 ) ;
  assign n19762 = ( n19693 & ~n19701 ) | ( n19693 & n19752 ) | ( ~n19701 & n19752 ) ;
  assign n19763 = ~n19761 & n19762 ;
  assign n19764 = n19757 | n19763 ;
  assign n19765 = n19674 &  n19702 ;
  assign n19758 = x68 | n19674 ;
  assign n19759 = x68 &  n19674 ;
  assign n19760 = ( n19758 & ~n19759 ) | ( n19758 & 1'b0 ) | ( ~n19759 & 1'b0 ) ;
  assign n19769 = ( n1104 & n19692 ) | ( n1104 & n19760 ) | ( n19692 & n19760 ) ;
  assign n19770 = ( n19692 & ~n19701 ) | ( n19692 & n19760 ) | ( ~n19701 & n19760 ) ;
  assign n19771 = ~n19769 & n19770 ;
  assign n19772 = n19765 | n19771 ;
  assign n19773 = n19679 &  n19702 ;
  assign n19766 = x67 | n19679 ;
  assign n19767 = x67 &  n19679 ;
  assign n19768 = ( n19766 & ~n19767 ) | ( n19766 & 1'b0 ) | ( ~n19767 & 1'b0 ) ;
  assign n19777 = ( n1104 & n19691 ) | ( n1104 & n19768 ) | ( n19691 & n19768 ) ;
  assign n19778 = ( n19691 & ~n19701 ) | ( n19691 & n19768 ) | ( ~n19701 & n19768 ) ;
  assign n19779 = ~n19777 & n19778 ;
  assign n19780 = n19773 | n19779 ;
  assign n19781 = n19685 &  n19702 ;
  assign n19774 = x66 | n19685 ;
  assign n19775 = x66 &  n19685 ;
  assign n19776 = ( n19774 & ~n19775 ) | ( n19774 & 1'b0 ) | ( ~n19775 & 1'b0 ) ;
  assign n19782 = ( n1104 & n19690 ) | ( n1104 & n19776 ) | ( n19690 & n19776 ) ;
  assign n19783 = ( n19690 & ~n19701 ) | ( n19690 & n19776 ) | ( ~n19701 & n19776 ) ;
  assign n19784 = ~n19782 & n19783 ;
  assign n19785 = n19781 | n19784 ;
  assign n19786 = n19689 &  n19702 ;
  assign n19787 = ( x65 & ~x52 ) | ( x65 & n19686 ) | ( ~x52 & n19686 ) ;
  assign n19788 = ( x52 & ~n19686 ) | ( x52 & x65 ) | ( ~n19686 & x65 ) ;
  assign n19789 = ( n19787 & ~x65 ) | ( n19787 & n19788 ) | ( ~x65 & n19788 ) ;
  assign n19790 = ( n1090 & ~n1104 ) | ( n1090 & n19789 ) | ( ~n1104 & n19789 ) ;
  assign n19791 = ( n1090 & n19701 ) | ( n1090 & n19789 ) | ( n19701 & n19789 ) ;
  assign n19792 = ( n19790 & ~n19791 ) | ( n19790 & 1'b0 ) | ( ~n19791 & 1'b0 ) ;
  assign n19793 = n19786 | n19792 ;
  assign n19794 = ( n1203 & ~n19701 ) | ( n1203 & 1'b0 ) | ( ~n19701 & 1'b0 ) ;
  assign n19795 = ( x51 & ~n19794 ) | ( x51 & 1'b0 ) | ( ~n19794 & 1'b0 ) ;
  assign n19796 = ( n1208 & ~n19701 ) | ( n1208 & 1'b0 ) | ( ~n19701 & 1'b0 ) ;
  assign n19797 = n19795 | n19796 ;
  assign n19798 = ( x65 & ~n19797 ) | ( x65 & n1211 ) | ( ~n19797 & n1211 ) ;
  assign n19799 = ( x66 & ~n19793 ) | ( x66 & n19798 ) | ( ~n19793 & n19798 ) ;
  assign n19800 = ( x67 & ~n19785 ) | ( x67 & n19799 ) | ( ~n19785 & n19799 ) ;
  assign n19801 = ( x68 & ~n19780 ) | ( x68 & n19800 ) | ( ~n19780 & n19800 ) ;
  assign n19802 = ( x69 & ~n19772 ) | ( x69 & n19801 ) | ( ~n19772 & n19801 ) ;
  assign n19803 = ( x70 & ~n19764 ) | ( x70 & n19802 ) | ( ~n19764 & n19802 ) ;
  assign n19804 = ( x71 & ~n19756 ) | ( x71 & n19803 ) | ( ~n19756 & n19803 ) ;
  assign n19805 = ( x72 & ~n19748 ) | ( x72 & n19804 ) | ( ~n19748 & n19804 ) ;
  assign n19806 = ( x73 & ~n19740 ) | ( x73 & n19805 ) | ( ~n19740 & n19805 ) ;
  assign n19807 = ( x74 & ~n19732 ) | ( x74 & n19806 ) | ( ~n19732 & n19806 ) ;
  assign n19808 = ( x75 & ~n19724 ) | ( x75 & n19807 ) | ( ~n19724 & n19807 ) ;
  assign n19809 = ( x76 & ~n19716 ) | ( x76 & n19808 ) | ( ~n19716 & n19808 ) ;
  assign n19810 = ( x77 & ~n19708 ) | ( x77 & n19809 ) | ( ~n19708 & n19809 ) ;
  assign n19811 = n1227 | n19810 ;
  assign n19812 = n19708 &  n19811 ;
  assign n19816 = ( n1227 & n19708 ) | ( n1227 & n19809 ) | ( n19708 & n19809 ) ;
  assign n19817 = ( x77 & ~n19816 ) | ( x77 & n19708 ) | ( ~n19816 & n19708 ) ;
  assign n19818 = ~x77 & n19817 ;
  assign n19819 = n19812 | n19818 ;
  assign n19820 = ~x78 & n19819 ;
  assign n19821 = n19716 &  n19811 ;
  assign n19813 = x76 | n19716 ;
  assign n19814 = x76 &  n19716 ;
  assign n19815 = ( n19813 & ~n19814 ) | ( n19813 & 1'b0 ) | ( ~n19814 & 1'b0 ) ;
  assign n19825 = ( n1227 & n19808 ) | ( n1227 & n19815 ) | ( n19808 & n19815 ) ;
  assign n19826 = ( n19808 & ~n19810 ) | ( n19808 & n19815 ) | ( ~n19810 & n19815 ) ;
  assign n19827 = ~n19825 & n19826 ;
  assign n19828 = n19821 | n19827 ;
  assign n19829 = n19724 &  n19811 ;
  assign n19822 = x75 | n19724 ;
  assign n19823 = x75 &  n19724 ;
  assign n19824 = ( n19822 & ~n19823 ) | ( n19822 & 1'b0 ) | ( ~n19823 & 1'b0 ) ;
  assign n19833 = ( n1227 & n19807 ) | ( n1227 & n19824 ) | ( n19807 & n19824 ) ;
  assign n19834 = ( n19807 & ~n19810 ) | ( n19807 & n19824 ) | ( ~n19810 & n19824 ) ;
  assign n19835 = ~n19833 & n19834 ;
  assign n19836 = n19829 | n19835 ;
  assign n19837 = n19732 &  n19811 ;
  assign n19830 = x74 | n19732 ;
  assign n19831 = x74 &  n19732 ;
  assign n19832 = ( n19830 & ~n19831 ) | ( n19830 & 1'b0 ) | ( ~n19831 & 1'b0 ) ;
  assign n19841 = ( n1227 & n19806 ) | ( n1227 & n19832 ) | ( n19806 & n19832 ) ;
  assign n19842 = ( n19806 & ~n19810 ) | ( n19806 & n19832 ) | ( ~n19810 & n19832 ) ;
  assign n19843 = ~n19841 & n19842 ;
  assign n19844 = n19837 | n19843 ;
  assign n19845 = n19740 &  n19811 ;
  assign n19838 = x73 | n19740 ;
  assign n19839 = x73 &  n19740 ;
  assign n19840 = ( n19838 & ~n19839 ) | ( n19838 & 1'b0 ) | ( ~n19839 & 1'b0 ) ;
  assign n19849 = ( n1227 & n19805 ) | ( n1227 & n19840 ) | ( n19805 & n19840 ) ;
  assign n19850 = ( n19805 & ~n19810 ) | ( n19805 & n19840 ) | ( ~n19810 & n19840 ) ;
  assign n19851 = ~n19849 & n19850 ;
  assign n19852 = n19845 | n19851 ;
  assign n19853 = n19748 &  n19811 ;
  assign n19846 = x72 | n19748 ;
  assign n19847 = x72 &  n19748 ;
  assign n19848 = ( n19846 & ~n19847 ) | ( n19846 & 1'b0 ) | ( ~n19847 & 1'b0 ) ;
  assign n19857 = ( n1227 & n19804 ) | ( n1227 & n19848 ) | ( n19804 & n19848 ) ;
  assign n19858 = ( n19804 & ~n19810 ) | ( n19804 & n19848 ) | ( ~n19810 & n19848 ) ;
  assign n19859 = ~n19857 & n19858 ;
  assign n19860 = n19853 | n19859 ;
  assign n19861 = n19756 &  n19811 ;
  assign n19854 = x71 | n19756 ;
  assign n19855 = x71 &  n19756 ;
  assign n19856 = ( n19854 & ~n19855 ) | ( n19854 & 1'b0 ) | ( ~n19855 & 1'b0 ) ;
  assign n19865 = ( n1227 & n19803 ) | ( n1227 & n19856 ) | ( n19803 & n19856 ) ;
  assign n19866 = ( n19803 & ~n19810 ) | ( n19803 & n19856 ) | ( ~n19810 & n19856 ) ;
  assign n19867 = ~n19865 & n19866 ;
  assign n19868 = n19861 | n19867 ;
  assign n19869 = n19764 &  n19811 ;
  assign n19862 = x70 | n19764 ;
  assign n19863 = x70 &  n19764 ;
  assign n19864 = ( n19862 & ~n19863 ) | ( n19862 & 1'b0 ) | ( ~n19863 & 1'b0 ) ;
  assign n19873 = ( n1227 & n19802 ) | ( n1227 & n19864 ) | ( n19802 & n19864 ) ;
  assign n19874 = ( n19802 & ~n19810 ) | ( n19802 & n19864 ) | ( ~n19810 & n19864 ) ;
  assign n19875 = ~n19873 & n19874 ;
  assign n19876 = n19869 | n19875 ;
  assign n19877 = n19772 &  n19811 ;
  assign n19870 = x69 | n19772 ;
  assign n19871 = x69 &  n19772 ;
  assign n19872 = ( n19870 & ~n19871 ) | ( n19870 & 1'b0 ) | ( ~n19871 & 1'b0 ) ;
  assign n19881 = ( n1227 & n19801 ) | ( n1227 & n19872 ) | ( n19801 & n19872 ) ;
  assign n19882 = ( n19801 & ~n19810 ) | ( n19801 & n19872 ) | ( ~n19810 & n19872 ) ;
  assign n19883 = ~n19881 & n19882 ;
  assign n19884 = n19877 | n19883 ;
  assign n19885 = n19780 &  n19811 ;
  assign n19878 = x68 | n19780 ;
  assign n19879 = x68 &  n19780 ;
  assign n19880 = ( n19878 & ~n19879 ) | ( n19878 & 1'b0 ) | ( ~n19879 & 1'b0 ) ;
  assign n19889 = ( n1227 & n19800 ) | ( n1227 & n19880 ) | ( n19800 & n19880 ) ;
  assign n19890 = ( n19800 & ~n19810 ) | ( n19800 & n19880 ) | ( ~n19810 & n19880 ) ;
  assign n19891 = ~n19889 & n19890 ;
  assign n19892 = n19885 | n19891 ;
  assign n19893 = n19785 &  n19811 ;
  assign n19886 = x67 | n19785 ;
  assign n19887 = x67 &  n19785 ;
  assign n19888 = ( n19886 & ~n19887 ) | ( n19886 & 1'b0 ) | ( ~n19887 & 1'b0 ) ;
  assign n19897 = ( n1227 & n19799 ) | ( n1227 & n19888 ) | ( n19799 & n19888 ) ;
  assign n19898 = ( n19799 & ~n19810 ) | ( n19799 & n19888 ) | ( ~n19810 & n19888 ) ;
  assign n19899 = ~n19897 & n19898 ;
  assign n19900 = n19893 | n19899 ;
  assign n19901 = n19793 &  n19811 ;
  assign n19894 = x66 | n19793 ;
  assign n19895 = x66 &  n19793 ;
  assign n19896 = ( n19894 & ~n19895 ) | ( n19894 & 1'b0 ) | ( ~n19895 & 1'b0 ) ;
  assign n19905 = ( n1227 & n19798 ) | ( n1227 & n19896 ) | ( n19798 & n19896 ) ;
  assign n19906 = ( n19798 & ~n19810 ) | ( n19798 & n19896 ) | ( ~n19810 & n19896 ) ;
  assign n19907 = ~n19905 & n19906 ;
  assign n19908 = n19901 | n19907 ;
  assign n19909 = n19797 &  n19811 ;
  assign n19902 = x65 &  n19797 ;
  assign n19903 = x65 | n19796 ;
  assign n19904 = n19795 | n19903 ;
  assign n19910 = ~n19902 & n19904 ;
  assign n19911 = ( n1211 & ~n1227 ) | ( n1211 & n19910 ) | ( ~n1227 & n19910 ) ;
  assign n19912 = ( n1211 & n19810 ) | ( n1211 & n19910 ) | ( n19810 & n19910 ) ;
  assign n19913 = ( n19911 & ~n19912 ) | ( n19911 & 1'b0 ) | ( ~n19912 & 1'b0 ) ;
  assign n19914 = n19909 | n19913 ;
  assign n19915 = ( n1315 & ~n19810 ) | ( n1315 & 1'b0 ) | ( ~n19810 & 1'b0 ) ;
  assign n19916 = ( x50 & ~n19915 ) | ( x50 & 1'b0 ) | ( ~n19915 & 1'b0 ) ;
  assign n19917 = ( n1321 & ~n19810 ) | ( n1321 & 1'b0 ) | ( ~n19810 & 1'b0 ) ;
  assign n19918 = n19916 | n19917 ;
  assign n19919 = ( x65 & ~n19918 ) | ( x65 & n1324 ) | ( ~n19918 & n1324 ) ;
  assign n19920 = ( x66 & ~n19914 ) | ( x66 & n19919 ) | ( ~n19914 & n19919 ) ;
  assign n19921 = ( x67 & ~n19908 ) | ( x67 & n19920 ) | ( ~n19908 & n19920 ) ;
  assign n19922 = ( x68 & ~n19900 ) | ( x68 & n19921 ) | ( ~n19900 & n19921 ) ;
  assign n19923 = ( x69 & ~n19892 ) | ( x69 & n19922 ) | ( ~n19892 & n19922 ) ;
  assign n19924 = ( x70 & ~n19884 ) | ( x70 & n19923 ) | ( ~n19884 & n19923 ) ;
  assign n19925 = ( x71 & ~n19876 ) | ( x71 & n19924 ) | ( ~n19876 & n19924 ) ;
  assign n19926 = ( x72 & ~n19868 ) | ( x72 & n19925 ) | ( ~n19868 & n19925 ) ;
  assign n19927 = ( x73 & ~n19860 ) | ( x73 & n19926 ) | ( ~n19860 & n19926 ) ;
  assign n19928 = ( x74 & ~n19852 ) | ( x74 & n19927 ) | ( ~n19852 & n19927 ) ;
  assign n19929 = ( x75 & ~n19844 ) | ( x75 & n19928 ) | ( ~n19844 & n19928 ) ;
  assign n19930 = ( x76 & ~n19836 ) | ( x76 & n19929 ) | ( ~n19836 & n19929 ) ;
  assign n19931 = ( x77 & ~n19828 ) | ( x77 & n19930 ) | ( ~n19828 & n19930 ) ;
  assign n19932 = ( x78 & ~n19812 ) | ( x78 & 1'b0 ) | ( ~n19812 & 1'b0 ) ;
  assign n19933 = ~n19818 & n19932 ;
  assign n19934 = ( n19931 & ~n19820 ) | ( n19931 & n19933 ) | ( ~n19820 & n19933 ) ;
  assign n19935 = ( n19820 & ~n1365 ) | ( n19820 & n19934 ) | ( ~n1365 & n19934 ) ;
  assign n19936 = n1365 | n19935 ;
  assign n19943 = n1227 &  n19708 ;
  assign n19944 = n19936 &  n19943 ;
  assign n19937 = ~n1227 & n19819 ;
  assign n19938 = ( n19936 & ~n19937 ) | ( n19936 & 1'b0 ) | ( ~n19937 & 1'b0 ) ;
  assign n19942 = n19820 | n19933 ;
  assign n19946 = ( n19931 & n19938 ) | ( n19931 & n19942 ) | ( n19938 & n19942 ) ;
  assign n19945 = n19931 | n19942 ;
  assign n19947 = ( n19944 & ~n19946 ) | ( n19944 & n19945 ) | ( ~n19946 & n19945 ) ;
  assign n19951 = ( n19828 & ~n19937 ) | ( n19828 & 1'b0 ) | ( ~n19937 & 1'b0 ) ;
  assign n19952 = n19936 &  n19951 ;
  assign n19939 = x77 | n19828 ;
  assign n19940 = x77 &  n19828 ;
  assign n19941 = ( n19939 & ~n19940 ) | ( n19939 & 1'b0 ) | ( ~n19940 & 1'b0 ) ;
  assign n19954 = ( n19930 & n19938 ) | ( n19930 & n19941 ) | ( n19938 & n19941 ) ;
  assign n19953 = n19930 | n19941 ;
  assign n19955 = ( n19952 & ~n19954 ) | ( n19952 & n19953 ) | ( ~n19954 & n19953 ) ;
  assign n19959 = ( n19836 & ~n19937 ) | ( n19836 & 1'b0 ) | ( ~n19937 & 1'b0 ) ;
  assign n19960 = n19936 &  n19959 ;
  assign n19948 = x76 | n19836 ;
  assign n19949 = x76 &  n19836 ;
  assign n19950 = ( n19948 & ~n19949 ) | ( n19948 & 1'b0 ) | ( ~n19949 & 1'b0 ) ;
  assign n19962 = ( n19929 & n19938 ) | ( n19929 & n19950 ) | ( n19938 & n19950 ) ;
  assign n19961 = n19929 | n19950 ;
  assign n19963 = ( n19960 & ~n19962 ) | ( n19960 & n19961 ) | ( ~n19962 & n19961 ) ;
  assign n19967 = ( n19844 & ~n19937 ) | ( n19844 & 1'b0 ) | ( ~n19937 & 1'b0 ) ;
  assign n19968 = n19936 &  n19967 ;
  assign n19956 = x75 | n19844 ;
  assign n19957 = x75 &  n19844 ;
  assign n19958 = ( n19956 & ~n19957 ) | ( n19956 & 1'b0 ) | ( ~n19957 & 1'b0 ) ;
  assign n19970 = ( n19928 & n19938 ) | ( n19928 & n19958 ) | ( n19938 & n19958 ) ;
  assign n19969 = n19928 | n19958 ;
  assign n19971 = ( n19968 & ~n19970 ) | ( n19968 & n19969 ) | ( ~n19970 & n19969 ) ;
  assign n19975 = ( n19852 & ~n19937 ) | ( n19852 & 1'b0 ) | ( ~n19937 & 1'b0 ) ;
  assign n19976 = n19936 &  n19975 ;
  assign n19964 = x74 | n19852 ;
  assign n19965 = x74 &  n19852 ;
  assign n19966 = ( n19964 & ~n19965 ) | ( n19964 & 1'b0 ) | ( ~n19965 & 1'b0 ) ;
  assign n19978 = ( n19927 & n19938 ) | ( n19927 & n19966 ) | ( n19938 & n19966 ) ;
  assign n19977 = n19927 | n19966 ;
  assign n19979 = ( n19976 & ~n19978 ) | ( n19976 & n19977 ) | ( ~n19978 & n19977 ) ;
  assign n19983 = ( n19860 & ~n19937 ) | ( n19860 & 1'b0 ) | ( ~n19937 & 1'b0 ) ;
  assign n19984 = n19936 &  n19983 ;
  assign n19972 = x73 | n19860 ;
  assign n19973 = x73 &  n19860 ;
  assign n19974 = ( n19972 & ~n19973 ) | ( n19972 & 1'b0 ) | ( ~n19973 & 1'b0 ) ;
  assign n19986 = ( n19926 & n19938 ) | ( n19926 & n19974 ) | ( n19938 & n19974 ) ;
  assign n19985 = n19926 | n19974 ;
  assign n19987 = ( n19984 & ~n19986 ) | ( n19984 & n19985 ) | ( ~n19986 & n19985 ) ;
  assign n19991 = ( n19868 & ~n19937 ) | ( n19868 & 1'b0 ) | ( ~n19937 & 1'b0 ) ;
  assign n19992 = n19936 &  n19991 ;
  assign n19980 = x72 | n19868 ;
  assign n19981 = x72 &  n19868 ;
  assign n19982 = ( n19980 & ~n19981 ) | ( n19980 & 1'b0 ) | ( ~n19981 & 1'b0 ) ;
  assign n19994 = ( n19925 & n19938 ) | ( n19925 & n19982 ) | ( n19938 & n19982 ) ;
  assign n19993 = n19925 | n19982 ;
  assign n19995 = ( n19992 & ~n19994 ) | ( n19992 & n19993 ) | ( ~n19994 & n19993 ) ;
  assign n19999 = ( n19876 & ~n19937 ) | ( n19876 & 1'b0 ) | ( ~n19937 & 1'b0 ) ;
  assign n20000 = n19936 &  n19999 ;
  assign n19988 = x71 | n19876 ;
  assign n19989 = x71 &  n19876 ;
  assign n19990 = ( n19988 & ~n19989 ) | ( n19988 & 1'b0 ) | ( ~n19989 & 1'b0 ) ;
  assign n20002 = ( n19924 & n19938 ) | ( n19924 & n19990 ) | ( n19938 & n19990 ) ;
  assign n20001 = n19924 | n19990 ;
  assign n20003 = ( n20000 & ~n20002 ) | ( n20000 & n20001 ) | ( ~n20002 & n20001 ) ;
  assign n20007 = ( n19884 & ~n19937 ) | ( n19884 & 1'b0 ) | ( ~n19937 & 1'b0 ) ;
  assign n20008 = n19936 &  n20007 ;
  assign n19996 = x70 | n19884 ;
  assign n19997 = x70 &  n19884 ;
  assign n19998 = ( n19996 & ~n19997 ) | ( n19996 & 1'b0 ) | ( ~n19997 & 1'b0 ) ;
  assign n20010 = ( n19923 & n19938 ) | ( n19923 & n19998 ) | ( n19938 & n19998 ) ;
  assign n20009 = n19923 | n19998 ;
  assign n20011 = ( n20008 & ~n20010 ) | ( n20008 & n20009 ) | ( ~n20010 & n20009 ) ;
  assign n20015 = ( n19892 & ~n19937 ) | ( n19892 & 1'b0 ) | ( ~n19937 & 1'b0 ) ;
  assign n20016 = n19936 &  n20015 ;
  assign n20004 = x69 | n19892 ;
  assign n20005 = x69 &  n19892 ;
  assign n20006 = ( n20004 & ~n20005 ) | ( n20004 & 1'b0 ) | ( ~n20005 & 1'b0 ) ;
  assign n20018 = ( n19922 & n19938 ) | ( n19922 & n20006 ) | ( n19938 & n20006 ) ;
  assign n20017 = n19922 | n20006 ;
  assign n20019 = ( n20016 & ~n20018 ) | ( n20016 & n20017 ) | ( ~n20018 & n20017 ) ;
  assign n20023 = ( n19900 & ~n19937 ) | ( n19900 & 1'b0 ) | ( ~n19937 & 1'b0 ) ;
  assign n20024 = n19936 &  n20023 ;
  assign n20012 = x68 | n19900 ;
  assign n20013 = x68 &  n19900 ;
  assign n20014 = ( n20012 & ~n20013 ) | ( n20012 & 1'b0 ) | ( ~n20013 & 1'b0 ) ;
  assign n20026 = ( n19921 & n19938 ) | ( n19921 & n20014 ) | ( n19938 & n20014 ) ;
  assign n20025 = n19921 | n20014 ;
  assign n20027 = ( n20024 & ~n20026 ) | ( n20024 & n20025 ) | ( ~n20026 & n20025 ) ;
  assign n20031 = ( n19908 & ~n19937 ) | ( n19908 & 1'b0 ) | ( ~n19937 & 1'b0 ) ;
  assign n20032 = n19936 &  n20031 ;
  assign n20020 = x67 | n19908 ;
  assign n20021 = x67 &  n19908 ;
  assign n20022 = ( n20020 & ~n20021 ) | ( n20020 & 1'b0 ) | ( ~n20021 & 1'b0 ) ;
  assign n20034 = ( n19920 & n19938 ) | ( n19920 & n20022 ) | ( n19938 & n20022 ) ;
  assign n20033 = n19920 | n20022 ;
  assign n20035 = ( n20032 & ~n20034 ) | ( n20032 & n20033 ) | ( ~n20034 & n20033 ) ;
  assign n20036 = ( n19914 & ~n19937 ) | ( n19914 & 1'b0 ) | ( ~n19937 & 1'b0 ) ;
  assign n20037 = n19936 &  n20036 ;
  assign n20028 = x66 | n19914 ;
  assign n20029 = x66 &  n19914 ;
  assign n20030 = ( n20028 & ~n20029 ) | ( n20028 & 1'b0 ) | ( ~n20029 & 1'b0 ) ;
  assign n20039 = ( n19919 & n19938 ) | ( n19919 & n20030 ) | ( n19938 & n20030 ) ;
  assign n20038 = n19919 | n20030 ;
  assign n20040 = ( n20037 & ~n20039 ) | ( n20037 & n20038 ) | ( ~n20039 & n20038 ) ;
  assign n20041 = ( x65 & ~n1324 ) | ( x65 & n19918 ) | ( ~n1324 & n19918 ) ;
  assign n20042 = ( n19919 & ~x65 ) | ( n19919 & n20041 ) | ( ~x65 & n20041 ) ;
  assign n20043 = ~n19938 & n20042 ;
  assign n20044 = ( n19918 & ~n19937 ) | ( n19918 & 1'b0 ) | ( ~n19937 & 1'b0 ) ;
  assign n20045 = n19936 &  n20044 ;
  assign n20046 = n20043 | n20045 ;
  assign n20047 = ( x64 & ~n19938 ) | ( x64 & 1'b0 ) | ( ~n19938 & 1'b0 ) ;
  assign n20048 = ( x49 & ~n20047 ) | ( x49 & 1'b0 ) | ( ~n20047 & 1'b0 ) ;
  assign n20049 = ( n1324 & ~n19938 ) | ( n1324 & 1'b0 ) | ( ~n19938 & 1'b0 ) ;
  assign n20050 = n20048 | n20049 ;
  assign n20051 = ( x65 & ~n20050 ) | ( x65 & n1479 ) | ( ~n20050 & n1479 ) ;
  assign n20052 = ( x66 & ~n20046 ) | ( x66 & n20051 ) | ( ~n20046 & n20051 ) ;
  assign n20053 = ( x67 & ~n20040 ) | ( x67 & n20052 ) | ( ~n20040 & n20052 ) ;
  assign n20054 = ( x68 & ~n20035 ) | ( x68 & n20053 ) | ( ~n20035 & n20053 ) ;
  assign n20055 = ( x69 & ~n20027 ) | ( x69 & n20054 ) | ( ~n20027 & n20054 ) ;
  assign n20056 = ( x70 & ~n20019 ) | ( x70 & n20055 ) | ( ~n20019 & n20055 ) ;
  assign n20057 = ( x71 & ~n20011 ) | ( x71 & n20056 ) | ( ~n20011 & n20056 ) ;
  assign n20058 = ( x72 & ~n20003 ) | ( x72 & n20057 ) | ( ~n20003 & n20057 ) ;
  assign n20059 = ( x73 & ~n19995 ) | ( x73 & n20058 ) | ( ~n19995 & n20058 ) ;
  assign n20060 = ( x74 & ~n19987 ) | ( x74 & n20059 ) | ( ~n19987 & n20059 ) ;
  assign n20061 = ( x75 & ~n19979 ) | ( x75 & n20060 ) | ( ~n19979 & n20060 ) ;
  assign n20062 = ( x76 & ~n19971 ) | ( x76 & n20061 ) | ( ~n19971 & n20061 ) ;
  assign n20063 = ( x77 & ~n19963 ) | ( x77 & n20062 ) | ( ~n19963 & n20062 ) ;
  assign n20064 = ( x78 & ~n19955 ) | ( x78 & n20063 ) | ( ~n19955 & n20063 ) ;
  assign n20071 = ( x79 & ~n282 ) | ( x79 & n20064 ) | ( ~n282 & n20064 ) ;
  assign n20070 = x79 &  n20064 ;
  assign n20072 = ( n19947 & ~n20071 ) | ( n19947 & n20070 ) | ( ~n20071 & n20070 ) ;
  assign n20065 = ( x79 & ~n19947 ) | ( x79 & n20064 ) | ( ~n19947 & n20064 ) ;
  assign n20066 = n282 | n20065 ;
  assign n20073 = n19955 &  n20066 ;
  assign n20067 = x78 | n19955 ;
  assign n20068 = x78 &  n19955 ;
  assign n20069 = ( n20067 & ~n20068 ) | ( n20067 & 1'b0 ) | ( ~n20068 & 1'b0 ) ;
  assign n20077 = ( n282 & n20063 ) | ( n282 & n20069 ) | ( n20063 & n20069 ) ;
  assign n20078 = ( n20063 & ~n20065 ) | ( n20063 & n20069 ) | ( ~n20065 & n20069 ) ;
  assign n20079 = ~n20077 & n20078 ;
  assign n20080 = n20073 | n20079 ;
  assign n20081 = n19963 &  n20066 ;
  assign n20074 = x77 | n19963 ;
  assign n20075 = x77 &  n19963 ;
  assign n20076 = ( n20074 & ~n20075 ) | ( n20074 & 1'b0 ) | ( ~n20075 & 1'b0 ) ;
  assign n20085 = ( n282 & n20062 ) | ( n282 & n20076 ) | ( n20062 & n20076 ) ;
  assign n20086 = ( n20062 & ~n20065 ) | ( n20062 & n20076 ) | ( ~n20065 & n20076 ) ;
  assign n20087 = ~n20085 & n20086 ;
  assign n20088 = n20081 | n20087 ;
  assign n20089 = n19971 &  n20066 ;
  assign n20082 = x76 | n19971 ;
  assign n20083 = x76 &  n19971 ;
  assign n20084 = ( n20082 & ~n20083 ) | ( n20082 & 1'b0 ) | ( ~n20083 & 1'b0 ) ;
  assign n20093 = ( n282 & n20061 ) | ( n282 & n20084 ) | ( n20061 & n20084 ) ;
  assign n20094 = ( n20061 & ~n20065 ) | ( n20061 & n20084 ) | ( ~n20065 & n20084 ) ;
  assign n20095 = ~n20093 & n20094 ;
  assign n20096 = n20089 | n20095 ;
  assign n20097 = n19979 &  n20066 ;
  assign n20090 = x75 | n19979 ;
  assign n20091 = x75 &  n19979 ;
  assign n20092 = ( n20090 & ~n20091 ) | ( n20090 & 1'b0 ) | ( ~n20091 & 1'b0 ) ;
  assign n20101 = ( n282 & n20060 ) | ( n282 & n20092 ) | ( n20060 & n20092 ) ;
  assign n20102 = ( n20060 & ~n20065 ) | ( n20060 & n20092 ) | ( ~n20065 & n20092 ) ;
  assign n20103 = ~n20101 & n20102 ;
  assign n20104 = n20097 | n20103 ;
  assign n20105 = n19987 &  n20066 ;
  assign n20098 = x74 | n19987 ;
  assign n20099 = x74 &  n19987 ;
  assign n20100 = ( n20098 & ~n20099 ) | ( n20098 & 1'b0 ) | ( ~n20099 & 1'b0 ) ;
  assign n20109 = ( n282 & n20059 ) | ( n282 & n20100 ) | ( n20059 & n20100 ) ;
  assign n20110 = ( n20059 & ~n20065 ) | ( n20059 & n20100 ) | ( ~n20065 & n20100 ) ;
  assign n20111 = ~n20109 & n20110 ;
  assign n20112 = n20105 | n20111 ;
  assign n20113 = n19995 &  n20066 ;
  assign n20106 = x73 | n19995 ;
  assign n20107 = x73 &  n19995 ;
  assign n20108 = ( n20106 & ~n20107 ) | ( n20106 & 1'b0 ) | ( ~n20107 & 1'b0 ) ;
  assign n20117 = ( n282 & n20058 ) | ( n282 & n20108 ) | ( n20058 & n20108 ) ;
  assign n20118 = ( n20058 & ~n20065 ) | ( n20058 & n20108 ) | ( ~n20065 & n20108 ) ;
  assign n20119 = ~n20117 & n20118 ;
  assign n20120 = n20113 | n20119 ;
  assign n20121 = n20003 &  n20066 ;
  assign n20114 = x72 | n20003 ;
  assign n20115 = x72 &  n20003 ;
  assign n20116 = ( n20114 & ~n20115 ) | ( n20114 & 1'b0 ) | ( ~n20115 & 1'b0 ) ;
  assign n20125 = ( n282 & n20057 ) | ( n282 & n20116 ) | ( n20057 & n20116 ) ;
  assign n20126 = ( n20057 & ~n20065 ) | ( n20057 & n20116 ) | ( ~n20065 & n20116 ) ;
  assign n20127 = ~n20125 & n20126 ;
  assign n20128 = n20121 | n20127 ;
  assign n20129 = n20011 &  n20066 ;
  assign n20122 = x71 | n20011 ;
  assign n20123 = x71 &  n20011 ;
  assign n20124 = ( n20122 & ~n20123 ) | ( n20122 & 1'b0 ) | ( ~n20123 & 1'b0 ) ;
  assign n20133 = ( n282 & n20056 ) | ( n282 & n20124 ) | ( n20056 & n20124 ) ;
  assign n20134 = ( n20056 & ~n20065 ) | ( n20056 & n20124 ) | ( ~n20065 & n20124 ) ;
  assign n20135 = ~n20133 & n20134 ;
  assign n20136 = n20129 | n20135 ;
  assign n20137 = n20019 &  n20066 ;
  assign n20130 = x70 | n20019 ;
  assign n20131 = x70 &  n20019 ;
  assign n20132 = ( n20130 & ~n20131 ) | ( n20130 & 1'b0 ) | ( ~n20131 & 1'b0 ) ;
  assign n20141 = ( n282 & n20055 ) | ( n282 & n20132 ) | ( n20055 & n20132 ) ;
  assign n20142 = ( n20055 & ~n20065 ) | ( n20055 & n20132 ) | ( ~n20065 & n20132 ) ;
  assign n20143 = ~n20141 & n20142 ;
  assign n20144 = n20137 | n20143 ;
  assign n20145 = n20027 &  n20066 ;
  assign n20138 = x69 | n20027 ;
  assign n20139 = x69 &  n20027 ;
  assign n20140 = ( n20138 & ~n20139 ) | ( n20138 & 1'b0 ) | ( ~n20139 & 1'b0 ) ;
  assign n20149 = ( n282 & n20054 ) | ( n282 & n20140 ) | ( n20054 & n20140 ) ;
  assign n20150 = ( n20054 & ~n20065 ) | ( n20054 & n20140 ) | ( ~n20065 & n20140 ) ;
  assign n20151 = ~n20149 & n20150 ;
  assign n20152 = n20145 | n20151 ;
  assign n20153 = n20035 &  n20066 ;
  assign n20146 = x68 | n20035 ;
  assign n20147 = x68 &  n20035 ;
  assign n20148 = ( n20146 & ~n20147 ) | ( n20146 & 1'b0 ) | ( ~n20147 & 1'b0 ) ;
  assign n20157 = ( n282 & n20053 ) | ( n282 & n20148 ) | ( n20053 & n20148 ) ;
  assign n20158 = ( n20053 & ~n20065 ) | ( n20053 & n20148 ) | ( ~n20065 & n20148 ) ;
  assign n20159 = ~n20157 & n20158 ;
  assign n20160 = n20153 | n20159 ;
  assign n20161 = n20040 &  n20066 ;
  assign n20154 = x67 | n20040 ;
  assign n20155 = x67 &  n20040 ;
  assign n20156 = ( n20154 & ~n20155 ) | ( n20154 & 1'b0 ) | ( ~n20155 & 1'b0 ) ;
  assign n20165 = ( n282 & n20052 ) | ( n282 & n20156 ) | ( n20052 & n20156 ) ;
  assign n20166 = ( n20052 & ~n20065 ) | ( n20052 & n20156 ) | ( ~n20065 & n20156 ) ;
  assign n20167 = ~n20165 & n20166 ;
  assign n20168 = n20161 | n20167 ;
  assign n20169 = n20046 &  n20066 ;
  assign n20162 = x66 | n20046 ;
  assign n20163 = x66 &  n20046 ;
  assign n20164 = ( n20162 & ~n20163 ) | ( n20162 & 1'b0 ) | ( ~n20163 & 1'b0 ) ;
  assign n20170 = ( n282 & n20051 ) | ( n282 & n20164 ) | ( n20051 & n20164 ) ;
  assign n20171 = ( n20051 & ~n20065 ) | ( n20051 & n20164 ) | ( ~n20065 & n20164 ) ;
  assign n20172 = ~n20170 & n20171 ;
  assign n20173 = n20169 | n20172 ;
  assign n20174 = n20050 &  n20066 ;
  assign n20175 = ( x65 & ~x49 ) | ( x65 & n20047 ) | ( ~x49 & n20047 ) ;
  assign n20176 = ( x49 & ~n20047 ) | ( x49 & x65 ) | ( ~n20047 & x65 ) ;
  assign n20177 = ( n20175 & ~x65 ) | ( n20175 & n20176 ) | ( ~x65 & n20176 ) ;
  assign n20178 = ( n1479 & ~n20065 ) | ( n1479 & n20177 ) | ( ~n20065 & n20177 ) ;
  assign n20179 = ( n282 & n1479 ) | ( n282 & n20177 ) | ( n1479 & n20177 ) ;
  assign n20180 = ( n20178 & ~n20179 ) | ( n20178 & 1'b0 ) | ( ~n20179 & 1'b0 ) ;
  assign n20181 = n20174 | n20180 ;
  assign n20182 = ( n1614 & ~n20065 ) | ( n1614 & 1'b0 ) | ( ~n20065 & 1'b0 ) ;
  assign n20183 = ( x48 & ~n20182 ) | ( x48 & 1'b0 ) | ( ~n20182 & 1'b0 ) ;
  assign n20184 = ( n1619 & ~n20065 ) | ( n1619 & 1'b0 ) | ( ~n20065 & 1'b0 ) ;
  assign n20185 = n20183 | n20184 ;
  assign n20186 = ( x65 & ~n20185 ) | ( x65 & n1622 ) | ( ~n20185 & n1622 ) ;
  assign n20187 = ( x66 & ~n20181 ) | ( x66 & n20186 ) | ( ~n20181 & n20186 ) ;
  assign n20188 = ( x67 & ~n20173 ) | ( x67 & n20187 ) | ( ~n20173 & n20187 ) ;
  assign n20189 = ( x68 & ~n20168 ) | ( x68 & n20188 ) | ( ~n20168 & n20188 ) ;
  assign n20190 = ( x69 & ~n20160 ) | ( x69 & n20189 ) | ( ~n20160 & n20189 ) ;
  assign n20191 = ( x70 & ~n20152 ) | ( x70 & n20190 ) | ( ~n20152 & n20190 ) ;
  assign n20192 = ( x71 & ~n20144 ) | ( x71 & n20191 ) | ( ~n20144 & n20191 ) ;
  assign n20193 = ( x72 & ~n20136 ) | ( x72 & n20192 ) | ( ~n20136 & n20192 ) ;
  assign n20194 = ( x73 & ~n20128 ) | ( x73 & n20193 ) | ( ~n20128 & n20193 ) ;
  assign n20195 = ( x74 & ~n20120 ) | ( x74 & n20194 ) | ( ~n20120 & n20194 ) ;
  assign n20196 = ( x75 & ~n20112 ) | ( x75 & n20195 ) | ( ~n20112 & n20195 ) ;
  assign n20197 = ( x76 & ~n20104 ) | ( x76 & n20196 ) | ( ~n20104 & n20196 ) ;
  assign n20198 = ( x77 & ~n20096 ) | ( x77 & n20197 ) | ( ~n20096 & n20197 ) ;
  assign n20199 = ( x78 & ~n20088 ) | ( x78 & n20198 ) | ( ~n20088 & n20198 ) ;
  assign n20200 = ( x79 & ~n20080 ) | ( x79 & n20199 ) | ( ~n20080 & n20199 ) ;
  assign n20201 = ( x80 & ~n20072 ) | ( x80 & n20200 ) | ( ~n20072 & n20200 ) ;
  assign n20202 = n317 | n20201 ;
  assign n20203 = n20072 &  n20202 ;
  assign n20207 = ( n317 & n20072 ) | ( n317 & n20200 ) | ( n20072 & n20200 ) ;
  assign n20208 = ( x80 & ~n20207 ) | ( x80 & n20072 ) | ( ~n20207 & n20072 ) ;
  assign n20209 = ~x80 & n20208 ;
  assign n20210 = n20203 | n20209 ;
  assign n20211 = ~x81 & n20210 ;
  assign n20212 = n20080 &  n20202 ;
  assign n20204 = x79 | n20080 ;
  assign n20205 = x79 &  n20080 ;
  assign n20206 = ( n20204 & ~n20205 ) | ( n20204 & 1'b0 ) | ( ~n20205 & 1'b0 ) ;
  assign n20216 = ( n317 & n20199 ) | ( n317 & n20206 ) | ( n20199 & n20206 ) ;
  assign n20217 = ( n20199 & ~n20201 ) | ( n20199 & n20206 ) | ( ~n20201 & n20206 ) ;
  assign n20218 = ~n20216 & n20217 ;
  assign n20219 = n20212 | n20218 ;
  assign n20220 = n20088 &  n20202 ;
  assign n20213 = x78 | n20088 ;
  assign n20214 = x78 &  n20088 ;
  assign n20215 = ( n20213 & ~n20214 ) | ( n20213 & 1'b0 ) | ( ~n20214 & 1'b0 ) ;
  assign n20224 = ( n317 & n20198 ) | ( n317 & n20215 ) | ( n20198 & n20215 ) ;
  assign n20225 = ( n20198 & ~n20201 ) | ( n20198 & n20215 ) | ( ~n20201 & n20215 ) ;
  assign n20226 = ~n20224 & n20225 ;
  assign n20227 = n20220 | n20226 ;
  assign n20228 = n20096 &  n20202 ;
  assign n20221 = x77 | n20096 ;
  assign n20222 = x77 &  n20096 ;
  assign n20223 = ( n20221 & ~n20222 ) | ( n20221 & 1'b0 ) | ( ~n20222 & 1'b0 ) ;
  assign n20232 = ( n317 & n20197 ) | ( n317 & n20223 ) | ( n20197 & n20223 ) ;
  assign n20233 = ( n20197 & ~n20201 ) | ( n20197 & n20223 ) | ( ~n20201 & n20223 ) ;
  assign n20234 = ~n20232 & n20233 ;
  assign n20235 = n20228 | n20234 ;
  assign n20236 = n20104 &  n20202 ;
  assign n20229 = x76 | n20104 ;
  assign n20230 = x76 &  n20104 ;
  assign n20231 = ( n20229 & ~n20230 ) | ( n20229 & 1'b0 ) | ( ~n20230 & 1'b0 ) ;
  assign n20240 = ( n317 & n20196 ) | ( n317 & n20231 ) | ( n20196 & n20231 ) ;
  assign n20241 = ( n20196 & ~n20201 ) | ( n20196 & n20231 ) | ( ~n20201 & n20231 ) ;
  assign n20242 = ~n20240 & n20241 ;
  assign n20243 = n20236 | n20242 ;
  assign n20244 = n20112 &  n20202 ;
  assign n20237 = x75 | n20112 ;
  assign n20238 = x75 &  n20112 ;
  assign n20239 = ( n20237 & ~n20238 ) | ( n20237 & 1'b0 ) | ( ~n20238 & 1'b0 ) ;
  assign n20248 = ( n317 & n20195 ) | ( n317 & n20239 ) | ( n20195 & n20239 ) ;
  assign n20249 = ( n20195 & ~n20201 ) | ( n20195 & n20239 ) | ( ~n20201 & n20239 ) ;
  assign n20250 = ~n20248 & n20249 ;
  assign n20251 = n20244 | n20250 ;
  assign n20252 = n20120 &  n20202 ;
  assign n20245 = x74 | n20120 ;
  assign n20246 = x74 &  n20120 ;
  assign n20247 = ( n20245 & ~n20246 ) | ( n20245 & 1'b0 ) | ( ~n20246 & 1'b0 ) ;
  assign n20256 = ( n317 & n20194 ) | ( n317 & n20247 ) | ( n20194 & n20247 ) ;
  assign n20257 = ( n20194 & ~n20201 ) | ( n20194 & n20247 ) | ( ~n20201 & n20247 ) ;
  assign n20258 = ~n20256 & n20257 ;
  assign n20259 = n20252 | n20258 ;
  assign n20260 = n20128 &  n20202 ;
  assign n20253 = x73 | n20128 ;
  assign n20254 = x73 &  n20128 ;
  assign n20255 = ( n20253 & ~n20254 ) | ( n20253 & 1'b0 ) | ( ~n20254 & 1'b0 ) ;
  assign n20264 = ( n317 & n20193 ) | ( n317 & n20255 ) | ( n20193 & n20255 ) ;
  assign n20265 = ( n20193 & ~n20201 ) | ( n20193 & n20255 ) | ( ~n20201 & n20255 ) ;
  assign n20266 = ~n20264 & n20265 ;
  assign n20267 = n20260 | n20266 ;
  assign n20268 = n20136 &  n20202 ;
  assign n20261 = x72 | n20136 ;
  assign n20262 = x72 &  n20136 ;
  assign n20263 = ( n20261 & ~n20262 ) | ( n20261 & 1'b0 ) | ( ~n20262 & 1'b0 ) ;
  assign n20272 = ( n317 & n20192 ) | ( n317 & n20263 ) | ( n20192 & n20263 ) ;
  assign n20273 = ( n20192 & ~n20201 ) | ( n20192 & n20263 ) | ( ~n20201 & n20263 ) ;
  assign n20274 = ~n20272 & n20273 ;
  assign n20275 = n20268 | n20274 ;
  assign n20276 = n20144 &  n20202 ;
  assign n20269 = x71 | n20144 ;
  assign n20270 = x71 &  n20144 ;
  assign n20271 = ( n20269 & ~n20270 ) | ( n20269 & 1'b0 ) | ( ~n20270 & 1'b0 ) ;
  assign n20280 = ( n317 & n20191 ) | ( n317 & n20271 ) | ( n20191 & n20271 ) ;
  assign n20281 = ( n20191 & ~n20201 ) | ( n20191 & n20271 ) | ( ~n20201 & n20271 ) ;
  assign n20282 = ~n20280 & n20281 ;
  assign n20283 = n20276 | n20282 ;
  assign n20284 = n20152 &  n20202 ;
  assign n20277 = x70 | n20152 ;
  assign n20278 = x70 &  n20152 ;
  assign n20279 = ( n20277 & ~n20278 ) | ( n20277 & 1'b0 ) | ( ~n20278 & 1'b0 ) ;
  assign n20288 = ( n317 & n20190 ) | ( n317 & n20279 ) | ( n20190 & n20279 ) ;
  assign n20289 = ( n20190 & ~n20201 ) | ( n20190 & n20279 ) | ( ~n20201 & n20279 ) ;
  assign n20290 = ~n20288 & n20289 ;
  assign n20291 = n20284 | n20290 ;
  assign n20292 = n20160 &  n20202 ;
  assign n20285 = x69 | n20160 ;
  assign n20286 = x69 &  n20160 ;
  assign n20287 = ( n20285 & ~n20286 ) | ( n20285 & 1'b0 ) | ( ~n20286 & 1'b0 ) ;
  assign n20296 = ( n317 & n20189 ) | ( n317 & n20287 ) | ( n20189 & n20287 ) ;
  assign n20297 = ( n20189 & ~n20201 ) | ( n20189 & n20287 ) | ( ~n20201 & n20287 ) ;
  assign n20298 = ~n20296 & n20297 ;
  assign n20299 = n20292 | n20298 ;
  assign n20300 = n20168 &  n20202 ;
  assign n20293 = x68 | n20168 ;
  assign n20294 = x68 &  n20168 ;
  assign n20295 = ( n20293 & ~n20294 ) | ( n20293 & 1'b0 ) | ( ~n20294 & 1'b0 ) ;
  assign n20304 = ( n317 & n20188 ) | ( n317 & n20295 ) | ( n20188 & n20295 ) ;
  assign n20305 = ( n20188 & ~n20201 ) | ( n20188 & n20295 ) | ( ~n20201 & n20295 ) ;
  assign n20306 = ~n20304 & n20305 ;
  assign n20307 = n20300 | n20306 ;
  assign n20308 = n20173 &  n20202 ;
  assign n20301 = x67 | n20173 ;
  assign n20302 = x67 &  n20173 ;
  assign n20303 = ( n20301 & ~n20302 ) | ( n20301 & 1'b0 ) | ( ~n20302 & 1'b0 ) ;
  assign n20312 = ( n317 & n20187 ) | ( n317 & n20303 ) | ( n20187 & n20303 ) ;
  assign n20313 = ( n20187 & ~n20201 ) | ( n20187 & n20303 ) | ( ~n20201 & n20303 ) ;
  assign n20314 = ~n20312 & n20313 ;
  assign n20315 = n20308 | n20314 ;
  assign n20316 = n20181 &  n20202 ;
  assign n20309 = x66 | n20181 ;
  assign n20310 = x66 &  n20181 ;
  assign n20311 = ( n20309 & ~n20310 ) | ( n20309 & 1'b0 ) | ( ~n20310 & 1'b0 ) ;
  assign n20320 = ( n317 & n20186 ) | ( n317 & n20311 ) | ( n20186 & n20311 ) ;
  assign n20321 = ( n20186 & ~n20201 ) | ( n20186 & n20311 ) | ( ~n20201 & n20311 ) ;
  assign n20322 = ~n20320 & n20321 ;
  assign n20323 = n20316 | n20322 ;
  assign n20324 = n20185 &  n20202 ;
  assign n20317 = x65 &  n20185 ;
  assign n20318 = x65 | n20184 ;
  assign n20319 = n20183 | n20318 ;
  assign n20325 = ~n20317 & n20319 ;
  assign n20326 = ( n1622 & ~n20201 ) | ( n1622 & n20325 ) | ( ~n20201 & n20325 ) ;
  assign n20327 = ( n317 & n1622 ) | ( n317 & n20325 ) | ( n1622 & n20325 ) ;
  assign n20328 = ( n20326 & ~n20327 ) | ( n20326 & 1'b0 ) | ( ~n20327 & 1'b0 ) ;
  assign n20329 = n20324 | n20328 ;
  assign n20330 = ( n1758 & ~n20201 ) | ( n1758 & 1'b0 ) | ( ~n20201 & 1'b0 ) ;
  assign n20331 = ( x47 & ~n20330 ) | ( x47 & 1'b0 ) | ( ~n20330 & 1'b0 ) ;
  assign n20332 = ( n1763 & ~n20201 ) | ( n1763 & 1'b0 ) | ( ~n20201 & 1'b0 ) ;
  assign n20333 = n20331 | n20332 ;
  assign n20334 = ( x65 & ~n20333 ) | ( x65 & n1766 ) | ( ~n20333 & n1766 ) ;
  assign n20335 = ( x66 & ~n20329 ) | ( x66 & n20334 ) | ( ~n20329 & n20334 ) ;
  assign n20336 = ( x67 & ~n20323 ) | ( x67 & n20335 ) | ( ~n20323 & n20335 ) ;
  assign n20337 = ( x68 & ~n20315 ) | ( x68 & n20336 ) | ( ~n20315 & n20336 ) ;
  assign n20338 = ( x69 & ~n20307 ) | ( x69 & n20337 ) | ( ~n20307 & n20337 ) ;
  assign n20339 = ( x70 & ~n20299 ) | ( x70 & n20338 ) | ( ~n20299 & n20338 ) ;
  assign n20340 = ( x71 & ~n20291 ) | ( x71 & n20339 ) | ( ~n20291 & n20339 ) ;
  assign n20341 = ( x72 & ~n20283 ) | ( x72 & n20340 ) | ( ~n20283 & n20340 ) ;
  assign n20342 = ( x73 & ~n20275 ) | ( x73 & n20341 ) | ( ~n20275 & n20341 ) ;
  assign n20343 = ( x74 & ~n20267 ) | ( x74 & n20342 ) | ( ~n20267 & n20342 ) ;
  assign n20344 = ( x75 & ~n20259 ) | ( x75 & n20343 ) | ( ~n20259 & n20343 ) ;
  assign n20345 = ( x76 & ~n20251 ) | ( x76 & n20344 ) | ( ~n20251 & n20344 ) ;
  assign n20346 = ( x77 & ~n20243 ) | ( x77 & n20345 ) | ( ~n20243 & n20345 ) ;
  assign n20347 = ( x78 & ~n20235 ) | ( x78 & n20346 ) | ( ~n20235 & n20346 ) ;
  assign n20348 = ( x79 & ~n20227 ) | ( x79 & n20347 ) | ( ~n20227 & n20347 ) ;
  assign n20349 = ( x80 & ~n20219 ) | ( x80 & n20348 ) | ( ~n20219 & n20348 ) ;
  assign n20350 = ( x81 & ~n20203 ) | ( x81 & 1'b0 ) | ( ~n20203 & 1'b0 ) ;
  assign n20351 = ~n20209 & n20350 ;
  assign n20352 = ( n20349 & ~n20211 ) | ( n20349 & n20351 ) | ( ~n20211 & n20351 ) ;
  assign n20353 = ( n20211 & ~n1803 ) | ( n20211 & n20352 ) | ( ~n1803 & n20352 ) ;
  assign n20354 = n1803 | n20353 ;
  assign n20361 = n317 &  n20072 ;
  assign n20362 = n20354 &  n20361 ;
  assign n20355 = ~n317 & n20210 ;
  assign n20356 = ( n20354 & ~n20355 ) | ( n20354 & 1'b0 ) | ( ~n20355 & 1'b0 ) ;
  assign n20360 = n20211 | n20351 ;
  assign n20364 = ( n20349 & n20356 ) | ( n20349 & n20360 ) | ( n20356 & n20360 ) ;
  assign n20363 = n20349 | n20360 ;
  assign n20365 = ( n20362 & ~n20364 ) | ( n20362 & n20363 ) | ( ~n20364 & n20363 ) ;
  assign n20369 = ( n20219 & ~n20355 ) | ( n20219 & 1'b0 ) | ( ~n20355 & 1'b0 ) ;
  assign n20370 = n20354 &  n20369 ;
  assign n20357 = x80 | n20219 ;
  assign n20358 = x80 &  n20219 ;
  assign n20359 = ( n20357 & ~n20358 ) | ( n20357 & 1'b0 ) | ( ~n20358 & 1'b0 ) ;
  assign n20372 = ( n20348 & n20356 ) | ( n20348 & n20359 ) | ( n20356 & n20359 ) ;
  assign n20371 = n20348 | n20359 ;
  assign n20373 = ( n20370 & ~n20372 ) | ( n20370 & n20371 ) | ( ~n20372 & n20371 ) ;
  assign n20377 = ( n20227 & ~n20355 ) | ( n20227 & 1'b0 ) | ( ~n20355 & 1'b0 ) ;
  assign n20378 = n20354 &  n20377 ;
  assign n20366 = x79 | n20227 ;
  assign n20367 = x79 &  n20227 ;
  assign n20368 = ( n20366 & ~n20367 ) | ( n20366 & 1'b0 ) | ( ~n20367 & 1'b0 ) ;
  assign n20380 = ( n20347 & n20356 ) | ( n20347 & n20368 ) | ( n20356 & n20368 ) ;
  assign n20379 = n20347 | n20368 ;
  assign n20381 = ( n20378 & ~n20380 ) | ( n20378 & n20379 ) | ( ~n20380 & n20379 ) ;
  assign n20385 = ( n20235 & ~n20355 ) | ( n20235 & 1'b0 ) | ( ~n20355 & 1'b0 ) ;
  assign n20386 = n20354 &  n20385 ;
  assign n20374 = x78 | n20235 ;
  assign n20375 = x78 &  n20235 ;
  assign n20376 = ( n20374 & ~n20375 ) | ( n20374 & 1'b0 ) | ( ~n20375 & 1'b0 ) ;
  assign n20388 = ( n20346 & n20356 ) | ( n20346 & n20376 ) | ( n20356 & n20376 ) ;
  assign n20387 = n20346 | n20376 ;
  assign n20389 = ( n20386 & ~n20388 ) | ( n20386 & n20387 ) | ( ~n20388 & n20387 ) ;
  assign n20393 = ( n20243 & ~n20355 ) | ( n20243 & 1'b0 ) | ( ~n20355 & 1'b0 ) ;
  assign n20394 = n20354 &  n20393 ;
  assign n20382 = x77 | n20243 ;
  assign n20383 = x77 &  n20243 ;
  assign n20384 = ( n20382 & ~n20383 ) | ( n20382 & 1'b0 ) | ( ~n20383 & 1'b0 ) ;
  assign n20396 = ( n20345 & n20356 ) | ( n20345 & n20384 ) | ( n20356 & n20384 ) ;
  assign n20395 = n20345 | n20384 ;
  assign n20397 = ( n20394 & ~n20396 ) | ( n20394 & n20395 ) | ( ~n20396 & n20395 ) ;
  assign n20401 = ( n20251 & ~n20355 ) | ( n20251 & 1'b0 ) | ( ~n20355 & 1'b0 ) ;
  assign n20402 = n20354 &  n20401 ;
  assign n20390 = x76 | n20251 ;
  assign n20391 = x76 &  n20251 ;
  assign n20392 = ( n20390 & ~n20391 ) | ( n20390 & 1'b0 ) | ( ~n20391 & 1'b0 ) ;
  assign n20404 = ( n20344 & n20356 ) | ( n20344 & n20392 ) | ( n20356 & n20392 ) ;
  assign n20403 = n20344 | n20392 ;
  assign n20405 = ( n20402 & ~n20404 ) | ( n20402 & n20403 ) | ( ~n20404 & n20403 ) ;
  assign n20409 = ( n20259 & ~n20355 ) | ( n20259 & 1'b0 ) | ( ~n20355 & 1'b0 ) ;
  assign n20410 = n20354 &  n20409 ;
  assign n20398 = x75 | n20259 ;
  assign n20399 = x75 &  n20259 ;
  assign n20400 = ( n20398 & ~n20399 ) | ( n20398 & 1'b0 ) | ( ~n20399 & 1'b0 ) ;
  assign n20412 = ( n20343 & n20356 ) | ( n20343 & n20400 ) | ( n20356 & n20400 ) ;
  assign n20411 = n20343 | n20400 ;
  assign n20413 = ( n20410 & ~n20412 ) | ( n20410 & n20411 ) | ( ~n20412 & n20411 ) ;
  assign n20417 = ( n20267 & ~n20355 ) | ( n20267 & 1'b0 ) | ( ~n20355 & 1'b0 ) ;
  assign n20418 = n20354 &  n20417 ;
  assign n20406 = x74 | n20267 ;
  assign n20407 = x74 &  n20267 ;
  assign n20408 = ( n20406 & ~n20407 ) | ( n20406 & 1'b0 ) | ( ~n20407 & 1'b0 ) ;
  assign n20420 = ( n20342 & n20356 ) | ( n20342 & n20408 ) | ( n20356 & n20408 ) ;
  assign n20419 = n20342 | n20408 ;
  assign n20421 = ( n20418 & ~n20420 ) | ( n20418 & n20419 ) | ( ~n20420 & n20419 ) ;
  assign n20425 = ( n20275 & ~n20355 ) | ( n20275 & 1'b0 ) | ( ~n20355 & 1'b0 ) ;
  assign n20426 = n20354 &  n20425 ;
  assign n20414 = x73 | n20275 ;
  assign n20415 = x73 &  n20275 ;
  assign n20416 = ( n20414 & ~n20415 ) | ( n20414 & 1'b0 ) | ( ~n20415 & 1'b0 ) ;
  assign n20428 = ( n20341 & n20356 ) | ( n20341 & n20416 ) | ( n20356 & n20416 ) ;
  assign n20427 = n20341 | n20416 ;
  assign n20429 = ( n20426 & ~n20428 ) | ( n20426 & n20427 ) | ( ~n20428 & n20427 ) ;
  assign n20433 = ( n20283 & ~n20355 ) | ( n20283 & 1'b0 ) | ( ~n20355 & 1'b0 ) ;
  assign n20434 = n20354 &  n20433 ;
  assign n20422 = x72 | n20283 ;
  assign n20423 = x72 &  n20283 ;
  assign n20424 = ( n20422 & ~n20423 ) | ( n20422 & 1'b0 ) | ( ~n20423 & 1'b0 ) ;
  assign n20436 = ( n20340 & n20356 ) | ( n20340 & n20424 ) | ( n20356 & n20424 ) ;
  assign n20435 = n20340 | n20424 ;
  assign n20437 = ( n20434 & ~n20436 ) | ( n20434 & n20435 ) | ( ~n20436 & n20435 ) ;
  assign n20441 = ( n20291 & ~n20355 ) | ( n20291 & 1'b0 ) | ( ~n20355 & 1'b0 ) ;
  assign n20442 = n20354 &  n20441 ;
  assign n20430 = x71 | n20291 ;
  assign n20431 = x71 &  n20291 ;
  assign n20432 = ( n20430 & ~n20431 ) | ( n20430 & 1'b0 ) | ( ~n20431 & 1'b0 ) ;
  assign n20444 = ( n20339 & n20356 ) | ( n20339 & n20432 ) | ( n20356 & n20432 ) ;
  assign n20443 = n20339 | n20432 ;
  assign n20445 = ( n20442 & ~n20444 ) | ( n20442 & n20443 ) | ( ~n20444 & n20443 ) ;
  assign n20449 = ( n20299 & ~n20355 ) | ( n20299 & 1'b0 ) | ( ~n20355 & 1'b0 ) ;
  assign n20450 = n20354 &  n20449 ;
  assign n20438 = x70 | n20299 ;
  assign n20439 = x70 &  n20299 ;
  assign n20440 = ( n20438 & ~n20439 ) | ( n20438 & 1'b0 ) | ( ~n20439 & 1'b0 ) ;
  assign n20452 = ( n20338 & n20356 ) | ( n20338 & n20440 ) | ( n20356 & n20440 ) ;
  assign n20451 = n20338 | n20440 ;
  assign n20453 = ( n20450 & ~n20452 ) | ( n20450 & n20451 ) | ( ~n20452 & n20451 ) ;
  assign n20457 = ( n20307 & ~n20355 ) | ( n20307 & 1'b0 ) | ( ~n20355 & 1'b0 ) ;
  assign n20458 = n20354 &  n20457 ;
  assign n20446 = x69 | n20307 ;
  assign n20447 = x69 &  n20307 ;
  assign n20448 = ( n20446 & ~n20447 ) | ( n20446 & 1'b0 ) | ( ~n20447 & 1'b0 ) ;
  assign n20460 = ( n20337 & n20356 ) | ( n20337 & n20448 ) | ( n20356 & n20448 ) ;
  assign n20459 = n20337 | n20448 ;
  assign n20461 = ( n20458 & ~n20460 ) | ( n20458 & n20459 ) | ( ~n20460 & n20459 ) ;
  assign n20465 = ( n20315 & ~n20355 ) | ( n20315 & 1'b0 ) | ( ~n20355 & 1'b0 ) ;
  assign n20466 = n20354 &  n20465 ;
  assign n20454 = x68 | n20315 ;
  assign n20455 = x68 &  n20315 ;
  assign n20456 = ( n20454 & ~n20455 ) | ( n20454 & 1'b0 ) | ( ~n20455 & 1'b0 ) ;
  assign n20468 = ( n20336 & n20356 ) | ( n20336 & n20456 ) | ( n20356 & n20456 ) ;
  assign n20467 = n20336 | n20456 ;
  assign n20469 = ( n20466 & ~n20468 ) | ( n20466 & n20467 ) | ( ~n20468 & n20467 ) ;
  assign n20473 = ( n20323 & ~n20355 ) | ( n20323 & 1'b0 ) | ( ~n20355 & 1'b0 ) ;
  assign n20474 = n20354 &  n20473 ;
  assign n20462 = x67 | n20323 ;
  assign n20463 = x67 &  n20323 ;
  assign n20464 = ( n20462 & ~n20463 ) | ( n20462 & 1'b0 ) | ( ~n20463 & 1'b0 ) ;
  assign n20476 = ( n20335 & n20356 ) | ( n20335 & n20464 ) | ( n20356 & n20464 ) ;
  assign n20475 = n20335 | n20464 ;
  assign n20477 = ( n20474 & ~n20476 ) | ( n20474 & n20475 ) | ( ~n20476 & n20475 ) ;
  assign n20478 = ( n20329 & ~n20355 ) | ( n20329 & 1'b0 ) | ( ~n20355 & 1'b0 ) ;
  assign n20479 = n20354 &  n20478 ;
  assign n20470 = x66 | n20329 ;
  assign n20471 = x66 &  n20329 ;
  assign n20472 = ( n20470 & ~n20471 ) | ( n20470 & 1'b0 ) | ( ~n20471 & 1'b0 ) ;
  assign n20481 = ( n20334 & n20356 ) | ( n20334 & n20472 ) | ( n20356 & n20472 ) ;
  assign n20480 = n20334 | n20472 ;
  assign n20482 = ( n20479 & ~n20481 ) | ( n20479 & n20480 ) | ( ~n20481 & n20480 ) ;
  assign n20483 = ( x65 & ~n1766 ) | ( x65 & n20333 ) | ( ~n1766 & n20333 ) ;
  assign n20484 = ( n20334 & ~x65 ) | ( n20334 & n20483 ) | ( ~x65 & n20483 ) ;
  assign n20485 = ~n20356 & n20484 ;
  assign n20486 = ( n20333 & ~n20355 ) | ( n20333 & 1'b0 ) | ( ~n20355 & 1'b0 ) ;
  assign n20487 = n20354 &  n20486 ;
  assign n20488 = n20485 | n20487 ;
  assign n20489 = ( x64 & ~n20356 ) | ( x64 & 1'b0 ) | ( ~n20356 & 1'b0 ) ;
  assign n20490 = ( x46 & ~n20489 ) | ( x46 & 1'b0 ) | ( ~n20489 & 1'b0 ) ;
  assign n20491 = ( n1766 & ~n20356 ) | ( n1766 & 1'b0 ) | ( ~n20356 & 1'b0 ) ;
  assign n20492 = n20490 | n20491 ;
  assign n20493 = ( x65 & ~n20492 ) | ( x65 & n1941 ) | ( ~n20492 & n1941 ) ;
  assign n20494 = ( x66 & ~n20488 ) | ( x66 & n20493 ) | ( ~n20488 & n20493 ) ;
  assign n20495 = ( x67 & ~n20482 ) | ( x67 & n20494 ) | ( ~n20482 & n20494 ) ;
  assign n20496 = ( x68 & ~n20477 ) | ( x68 & n20495 ) | ( ~n20477 & n20495 ) ;
  assign n20497 = ( x69 & ~n20469 ) | ( x69 & n20496 ) | ( ~n20469 & n20496 ) ;
  assign n20498 = ( x70 & ~n20461 ) | ( x70 & n20497 ) | ( ~n20461 & n20497 ) ;
  assign n20499 = ( x71 & ~n20453 ) | ( x71 & n20498 ) | ( ~n20453 & n20498 ) ;
  assign n20500 = ( x72 & ~n20445 ) | ( x72 & n20499 ) | ( ~n20445 & n20499 ) ;
  assign n20501 = ( x73 & ~n20437 ) | ( x73 & n20500 ) | ( ~n20437 & n20500 ) ;
  assign n20502 = ( x74 & ~n20429 ) | ( x74 & n20501 ) | ( ~n20429 & n20501 ) ;
  assign n20503 = ( x75 & ~n20421 ) | ( x75 & n20502 ) | ( ~n20421 & n20502 ) ;
  assign n20504 = ( x76 & ~n20413 ) | ( x76 & n20503 ) | ( ~n20413 & n20503 ) ;
  assign n20505 = ( x77 & ~n20405 ) | ( x77 & n20504 ) | ( ~n20405 & n20504 ) ;
  assign n20506 = ( x78 & ~n20397 ) | ( x78 & n20505 ) | ( ~n20397 & n20505 ) ;
  assign n20507 = ( x79 & ~n20389 ) | ( x79 & n20506 ) | ( ~n20389 & n20506 ) ;
  assign n20508 = ( x80 & ~n20381 ) | ( x80 & n20507 ) | ( ~n20381 & n20507 ) ;
  assign n20509 = ( x81 & ~n20373 ) | ( x81 & n20508 ) | ( ~n20373 & n20508 ) ;
  assign n20516 = ( x82 & ~n1963 ) | ( x82 & n20509 ) | ( ~n1963 & n20509 ) ;
  assign n20515 = x82 &  n20509 ;
  assign n20517 = ( n20365 & ~n20516 ) | ( n20365 & n20515 ) | ( ~n20516 & n20515 ) ;
  assign n20510 = ( x82 & ~n20365 ) | ( x82 & n20509 ) | ( ~n20365 & n20509 ) ;
  assign n20511 = n1963 | n20510 ;
  assign n20518 = n20373 &  n20511 ;
  assign n20512 = x81 | n20373 ;
  assign n20513 = x81 &  n20373 ;
  assign n20514 = ( n20512 & ~n20513 ) | ( n20512 & 1'b0 ) | ( ~n20513 & 1'b0 ) ;
  assign n20522 = ( n1963 & n20508 ) | ( n1963 & n20514 ) | ( n20508 & n20514 ) ;
  assign n20523 = ( n20508 & ~n20510 ) | ( n20508 & n20514 ) | ( ~n20510 & n20514 ) ;
  assign n20524 = ~n20522 & n20523 ;
  assign n20525 = n20518 | n20524 ;
  assign n20526 = n20381 &  n20511 ;
  assign n20519 = x80 | n20381 ;
  assign n20520 = x80 &  n20381 ;
  assign n20521 = ( n20519 & ~n20520 ) | ( n20519 & 1'b0 ) | ( ~n20520 & 1'b0 ) ;
  assign n20530 = ( n1963 & n20507 ) | ( n1963 & n20521 ) | ( n20507 & n20521 ) ;
  assign n20531 = ( n20507 & ~n20510 ) | ( n20507 & n20521 ) | ( ~n20510 & n20521 ) ;
  assign n20532 = ~n20530 & n20531 ;
  assign n20533 = n20526 | n20532 ;
  assign n20534 = n20389 &  n20511 ;
  assign n20527 = x79 | n20389 ;
  assign n20528 = x79 &  n20389 ;
  assign n20529 = ( n20527 & ~n20528 ) | ( n20527 & 1'b0 ) | ( ~n20528 & 1'b0 ) ;
  assign n20538 = ( n1963 & n20506 ) | ( n1963 & n20529 ) | ( n20506 & n20529 ) ;
  assign n20539 = ( n20506 & ~n20510 ) | ( n20506 & n20529 ) | ( ~n20510 & n20529 ) ;
  assign n20540 = ~n20538 & n20539 ;
  assign n20541 = n20534 | n20540 ;
  assign n20542 = n20397 &  n20511 ;
  assign n20535 = x78 | n20397 ;
  assign n20536 = x78 &  n20397 ;
  assign n20537 = ( n20535 & ~n20536 ) | ( n20535 & 1'b0 ) | ( ~n20536 & 1'b0 ) ;
  assign n20546 = ( n1963 & n20505 ) | ( n1963 & n20537 ) | ( n20505 & n20537 ) ;
  assign n20547 = ( n20505 & ~n20510 ) | ( n20505 & n20537 ) | ( ~n20510 & n20537 ) ;
  assign n20548 = ~n20546 & n20547 ;
  assign n20549 = n20542 | n20548 ;
  assign n20550 = n20405 &  n20511 ;
  assign n20543 = x77 | n20405 ;
  assign n20544 = x77 &  n20405 ;
  assign n20545 = ( n20543 & ~n20544 ) | ( n20543 & 1'b0 ) | ( ~n20544 & 1'b0 ) ;
  assign n20554 = ( n1963 & n20504 ) | ( n1963 & n20545 ) | ( n20504 & n20545 ) ;
  assign n20555 = ( n20504 & ~n20510 ) | ( n20504 & n20545 ) | ( ~n20510 & n20545 ) ;
  assign n20556 = ~n20554 & n20555 ;
  assign n20557 = n20550 | n20556 ;
  assign n20558 = n20413 &  n20511 ;
  assign n20551 = x76 | n20413 ;
  assign n20552 = x76 &  n20413 ;
  assign n20553 = ( n20551 & ~n20552 ) | ( n20551 & 1'b0 ) | ( ~n20552 & 1'b0 ) ;
  assign n20562 = ( n1963 & n20503 ) | ( n1963 & n20553 ) | ( n20503 & n20553 ) ;
  assign n20563 = ( n20503 & ~n20510 ) | ( n20503 & n20553 ) | ( ~n20510 & n20553 ) ;
  assign n20564 = ~n20562 & n20563 ;
  assign n20565 = n20558 | n20564 ;
  assign n20566 = n20421 &  n20511 ;
  assign n20559 = x75 | n20421 ;
  assign n20560 = x75 &  n20421 ;
  assign n20561 = ( n20559 & ~n20560 ) | ( n20559 & 1'b0 ) | ( ~n20560 & 1'b0 ) ;
  assign n20570 = ( n1963 & n20502 ) | ( n1963 & n20561 ) | ( n20502 & n20561 ) ;
  assign n20571 = ( n20502 & ~n20510 ) | ( n20502 & n20561 ) | ( ~n20510 & n20561 ) ;
  assign n20572 = ~n20570 & n20571 ;
  assign n20573 = n20566 | n20572 ;
  assign n20574 = n20429 &  n20511 ;
  assign n20567 = x74 | n20429 ;
  assign n20568 = x74 &  n20429 ;
  assign n20569 = ( n20567 & ~n20568 ) | ( n20567 & 1'b0 ) | ( ~n20568 & 1'b0 ) ;
  assign n20578 = ( n1963 & n20501 ) | ( n1963 & n20569 ) | ( n20501 & n20569 ) ;
  assign n20579 = ( n20501 & ~n20510 ) | ( n20501 & n20569 ) | ( ~n20510 & n20569 ) ;
  assign n20580 = ~n20578 & n20579 ;
  assign n20581 = n20574 | n20580 ;
  assign n20582 = n20437 &  n20511 ;
  assign n20575 = x73 | n20437 ;
  assign n20576 = x73 &  n20437 ;
  assign n20577 = ( n20575 & ~n20576 ) | ( n20575 & 1'b0 ) | ( ~n20576 & 1'b0 ) ;
  assign n20586 = ( n1963 & n20500 ) | ( n1963 & n20577 ) | ( n20500 & n20577 ) ;
  assign n20587 = ( n20500 & ~n20510 ) | ( n20500 & n20577 ) | ( ~n20510 & n20577 ) ;
  assign n20588 = ~n20586 & n20587 ;
  assign n20589 = n20582 | n20588 ;
  assign n20590 = n20445 &  n20511 ;
  assign n20583 = x72 | n20445 ;
  assign n20584 = x72 &  n20445 ;
  assign n20585 = ( n20583 & ~n20584 ) | ( n20583 & 1'b0 ) | ( ~n20584 & 1'b0 ) ;
  assign n20594 = ( n1963 & n20499 ) | ( n1963 & n20585 ) | ( n20499 & n20585 ) ;
  assign n20595 = ( n20499 & ~n20510 ) | ( n20499 & n20585 ) | ( ~n20510 & n20585 ) ;
  assign n20596 = ~n20594 & n20595 ;
  assign n20597 = n20590 | n20596 ;
  assign n20598 = n20453 &  n20511 ;
  assign n20591 = x71 | n20453 ;
  assign n20592 = x71 &  n20453 ;
  assign n20593 = ( n20591 & ~n20592 ) | ( n20591 & 1'b0 ) | ( ~n20592 & 1'b0 ) ;
  assign n20602 = ( n1963 & n20498 ) | ( n1963 & n20593 ) | ( n20498 & n20593 ) ;
  assign n20603 = ( n20498 & ~n20510 ) | ( n20498 & n20593 ) | ( ~n20510 & n20593 ) ;
  assign n20604 = ~n20602 & n20603 ;
  assign n20605 = n20598 | n20604 ;
  assign n20606 = n20461 &  n20511 ;
  assign n20599 = x70 | n20461 ;
  assign n20600 = x70 &  n20461 ;
  assign n20601 = ( n20599 & ~n20600 ) | ( n20599 & 1'b0 ) | ( ~n20600 & 1'b0 ) ;
  assign n20610 = ( n1963 & n20497 ) | ( n1963 & n20601 ) | ( n20497 & n20601 ) ;
  assign n20611 = ( n20497 & ~n20510 ) | ( n20497 & n20601 ) | ( ~n20510 & n20601 ) ;
  assign n20612 = ~n20610 & n20611 ;
  assign n20613 = n20606 | n20612 ;
  assign n20614 = n20469 &  n20511 ;
  assign n20607 = x69 | n20469 ;
  assign n20608 = x69 &  n20469 ;
  assign n20609 = ( n20607 & ~n20608 ) | ( n20607 & 1'b0 ) | ( ~n20608 & 1'b0 ) ;
  assign n20618 = ( n1963 & n20496 ) | ( n1963 & n20609 ) | ( n20496 & n20609 ) ;
  assign n20619 = ( n20496 & ~n20510 ) | ( n20496 & n20609 ) | ( ~n20510 & n20609 ) ;
  assign n20620 = ~n20618 & n20619 ;
  assign n20621 = n20614 | n20620 ;
  assign n20622 = n20477 &  n20511 ;
  assign n20615 = x68 | n20477 ;
  assign n20616 = x68 &  n20477 ;
  assign n20617 = ( n20615 & ~n20616 ) | ( n20615 & 1'b0 ) | ( ~n20616 & 1'b0 ) ;
  assign n20626 = ( n1963 & n20495 ) | ( n1963 & n20617 ) | ( n20495 & n20617 ) ;
  assign n20627 = ( n20495 & ~n20510 ) | ( n20495 & n20617 ) | ( ~n20510 & n20617 ) ;
  assign n20628 = ~n20626 & n20627 ;
  assign n20629 = n20622 | n20628 ;
  assign n20630 = n20482 &  n20511 ;
  assign n20623 = x67 | n20482 ;
  assign n20624 = x67 &  n20482 ;
  assign n20625 = ( n20623 & ~n20624 ) | ( n20623 & 1'b0 ) | ( ~n20624 & 1'b0 ) ;
  assign n20634 = ( n1963 & n20494 ) | ( n1963 & n20625 ) | ( n20494 & n20625 ) ;
  assign n20635 = ( n20494 & ~n20510 ) | ( n20494 & n20625 ) | ( ~n20510 & n20625 ) ;
  assign n20636 = ~n20634 & n20635 ;
  assign n20637 = n20630 | n20636 ;
  assign n20638 = n20488 &  n20511 ;
  assign n20631 = x66 | n20488 ;
  assign n20632 = x66 &  n20488 ;
  assign n20633 = ( n20631 & ~n20632 ) | ( n20631 & 1'b0 ) | ( ~n20632 & 1'b0 ) ;
  assign n20639 = ( n1963 & n20493 ) | ( n1963 & n20633 ) | ( n20493 & n20633 ) ;
  assign n20640 = ( n20493 & ~n20510 ) | ( n20493 & n20633 ) | ( ~n20510 & n20633 ) ;
  assign n20641 = ~n20639 & n20640 ;
  assign n20642 = n20638 | n20641 ;
  assign n20643 = n20492 &  n20511 ;
  assign n20644 = ( x65 & ~x46 ) | ( x65 & n20489 ) | ( ~x46 & n20489 ) ;
  assign n20645 = ( x46 & ~n20489 ) | ( x46 & x65 ) | ( ~n20489 & x65 ) ;
  assign n20646 = ( n20644 & ~x65 ) | ( n20644 & n20645 ) | ( ~x65 & n20645 ) ;
  assign n20647 = ( n1941 & ~n1963 ) | ( n1941 & n20646 ) | ( ~n1963 & n20646 ) ;
  assign n20648 = ( n1941 & n20510 ) | ( n1941 & n20646 ) | ( n20510 & n20646 ) ;
  assign n20649 = ( n20647 & ~n20648 ) | ( n20647 & 1'b0 ) | ( ~n20648 & 1'b0 ) ;
  assign n20650 = n20643 | n20649 ;
  assign n20651 = ( n2110 & ~n20510 ) | ( n2110 & 1'b0 ) | ( ~n20510 & 1'b0 ) ;
  assign n20652 = ( x45 & ~n20651 ) | ( x45 & 1'b0 ) | ( ~n20651 & 1'b0 ) ;
  assign n20653 = ( n2117 & ~n20510 ) | ( n2117 & 1'b0 ) | ( ~n20510 & 1'b0 ) ;
  assign n20654 = n20652 | n20653 ;
  assign n20655 = ( x65 & ~n20654 ) | ( x65 & n2120 ) | ( ~n20654 & n2120 ) ;
  assign n20656 = ( x66 & ~n20650 ) | ( x66 & n20655 ) | ( ~n20650 & n20655 ) ;
  assign n20657 = ( x67 & ~n20642 ) | ( x67 & n20656 ) | ( ~n20642 & n20656 ) ;
  assign n20658 = ( x68 & ~n20637 ) | ( x68 & n20657 ) | ( ~n20637 & n20657 ) ;
  assign n20659 = ( x69 & ~n20629 ) | ( x69 & n20658 ) | ( ~n20629 & n20658 ) ;
  assign n20660 = ( x70 & ~n20621 ) | ( x70 & n20659 ) | ( ~n20621 & n20659 ) ;
  assign n20661 = ( x71 & ~n20613 ) | ( x71 & n20660 ) | ( ~n20613 & n20660 ) ;
  assign n20662 = ( x72 & ~n20605 ) | ( x72 & n20661 ) | ( ~n20605 & n20661 ) ;
  assign n20663 = ( x73 & ~n20597 ) | ( x73 & n20662 ) | ( ~n20597 & n20662 ) ;
  assign n20664 = ( x74 & ~n20589 ) | ( x74 & n20663 ) | ( ~n20589 & n20663 ) ;
  assign n20665 = ( x75 & ~n20581 ) | ( x75 & n20664 ) | ( ~n20581 & n20664 ) ;
  assign n20666 = ( x76 & ~n20573 ) | ( x76 & n20665 ) | ( ~n20573 & n20665 ) ;
  assign n20667 = ( x77 & ~n20565 ) | ( x77 & n20666 ) | ( ~n20565 & n20666 ) ;
  assign n20668 = ( x78 & ~n20557 ) | ( x78 & n20667 ) | ( ~n20557 & n20667 ) ;
  assign n20669 = ( x79 & ~n20549 ) | ( x79 & n20668 ) | ( ~n20549 & n20668 ) ;
  assign n20670 = ( x80 & ~n20541 ) | ( x80 & n20669 ) | ( ~n20541 & n20669 ) ;
  assign n20671 = ( x81 & ~n20533 ) | ( x81 & n20670 ) | ( ~n20533 & n20670 ) ;
  assign n20672 = ( x82 & ~n20525 ) | ( x82 & n20671 ) | ( ~n20525 & n20671 ) ;
  assign n20673 = ( x83 & ~n20517 ) | ( x83 & n20672 ) | ( ~n20517 & n20672 ) ;
  assign n20674 = n192 | n20673 ;
  assign n20675 = n20517 &  n20674 ;
  assign n20679 = ( n192 & n20517 ) | ( n192 & n20672 ) | ( n20517 & n20672 ) ;
  assign n20680 = ( x83 & ~n20679 ) | ( x83 & n20517 ) | ( ~n20679 & n20517 ) ;
  assign n20681 = ~x83 & n20680 ;
  assign n20682 = n20675 | n20681 ;
  assign n20683 = ~x84 & n20682 ;
  assign n20684 = n20525 &  n20674 ;
  assign n20676 = x82 | n20525 ;
  assign n20677 = x82 &  n20525 ;
  assign n20678 = ( n20676 & ~n20677 ) | ( n20676 & 1'b0 ) | ( ~n20677 & 1'b0 ) ;
  assign n20688 = ( n192 & n20671 ) | ( n192 & n20678 ) | ( n20671 & n20678 ) ;
  assign n20689 = ( n20671 & ~n20673 ) | ( n20671 & n20678 ) | ( ~n20673 & n20678 ) ;
  assign n20690 = ~n20688 & n20689 ;
  assign n20691 = n20684 | n20690 ;
  assign n20692 = n20533 &  n20674 ;
  assign n20685 = x81 | n20533 ;
  assign n20686 = x81 &  n20533 ;
  assign n20687 = ( n20685 & ~n20686 ) | ( n20685 & 1'b0 ) | ( ~n20686 & 1'b0 ) ;
  assign n20696 = ( n192 & n20670 ) | ( n192 & n20687 ) | ( n20670 & n20687 ) ;
  assign n20697 = ( n20670 & ~n20673 ) | ( n20670 & n20687 ) | ( ~n20673 & n20687 ) ;
  assign n20698 = ~n20696 & n20697 ;
  assign n20699 = n20692 | n20698 ;
  assign n20700 = n20541 &  n20674 ;
  assign n20693 = x80 | n20541 ;
  assign n20694 = x80 &  n20541 ;
  assign n20695 = ( n20693 & ~n20694 ) | ( n20693 & 1'b0 ) | ( ~n20694 & 1'b0 ) ;
  assign n20704 = ( n192 & n20669 ) | ( n192 & n20695 ) | ( n20669 & n20695 ) ;
  assign n20705 = ( n20669 & ~n20673 ) | ( n20669 & n20695 ) | ( ~n20673 & n20695 ) ;
  assign n20706 = ~n20704 & n20705 ;
  assign n20707 = n20700 | n20706 ;
  assign n20708 = n20549 &  n20674 ;
  assign n20701 = x79 | n20549 ;
  assign n20702 = x79 &  n20549 ;
  assign n20703 = ( n20701 & ~n20702 ) | ( n20701 & 1'b0 ) | ( ~n20702 & 1'b0 ) ;
  assign n20712 = ( n192 & n20668 ) | ( n192 & n20703 ) | ( n20668 & n20703 ) ;
  assign n20713 = ( n20668 & ~n20673 ) | ( n20668 & n20703 ) | ( ~n20673 & n20703 ) ;
  assign n20714 = ~n20712 & n20713 ;
  assign n20715 = n20708 | n20714 ;
  assign n20716 = n20557 &  n20674 ;
  assign n20709 = x78 | n20557 ;
  assign n20710 = x78 &  n20557 ;
  assign n20711 = ( n20709 & ~n20710 ) | ( n20709 & 1'b0 ) | ( ~n20710 & 1'b0 ) ;
  assign n20720 = ( n192 & n20667 ) | ( n192 & n20711 ) | ( n20667 & n20711 ) ;
  assign n20721 = ( n20667 & ~n20673 ) | ( n20667 & n20711 ) | ( ~n20673 & n20711 ) ;
  assign n20722 = ~n20720 & n20721 ;
  assign n20723 = n20716 | n20722 ;
  assign n20724 = n20565 &  n20674 ;
  assign n20717 = x77 | n20565 ;
  assign n20718 = x77 &  n20565 ;
  assign n20719 = ( n20717 & ~n20718 ) | ( n20717 & 1'b0 ) | ( ~n20718 & 1'b0 ) ;
  assign n20728 = ( n192 & n20666 ) | ( n192 & n20719 ) | ( n20666 & n20719 ) ;
  assign n20729 = ( n20666 & ~n20673 ) | ( n20666 & n20719 ) | ( ~n20673 & n20719 ) ;
  assign n20730 = ~n20728 & n20729 ;
  assign n20731 = n20724 | n20730 ;
  assign n20732 = n20573 &  n20674 ;
  assign n20725 = x76 | n20573 ;
  assign n20726 = x76 &  n20573 ;
  assign n20727 = ( n20725 & ~n20726 ) | ( n20725 & 1'b0 ) | ( ~n20726 & 1'b0 ) ;
  assign n20736 = ( n192 & n20665 ) | ( n192 & n20727 ) | ( n20665 & n20727 ) ;
  assign n20737 = ( n20665 & ~n20673 ) | ( n20665 & n20727 ) | ( ~n20673 & n20727 ) ;
  assign n20738 = ~n20736 & n20737 ;
  assign n20739 = n20732 | n20738 ;
  assign n20740 = n20581 &  n20674 ;
  assign n20733 = x75 | n20581 ;
  assign n20734 = x75 &  n20581 ;
  assign n20735 = ( n20733 & ~n20734 ) | ( n20733 & 1'b0 ) | ( ~n20734 & 1'b0 ) ;
  assign n20744 = ( n192 & n20664 ) | ( n192 & n20735 ) | ( n20664 & n20735 ) ;
  assign n20745 = ( n20664 & ~n20673 ) | ( n20664 & n20735 ) | ( ~n20673 & n20735 ) ;
  assign n20746 = ~n20744 & n20745 ;
  assign n20747 = n20740 | n20746 ;
  assign n20748 = n20589 &  n20674 ;
  assign n20741 = x74 | n20589 ;
  assign n20742 = x74 &  n20589 ;
  assign n20743 = ( n20741 & ~n20742 ) | ( n20741 & 1'b0 ) | ( ~n20742 & 1'b0 ) ;
  assign n20752 = ( n192 & n20663 ) | ( n192 & n20743 ) | ( n20663 & n20743 ) ;
  assign n20753 = ( n20663 & ~n20673 ) | ( n20663 & n20743 ) | ( ~n20673 & n20743 ) ;
  assign n20754 = ~n20752 & n20753 ;
  assign n20755 = n20748 | n20754 ;
  assign n20756 = n20597 &  n20674 ;
  assign n20749 = x73 | n20597 ;
  assign n20750 = x73 &  n20597 ;
  assign n20751 = ( n20749 & ~n20750 ) | ( n20749 & 1'b0 ) | ( ~n20750 & 1'b0 ) ;
  assign n20760 = ( n192 & n20662 ) | ( n192 & n20751 ) | ( n20662 & n20751 ) ;
  assign n20761 = ( n20662 & ~n20673 ) | ( n20662 & n20751 ) | ( ~n20673 & n20751 ) ;
  assign n20762 = ~n20760 & n20761 ;
  assign n20763 = n20756 | n20762 ;
  assign n20764 = n20605 &  n20674 ;
  assign n20757 = x72 | n20605 ;
  assign n20758 = x72 &  n20605 ;
  assign n20759 = ( n20757 & ~n20758 ) | ( n20757 & 1'b0 ) | ( ~n20758 & 1'b0 ) ;
  assign n20768 = ( n192 & n20661 ) | ( n192 & n20759 ) | ( n20661 & n20759 ) ;
  assign n20769 = ( n20661 & ~n20673 ) | ( n20661 & n20759 ) | ( ~n20673 & n20759 ) ;
  assign n20770 = ~n20768 & n20769 ;
  assign n20771 = n20764 | n20770 ;
  assign n20772 = n20613 &  n20674 ;
  assign n20765 = x71 | n20613 ;
  assign n20766 = x71 &  n20613 ;
  assign n20767 = ( n20765 & ~n20766 ) | ( n20765 & 1'b0 ) | ( ~n20766 & 1'b0 ) ;
  assign n20776 = ( n192 & n20660 ) | ( n192 & n20767 ) | ( n20660 & n20767 ) ;
  assign n20777 = ( n20660 & ~n20673 ) | ( n20660 & n20767 ) | ( ~n20673 & n20767 ) ;
  assign n20778 = ~n20776 & n20777 ;
  assign n20779 = n20772 | n20778 ;
  assign n20780 = n20621 &  n20674 ;
  assign n20773 = x70 | n20621 ;
  assign n20774 = x70 &  n20621 ;
  assign n20775 = ( n20773 & ~n20774 ) | ( n20773 & 1'b0 ) | ( ~n20774 & 1'b0 ) ;
  assign n20784 = ( n192 & n20659 ) | ( n192 & n20775 ) | ( n20659 & n20775 ) ;
  assign n20785 = ( n20659 & ~n20673 ) | ( n20659 & n20775 ) | ( ~n20673 & n20775 ) ;
  assign n20786 = ~n20784 & n20785 ;
  assign n20787 = n20780 | n20786 ;
  assign n20788 = n20629 &  n20674 ;
  assign n20781 = x69 | n20629 ;
  assign n20782 = x69 &  n20629 ;
  assign n20783 = ( n20781 & ~n20782 ) | ( n20781 & 1'b0 ) | ( ~n20782 & 1'b0 ) ;
  assign n20792 = ( n192 & n20658 ) | ( n192 & n20783 ) | ( n20658 & n20783 ) ;
  assign n20793 = ( n20658 & ~n20673 ) | ( n20658 & n20783 ) | ( ~n20673 & n20783 ) ;
  assign n20794 = ~n20792 & n20793 ;
  assign n20795 = n20788 | n20794 ;
  assign n20796 = n20637 &  n20674 ;
  assign n20789 = x68 | n20637 ;
  assign n20790 = x68 &  n20637 ;
  assign n20791 = ( n20789 & ~n20790 ) | ( n20789 & 1'b0 ) | ( ~n20790 & 1'b0 ) ;
  assign n20800 = ( n192 & n20657 ) | ( n192 & n20791 ) | ( n20657 & n20791 ) ;
  assign n20801 = ( n20657 & ~n20673 ) | ( n20657 & n20791 ) | ( ~n20673 & n20791 ) ;
  assign n20802 = ~n20800 & n20801 ;
  assign n20803 = n20796 | n20802 ;
  assign n20804 = n20642 &  n20674 ;
  assign n20797 = x67 | n20642 ;
  assign n20798 = x67 &  n20642 ;
  assign n20799 = ( n20797 & ~n20798 ) | ( n20797 & 1'b0 ) | ( ~n20798 & 1'b0 ) ;
  assign n20808 = ( n192 & n20656 ) | ( n192 & n20799 ) | ( n20656 & n20799 ) ;
  assign n20809 = ( n20656 & ~n20673 ) | ( n20656 & n20799 ) | ( ~n20673 & n20799 ) ;
  assign n20810 = ~n20808 & n20809 ;
  assign n20811 = n20804 | n20810 ;
  assign n20812 = n20650 &  n20674 ;
  assign n20805 = x66 | n20650 ;
  assign n20806 = x66 &  n20650 ;
  assign n20807 = ( n20805 & ~n20806 ) | ( n20805 & 1'b0 ) | ( ~n20806 & 1'b0 ) ;
  assign n20816 = ( n192 & n20655 ) | ( n192 & n20807 ) | ( n20655 & n20807 ) ;
  assign n20817 = ( n20655 & ~n20673 ) | ( n20655 & n20807 ) | ( ~n20673 & n20807 ) ;
  assign n20818 = ~n20816 & n20817 ;
  assign n20819 = n20812 | n20818 ;
  assign n20820 = n20654 &  n20674 ;
  assign n20813 = x65 &  n20654 ;
  assign n20814 = x65 | n20653 ;
  assign n20815 = n20652 | n20814 ;
  assign n20821 = ~n20813 & n20815 ;
  assign n20822 = ( n2120 & ~n20673 ) | ( n2120 & n20821 ) | ( ~n20673 & n20821 ) ;
  assign n20823 = ( n192 & n2120 ) | ( n192 & n20821 ) | ( n2120 & n20821 ) ;
  assign n20824 = ( n20822 & ~n20823 ) | ( n20822 & 1'b0 ) | ( ~n20823 & 1'b0 ) ;
  assign n20825 = n20820 | n20824 ;
  assign n20826 = ( n2290 & ~n20673 ) | ( n2290 & 1'b0 ) | ( ~n20673 & 1'b0 ) ;
  assign n20827 = ( x44 & ~n20826 ) | ( x44 & 1'b0 ) | ( ~n20826 & 1'b0 ) ;
  assign n20828 = ( n2296 & ~n20673 ) | ( n2296 & 1'b0 ) | ( ~n20673 & 1'b0 ) ;
  assign n20829 = n20827 | n20828 ;
  assign n20830 = ( x65 & ~n20829 ) | ( x65 & n2299 ) | ( ~n20829 & n2299 ) ;
  assign n20831 = ( x66 & ~n20825 ) | ( x66 & n20830 ) | ( ~n20825 & n20830 ) ;
  assign n20832 = ( x67 & ~n20819 ) | ( x67 & n20831 ) | ( ~n20819 & n20831 ) ;
  assign n20833 = ( x68 & ~n20811 ) | ( x68 & n20832 ) | ( ~n20811 & n20832 ) ;
  assign n20834 = ( x69 & ~n20803 ) | ( x69 & n20833 ) | ( ~n20803 & n20833 ) ;
  assign n20835 = ( x70 & ~n20795 ) | ( x70 & n20834 ) | ( ~n20795 & n20834 ) ;
  assign n20836 = ( x71 & ~n20787 ) | ( x71 & n20835 ) | ( ~n20787 & n20835 ) ;
  assign n20837 = ( x72 & ~n20779 ) | ( x72 & n20836 ) | ( ~n20779 & n20836 ) ;
  assign n20838 = ( x73 & ~n20771 ) | ( x73 & n20837 ) | ( ~n20771 & n20837 ) ;
  assign n20839 = ( x74 & ~n20763 ) | ( x74 & n20838 ) | ( ~n20763 & n20838 ) ;
  assign n20840 = ( x75 & ~n20755 ) | ( x75 & n20839 ) | ( ~n20755 & n20839 ) ;
  assign n20841 = ( x76 & ~n20747 ) | ( x76 & n20840 ) | ( ~n20747 & n20840 ) ;
  assign n20842 = ( x77 & ~n20739 ) | ( x77 & n20841 ) | ( ~n20739 & n20841 ) ;
  assign n20843 = ( x78 & ~n20731 ) | ( x78 & n20842 ) | ( ~n20731 & n20842 ) ;
  assign n20844 = ( x79 & ~n20723 ) | ( x79 & n20843 ) | ( ~n20723 & n20843 ) ;
  assign n20845 = ( x80 & ~n20715 ) | ( x80 & n20844 ) | ( ~n20715 & n20844 ) ;
  assign n20846 = ( x81 & ~n20707 ) | ( x81 & n20845 ) | ( ~n20707 & n20845 ) ;
  assign n20847 = ( x82 & ~n20699 ) | ( x82 & n20846 ) | ( ~n20699 & n20846 ) ;
  assign n20848 = ( x83 & ~n20691 ) | ( x83 & n20847 ) | ( ~n20691 & n20847 ) ;
  assign n20849 = ( x84 & ~n20675 ) | ( x84 & 1'b0 ) | ( ~n20675 & 1'b0 ) ;
  assign n20850 = ~n20681 & n20849 ;
  assign n20851 = ( n20848 & ~n20683 ) | ( n20848 & n20850 ) | ( ~n20683 & n20850 ) ;
  assign n20852 = ( n20683 & ~n462 ) | ( n20683 & n20851 ) | ( ~n462 & n20851 ) ;
  assign n20853 = n462 | n20852 ;
  assign n20860 = n192 &  n20517 ;
  assign n20861 = n20853 &  n20860 ;
  assign n20854 = ~n192 & n20682 ;
  assign n20855 = ( n20853 & ~n20854 ) | ( n20853 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20859 = n20683 | n20850 ;
  assign n20863 = ( n20848 & n20855 ) | ( n20848 & n20859 ) | ( n20855 & n20859 ) ;
  assign n20862 = n20848 | n20859 ;
  assign n20864 = ( n20861 & ~n20863 ) | ( n20861 & n20862 ) | ( ~n20863 & n20862 ) ;
  assign n20868 = ( n20691 & ~n20854 ) | ( n20691 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20869 = n20853 &  n20868 ;
  assign n20856 = x83 | n20691 ;
  assign n20857 = x83 &  n20691 ;
  assign n20858 = ( n20856 & ~n20857 ) | ( n20856 & 1'b0 ) | ( ~n20857 & 1'b0 ) ;
  assign n20871 = ( n20847 & n20855 ) | ( n20847 & n20858 ) | ( n20855 & n20858 ) ;
  assign n20870 = n20847 | n20858 ;
  assign n20872 = ( n20869 & ~n20871 ) | ( n20869 & n20870 ) | ( ~n20871 & n20870 ) ;
  assign n20876 = ( n20699 & ~n20854 ) | ( n20699 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20877 = n20853 &  n20876 ;
  assign n20865 = x82 | n20699 ;
  assign n20866 = x82 &  n20699 ;
  assign n20867 = ( n20865 & ~n20866 ) | ( n20865 & 1'b0 ) | ( ~n20866 & 1'b0 ) ;
  assign n20879 = ( n20846 & n20855 ) | ( n20846 & n20867 ) | ( n20855 & n20867 ) ;
  assign n20878 = n20846 | n20867 ;
  assign n20880 = ( n20877 & ~n20879 ) | ( n20877 & n20878 ) | ( ~n20879 & n20878 ) ;
  assign n20884 = ( n20707 & ~n20854 ) | ( n20707 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20885 = n20853 &  n20884 ;
  assign n20873 = x81 | n20707 ;
  assign n20874 = x81 &  n20707 ;
  assign n20875 = ( n20873 & ~n20874 ) | ( n20873 & 1'b0 ) | ( ~n20874 & 1'b0 ) ;
  assign n20887 = ( n20845 & n20855 ) | ( n20845 & n20875 ) | ( n20855 & n20875 ) ;
  assign n20886 = n20845 | n20875 ;
  assign n20888 = ( n20885 & ~n20887 ) | ( n20885 & n20886 ) | ( ~n20887 & n20886 ) ;
  assign n20892 = ( n20715 & ~n20854 ) | ( n20715 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20893 = n20853 &  n20892 ;
  assign n20881 = x80 | n20715 ;
  assign n20882 = x80 &  n20715 ;
  assign n20883 = ( n20881 & ~n20882 ) | ( n20881 & 1'b0 ) | ( ~n20882 & 1'b0 ) ;
  assign n20895 = ( n20844 & n20855 ) | ( n20844 & n20883 ) | ( n20855 & n20883 ) ;
  assign n20894 = n20844 | n20883 ;
  assign n20896 = ( n20893 & ~n20895 ) | ( n20893 & n20894 ) | ( ~n20895 & n20894 ) ;
  assign n20900 = ( n20723 & ~n20854 ) | ( n20723 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20901 = n20853 &  n20900 ;
  assign n20889 = x79 | n20723 ;
  assign n20890 = x79 &  n20723 ;
  assign n20891 = ( n20889 & ~n20890 ) | ( n20889 & 1'b0 ) | ( ~n20890 & 1'b0 ) ;
  assign n20903 = ( n20843 & n20855 ) | ( n20843 & n20891 ) | ( n20855 & n20891 ) ;
  assign n20902 = n20843 | n20891 ;
  assign n20904 = ( n20901 & ~n20903 ) | ( n20901 & n20902 ) | ( ~n20903 & n20902 ) ;
  assign n20908 = ( n20731 & ~n20854 ) | ( n20731 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20909 = n20853 &  n20908 ;
  assign n20897 = x78 | n20731 ;
  assign n20898 = x78 &  n20731 ;
  assign n20899 = ( n20897 & ~n20898 ) | ( n20897 & 1'b0 ) | ( ~n20898 & 1'b0 ) ;
  assign n20911 = ( n20842 & n20855 ) | ( n20842 & n20899 ) | ( n20855 & n20899 ) ;
  assign n20910 = n20842 | n20899 ;
  assign n20912 = ( n20909 & ~n20911 ) | ( n20909 & n20910 ) | ( ~n20911 & n20910 ) ;
  assign n20916 = ( n20739 & ~n20854 ) | ( n20739 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20917 = n20853 &  n20916 ;
  assign n20905 = x77 | n20739 ;
  assign n20906 = x77 &  n20739 ;
  assign n20907 = ( n20905 & ~n20906 ) | ( n20905 & 1'b0 ) | ( ~n20906 & 1'b0 ) ;
  assign n20919 = ( n20841 & n20855 ) | ( n20841 & n20907 ) | ( n20855 & n20907 ) ;
  assign n20918 = n20841 | n20907 ;
  assign n20920 = ( n20917 & ~n20919 ) | ( n20917 & n20918 ) | ( ~n20919 & n20918 ) ;
  assign n20924 = ( n20747 & ~n20854 ) | ( n20747 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20925 = n20853 &  n20924 ;
  assign n20913 = x76 | n20747 ;
  assign n20914 = x76 &  n20747 ;
  assign n20915 = ( n20913 & ~n20914 ) | ( n20913 & 1'b0 ) | ( ~n20914 & 1'b0 ) ;
  assign n20927 = ( n20840 & n20855 ) | ( n20840 & n20915 ) | ( n20855 & n20915 ) ;
  assign n20926 = n20840 | n20915 ;
  assign n20928 = ( n20925 & ~n20927 ) | ( n20925 & n20926 ) | ( ~n20927 & n20926 ) ;
  assign n20932 = ( n20755 & ~n20854 ) | ( n20755 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20933 = n20853 &  n20932 ;
  assign n20921 = x75 | n20755 ;
  assign n20922 = x75 &  n20755 ;
  assign n20923 = ( n20921 & ~n20922 ) | ( n20921 & 1'b0 ) | ( ~n20922 & 1'b0 ) ;
  assign n20935 = ( n20839 & n20855 ) | ( n20839 & n20923 ) | ( n20855 & n20923 ) ;
  assign n20934 = n20839 | n20923 ;
  assign n20936 = ( n20933 & ~n20935 ) | ( n20933 & n20934 ) | ( ~n20935 & n20934 ) ;
  assign n20940 = ( n20763 & ~n20854 ) | ( n20763 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20941 = n20853 &  n20940 ;
  assign n20929 = x74 | n20763 ;
  assign n20930 = x74 &  n20763 ;
  assign n20931 = ( n20929 & ~n20930 ) | ( n20929 & 1'b0 ) | ( ~n20930 & 1'b0 ) ;
  assign n20943 = ( n20838 & n20855 ) | ( n20838 & n20931 ) | ( n20855 & n20931 ) ;
  assign n20942 = n20838 | n20931 ;
  assign n20944 = ( n20941 & ~n20943 ) | ( n20941 & n20942 ) | ( ~n20943 & n20942 ) ;
  assign n20948 = ( n20771 & ~n20854 ) | ( n20771 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20949 = n20853 &  n20948 ;
  assign n20937 = x73 | n20771 ;
  assign n20938 = x73 &  n20771 ;
  assign n20939 = ( n20937 & ~n20938 ) | ( n20937 & 1'b0 ) | ( ~n20938 & 1'b0 ) ;
  assign n20951 = ( n20837 & n20855 ) | ( n20837 & n20939 ) | ( n20855 & n20939 ) ;
  assign n20950 = n20837 | n20939 ;
  assign n20952 = ( n20949 & ~n20951 ) | ( n20949 & n20950 ) | ( ~n20951 & n20950 ) ;
  assign n20956 = ( n20779 & ~n20854 ) | ( n20779 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20957 = n20853 &  n20956 ;
  assign n20945 = x72 | n20779 ;
  assign n20946 = x72 &  n20779 ;
  assign n20947 = ( n20945 & ~n20946 ) | ( n20945 & 1'b0 ) | ( ~n20946 & 1'b0 ) ;
  assign n20959 = ( n20836 & n20855 ) | ( n20836 & n20947 ) | ( n20855 & n20947 ) ;
  assign n20958 = n20836 | n20947 ;
  assign n20960 = ( n20957 & ~n20959 ) | ( n20957 & n20958 ) | ( ~n20959 & n20958 ) ;
  assign n20964 = ( n20787 & ~n20854 ) | ( n20787 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20965 = n20853 &  n20964 ;
  assign n20953 = x71 | n20787 ;
  assign n20954 = x71 &  n20787 ;
  assign n20955 = ( n20953 & ~n20954 ) | ( n20953 & 1'b0 ) | ( ~n20954 & 1'b0 ) ;
  assign n20967 = ( n20835 & n20855 ) | ( n20835 & n20955 ) | ( n20855 & n20955 ) ;
  assign n20966 = n20835 | n20955 ;
  assign n20968 = ( n20965 & ~n20967 ) | ( n20965 & n20966 ) | ( ~n20967 & n20966 ) ;
  assign n20972 = ( n20795 & ~n20854 ) | ( n20795 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20973 = n20853 &  n20972 ;
  assign n20961 = x70 | n20795 ;
  assign n20962 = x70 &  n20795 ;
  assign n20963 = ( n20961 & ~n20962 ) | ( n20961 & 1'b0 ) | ( ~n20962 & 1'b0 ) ;
  assign n20975 = ( n20834 & n20855 ) | ( n20834 & n20963 ) | ( n20855 & n20963 ) ;
  assign n20974 = n20834 | n20963 ;
  assign n20976 = ( n20973 & ~n20975 ) | ( n20973 & n20974 ) | ( ~n20975 & n20974 ) ;
  assign n20980 = ( n20803 & ~n20854 ) | ( n20803 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20981 = n20853 &  n20980 ;
  assign n20969 = x69 | n20803 ;
  assign n20970 = x69 &  n20803 ;
  assign n20971 = ( n20969 & ~n20970 ) | ( n20969 & 1'b0 ) | ( ~n20970 & 1'b0 ) ;
  assign n20983 = ( n20833 & n20855 ) | ( n20833 & n20971 ) | ( n20855 & n20971 ) ;
  assign n20982 = n20833 | n20971 ;
  assign n20984 = ( n20981 & ~n20983 ) | ( n20981 & n20982 ) | ( ~n20983 & n20982 ) ;
  assign n20988 = ( n20811 & ~n20854 ) | ( n20811 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20989 = n20853 &  n20988 ;
  assign n20977 = x68 | n20811 ;
  assign n20978 = x68 &  n20811 ;
  assign n20979 = ( n20977 & ~n20978 ) | ( n20977 & 1'b0 ) | ( ~n20978 & 1'b0 ) ;
  assign n20991 = ( n20832 & n20855 ) | ( n20832 & n20979 ) | ( n20855 & n20979 ) ;
  assign n20990 = n20832 | n20979 ;
  assign n20992 = ( n20989 & ~n20991 ) | ( n20989 & n20990 ) | ( ~n20991 & n20990 ) ;
  assign n20996 = ( n20819 & ~n20854 ) | ( n20819 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n20997 = n20853 &  n20996 ;
  assign n20985 = x67 | n20819 ;
  assign n20986 = x67 &  n20819 ;
  assign n20987 = ( n20985 & ~n20986 ) | ( n20985 & 1'b0 ) | ( ~n20986 & 1'b0 ) ;
  assign n20999 = ( n20831 & n20855 ) | ( n20831 & n20987 ) | ( n20855 & n20987 ) ;
  assign n20998 = n20831 | n20987 ;
  assign n21000 = ( n20997 & ~n20999 ) | ( n20997 & n20998 ) | ( ~n20999 & n20998 ) ;
  assign n21001 = ( n20825 & ~n20854 ) | ( n20825 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n21002 = n20853 &  n21001 ;
  assign n20993 = x66 | n20825 ;
  assign n20994 = x66 &  n20825 ;
  assign n20995 = ( n20993 & ~n20994 ) | ( n20993 & 1'b0 ) | ( ~n20994 & 1'b0 ) ;
  assign n21004 = ( n20830 & n20855 ) | ( n20830 & n20995 ) | ( n20855 & n20995 ) ;
  assign n21003 = n20830 | n20995 ;
  assign n21005 = ( n21002 & ~n21004 ) | ( n21002 & n21003 ) | ( ~n21004 & n21003 ) ;
  assign n21006 = ( x65 & ~n2299 ) | ( x65 & n20829 ) | ( ~n2299 & n20829 ) ;
  assign n21007 = ( n20830 & ~x65 ) | ( n20830 & n21006 ) | ( ~x65 & n21006 ) ;
  assign n21008 = ~n20855 & n21007 ;
  assign n21009 = ( n20829 & ~n20854 ) | ( n20829 & 1'b0 ) | ( ~n20854 & 1'b0 ) ;
  assign n21010 = n20853 &  n21009 ;
  assign n21011 = n21008 | n21010 ;
  assign n21012 = ( x64 & ~n20855 ) | ( x64 & 1'b0 ) | ( ~n20855 & 1'b0 ) ;
  assign n21013 = ( x43 & ~n21012 ) | ( x43 & 1'b0 ) | ( ~n21012 & 1'b0 ) ;
  assign n21014 = ( n2299 & ~n20855 ) | ( n2299 & 1'b0 ) | ( ~n20855 & 1'b0 ) ;
  assign n21015 = n21013 | n21014 ;
  assign n21016 = ( x65 & ~n21015 ) | ( x65 & n2492 ) | ( ~n21015 & n2492 ) ;
  assign n21017 = ( x66 & ~n21011 ) | ( x66 & n21016 ) | ( ~n21011 & n21016 ) ;
  assign n21018 = ( x67 & ~n21005 ) | ( x67 & n21017 ) | ( ~n21005 & n21017 ) ;
  assign n21019 = ( x68 & ~n21000 ) | ( x68 & n21018 ) | ( ~n21000 & n21018 ) ;
  assign n21020 = ( x69 & ~n20992 ) | ( x69 & n21019 ) | ( ~n20992 & n21019 ) ;
  assign n21021 = ( x70 & ~n20984 ) | ( x70 & n21020 ) | ( ~n20984 & n21020 ) ;
  assign n21022 = ( x71 & ~n20976 ) | ( x71 & n21021 ) | ( ~n20976 & n21021 ) ;
  assign n21023 = ( x72 & ~n20968 ) | ( x72 & n21022 ) | ( ~n20968 & n21022 ) ;
  assign n21024 = ( x73 & ~n20960 ) | ( x73 & n21023 ) | ( ~n20960 & n21023 ) ;
  assign n21025 = ( x74 & ~n20952 ) | ( x74 & n21024 ) | ( ~n20952 & n21024 ) ;
  assign n21026 = ( x75 & ~n20944 ) | ( x75 & n21025 ) | ( ~n20944 & n21025 ) ;
  assign n21027 = ( x76 & ~n20936 ) | ( x76 & n21026 ) | ( ~n20936 & n21026 ) ;
  assign n21028 = ( x77 & ~n20928 ) | ( x77 & n21027 ) | ( ~n20928 & n21027 ) ;
  assign n21029 = ( x78 & ~n20920 ) | ( x78 & n21028 ) | ( ~n20920 & n21028 ) ;
  assign n21030 = ( x79 & ~n20912 ) | ( x79 & n21029 ) | ( ~n20912 & n21029 ) ;
  assign n21031 = ( x80 & ~n20904 ) | ( x80 & n21030 ) | ( ~n20904 & n21030 ) ;
  assign n21032 = ( x81 & ~n20896 ) | ( x81 & n21031 ) | ( ~n20896 & n21031 ) ;
  assign n21033 = ( x82 & ~n20888 ) | ( x82 & n21032 ) | ( ~n20888 & n21032 ) ;
  assign n21034 = ( x83 & ~n20880 ) | ( x83 & n21033 ) | ( ~n20880 & n21033 ) ;
  assign n21035 = ( x84 & ~n20872 ) | ( x84 & n21034 ) | ( ~n20872 & n21034 ) ;
  assign n21042 = ( x85 & ~n2517 ) | ( x85 & n21035 ) | ( ~n2517 & n21035 ) ;
  assign n21041 = x85 &  n21035 ;
  assign n21043 = ( n20864 & ~n21042 ) | ( n20864 & n21041 ) | ( ~n21042 & n21041 ) ;
  assign n21036 = ( x85 & ~n20864 ) | ( x85 & n21035 ) | ( ~n20864 & n21035 ) ;
  assign n21037 = n2517 | n21036 ;
  assign n21044 = n20872 &  n21037 ;
  assign n21038 = x84 | n20872 ;
  assign n21039 = x84 &  n20872 ;
  assign n21040 = ( n21038 & ~n21039 ) | ( n21038 & 1'b0 ) | ( ~n21039 & 1'b0 ) ;
  assign n21048 = ( n2517 & n21034 ) | ( n2517 & n21040 ) | ( n21034 & n21040 ) ;
  assign n21049 = ( n21034 & ~n21036 ) | ( n21034 & n21040 ) | ( ~n21036 & n21040 ) ;
  assign n21050 = ~n21048 & n21049 ;
  assign n21051 = n21044 | n21050 ;
  assign n21052 = n20880 &  n21037 ;
  assign n21045 = x83 | n20880 ;
  assign n21046 = x83 &  n20880 ;
  assign n21047 = ( n21045 & ~n21046 ) | ( n21045 & 1'b0 ) | ( ~n21046 & 1'b0 ) ;
  assign n21056 = ( n2517 & n21033 ) | ( n2517 & n21047 ) | ( n21033 & n21047 ) ;
  assign n21057 = ( n21033 & ~n21036 ) | ( n21033 & n21047 ) | ( ~n21036 & n21047 ) ;
  assign n21058 = ~n21056 & n21057 ;
  assign n21059 = n21052 | n21058 ;
  assign n21060 = n20888 &  n21037 ;
  assign n21053 = x82 | n20888 ;
  assign n21054 = x82 &  n20888 ;
  assign n21055 = ( n21053 & ~n21054 ) | ( n21053 & 1'b0 ) | ( ~n21054 & 1'b0 ) ;
  assign n21064 = ( n2517 & n21032 ) | ( n2517 & n21055 ) | ( n21032 & n21055 ) ;
  assign n21065 = ( n21032 & ~n21036 ) | ( n21032 & n21055 ) | ( ~n21036 & n21055 ) ;
  assign n21066 = ~n21064 & n21065 ;
  assign n21067 = n21060 | n21066 ;
  assign n21068 = n20896 &  n21037 ;
  assign n21061 = x81 | n20896 ;
  assign n21062 = x81 &  n20896 ;
  assign n21063 = ( n21061 & ~n21062 ) | ( n21061 & 1'b0 ) | ( ~n21062 & 1'b0 ) ;
  assign n21072 = ( n2517 & n21031 ) | ( n2517 & n21063 ) | ( n21031 & n21063 ) ;
  assign n21073 = ( n21031 & ~n21036 ) | ( n21031 & n21063 ) | ( ~n21036 & n21063 ) ;
  assign n21074 = ~n21072 & n21073 ;
  assign n21075 = n21068 | n21074 ;
  assign n21076 = n20904 &  n21037 ;
  assign n21069 = x80 | n20904 ;
  assign n21070 = x80 &  n20904 ;
  assign n21071 = ( n21069 & ~n21070 ) | ( n21069 & 1'b0 ) | ( ~n21070 & 1'b0 ) ;
  assign n21080 = ( n2517 & n21030 ) | ( n2517 & n21071 ) | ( n21030 & n21071 ) ;
  assign n21081 = ( n21030 & ~n21036 ) | ( n21030 & n21071 ) | ( ~n21036 & n21071 ) ;
  assign n21082 = ~n21080 & n21081 ;
  assign n21083 = n21076 | n21082 ;
  assign n21084 = n20912 &  n21037 ;
  assign n21077 = x79 | n20912 ;
  assign n21078 = x79 &  n20912 ;
  assign n21079 = ( n21077 & ~n21078 ) | ( n21077 & 1'b0 ) | ( ~n21078 & 1'b0 ) ;
  assign n21088 = ( n2517 & n21029 ) | ( n2517 & n21079 ) | ( n21029 & n21079 ) ;
  assign n21089 = ( n21029 & ~n21036 ) | ( n21029 & n21079 ) | ( ~n21036 & n21079 ) ;
  assign n21090 = ~n21088 & n21089 ;
  assign n21091 = n21084 | n21090 ;
  assign n21092 = n20920 &  n21037 ;
  assign n21085 = x78 | n20920 ;
  assign n21086 = x78 &  n20920 ;
  assign n21087 = ( n21085 & ~n21086 ) | ( n21085 & 1'b0 ) | ( ~n21086 & 1'b0 ) ;
  assign n21096 = ( n2517 & n21028 ) | ( n2517 & n21087 ) | ( n21028 & n21087 ) ;
  assign n21097 = ( n21028 & ~n21036 ) | ( n21028 & n21087 ) | ( ~n21036 & n21087 ) ;
  assign n21098 = ~n21096 & n21097 ;
  assign n21099 = n21092 | n21098 ;
  assign n21100 = n20928 &  n21037 ;
  assign n21093 = x77 | n20928 ;
  assign n21094 = x77 &  n20928 ;
  assign n21095 = ( n21093 & ~n21094 ) | ( n21093 & 1'b0 ) | ( ~n21094 & 1'b0 ) ;
  assign n21104 = ( n2517 & n21027 ) | ( n2517 & n21095 ) | ( n21027 & n21095 ) ;
  assign n21105 = ( n21027 & ~n21036 ) | ( n21027 & n21095 ) | ( ~n21036 & n21095 ) ;
  assign n21106 = ~n21104 & n21105 ;
  assign n21107 = n21100 | n21106 ;
  assign n21108 = n20936 &  n21037 ;
  assign n21101 = x76 | n20936 ;
  assign n21102 = x76 &  n20936 ;
  assign n21103 = ( n21101 & ~n21102 ) | ( n21101 & 1'b0 ) | ( ~n21102 & 1'b0 ) ;
  assign n21112 = ( n2517 & n21026 ) | ( n2517 & n21103 ) | ( n21026 & n21103 ) ;
  assign n21113 = ( n21026 & ~n21036 ) | ( n21026 & n21103 ) | ( ~n21036 & n21103 ) ;
  assign n21114 = ~n21112 & n21113 ;
  assign n21115 = n21108 | n21114 ;
  assign n21116 = n20944 &  n21037 ;
  assign n21109 = x75 | n20944 ;
  assign n21110 = x75 &  n20944 ;
  assign n21111 = ( n21109 & ~n21110 ) | ( n21109 & 1'b0 ) | ( ~n21110 & 1'b0 ) ;
  assign n21120 = ( n2517 & n21025 ) | ( n2517 & n21111 ) | ( n21025 & n21111 ) ;
  assign n21121 = ( n21025 & ~n21036 ) | ( n21025 & n21111 ) | ( ~n21036 & n21111 ) ;
  assign n21122 = ~n21120 & n21121 ;
  assign n21123 = n21116 | n21122 ;
  assign n21124 = n20952 &  n21037 ;
  assign n21117 = x74 | n20952 ;
  assign n21118 = x74 &  n20952 ;
  assign n21119 = ( n21117 & ~n21118 ) | ( n21117 & 1'b0 ) | ( ~n21118 & 1'b0 ) ;
  assign n21128 = ( n2517 & n21024 ) | ( n2517 & n21119 ) | ( n21024 & n21119 ) ;
  assign n21129 = ( n21024 & ~n21036 ) | ( n21024 & n21119 ) | ( ~n21036 & n21119 ) ;
  assign n21130 = ~n21128 & n21129 ;
  assign n21131 = n21124 | n21130 ;
  assign n21132 = n20960 &  n21037 ;
  assign n21125 = x73 | n20960 ;
  assign n21126 = x73 &  n20960 ;
  assign n21127 = ( n21125 & ~n21126 ) | ( n21125 & 1'b0 ) | ( ~n21126 & 1'b0 ) ;
  assign n21136 = ( n2517 & n21023 ) | ( n2517 & n21127 ) | ( n21023 & n21127 ) ;
  assign n21137 = ( n21023 & ~n21036 ) | ( n21023 & n21127 ) | ( ~n21036 & n21127 ) ;
  assign n21138 = ~n21136 & n21137 ;
  assign n21139 = n21132 | n21138 ;
  assign n21140 = n20968 &  n21037 ;
  assign n21133 = x72 | n20968 ;
  assign n21134 = x72 &  n20968 ;
  assign n21135 = ( n21133 & ~n21134 ) | ( n21133 & 1'b0 ) | ( ~n21134 & 1'b0 ) ;
  assign n21144 = ( n2517 & n21022 ) | ( n2517 & n21135 ) | ( n21022 & n21135 ) ;
  assign n21145 = ( n21022 & ~n21036 ) | ( n21022 & n21135 ) | ( ~n21036 & n21135 ) ;
  assign n21146 = ~n21144 & n21145 ;
  assign n21147 = n21140 | n21146 ;
  assign n21148 = n20976 &  n21037 ;
  assign n21141 = x71 | n20976 ;
  assign n21142 = x71 &  n20976 ;
  assign n21143 = ( n21141 & ~n21142 ) | ( n21141 & 1'b0 ) | ( ~n21142 & 1'b0 ) ;
  assign n21152 = ( n2517 & n21021 ) | ( n2517 & n21143 ) | ( n21021 & n21143 ) ;
  assign n21153 = ( n21021 & ~n21036 ) | ( n21021 & n21143 ) | ( ~n21036 & n21143 ) ;
  assign n21154 = ~n21152 & n21153 ;
  assign n21155 = n21148 | n21154 ;
  assign n21156 = n20984 &  n21037 ;
  assign n21149 = x70 | n20984 ;
  assign n21150 = x70 &  n20984 ;
  assign n21151 = ( n21149 & ~n21150 ) | ( n21149 & 1'b0 ) | ( ~n21150 & 1'b0 ) ;
  assign n21160 = ( n2517 & n21020 ) | ( n2517 & n21151 ) | ( n21020 & n21151 ) ;
  assign n21161 = ( n21020 & ~n21036 ) | ( n21020 & n21151 ) | ( ~n21036 & n21151 ) ;
  assign n21162 = ~n21160 & n21161 ;
  assign n21163 = n21156 | n21162 ;
  assign n21164 = n20992 &  n21037 ;
  assign n21157 = x69 | n20992 ;
  assign n21158 = x69 &  n20992 ;
  assign n21159 = ( n21157 & ~n21158 ) | ( n21157 & 1'b0 ) | ( ~n21158 & 1'b0 ) ;
  assign n21168 = ( n2517 & n21019 ) | ( n2517 & n21159 ) | ( n21019 & n21159 ) ;
  assign n21169 = ( n21019 & ~n21036 ) | ( n21019 & n21159 ) | ( ~n21036 & n21159 ) ;
  assign n21170 = ~n21168 & n21169 ;
  assign n21171 = n21164 | n21170 ;
  assign n21172 = n21000 &  n21037 ;
  assign n21165 = x68 | n21000 ;
  assign n21166 = x68 &  n21000 ;
  assign n21167 = ( n21165 & ~n21166 ) | ( n21165 & 1'b0 ) | ( ~n21166 & 1'b0 ) ;
  assign n21176 = ( n2517 & n21018 ) | ( n2517 & n21167 ) | ( n21018 & n21167 ) ;
  assign n21177 = ( n21018 & ~n21036 ) | ( n21018 & n21167 ) | ( ~n21036 & n21167 ) ;
  assign n21178 = ~n21176 & n21177 ;
  assign n21179 = n21172 | n21178 ;
  assign n21180 = n21005 &  n21037 ;
  assign n21173 = x67 | n21005 ;
  assign n21174 = x67 &  n21005 ;
  assign n21175 = ( n21173 & ~n21174 ) | ( n21173 & 1'b0 ) | ( ~n21174 & 1'b0 ) ;
  assign n21184 = ( n2517 & n21017 ) | ( n2517 & n21175 ) | ( n21017 & n21175 ) ;
  assign n21185 = ( n21017 & ~n21036 ) | ( n21017 & n21175 ) | ( ~n21036 & n21175 ) ;
  assign n21186 = ~n21184 & n21185 ;
  assign n21187 = n21180 | n21186 ;
  assign n21188 = n21011 &  n21037 ;
  assign n21181 = x66 | n21011 ;
  assign n21182 = x66 &  n21011 ;
  assign n21183 = ( n21181 & ~n21182 ) | ( n21181 & 1'b0 ) | ( ~n21182 & 1'b0 ) ;
  assign n21189 = ( n2517 & n21016 ) | ( n2517 & n21183 ) | ( n21016 & n21183 ) ;
  assign n21190 = ( n21016 & ~n21036 ) | ( n21016 & n21183 ) | ( ~n21036 & n21183 ) ;
  assign n21191 = ~n21189 & n21190 ;
  assign n21192 = n21188 | n21191 ;
  assign n21193 = n21015 &  n21037 ;
  assign n21194 = ( x65 & ~x43 ) | ( x65 & n21012 ) | ( ~x43 & n21012 ) ;
  assign n21195 = ( x43 & ~n21012 ) | ( x43 & x65 ) | ( ~n21012 & x65 ) ;
  assign n21196 = ( n21194 & ~x65 ) | ( n21194 & n21195 ) | ( ~x65 & n21195 ) ;
  assign n21197 = ( n2492 & ~n2517 ) | ( n2492 & n21196 ) | ( ~n2517 & n21196 ) ;
  assign n21198 = ( n2492 & n21036 ) | ( n2492 & n21196 ) | ( n21036 & n21196 ) ;
  assign n21199 = ( n21197 & ~n21198 ) | ( n21197 & 1'b0 ) | ( ~n21198 & 1'b0 ) ;
  assign n21200 = n21193 | n21199 ;
  assign n21201 = ( n2689 & ~n21036 ) | ( n2689 & 1'b0 ) | ( ~n21036 & 1'b0 ) ;
  assign n21202 = ( x42 & ~n21201 ) | ( x42 & 1'b0 ) | ( ~n21201 & 1'b0 ) ;
  assign n21203 = ( n2696 & ~n21036 ) | ( n2696 & 1'b0 ) | ( ~n21036 & 1'b0 ) ;
  assign n21204 = n21202 | n21203 ;
  assign n21205 = ( x65 & ~n21204 ) | ( x65 & n2699 ) | ( ~n21204 & n2699 ) ;
  assign n21206 = ( x66 & ~n21200 ) | ( x66 & n21205 ) | ( ~n21200 & n21205 ) ;
  assign n21207 = ( x67 & ~n21192 ) | ( x67 & n21206 ) | ( ~n21192 & n21206 ) ;
  assign n21208 = ( x68 & ~n21187 ) | ( x68 & n21207 ) | ( ~n21187 & n21207 ) ;
  assign n21209 = ( x69 & ~n21179 ) | ( x69 & n21208 ) | ( ~n21179 & n21208 ) ;
  assign n21210 = ( x70 & ~n21171 ) | ( x70 & n21209 ) | ( ~n21171 & n21209 ) ;
  assign n21211 = ( x71 & ~n21163 ) | ( x71 & n21210 ) | ( ~n21163 & n21210 ) ;
  assign n21212 = ( x72 & ~n21155 ) | ( x72 & n21211 ) | ( ~n21155 & n21211 ) ;
  assign n21213 = ( x73 & ~n21147 ) | ( x73 & n21212 ) | ( ~n21147 & n21212 ) ;
  assign n21214 = ( x74 & ~n21139 ) | ( x74 & n21213 ) | ( ~n21139 & n21213 ) ;
  assign n21215 = ( x75 & ~n21131 ) | ( x75 & n21214 ) | ( ~n21131 & n21214 ) ;
  assign n21216 = ( x76 & ~n21123 ) | ( x76 & n21215 ) | ( ~n21123 & n21215 ) ;
  assign n21217 = ( x77 & ~n21115 ) | ( x77 & n21216 ) | ( ~n21115 & n21216 ) ;
  assign n21218 = ( x78 & ~n21107 ) | ( x78 & n21217 ) | ( ~n21107 & n21217 ) ;
  assign n21219 = ( x79 & ~n21099 ) | ( x79 & n21218 ) | ( ~n21099 & n21218 ) ;
  assign n21220 = ( x80 & ~n21091 ) | ( x80 & n21219 ) | ( ~n21091 & n21219 ) ;
  assign n21221 = ( x81 & ~n21083 ) | ( x81 & n21220 ) | ( ~n21083 & n21220 ) ;
  assign n21222 = ( x82 & ~n21075 ) | ( x82 & n21221 ) | ( ~n21075 & n21221 ) ;
  assign n21223 = ( x83 & ~n21067 ) | ( x83 & n21222 ) | ( ~n21067 & n21222 ) ;
  assign n21224 = ( x84 & ~n21059 ) | ( x84 & n21223 ) | ( ~n21059 & n21223 ) ;
  assign n21225 = ( x85 & ~n21051 ) | ( x85 & n21224 ) | ( ~n21051 & n21224 ) ;
  assign n21226 = ( x86 & ~n21043 ) | ( x86 & n21225 ) | ( ~n21043 & n21225 ) ;
  assign n21227 = n2741 | n21226 ;
  assign n21228 = n21043 &  n21227 ;
  assign n21232 = ( n2741 & n21043 ) | ( n2741 & n21225 ) | ( n21043 & n21225 ) ;
  assign n21233 = ( x86 & ~n21232 ) | ( x86 & n21043 ) | ( ~n21232 & n21043 ) ;
  assign n21234 = ~x86 & n21233 ;
  assign n21235 = n21228 | n21234 ;
  assign n21236 = ~x87 & n21235 ;
  assign n21237 = n21051 &  n21227 ;
  assign n21229 = x85 | n21051 ;
  assign n21230 = x85 &  n21051 ;
  assign n21231 = ( n21229 & ~n21230 ) | ( n21229 & 1'b0 ) | ( ~n21230 & 1'b0 ) ;
  assign n21241 = ( n2741 & n21224 ) | ( n2741 & n21231 ) | ( n21224 & n21231 ) ;
  assign n21242 = ( n21224 & ~n21226 ) | ( n21224 & n21231 ) | ( ~n21226 & n21231 ) ;
  assign n21243 = ~n21241 & n21242 ;
  assign n21244 = n21237 | n21243 ;
  assign n21245 = n21059 &  n21227 ;
  assign n21238 = x84 | n21059 ;
  assign n21239 = x84 &  n21059 ;
  assign n21240 = ( n21238 & ~n21239 ) | ( n21238 & 1'b0 ) | ( ~n21239 & 1'b0 ) ;
  assign n21249 = ( n2741 & n21223 ) | ( n2741 & n21240 ) | ( n21223 & n21240 ) ;
  assign n21250 = ( n21223 & ~n21226 ) | ( n21223 & n21240 ) | ( ~n21226 & n21240 ) ;
  assign n21251 = ~n21249 & n21250 ;
  assign n21252 = n21245 | n21251 ;
  assign n21253 = n21067 &  n21227 ;
  assign n21246 = x83 | n21067 ;
  assign n21247 = x83 &  n21067 ;
  assign n21248 = ( n21246 & ~n21247 ) | ( n21246 & 1'b0 ) | ( ~n21247 & 1'b0 ) ;
  assign n21257 = ( n2741 & n21222 ) | ( n2741 & n21248 ) | ( n21222 & n21248 ) ;
  assign n21258 = ( n21222 & ~n21226 ) | ( n21222 & n21248 ) | ( ~n21226 & n21248 ) ;
  assign n21259 = ~n21257 & n21258 ;
  assign n21260 = n21253 | n21259 ;
  assign n21261 = n21075 &  n21227 ;
  assign n21254 = x82 | n21075 ;
  assign n21255 = x82 &  n21075 ;
  assign n21256 = ( n21254 & ~n21255 ) | ( n21254 & 1'b0 ) | ( ~n21255 & 1'b0 ) ;
  assign n21265 = ( n2741 & n21221 ) | ( n2741 & n21256 ) | ( n21221 & n21256 ) ;
  assign n21266 = ( n21221 & ~n21226 ) | ( n21221 & n21256 ) | ( ~n21226 & n21256 ) ;
  assign n21267 = ~n21265 & n21266 ;
  assign n21268 = n21261 | n21267 ;
  assign n21269 = n21083 &  n21227 ;
  assign n21262 = x81 | n21083 ;
  assign n21263 = x81 &  n21083 ;
  assign n21264 = ( n21262 & ~n21263 ) | ( n21262 & 1'b0 ) | ( ~n21263 & 1'b0 ) ;
  assign n21273 = ( n2741 & n21220 ) | ( n2741 & n21264 ) | ( n21220 & n21264 ) ;
  assign n21274 = ( n21220 & ~n21226 ) | ( n21220 & n21264 ) | ( ~n21226 & n21264 ) ;
  assign n21275 = ~n21273 & n21274 ;
  assign n21276 = n21269 | n21275 ;
  assign n21277 = n21091 &  n21227 ;
  assign n21270 = x80 | n21091 ;
  assign n21271 = x80 &  n21091 ;
  assign n21272 = ( n21270 & ~n21271 ) | ( n21270 & 1'b0 ) | ( ~n21271 & 1'b0 ) ;
  assign n21281 = ( n2741 & n21219 ) | ( n2741 & n21272 ) | ( n21219 & n21272 ) ;
  assign n21282 = ( n21219 & ~n21226 ) | ( n21219 & n21272 ) | ( ~n21226 & n21272 ) ;
  assign n21283 = ~n21281 & n21282 ;
  assign n21284 = n21277 | n21283 ;
  assign n21285 = n21099 &  n21227 ;
  assign n21278 = x79 | n21099 ;
  assign n21279 = x79 &  n21099 ;
  assign n21280 = ( n21278 & ~n21279 ) | ( n21278 & 1'b0 ) | ( ~n21279 & 1'b0 ) ;
  assign n21289 = ( n2741 & n21218 ) | ( n2741 & n21280 ) | ( n21218 & n21280 ) ;
  assign n21290 = ( n21218 & ~n21226 ) | ( n21218 & n21280 ) | ( ~n21226 & n21280 ) ;
  assign n21291 = ~n21289 & n21290 ;
  assign n21292 = n21285 | n21291 ;
  assign n21293 = n21107 &  n21227 ;
  assign n21286 = x78 | n21107 ;
  assign n21287 = x78 &  n21107 ;
  assign n21288 = ( n21286 & ~n21287 ) | ( n21286 & 1'b0 ) | ( ~n21287 & 1'b0 ) ;
  assign n21297 = ( n2741 & n21217 ) | ( n2741 & n21288 ) | ( n21217 & n21288 ) ;
  assign n21298 = ( n21217 & ~n21226 ) | ( n21217 & n21288 ) | ( ~n21226 & n21288 ) ;
  assign n21299 = ~n21297 & n21298 ;
  assign n21300 = n21293 | n21299 ;
  assign n21301 = n21115 &  n21227 ;
  assign n21294 = x77 | n21115 ;
  assign n21295 = x77 &  n21115 ;
  assign n21296 = ( n21294 & ~n21295 ) | ( n21294 & 1'b0 ) | ( ~n21295 & 1'b0 ) ;
  assign n21305 = ( n2741 & n21216 ) | ( n2741 & n21296 ) | ( n21216 & n21296 ) ;
  assign n21306 = ( n21216 & ~n21226 ) | ( n21216 & n21296 ) | ( ~n21226 & n21296 ) ;
  assign n21307 = ~n21305 & n21306 ;
  assign n21308 = n21301 | n21307 ;
  assign n21309 = n21123 &  n21227 ;
  assign n21302 = x76 | n21123 ;
  assign n21303 = x76 &  n21123 ;
  assign n21304 = ( n21302 & ~n21303 ) | ( n21302 & 1'b0 ) | ( ~n21303 & 1'b0 ) ;
  assign n21313 = ( n2741 & n21215 ) | ( n2741 & n21304 ) | ( n21215 & n21304 ) ;
  assign n21314 = ( n21215 & ~n21226 ) | ( n21215 & n21304 ) | ( ~n21226 & n21304 ) ;
  assign n21315 = ~n21313 & n21314 ;
  assign n21316 = n21309 | n21315 ;
  assign n21317 = n21131 &  n21227 ;
  assign n21310 = x75 | n21131 ;
  assign n21311 = x75 &  n21131 ;
  assign n21312 = ( n21310 & ~n21311 ) | ( n21310 & 1'b0 ) | ( ~n21311 & 1'b0 ) ;
  assign n21321 = ( n2741 & n21214 ) | ( n2741 & n21312 ) | ( n21214 & n21312 ) ;
  assign n21322 = ( n21214 & ~n21226 ) | ( n21214 & n21312 ) | ( ~n21226 & n21312 ) ;
  assign n21323 = ~n21321 & n21322 ;
  assign n21324 = n21317 | n21323 ;
  assign n21325 = n21139 &  n21227 ;
  assign n21318 = x74 | n21139 ;
  assign n21319 = x74 &  n21139 ;
  assign n21320 = ( n21318 & ~n21319 ) | ( n21318 & 1'b0 ) | ( ~n21319 & 1'b0 ) ;
  assign n21329 = ( n2741 & n21213 ) | ( n2741 & n21320 ) | ( n21213 & n21320 ) ;
  assign n21330 = ( n21213 & ~n21226 ) | ( n21213 & n21320 ) | ( ~n21226 & n21320 ) ;
  assign n21331 = ~n21329 & n21330 ;
  assign n21332 = n21325 | n21331 ;
  assign n21333 = n21147 &  n21227 ;
  assign n21326 = x73 | n21147 ;
  assign n21327 = x73 &  n21147 ;
  assign n21328 = ( n21326 & ~n21327 ) | ( n21326 & 1'b0 ) | ( ~n21327 & 1'b0 ) ;
  assign n21337 = ( n2741 & n21212 ) | ( n2741 & n21328 ) | ( n21212 & n21328 ) ;
  assign n21338 = ( n21212 & ~n21226 ) | ( n21212 & n21328 ) | ( ~n21226 & n21328 ) ;
  assign n21339 = ~n21337 & n21338 ;
  assign n21340 = n21333 | n21339 ;
  assign n21341 = n21155 &  n21227 ;
  assign n21334 = x72 | n21155 ;
  assign n21335 = x72 &  n21155 ;
  assign n21336 = ( n21334 & ~n21335 ) | ( n21334 & 1'b0 ) | ( ~n21335 & 1'b0 ) ;
  assign n21345 = ( n2741 & n21211 ) | ( n2741 & n21336 ) | ( n21211 & n21336 ) ;
  assign n21346 = ( n21211 & ~n21226 ) | ( n21211 & n21336 ) | ( ~n21226 & n21336 ) ;
  assign n21347 = ~n21345 & n21346 ;
  assign n21348 = n21341 | n21347 ;
  assign n21349 = n21163 &  n21227 ;
  assign n21342 = x71 | n21163 ;
  assign n21343 = x71 &  n21163 ;
  assign n21344 = ( n21342 & ~n21343 ) | ( n21342 & 1'b0 ) | ( ~n21343 & 1'b0 ) ;
  assign n21353 = ( n2741 & n21210 ) | ( n2741 & n21344 ) | ( n21210 & n21344 ) ;
  assign n21354 = ( n21210 & ~n21226 ) | ( n21210 & n21344 ) | ( ~n21226 & n21344 ) ;
  assign n21355 = ~n21353 & n21354 ;
  assign n21356 = n21349 | n21355 ;
  assign n21357 = n21171 &  n21227 ;
  assign n21350 = x70 | n21171 ;
  assign n21351 = x70 &  n21171 ;
  assign n21352 = ( n21350 & ~n21351 ) | ( n21350 & 1'b0 ) | ( ~n21351 & 1'b0 ) ;
  assign n21361 = ( n2741 & n21209 ) | ( n2741 & n21352 ) | ( n21209 & n21352 ) ;
  assign n21362 = ( n21209 & ~n21226 ) | ( n21209 & n21352 ) | ( ~n21226 & n21352 ) ;
  assign n21363 = ~n21361 & n21362 ;
  assign n21364 = n21357 | n21363 ;
  assign n21365 = n21179 &  n21227 ;
  assign n21358 = x69 | n21179 ;
  assign n21359 = x69 &  n21179 ;
  assign n21360 = ( n21358 & ~n21359 ) | ( n21358 & 1'b0 ) | ( ~n21359 & 1'b0 ) ;
  assign n21369 = ( n2741 & n21208 ) | ( n2741 & n21360 ) | ( n21208 & n21360 ) ;
  assign n21370 = ( n21208 & ~n21226 ) | ( n21208 & n21360 ) | ( ~n21226 & n21360 ) ;
  assign n21371 = ~n21369 & n21370 ;
  assign n21372 = n21365 | n21371 ;
  assign n21373 = n21187 &  n21227 ;
  assign n21366 = x68 | n21187 ;
  assign n21367 = x68 &  n21187 ;
  assign n21368 = ( n21366 & ~n21367 ) | ( n21366 & 1'b0 ) | ( ~n21367 & 1'b0 ) ;
  assign n21377 = ( n2741 & n21207 ) | ( n2741 & n21368 ) | ( n21207 & n21368 ) ;
  assign n21378 = ( n21207 & ~n21226 ) | ( n21207 & n21368 ) | ( ~n21226 & n21368 ) ;
  assign n21379 = ~n21377 & n21378 ;
  assign n21380 = n21373 | n21379 ;
  assign n21381 = n21192 &  n21227 ;
  assign n21374 = x67 | n21192 ;
  assign n21375 = x67 &  n21192 ;
  assign n21376 = ( n21374 & ~n21375 ) | ( n21374 & 1'b0 ) | ( ~n21375 & 1'b0 ) ;
  assign n21385 = ( n2741 & n21206 ) | ( n2741 & n21376 ) | ( n21206 & n21376 ) ;
  assign n21386 = ( n21206 & ~n21226 ) | ( n21206 & n21376 ) | ( ~n21226 & n21376 ) ;
  assign n21387 = ~n21385 & n21386 ;
  assign n21388 = n21381 | n21387 ;
  assign n21389 = n21200 &  n21227 ;
  assign n21382 = x66 | n21200 ;
  assign n21383 = x66 &  n21200 ;
  assign n21384 = ( n21382 & ~n21383 ) | ( n21382 & 1'b0 ) | ( ~n21383 & 1'b0 ) ;
  assign n21393 = ( n2741 & n21205 ) | ( n2741 & n21384 ) | ( n21205 & n21384 ) ;
  assign n21394 = ( n21205 & ~n21226 ) | ( n21205 & n21384 ) | ( ~n21226 & n21384 ) ;
  assign n21395 = ~n21393 & n21394 ;
  assign n21396 = n21389 | n21395 ;
  assign n21397 = n21204 &  n21227 ;
  assign n21390 = x65 &  n21204 ;
  assign n21391 = x65 | n21203 ;
  assign n21392 = n21202 | n21391 ;
  assign n21398 = ~n21390 & n21392 ;
  assign n21399 = ( n2699 & ~n2741 ) | ( n2699 & n21398 ) | ( ~n2741 & n21398 ) ;
  assign n21400 = ( n2699 & n21226 ) | ( n2699 & n21398 ) | ( n21226 & n21398 ) ;
  assign n21401 = ( n21399 & ~n21400 ) | ( n21399 & 1'b0 ) | ( ~n21400 & 1'b0 ) ;
  assign n21402 = n21397 | n21401 ;
  assign n21403 = ( n2726 & ~n21226 ) | ( n2726 & 1'b0 ) | ( ~n21226 & 1'b0 ) ;
  assign n21404 = ( x41 & ~n21403 ) | ( x41 & 1'b0 ) | ( ~n21403 & 1'b0 ) ;
  assign n21405 = ( n2733 & ~n21226 ) | ( n2733 & 1'b0 ) | ( ~n21226 & 1'b0 ) ;
  assign n21406 = n21404 | n21405 ;
  assign n21407 = ( x65 & ~n21406 ) | ( x65 & n2736 ) | ( ~n21406 & n2736 ) ;
  assign n21408 = ( x66 & ~n21402 ) | ( x66 & n21407 ) | ( ~n21402 & n21407 ) ;
  assign n21409 = ( x67 & ~n21396 ) | ( x67 & n21408 ) | ( ~n21396 & n21408 ) ;
  assign n21410 = ( x68 & ~n21388 ) | ( x68 & n21409 ) | ( ~n21388 & n21409 ) ;
  assign n21411 = ( x69 & ~n21380 ) | ( x69 & n21410 ) | ( ~n21380 & n21410 ) ;
  assign n21412 = ( x70 & ~n21372 ) | ( x70 & n21411 ) | ( ~n21372 & n21411 ) ;
  assign n21413 = ( x71 & ~n21364 ) | ( x71 & n21412 ) | ( ~n21364 & n21412 ) ;
  assign n21414 = ( x72 & ~n21356 ) | ( x72 & n21413 ) | ( ~n21356 & n21413 ) ;
  assign n21415 = ( x73 & ~n21348 ) | ( x73 & n21414 ) | ( ~n21348 & n21414 ) ;
  assign n21416 = ( x74 & ~n21340 ) | ( x74 & n21415 ) | ( ~n21340 & n21415 ) ;
  assign n21417 = ( x75 & ~n21332 ) | ( x75 & n21416 ) | ( ~n21332 & n21416 ) ;
  assign n21418 = ( x76 & ~n21324 ) | ( x76 & n21417 ) | ( ~n21324 & n21417 ) ;
  assign n21419 = ( x77 & ~n21316 ) | ( x77 & n21418 ) | ( ~n21316 & n21418 ) ;
  assign n21420 = ( x78 & ~n21308 ) | ( x78 & n21419 ) | ( ~n21308 & n21419 ) ;
  assign n21421 = ( x79 & ~n21300 ) | ( x79 & n21420 ) | ( ~n21300 & n21420 ) ;
  assign n21422 = ( x80 & ~n21292 ) | ( x80 & n21421 ) | ( ~n21292 & n21421 ) ;
  assign n21423 = ( x81 & ~n21284 ) | ( x81 & n21422 ) | ( ~n21284 & n21422 ) ;
  assign n21424 = ( x82 & ~n21276 ) | ( x82 & n21423 ) | ( ~n21276 & n21423 ) ;
  assign n21425 = ( x83 & ~n21268 ) | ( x83 & n21424 ) | ( ~n21268 & n21424 ) ;
  assign n21426 = ( x84 & ~n21260 ) | ( x84 & n21425 ) | ( ~n21260 & n21425 ) ;
  assign n21427 = ( x85 & ~n21252 ) | ( x85 & n21426 ) | ( ~n21252 & n21426 ) ;
  assign n21428 = ( x86 & ~n21244 ) | ( x86 & n21427 ) | ( ~n21244 & n21427 ) ;
  assign n21429 = ( x87 & ~n21228 ) | ( x87 & 1'b0 ) | ( ~n21228 & 1'b0 ) ;
  assign n21430 = ~n21234 & n21429 ;
  assign n21431 = ( n21428 & ~n21236 ) | ( n21428 & n21430 ) | ( ~n21236 & n21430 ) ;
  assign n21432 = ( n21236 & ~n2941 ) | ( n21236 & n21431 ) | ( ~n2941 & n21431 ) ;
  assign n21433 = n2941 | n21432 ;
  assign n21440 = n2741 &  n21043 ;
  assign n21441 = n21433 &  n21440 ;
  assign n21434 = ~n21235 |  n2741 ;
  assign n21435 = n21433 &  n21434 ;
  assign n21439 = n21236 | n21430 ;
  assign n21443 = ( n21428 & n21435 ) | ( n21428 & n21439 ) | ( n21435 & n21439 ) ;
  assign n21442 = n21428 | n21439 ;
  assign n21444 = ( n21441 & ~n21443 ) | ( n21441 & n21442 ) | ( ~n21443 & n21442 ) ;
  assign n21448 = n21244 &  n21434 ;
  assign n21449 = n21433 &  n21448 ;
  assign n21436 = x86 | n21244 ;
  assign n21437 = x86 &  n21244 ;
  assign n21438 = ( n21436 & ~n21437 ) | ( n21436 & 1'b0 ) | ( ~n21437 & 1'b0 ) ;
  assign n21451 = ( n21427 & n21435 ) | ( n21427 & n21438 ) | ( n21435 & n21438 ) ;
  assign n21450 = n21427 | n21438 ;
  assign n21452 = ( n21449 & ~n21451 ) | ( n21449 & n21450 ) | ( ~n21451 & n21450 ) ;
  assign n21456 = n21252 &  n21434 ;
  assign n21457 = n21433 &  n21456 ;
  assign n21445 = x85 | n21252 ;
  assign n21446 = x85 &  n21252 ;
  assign n21447 = ( n21445 & ~n21446 ) | ( n21445 & 1'b0 ) | ( ~n21446 & 1'b0 ) ;
  assign n21459 = ( n21426 & n21435 ) | ( n21426 & n21447 ) | ( n21435 & n21447 ) ;
  assign n21458 = n21426 | n21447 ;
  assign n21460 = ( n21457 & ~n21459 ) | ( n21457 & n21458 ) | ( ~n21459 & n21458 ) ;
  assign n21464 = n21260 &  n21434 ;
  assign n21465 = n21433 &  n21464 ;
  assign n21453 = x84 | n21260 ;
  assign n21454 = x84 &  n21260 ;
  assign n21455 = ( n21453 & ~n21454 ) | ( n21453 & 1'b0 ) | ( ~n21454 & 1'b0 ) ;
  assign n21467 = ( n21425 & n21435 ) | ( n21425 & n21455 ) | ( n21435 & n21455 ) ;
  assign n21466 = n21425 | n21455 ;
  assign n21468 = ( n21465 & ~n21467 ) | ( n21465 & n21466 ) | ( ~n21467 & n21466 ) ;
  assign n21472 = n21268 &  n21434 ;
  assign n21473 = n21433 &  n21472 ;
  assign n21461 = x83 | n21268 ;
  assign n21462 = x83 &  n21268 ;
  assign n21463 = ( n21461 & ~n21462 ) | ( n21461 & 1'b0 ) | ( ~n21462 & 1'b0 ) ;
  assign n21475 = ( n21424 & n21435 ) | ( n21424 & n21463 ) | ( n21435 & n21463 ) ;
  assign n21474 = n21424 | n21463 ;
  assign n21476 = ( n21473 & ~n21475 ) | ( n21473 & n21474 ) | ( ~n21475 & n21474 ) ;
  assign n21480 = n21276 &  n21434 ;
  assign n21481 = n21433 &  n21480 ;
  assign n21469 = x82 | n21276 ;
  assign n21470 = x82 &  n21276 ;
  assign n21471 = ( n21469 & ~n21470 ) | ( n21469 & 1'b0 ) | ( ~n21470 & 1'b0 ) ;
  assign n21483 = ( n21423 & n21435 ) | ( n21423 & n21471 ) | ( n21435 & n21471 ) ;
  assign n21482 = n21423 | n21471 ;
  assign n21484 = ( n21481 & ~n21483 ) | ( n21481 & n21482 ) | ( ~n21483 & n21482 ) ;
  assign n21488 = n21284 &  n21434 ;
  assign n21489 = n21433 &  n21488 ;
  assign n21477 = x81 | n21284 ;
  assign n21478 = x81 &  n21284 ;
  assign n21479 = ( n21477 & ~n21478 ) | ( n21477 & 1'b0 ) | ( ~n21478 & 1'b0 ) ;
  assign n21491 = ( n21422 & n21435 ) | ( n21422 & n21479 ) | ( n21435 & n21479 ) ;
  assign n21490 = n21422 | n21479 ;
  assign n21492 = ( n21489 & ~n21491 ) | ( n21489 & n21490 ) | ( ~n21491 & n21490 ) ;
  assign n21496 = n21292 &  n21434 ;
  assign n21497 = n21433 &  n21496 ;
  assign n21485 = x80 | n21292 ;
  assign n21486 = x80 &  n21292 ;
  assign n21487 = ( n21485 & ~n21486 ) | ( n21485 & 1'b0 ) | ( ~n21486 & 1'b0 ) ;
  assign n21499 = ( n21421 & n21435 ) | ( n21421 & n21487 ) | ( n21435 & n21487 ) ;
  assign n21498 = n21421 | n21487 ;
  assign n21500 = ( n21497 & ~n21499 ) | ( n21497 & n21498 ) | ( ~n21499 & n21498 ) ;
  assign n21504 = n21300 &  n21434 ;
  assign n21505 = n21433 &  n21504 ;
  assign n21493 = x79 | n21300 ;
  assign n21494 = x79 &  n21300 ;
  assign n21495 = ( n21493 & ~n21494 ) | ( n21493 & 1'b0 ) | ( ~n21494 & 1'b0 ) ;
  assign n21507 = ( n21420 & n21435 ) | ( n21420 & n21495 ) | ( n21435 & n21495 ) ;
  assign n21506 = n21420 | n21495 ;
  assign n21508 = ( n21505 & ~n21507 ) | ( n21505 & n21506 ) | ( ~n21507 & n21506 ) ;
  assign n21512 = n21308 &  n21434 ;
  assign n21513 = n21433 &  n21512 ;
  assign n21501 = x78 | n21308 ;
  assign n21502 = x78 &  n21308 ;
  assign n21503 = ( n21501 & ~n21502 ) | ( n21501 & 1'b0 ) | ( ~n21502 & 1'b0 ) ;
  assign n21515 = ( n21419 & n21435 ) | ( n21419 & n21503 ) | ( n21435 & n21503 ) ;
  assign n21514 = n21419 | n21503 ;
  assign n21516 = ( n21513 & ~n21515 ) | ( n21513 & n21514 ) | ( ~n21515 & n21514 ) ;
  assign n21520 = n21316 &  n21434 ;
  assign n21521 = n21433 &  n21520 ;
  assign n21509 = x77 | n21316 ;
  assign n21510 = x77 &  n21316 ;
  assign n21511 = ( n21509 & ~n21510 ) | ( n21509 & 1'b0 ) | ( ~n21510 & 1'b0 ) ;
  assign n21523 = ( n21418 & n21435 ) | ( n21418 & n21511 ) | ( n21435 & n21511 ) ;
  assign n21522 = n21418 | n21511 ;
  assign n21524 = ( n21521 & ~n21523 ) | ( n21521 & n21522 ) | ( ~n21523 & n21522 ) ;
  assign n21528 = n21324 &  n21434 ;
  assign n21529 = n21433 &  n21528 ;
  assign n21517 = x76 | n21324 ;
  assign n21518 = x76 &  n21324 ;
  assign n21519 = ( n21517 & ~n21518 ) | ( n21517 & 1'b0 ) | ( ~n21518 & 1'b0 ) ;
  assign n21531 = ( n21417 & n21435 ) | ( n21417 & n21519 ) | ( n21435 & n21519 ) ;
  assign n21530 = n21417 | n21519 ;
  assign n21532 = ( n21529 & ~n21531 ) | ( n21529 & n21530 ) | ( ~n21531 & n21530 ) ;
  assign n21536 = n21332 &  n21434 ;
  assign n21537 = n21433 &  n21536 ;
  assign n21525 = x75 | n21332 ;
  assign n21526 = x75 &  n21332 ;
  assign n21527 = ( n21525 & ~n21526 ) | ( n21525 & 1'b0 ) | ( ~n21526 & 1'b0 ) ;
  assign n21539 = ( n21416 & n21435 ) | ( n21416 & n21527 ) | ( n21435 & n21527 ) ;
  assign n21538 = n21416 | n21527 ;
  assign n21540 = ( n21537 & ~n21539 ) | ( n21537 & n21538 ) | ( ~n21539 & n21538 ) ;
  assign n21544 = n21340 &  n21434 ;
  assign n21545 = n21433 &  n21544 ;
  assign n21533 = x74 | n21340 ;
  assign n21534 = x74 &  n21340 ;
  assign n21535 = ( n21533 & ~n21534 ) | ( n21533 & 1'b0 ) | ( ~n21534 & 1'b0 ) ;
  assign n21547 = ( n21415 & n21435 ) | ( n21415 & n21535 ) | ( n21435 & n21535 ) ;
  assign n21546 = n21415 | n21535 ;
  assign n21548 = ( n21545 & ~n21547 ) | ( n21545 & n21546 ) | ( ~n21547 & n21546 ) ;
  assign n21552 = n21348 &  n21434 ;
  assign n21553 = n21433 &  n21552 ;
  assign n21541 = x73 | n21348 ;
  assign n21542 = x73 &  n21348 ;
  assign n21543 = ( n21541 & ~n21542 ) | ( n21541 & 1'b0 ) | ( ~n21542 & 1'b0 ) ;
  assign n21555 = ( n21414 & n21435 ) | ( n21414 & n21543 ) | ( n21435 & n21543 ) ;
  assign n21554 = n21414 | n21543 ;
  assign n21556 = ( n21553 & ~n21555 ) | ( n21553 & n21554 ) | ( ~n21555 & n21554 ) ;
  assign n21560 = n21356 &  n21434 ;
  assign n21561 = n21433 &  n21560 ;
  assign n21549 = x72 | n21356 ;
  assign n21550 = x72 &  n21356 ;
  assign n21551 = ( n21549 & ~n21550 ) | ( n21549 & 1'b0 ) | ( ~n21550 & 1'b0 ) ;
  assign n21563 = ( n21413 & n21435 ) | ( n21413 & n21551 ) | ( n21435 & n21551 ) ;
  assign n21562 = n21413 | n21551 ;
  assign n21564 = ( n21561 & ~n21563 ) | ( n21561 & n21562 ) | ( ~n21563 & n21562 ) ;
  assign n21568 = n21364 &  n21434 ;
  assign n21569 = n21433 &  n21568 ;
  assign n21557 = x71 | n21364 ;
  assign n21558 = x71 &  n21364 ;
  assign n21559 = ( n21557 & ~n21558 ) | ( n21557 & 1'b0 ) | ( ~n21558 & 1'b0 ) ;
  assign n21571 = ( n21412 & n21435 ) | ( n21412 & n21559 ) | ( n21435 & n21559 ) ;
  assign n21570 = n21412 | n21559 ;
  assign n21572 = ( n21569 & ~n21571 ) | ( n21569 & n21570 ) | ( ~n21571 & n21570 ) ;
  assign n21576 = n21372 &  n21434 ;
  assign n21577 = n21433 &  n21576 ;
  assign n21565 = x70 | n21372 ;
  assign n21566 = x70 &  n21372 ;
  assign n21567 = ( n21565 & ~n21566 ) | ( n21565 & 1'b0 ) | ( ~n21566 & 1'b0 ) ;
  assign n21579 = ( n21411 & n21435 ) | ( n21411 & n21567 ) | ( n21435 & n21567 ) ;
  assign n21578 = n21411 | n21567 ;
  assign n21580 = ( n21577 & ~n21579 ) | ( n21577 & n21578 ) | ( ~n21579 & n21578 ) ;
  assign n21584 = n21380 &  n21434 ;
  assign n21585 = n21433 &  n21584 ;
  assign n21573 = x69 | n21380 ;
  assign n21574 = x69 &  n21380 ;
  assign n21575 = ( n21573 & ~n21574 ) | ( n21573 & 1'b0 ) | ( ~n21574 & 1'b0 ) ;
  assign n21587 = ( n21410 & n21435 ) | ( n21410 & n21575 ) | ( n21435 & n21575 ) ;
  assign n21586 = n21410 | n21575 ;
  assign n21588 = ( n21585 & ~n21587 ) | ( n21585 & n21586 ) | ( ~n21587 & n21586 ) ;
  assign n21592 = n21388 &  n21434 ;
  assign n21593 = n21433 &  n21592 ;
  assign n21581 = x68 | n21388 ;
  assign n21582 = x68 &  n21388 ;
  assign n21583 = ( n21581 & ~n21582 ) | ( n21581 & 1'b0 ) | ( ~n21582 & 1'b0 ) ;
  assign n21595 = ( n21409 & n21435 ) | ( n21409 & n21583 ) | ( n21435 & n21583 ) ;
  assign n21594 = n21409 | n21583 ;
  assign n21596 = ( n21593 & ~n21595 ) | ( n21593 & n21594 ) | ( ~n21595 & n21594 ) ;
  assign n21600 = n21396 &  n21434 ;
  assign n21601 = n21433 &  n21600 ;
  assign n21589 = x67 | n21396 ;
  assign n21590 = x67 &  n21396 ;
  assign n21591 = ( n21589 & ~n21590 ) | ( n21589 & 1'b0 ) | ( ~n21590 & 1'b0 ) ;
  assign n21603 = ( n21408 & n21435 ) | ( n21408 & n21591 ) | ( n21435 & n21591 ) ;
  assign n21602 = n21408 | n21591 ;
  assign n21604 = ( n21601 & ~n21603 ) | ( n21601 & n21602 ) | ( ~n21603 & n21602 ) ;
  assign n21605 = n21402 &  n21434 ;
  assign n21606 = n21433 &  n21605 ;
  assign n21597 = x66 | n21402 ;
  assign n21598 = x66 &  n21402 ;
  assign n21599 = ( n21597 & ~n21598 ) | ( n21597 & 1'b0 ) | ( ~n21598 & 1'b0 ) ;
  assign n21608 = ( n21407 & n21435 ) | ( n21407 & n21599 ) | ( n21435 & n21599 ) ;
  assign n21607 = n21407 | n21599 ;
  assign n21609 = ( n21606 & ~n21608 ) | ( n21606 & n21607 ) | ( ~n21608 & n21607 ) ;
  assign n21610 = ( x65 & ~n2736 ) | ( x65 & n21406 ) | ( ~n2736 & n21406 ) ;
  assign n21611 = ( n21407 & ~x65 ) | ( n21407 & n21610 ) | ( ~x65 & n21610 ) ;
  assign n21612 = ~n21435 & n21611 ;
  assign n21613 = n21406 &  n21434 ;
  assign n21614 = n21433 &  n21613 ;
  assign n21615 = n21612 | n21614 ;
  assign n21616 = ( x64 & ~n21435 ) | ( x64 & 1'b0 ) | ( ~n21435 & 1'b0 ) ;
  assign n21617 = ( x40 & ~n21616 ) | ( x40 & 1'b0 ) | ( ~n21616 & 1'b0 ) ;
  assign n21618 = ( n2736 & ~n21435 ) | ( n2736 & 1'b0 ) | ( ~n21435 & 1'b0 ) ;
  assign n21619 = n21617 | n21618 ;
  assign n21620 = ( x65 & ~n21619 ) | ( x65 & n3130 ) | ( ~n21619 & n3130 ) ;
  assign n21621 = ( x66 & ~n21615 ) | ( x66 & n21620 ) | ( ~n21615 & n21620 ) ;
  assign n21622 = ( x67 & ~n21609 ) | ( x67 & n21621 ) | ( ~n21609 & n21621 ) ;
  assign n21623 = ( x68 & ~n21604 ) | ( x68 & n21622 ) | ( ~n21604 & n21622 ) ;
  assign n21624 = ( x69 & ~n21596 ) | ( x69 & n21623 ) | ( ~n21596 & n21623 ) ;
  assign n21625 = ( x70 & ~n21588 ) | ( x70 & n21624 ) | ( ~n21588 & n21624 ) ;
  assign n21626 = ( x71 & ~n21580 ) | ( x71 & n21625 ) | ( ~n21580 & n21625 ) ;
  assign n21627 = ( x72 & ~n21572 ) | ( x72 & n21626 ) | ( ~n21572 & n21626 ) ;
  assign n21628 = ( x73 & ~n21564 ) | ( x73 & n21627 ) | ( ~n21564 & n21627 ) ;
  assign n21629 = ( x74 & ~n21556 ) | ( x74 & n21628 ) | ( ~n21556 & n21628 ) ;
  assign n21630 = ( x75 & ~n21548 ) | ( x75 & n21629 ) | ( ~n21548 & n21629 ) ;
  assign n21631 = ( x76 & ~n21540 ) | ( x76 & n21630 ) | ( ~n21540 & n21630 ) ;
  assign n21632 = ( x77 & ~n21532 ) | ( x77 & n21631 ) | ( ~n21532 & n21631 ) ;
  assign n21633 = ( x78 & ~n21524 ) | ( x78 & n21632 ) | ( ~n21524 & n21632 ) ;
  assign n21634 = ( x79 & ~n21516 ) | ( x79 & n21633 ) | ( ~n21516 & n21633 ) ;
  assign n21635 = ( x80 & ~n21508 ) | ( x80 & n21634 ) | ( ~n21508 & n21634 ) ;
  assign n21636 = ( x81 & ~n21500 ) | ( x81 & n21635 ) | ( ~n21500 & n21635 ) ;
  assign n21637 = ( x82 & ~n21492 ) | ( x82 & n21636 ) | ( ~n21492 & n21636 ) ;
  assign n21638 = ( x83 & ~n21484 ) | ( x83 & n21637 ) | ( ~n21484 & n21637 ) ;
  assign n21639 = ( x84 & ~n21476 ) | ( x84 & n21638 ) | ( ~n21476 & n21638 ) ;
  assign n21640 = ( x85 & ~n21468 ) | ( x85 & n21639 ) | ( ~n21468 & n21639 ) ;
  assign n21641 = ( x86 & ~n21460 ) | ( x86 & n21640 ) | ( ~n21460 & n21640 ) ;
  assign n21642 = ( x87 & ~n21452 ) | ( x87 & n21641 ) | ( ~n21452 & n21641 ) ;
  assign n21649 = ( x88 & ~n3156 ) | ( x88 & n21642 ) | ( ~n3156 & n21642 ) ;
  assign n21648 = x88 &  n21642 ;
  assign n21650 = ( n21444 & ~n21649 ) | ( n21444 & n21648 ) | ( ~n21649 & n21648 ) ;
  assign n21643 = ( x88 & ~n21444 ) | ( x88 & n21642 ) | ( ~n21444 & n21642 ) ;
  assign n21644 = n3156 | n21643 ;
  assign n21651 = n21452 &  n21644 ;
  assign n21645 = x87 | n21452 ;
  assign n21646 = x87 &  n21452 ;
  assign n21647 = ( n21645 & ~n21646 ) | ( n21645 & 1'b0 ) | ( ~n21646 & 1'b0 ) ;
  assign n21655 = ( n3156 & n21641 ) | ( n3156 & n21647 ) | ( n21641 & n21647 ) ;
  assign n21656 = ( n21641 & ~n21643 ) | ( n21641 & n21647 ) | ( ~n21643 & n21647 ) ;
  assign n21657 = ~n21655 & n21656 ;
  assign n21658 = n21651 | n21657 ;
  assign n21659 = n21460 &  n21644 ;
  assign n21652 = x86 | n21460 ;
  assign n21653 = x86 &  n21460 ;
  assign n21654 = ( n21652 & ~n21653 ) | ( n21652 & 1'b0 ) | ( ~n21653 & 1'b0 ) ;
  assign n21663 = ( n3156 & n21640 ) | ( n3156 & n21654 ) | ( n21640 & n21654 ) ;
  assign n21664 = ( n21640 & ~n21643 ) | ( n21640 & n21654 ) | ( ~n21643 & n21654 ) ;
  assign n21665 = ~n21663 & n21664 ;
  assign n21666 = n21659 | n21665 ;
  assign n21667 = n21468 &  n21644 ;
  assign n21660 = x85 | n21468 ;
  assign n21661 = x85 &  n21468 ;
  assign n21662 = ( n21660 & ~n21661 ) | ( n21660 & 1'b0 ) | ( ~n21661 & 1'b0 ) ;
  assign n21671 = ( n3156 & n21639 ) | ( n3156 & n21662 ) | ( n21639 & n21662 ) ;
  assign n21672 = ( n21639 & ~n21643 ) | ( n21639 & n21662 ) | ( ~n21643 & n21662 ) ;
  assign n21673 = ~n21671 & n21672 ;
  assign n21674 = n21667 | n21673 ;
  assign n21675 = n21476 &  n21644 ;
  assign n21668 = x84 | n21476 ;
  assign n21669 = x84 &  n21476 ;
  assign n21670 = ( n21668 & ~n21669 ) | ( n21668 & 1'b0 ) | ( ~n21669 & 1'b0 ) ;
  assign n21679 = ( n3156 & n21638 ) | ( n3156 & n21670 ) | ( n21638 & n21670 ) ;
  assign n21680 = ( n21638 & ~n21643 ) | ( n21638 & n21670 ) | ( ~n21643 & n21670 ) ;
  assign n21681 = ~n21679 & n21680 ;
  assign n21682 = n21675 | n21681 ;
  assign n21683 = n21484 &  n21644 ;
  assign n21676 = x83 | n21484 ;
  assign n21677 = x83 &  n21484 ;
  assign n21678 = ( n21676 & ~n21677 ) | ( n21676 & 1'b0 ) | ( ~n21677 & 1'b0 ) ;
  assign n21687 = ( n3156 & n21637 ) | ( n3156 & n21678 ) | ( n21637 & n21678 ) ;
  assign n21688 = ( n21637 & ~n21643 ) | ( n21637 & n21678 ) | ( ~n21643 & n21678 ) ;
  assign n21689 = ~n21687 & n21688 ;
  assign n21690 = n21683 | n21689 ;
  assign n21691 = n21492 &  n21644 ;
  assign n21684 = x82 | n21492 ;
  assign n21685 = x82 &  n21492 ;
  assign n21686 = ( n21684 & ~n21685 ) | ( n21684 & 1'b0 ) | ( ~n21685 & 1'b0 ) ;
  assign n21695 = ( n3156 & n21636 ) | ( n3156 & n21686 ) | ( n21636 & n21686 ) ;
  assign n21696 = ( n21636 & ~n21643 ) | ( n21636 & n21686 ) | ( ~n21643 & n21686 ) ;
  assign n21697 = ~n21695 & n21696 ;
  assign n21698 = n21691 | n21697 ;
  assign n21699 = n21500 &  n21644 ;
  assign n21692 = x81 | n21500 ;
  assign n21693 = x81 &  n21500 ;
  assign n21694 = ( n21692 & ~n21693 ) | ( n21692 & 1'b0 ) | ( ~n21693 & 1'b0 ) ;
  assign n21703 = ( n3156 & n21635 ) | ( n3156 & n21694 ) | ( n21635 & n21694 ) ;
  assign n21704 = ( n21635 & ~n21643 ) | ( n21635 & n21694 ) | ( ~n21643 & n21694 ) ;
  assign n21705 = ~n21703 & n21704 ;
  assign n21706 = n21699 | n21705 ;
  assign n21707 = n21508 &  n21644 ;
  assign n21700 = x80 | n21508 ;
  assign n21701 = x80 &  n21508 ;
  assign n21702 = ( n21700 & ~n21701 ) | ( n21700 & 1'b0 ) | ( ~n21701 & 1'b0 ) ;
  assign n21711 = ( n3156 & n21634 ) | ( n3156 & n21702 ) | ( n21634 & n21702 ) ;
  assign n21712 = ( n21634 & ~n21643 ) | ( n21634 & n21702 ) | ( ~n21643 & n21702 ) ;
  assign n21713 = ~n21711 & n21712 ;
  assign n21714 = n21707 | n21713 ;
  assign n21715 = n21516 &  n21644 ;
  assign n21708 = x79 | n21516 ;
  assign n21709 = x79 &  n21516 ;
  assign n21710 = ( n21708 & ~n21709 ) | ( n21708 & 1'b0 ) | ( ~n21709 & 1'b0 ) ;
  assign n21719 = ( n3156 & n21633 ) | ( n3156 & n21710 ) | ( n21633 & n21710 ) ;
  assign n21720 = ( n21633 & ~n21643 ) | ( n21633 & n21710 ) | ( ~n21643 & n21710 ) ;
  assign n21721 = ~n21719 & n21720 ;
  assign n21722 = n21715 | n21721 ;
  assign n21723 = n21524 &  n21644 ;
  assign n21716 = x78 | n21524 ;
  assign n21717 = x78 &  n21524 ;
  assign n21718 = ( n21716 & ~n21717 ) | ( n21716 & 1'b0 ) | ( ~n21717 & 1'b0 ) ;
  assign n21727 = ( n3156 & n21632 ) | ( n3156 & n21718 ) | ( n21632 & n21718 ) ;
  assign n21728 = ( n21632 & ~n21643 ) | ( n21632 & n21718 ) | ( ~n21643 & n21718 ) ;
  assign n21729 = ~n21727 & n21728 ;
  assign n21730 = n21723 | n21729 ;
  assign n21731 = n21532 &  n21644 ;
  assign n21724 = x77 | n21532 ;
  assign n21725 = x77 &  n21532 ;
  assign n21726 = ( n21724 & ~n21725 ) | ( n21724 & 1'b0 ) | ( ~n21725 & 1'b0 ) ;
  assign n21735 = ( n3156 & n21631 ) | ( n3156 & n21726 ) | ( n21631 & n21726 ) ;
  assign n21736 = ( n21631 & ~n21643 ) | ( n21631 & n21726 ) | ( ~n21643 & n21726 ) ;
  assign n21737 = ~n21735 & n21736 ;
  assign n21738 = n21731 | n21737 ;
  assign n21739 = n21540 &  n21644 ;
  assign n21732 = x76 | n21540 ;
  assign n21733 = x76 &  n21540 ;
  assign n21734 = ( n21732 & ~n21733 ) | ( n21732 & 1'b0 ) | ( ~n21733 & 1'b0 ) ;
  assign n21743 = ( n3156 & n21630 ) | ( n3156 & n21734 ) | ( n21630 & n21734 ) ;
  assign n21744 = ( n21630 & ~n21643 ) | ( n21630 & n21734 ) | ( ~n21643 & n21734 ) ;
  assign n21745 = ~n21743 & n21744 ;
  assign n21746 = n21739 | n21745 ;
  assign n21747 = n21548 &  n21644 ;
  assign n21740 = x75 | n21548 ;
  assign n21741 = x75 &  n21548 ;
  assign n21742 = ( n21740 & ~n21741 ) | ( n21740 & 1'b0 ) | ( ~n21741 & 1'b0 ) ;
  assign n21751 = ( n3156 & n21629 ) | ( n3156 & n21742 ) | ( n21629 & n21742 ) ;
  assign n21752 = ( n21629 & ~n21643 ) | ( n21629 & n21742 ) | ( ~n21643 & n21742 ) ;
  assign n21753 = ~n21751 & n21752 ;
  assign n21754 = n21747 | n21753 ;
  assign n21755 = n21556 &  n21644 ;
  assign n21748 = x74 | n21556 ;
  assign n21749 = x74 &  n21556 ;
  assign n21750 = ( n21748 & ~n21749 ) | ( n21748 & 1'b0 ) | ( ~n21749 & 1'b0 ) ;
  assign n21759 = ( n3156 & n21628 ) | ( n3156 & n21750 ) | ( n21628 & n21750 ) ;
  assign n21760 = ( n21628 & ~n21643 ) | ( n21628 & n21750 ) | ( ~n21643 & n21750 ) ;
  assign n21761 = ~n21759 & n21760 ;
  assign n21762 = n21755 | n21761 ;
  assign n21763 = n21564 &  n21644 ;
  assign n21756 = x73 | n21564 ;
  assign n21757 = x73 &  n21564 ;
  assign n21758 = ( n21756 & ~n21757 ) | ( n21756 & 1'b0 ) | ( ~n21757 & 1'b0 ) ;
  assign n21767 = ( n3156 & n21627 ) | ( n3156 & n21758 ) | ( n21627 & n21758 ) ;
  assign n21768 = ( n21627 & ~n21643 ) | ( n21627 & n21758 ) | ( ~n21643 & n21758 ) ;
  assign n21769 = ~n21767 & n21768 ;
  assign n21770 = n21763 | n21769 ;
  assign n21771 = n21572 &  n21644 ;
  assign n21764 = x72 | n21572 ;
  assign n21765 = x72 &  n21572 ;
  assign n21766 = ( n21764 & ~n21765 ) | ( n21764 & 1'b0 ) | ( ~n21765 & 1'b0 ) ;
  assign n21775 = ( n3156 & n21626 ) | ( n3156 & n21766 ) | ( n21626 & n21766 ) ;
  assign n21776 = ( n21626 & ~n21643 ) | ( n21626 & n21766 ) | ( ~n21643 & n21766 ) ;
  assign n21777 = ~n21775 & n21776 ;
  assign n21778 = n21771 | n21777 ;
  assign n21779 = n21580 &  n21644 ;
  assign n21772 = x71 | n21580 ;
  assign n21773 = x71 &  n21580 ;
  assign n21774 = ( n21772 & ~n21773 ) | ( n21772 & 1'b0 ) | ( ~n21773 & 1'b0 ) ;
  assign n21783 = ( n3156 & n21625 ) | ( n3156 & n21774 ) | ( n21625 & n21774 ) ;
  assign n21784 = ( n21625 & ~n21643 ) | ( n21625 & n21774 ) | ( ~n21643 & n21774 ) ;
  assign n21785 = ~n21783 & n21784 ;
  assign n21786 = n21779 | n21785 ;
  assign n21787 = n21588 &  n21644 ;
  assign n21780 = x70 | n21588 ;
  assign n21781 = x70 &  n21588 ;
  assign n21782 = ( n21780 & ~n21781 ) | ( n21780 & 1'b0 ) | ( ~n21781 & 1'b0 ) ;
  assign n21791 = ( n3156 & n21624 ) | ( n3156 & n21782 ) | ( n21624 & n21782 ) ;
  assign n21792 = ( n21624 & ~n21643 ) | ( n21624 & n21782 ) | ( ~n21643 & n21782 ) ;
  assign n21793 = ~n21791 & n21792 ;
  assign n21794 = n21787 | n21793 ;
  assign n21795 = n21596 &  n21644 ;
  assign n21788 = x69 | n21596 ;
  assign n21789 = x69 &  n21596 ;
  assign n21790 = ( n21788 & ~n21789 ) | ( n21788 & 1'b0 ) | ( ~n21789 & 1'b0 ) ;
  assign n21799 = ( n3156 & n21623 ) | ( n3156 & n21790 ) | ( n21623 & n21790 ) ;
  assign n21800 = ( n21623 & ~n21643 ) | ( n21623 & n21790 ) | ( ~n21643 & n21790 ) ;
  assign n21801 = ~n21799 & n21800 ;
  assign n21802 = n21795 | n21801 ;
  assign n21803 = n21604 &  n21644 ;
  assign n21796 = x68 | n21604 ;
  assign n21797 = x68 &  n21604 ;
  assign n21798 = ( n21796 & ~n21797 ) | ( n21796 & 1'b0 ) | ( ~n21797 & 1'b0 ) ;
  assign n21807 = ( n3156 & n21622 ) | ( n3156 & n21798 ) | ( n21622 & n21798 ) ;
  assign n21808 = ( n21622 & ~n21643 ) | ( n21622 & n21798 ) | ( ~n21643 & n21798 ) ;
  assign n21809 = ~n21807 & n21808 ;
  assign n21810 = n21803 | n21809 ;
  assign n21811 = n21609 &  n21644 ;
  assign n21804 = x67 | n21609 ;
  assign n21805 = x67 &  n21609 ;
  assign n21806 = ( n21804 & ~n21805 ) | ( n21804 & 1'b0 ) | ( ~n21805 & 1'b0 ) ;
  assign n21815 = ( n3156 & n21621 ) | ( n3156 & n21806 ) | ( n21621 & n21806 ) ;
  assign n21816 = ( n21621 & ~n21643 ) | ( n21621 & n21806 ) | ( ~n21643 & n21806 ) ;
  assign n21817 = ~n21815 & n21816 ;
  assign n21818 = n21811 | n21817 ;
  assign n21819 = n21615 &  n21644 ;
  assign n21812 = x66 | n21615 ;
  assign n21813 = x66 &  n21615 ;
  assign n21814 = ( n21812 & ~n21813 ) | ( n21812 & 1'b0 ) | ( ~n21813 & 1'b0 ) ;
  assign n21820 = ( n3156 & n21620 ) | ( n3156 & n21814 ) | ( n21620 & n21814 ) ;
  assign n21821 = ( n21620 & ~n21643 ) | ( n21620 & n21814 ) | ( ~n21643 & n21814 ) ;
  assign n21822 = ~n21820 & n21821 ;
  assign n21823 = n21819 | n21822 ;
  assign n21824 = n21619 &  n21644 ;
  assign n21825 = ( x65 & ~x40 ) | ( x65 & n21616 ) | ( ~x40 & n21616 ) ;
  assign n21826 = ( x40 & ~n21616 ) | ( x40 & x65 ) | ( ~n21616 & x65 ) ;
  assign n21827 = ( n21825 & ~x65 ) | ( n21825 & n21826 ) | ( ~x65 & n21826 ) ;
  assign n21828 = ( n3130 & ~n3156 ) | ( n3130 & n21827 ) | ( ~n3156 & n21827 ) ;
  assign n21829 = ( n3130 & n21643 ) | ( n3130 & n21827 ) | ( n21643 & n21827 ) ;
  assign n21830 = ( n21828 & ~n21829 ) | ( n21828 & 1'b0 ) | ( ~n21829 & 1'b0 ) ;
  assign n21831 = n21824 | n21830 ;
  assign n21832 = ( n3351 & ~n21643 ) | ( n3351 & 1'b0 ) | ( ~n21643 & 1'b0 ) ;
  assign n21833 = ( x39 & ~n21832 ) | ( x39 & 1'b0 ) | ( ~n21832 & 1'b0 ) ;
  assign n21834 = ( n3357 & ~n21643 ) | ( n3357 & 1'b0 ) | ( ~n21643 & 1'b0 ) ;
  assign n21835 = n21833 | n21834 ;
  assign n21836 = ( x65 & ~n21835 ) | ( x65 & n3360 ) | ( ~n21835 & n3360 ) ;
  assign n21837 = ( x66 & ~n21831 ) | ( x66 & n21836 ) | ( ~n21831 & n21836 ) ;
  assign n21838 = ( x67 & ~n21823 ) | ( x67 & n21837 ) | ( ~n21823 & n21837 ) ;
  assign n21839 = ( x68 & ~n21818 ) | ( x68 & n21838 ) | ( ~n21818 & n21838 ) ;
  assign n21840 = ( x69 & ~n21810 ) | ( x69 & n21839 ) | ( ~n21810 & n21839 ) ;
  assign n21841 = ( x70 & ~n21802 ) | ( x70 & n21840 ) | ( ~n21802 & n21840 ) ;
  assign n21842 = ( x71 & ~n21794 ) | ( x71 & n21841 ) | ( ~n21794 & n21841 ) ;
  assign n21843 = ( x72 & ~n21786 ) | ( x72 & n21842 ) | ( ~n21786 & n21842 ) ;
  assign n21844 = ( x73 & ~n21778 ) | ( x73 & n21843 ) | ( ~n21778 & n21843 ) ;
  assign n21845 = ( x74 & ~n21770 ) | ( x74 & n21844 ) | ( ~n21770 & n21844 ) ;
  assign n21846 = ( x75 & ~n21762 ) | ( x75 & n21845 ) | ( ~n21762 & n21845 ) ;
  assign n21847 = ( x76 & ~n21754 ) | ( x76 & n21846 ) | ( ~n21754 & n21846 ) ;
  assign n21848 = ( x77 & ~n21746 ) | ( x77 & n21847 ) | ( ~n21746 & n21847 ) ;
  assign n21849 = ( x78 & ~n21738 ) | ( x78 & n21848 ) | ( ~n21738 & n21848 ) ;
  assign n21850 = ( x79 & ~n21730 ) | ( x79 & n21849 ) | ( ~n21730 & n21849 ) ;
  assign n21851 = ( x80 & ~n21722 ) | ( x80 & n21850 ) | ( ~n21722 & n21850 ) ;
  assign n21852 = ( x81 & ~n21714 ) | ( x81 & n21851 ) | ( ~n21714 & n21851 ) ;
  assign n21853 = ( x82 & ~n21706 ) | ( x82 & n21852 ) | ( ~n21706 & n21852 ) ;
  assign n21854 = ( x83 & ~n21698 ) | ( x83 & n21853 ) | ( ~n21698 & n21853 ) ;
  assign n21855 = ( x84 & ~n21690 ) | ( x84 & n21854 ) | ( ~n21690 & n21854 ) ;
  assign n21856 = ( x85 & ~n21682 ) | ( x85 & n21855 ) | ( ~n21682 & n21855 ) ;
  assign n21857 = ( x86 & ~n21674 ) | ( x86 & n21856 ) | ( ~n21674 & n21856 ) ;
  assign n21858 = ( x87 & ~n21666 ) | ( x87 & n21857 ) | ( ~n21666 & n21857 ) ;
  assign n21859 = ( x88 & ~n21658 ) | ( x88 & n21858 ) | ( ~n21658 & n21858 ) ;
  assign n21860 = ( x89 & ~n21650 ) | ( x89 & n21859 ) | ( ~n21650 & n21859 ) ;
  assign n21861 = n3388 | n21860 ;
  assign n21862 = n21650 &  n21861 ;
  assign n21866 = ( n3388 & n21650 ) | ( n3388 & n21859 ) | ( n21650 & n21859 ) ;
  assign n21867 = ( x89 & ~n21866 ) | ( x89 & n21650 ) | ( ~n21866 & n21650 ) ;
  assign n21868 = ~x89 & n21867 ;
  assign n21869 = n21862 | n21868 ;
  assign n21870 = ~x90 & n21869 ;
  assign n21871 = n21658 &  n21861 ;
  assign n21863 = x88 | n21658 ;
  assign n21864 = x88 &  n21658 ;
  assign n21865 = ( n21863 & ~n21864 ) | ( n21863 & 1'b0 ) | ( ~n21864 & 1'b0 ) ;
  assign n21875 = ( n3388 & n21858 ) | ( n3388 & n21865 ) | ( n21858 & n21865 ) ;
  assign n21876 = ( n21858 & ~n21860 ) | ( n21858 & n21865 ) | ( ~n21860 & n21865 ) ;
  assign n21877 = ~n21875 & n21876 ;
  assign n21878 = n21871 | n21877 ;
  assign n21879 = n21666 &  n21861 ;
  assign n21872 = x87 | n21666 ;
  assign n21873 = x87 &  n21666 ;
  assign n21874 = ( n21872 & ~n21873 ) | ( n21872 & 1'b0 ) | ( ~n21873 & 1'b0 ) ;
  assign n21883 = ( n3388 & n21857 ) | ( n3388 & n21874 ) | ( n21857 & n21874 ) ;
  assign n21884 = ( n21857 & ~n21860 ) | ( n21857 & n21874 ) | ( ~n21860 & n21874 ) ;
  assign n21885 = ~n21883 & n21884 ;
  assign n21886 = n21879 | n21885 ;
  assign n21887 = n21674 &  n21861 ;
  assign n21880 = x86 | n21674 ;
  assign n21881 = x86 &  n21674 ;
  assign n21882 = ( n21880 & ~n21881 ) | ( n21880 & 1'b0 ) | ( ~n21881 & 1'b0 ) ;
  assign n21891 = ( n3388 & n21856 ) | ( n3388 & n21882 ) | ( n21856 & n21882 ) ;
  assign n21892 = ( n21856 & ~n21860 ) | ( n21856 & n21882 ) | ( ~n21860 & n21882 ) ;
  assign n21893 = ~n21891 & n21892 ;
  assign n21894 = n21887 | n21893 ;
  assign n21895 = n21682 &  n21861 ;
  assign n21888 = x85 | n21682 ;
  assign n21889 = x85 &  n21682 ;
  assign n21890 = ( n21888 & ~n21889 ) | ( n21888 & 1'b0 ) | ( ~n21889 & 1'b0 ) ;
  assign n21899 = ( n3388 & n21855 ) | ( n3388 & n21890 ) | ( n21855 & n21890 ) ;
  assign n21900 = ( n21855 & ~n21860 ) | ( n21855 & n21890 ) | ( ~n21860 & n21890 ) ;
  assign n21901 = ~n21899 & n21900 ;
  assign n21902 = n21895 | n21901 ;
  assign n21903 = n21690 &  n21861 ;
  assign n21896 = x84 | n21690 ;
  assign n21897 = x84 &  n21690 ;
  assign n21898 = ( n21896 & ~n21897 ) | ( n21896 & 1'b0 ) | ( ~n21897 & 1'b0 ) ;
  assign n21907 = ( n3388 & n21854 ) | ( n3388 & n21898 ) | ( n21854 & n21898 ) ;
  assign n21908 = ( n21854 & ~n21860 ) | ( n21854 & n21898 ) | ( ~n21860 & n21898 ) ;
  assign n21909 = ~n21907 & n21908 ;
  assign n21910 = n21903 | n21909 ;
  assign n21911 = n21698 &  n21861 ;
  assign n21904 = x83 | n21698 ;
  assign n21905 = x83 &  n21698 ;
  assign n21906 = ( n21904 & ~n21905 ) | ( n21904 & 1'b0 ) | ( ~n21905 & 1'b0 ) ;
  assign n21915 = ( n3388 & n21853 ) | ( n3388 & n21906 ) | ( n21853 & n21906 ) ;
  assign n21916 = ( n21853 & ~n21860 ) | ( n21853 & n21906 ) | ( ~n21860 & n21906 ) ;
  assign n21917 = ~n21915 & n21916 ;
  assign n21918 = n21911 | n21917 ;
  assign n21919 = n21706 &  n21861 ;
  assign n21912 = x82 | n21706 ;
  assign n21913 = x82 &  n21706 ;
  assign n21914 = ( n21912 & ~n21913 ) | ( n21912 & 1'b0 ) | ( ~n21913 & 1'b0 ) ;
  assign n21923 = ( n3388 & n21852 ) | ( n3388 & n21914 ) | ( n21852 & n21914 ) ;
  assign n21924 = ( n21852 & ~n21860 ) | ( n21852 & n21914 ) | ( ~n21860 & n21914 ) ;
  assign n21925 = ~n21923 & n21924 ;
  assign n21926 = n21919 | n21925 ;
  assign n21927 = n21714 &  n21861 ;
  assign n21920 = x81 | n21714 ;
  assign n21921 = x81 &  n21714 ;
  assign n21922 = ( n21920 & ~n21921 ) | ( n21920 & 1'b0 ) | ( ~n21921 & 1'b0 ) ;
  assign n21931 = ( n3388 & n21851 ) | ( n3388 & n21922 ) | ( n21851 & n21922 ) ;
  assign n21932 = ( n21851 & ~n21860 ) | ( n21851 & n21922 ) | ( ~n21860 & n21922 ) ;
  assign n21933 = ~n21931 & n21932 ;
  assign n21934 = n21927 | n21933 ;
  assign n21935 = n21722 &  n21861 ;
  assign n21928 = x80 | n21722 ;
  assign n21929 = x80 &  n21722 ;
  assign n21930 = ( n21928 & ~n21929 ) | ( n21928 & 1'b0 ) | ( ~n21929 & 1'b0 ) ;
  assign n21939 = ( n3388 & n21850 ) | ( n3388 & n21930 ) | ( n21850 & n21930 ) ;
  assign n21940 = ( n21850 & ~n21860 ) | ( n21850 & n21930 ) | ( ~n21860 & n21930 ) ;
  assign n21941 = ~n21939 & n21940 ;
  assign n21942 = n21935 | n21941 ;
  assign n21943 = n21730 &  n21861 ;
  assign n21936 = x79 | n21730 ;
  assign n21937 = x79 &  n21730 ;
  assign n21938 = ( n21936 & ~n21937 ) | ( n21936 & 1'b0 ) | ( ~n21937 & 1'b0 ) ;
  assign n21947 = ( n3388 & n21849 ) | ( n3388 & n21938 ) | ( n21849 & n21938 ) ;
  assign n21948 = ( n21849 & ~n21860 ) | ( n21849 & n21938 ) | ( ~n21860 & n21938 ) ;
  assign n21949 = ~n21947 & n21948 ;
  assign n21950 = n21943 | n21949 ;
  assign n21951 = n21738 &  n21861 ;
  assign n21944 = x78 | n21738 ;
  assign n21945 = x78 &  n21738 ;
  assign n21946 = ( n21944 & ~n21945 ) | ( n21944 & 1'b0 ) | ( ~n21945 & 1'b0 ) ;
  assign n21955 = ( n3388 & n21848 ) | ( n3388 & n21946 ) | ( n21848 & n21946 ) ;
  assign n21956 = ( n21848 & ~n21860 ) | ( n21848 & n21946 ) | ( ~n21860 & n21946 ) ;
  assign n21957 = ~n21955 & n21956 ;
  assign n21958 = n21951 | n21957 ;
  assign n21959 = n21746 &  n21861 ;
  assign n21952 = x77 | n21746 ;
  assign n21953 = x77 &  n21746 ;
  assign n21954 = ( n21952 & ~n21953 ) | ( n21952 & 1'b0 ) | ( ~n21953 & 1'b0 ) ;
  assign n21963 = ( n3388 & n21847 ) | ( n3388 & n21954 ) | ( n21847 & n21954 ) ;
  assign n21964 = ( n21847 & ~n21860 ) | ( n21847 & n21954 ) | ( ~n21860 & n21954 ) ;
  assign n21965 = ~n21963 & n21964 ;
  assign n21966 = n21959 | n21965 ;
  assign n21967 = n21754 &  n21861 ;
  assign n21960 = x76 | n21754 ;
  assign n21961 = x76 &  n21754 ;
  assign n21962 = ( n21960 & ~n21961 ) | ( n21960 & 1'b0 ) | ( ~n21961 & 1'b0 ) ;
  assign n21971 = ( n3388 & n21846 ) | ( n3388 & n21962 ) | ( n21846 & n21962 ) ;
  assign n21972 = ( n21846 & ~n21860 ) | ( n21846 & n21962 ) | ( ~n21860 & n21962 ) ;
  assign n21973 = ~n21971 & n21972 ;
  assign n21974 = n21967 | n21973 ;
  assign n21975 = n21762 &  n21861 ;
  assign n21968 = x75 | n21762 ;
  assign n21969 = x75 &  n21762 ;
  assign n21970 = ( n21968 & ~n21969 ) | ( n21968 & 1'b0 ) | ( ~n21969 & 1'b0 ) ;
  assign n21979 = ( n3388 & n21845 ) | ( n3388 & n21970 ) | ( n21845 & n21970 ) ;
  assign n21980 = ( n21845 & ~n21860 ) | ( n21845 & n21970 ) | ( ~n21860 & n21970 ) ;
  assign n21981 = ~n21979 & n21980 ;
  assign n21982 = n21975 | n21981 ;
  assign n21983 = n21770 &  n21861 ;
  assign n21976 = x74 | n21770 ;
  assign n21977 = x74 &  n21770 ;
  assign n21978 = ( n21976 & ~n21977 ) | ( n21976 & 1'b0 ) | ( ~n21977 & 1'b0 ) ;
  assign n21987 = ( n3388 & n21844 ) | ( n3388 & n21978 ) | ( n21844 & n21978 ) ;
  assign n21988 = ( n21844 & ~n21860 ) | ( n21844 & n21978 ) | ( ~n21860 & n21978 ) ;
  assign n21989 = ~n21987 & n21988 ;
  assign n21990 = n21983 | n21989 ;
  assign n21991 = n21778 &  n21861 ;
  assign n21984 = x73 | n21778 ;
  assign n21985 = x73 &  n21778 ;
  assign n21986 = ( n21984 & ~n21985 ) | ( n21984 & 1'b0 ) | ( ~n21985 & 1'b0 ) ;
  assign n21995 = ( n3388 & n21843 ) | ( n3388 & n21986 ) | ( n21843 & n21986 ) ;
  assign n21996 = ( n21843 & ~n21860 ) | ( n21843 & n21986 ) | ( ~n21860 & n21986 ) ;
  assign n21997 = ~n21995 & n21996 ;
  assign n21998 = n21991 | n21997 ;
  assign n21999 = n21786 &  n21861 ;
  assign n21992 = x72 | n21786 ;
  assign n21993 = x72 &  n21786 ;
  assign n21994 = ( n21992 & ~n21993 ) | ( n21992 & 1'b0 ) | ( ~n21993 & 1'b0 ) ;
  assign n22003 = ( n3388 & n21842 ) | ( n3388 & n21994 ) | ( n21842 & n21994 ) ;
  assign n22004 = ( n21842 & ~n21860 ) | ( n21842 & n21994 ) | ( ~n21860 & n21994 ) ;
  assign n22005 = ~n22003 & n22004 ;
  assign n22006 = n21999 | n22005 ;
  assign n22007 = n21794 &  n21861 ;
  assign n22000 = x71 | n21794 ;
  assign n22001 = x71 &  n21794 ;
  assign n22002 = ( n22000 & ~n22001 ) | ( n22000 & 1'b0 ) | ( ~n22001 & 1'b0 ) ;
  assign n22011 = ( n3388 & n21841 ) | ( n3388 & n22002 ) | ( n21841 & n22002 ) ;
  assign n22012 = ( n21841 & ~n21860 ) | ( n21841 & n22002 ) | ( ~n21860 & n22002 ) ;
  assign n22013 = ~n22011 & n22012 ;
  assign n22014 = n22007 | n22013 ;
  assign n22015 = n21802 &  n21861 ;
  assign n22008 = x70 | n21802 ;
  assign n22009 = x70 &  n21802 ;
  assign n22010 = ( n22008 & ~n22009 ) | ( n22008 & 1'b0 ) | ( ~n22009 & 1'b0 ) ;
  assign n22019 = ( n3388 & n21840 ) | ( n3388 & n22010 ) | ( n21840 & n22010 ) ;
  assign n22020 = ( n21840 & ~n21860 ) | ( n21840 & n22010 ) | ( ~n21860 & n22010 ) ;
  assign n22021 = ~n22019 & n22020 ;
  assign n22022 = n22015 | n22021 ;
  assign n22023 = n21810 &  n21861 ;
  assign n22016 = x69 | n21810 ;
  assign n22017 = x69 &  n21810 ;
  assign n22018 = ( n22016 & ~n22017 ) | ( n22016 & 1'b0 ) | ( ~n22017 & 1'b0 ) ;
  assign n22027 = ( n3388 & n21839 ) | ( n3388 & n22018 ) | ( n21839 & n22018 ) ;
  assign n22028 = ( n21839 & ~n21860 ) | ( n21839 & n22018 ) | ( ~n21860 & n22018 ) ;
  assign n22029 = ~n22027 & n22028 ;
  assign n22030 = n22023 | n22029 ;
  assign n22031 = n21818 &  n21861 ;
  assign n22024 = x68 | n21818 ;
  assign n22025 = x68 &  n21818 ;
  assign n22026 = ( n22024 & ~n22025 ) | ( n22024 & 1'b0 ) | ( ~n22025 & 1'b0 ) ;
  assign n22035 = ( n3388 & n21838 ) | ( n3388 & n22026 ) | ( n21838 & n22026 ) ;
  assign n22036 = ( n21838 & ~n21860 ) | ( n21838 & n22026 ) | ( ~n21860 & n22026 ) ;
  assign n22037 = ~n22035 & n22036 ;
  assign n22038 = n22031 | n22037 ;
  assign n22039 = n21823 &  n21861 ;
  assign n22032 = x67 | n21823 ;
  assign n22033 = x67 &  n21823 ;
  assign n22034 = ( n22032 & ~n22033 ) | ( n22032 & 1'b0 ) | ( ~n22033 & 1'b0 ) ;
  assign n22043 = ( n3388 & n21837 ) | ( n3388 & n22034 ) | ( n21837 & n22034 ) ;
  assign n22044 = ( n21837 & ~n21860 ) | ( n21837 & n22034 ) | ( ~n21860 & n22034 ) ;
  assign n22045 = ~n22043 & n22044 ;
  assign n22046 = n22039 | n22045 ;
  assign n22047 = n21831 &  n21861 ;
  assign n22040 = x66 | n21831 ;
  assign n22041 = x66 &  n21831 ;
  assign n22042 = ( n22040 & ~n22041 ) | ( n22040 & 1'b0 ) | ( ~n22041 & 1'b0 ) ;
  assign n22051 = ( n3388 & n21836 ) | ( n3388 & n22042 ) | ( n21836 & n22042 ) ;
  assign n22052 = ( n21836 & ~n21860 ) | ( n21836 & n22042 ) | ( ~n21860 & n22042 ) ;
  assign n22053 = ~n22051 & n22052 ;
  assign n22054 = n22047 | n22053 ;
  assign n22055 = n21835 &  n21861 ;
  assign n22048 = x65 &  n21835 ;
  assign n22049 = x65 | n21834 ;
  assign n22050 = n21833 | n22049 ;
  assign n22056 = ~n22048 & n22050 ;
  assign n22057 = ( n3360 & ~n3388 ) | ( n3360 & n22056 ) | ( ~n3388 & n22056 ) ;
  assign n22058 = ( n3360 & n21860 ) | ( n3360 & n22056 ) | ( n21860 & n22056 ) ;
  assign n22059 = ( n22057 & ~n22058 ) | ( n22057 & 1'b0 ) | ( ~n22058 & 1'b0 ) ;
  assign n22060 = n22055 | n22059 ;
  assign n22061 = ( n3428 & ~n21860 ) | ( n3428 & 1'b0 ) | ( ~n21860 & 1'b0 ) ;
  assign n22062 = ( x38 & ~n22061 ) | ( x38 & 1'b0 ) | ( ~n22061 & 1'b0 ) ;
  assign n22063 = ( n3434 & ~n21860 ) | ( n3434 & 1'b0 ) | ( ~n21860 & 1'b0 ) ;
  assign n22064 = n22062 | n22063 ;
  assign n22065 = ( x65 & ~n22064 ) | ( x65 & n3437 ) | ( ~n22064 & n3437 ) ;
  assign n22066 = ( x66 & ~n22060 ) | ( x66 & n22065 ) | ( ~n22060 & n22065 ) ;
  assign n22067 = ( x67 & ~n22054 ) | ( x67 & n22066 ) | ( ~n22054 & n22066 ) ;
  assign n22068 = ( x68 & ~n22046 ) | ( x68 & n22067 ) | ( ~n22046 & n22067 ) ;
  assign n22069 = ( x69 & ~n22038 ) | ( x69 & n22068 ) | ( ~n22038 & n22068 ) ;
  assign n22070 = ( x70 & ~n22030 ) | ( x70 & n22069 ) | ( ~n22030 & n22069 ) ;
  assign n22071 = ( x71 & ~n22022 ) | ( x71 & n22070 ) | ( ~n22022 & n22070 ) ;
  assign n22072 = ( x72 & ~n22014 ) | ( x72 & n22071 ) | ( ~n22014 & n22071 ) ;
  assign n22073 = ( x73 & ~n22006 ) | ( x73 & n22072 ) | ( ~n22006 & n22072 ) ;
  assign n22074 = ( x74 & ~n21998 ) | ( x74 & n22073 ) | ( ~n21998 & n22073 ) ;
  assign n22075 = ( x75 & ~n21990 ) | ( x75 & n22074 ) | ( ~n21990 & n22074 ) ;
  assign n22076 = ( x76 & ~n21982 ) | ( x76 & n22075 ) | ( ~n21982 & n22075 ) ;
  assign n22077 = ( x77 & ~n21974 ) | ( x77 & n22076 ) | ( ~n21974 & n22076 ) ;
  assign n22078 = ( x78 & ~n21966 ) | ( x78 & n22077 ) | ( ~n21966 & n22077 ) ;
  assign n22079 = ( x79 & ~n21958 ) | ( x79 & n22078 ) | ( ~n21958 & n22078 ) ;
  assign n22080 = ( x80 & ~n21950 ) | ( x80 & n22079 ) | ( ~n21950 & n22079 ) ;
  assign n22081 = ( x81 & ~n21942 ) | ( x81 & n22080 ) | ( ~n21942 & n22080 ) ;
  assign n22082 = ( x82 & ~n21934 ) | ( x82 & n22081 ) | ( ~n21934 & n22081 ) ;
  assign n22083 = ( x83 & ~n21926 ) | ( x83 & n22082 ) | ( ~n21926 & n22082 ) ;
  assign n22084 = ( x84 & ~n21918 ) | ( x84 & n22083 ) | ( ~n21918 & n22083 ) ;
  assign n22085 = ( x85 & ~n21910 ) | ( x85 & n22084 ) | ( ~n21910 & n22084 ) ;
  assign n22086 = ( x86 & ~n21902 ) | ( x86 & n22085 ) | ( ~n21902 & n22085 ) ;
  assign n22087 = ( x87 & ~n21894 ) | ( x87 & n22086 ) | ( ~n21894 & n22086 ) ;
  assign n22088 = ( x88 & ~n21886 ) | ( x88 & n22087 ) | ( ~n21886 & n22087 ) ;
  assign n22089 = ( x89 & ~n21878 ) | ( x89 & n22088 ) | ( ~n21878 & n22088 ) ;
  assign n22090 = ( x90 & ~n21862 ) | ( x90 & 1'b0 ) | ( ~n21862 & 1'b0 ) ;
  assign n22091 = ~n21868 & n22090 ;
  assign n22092 = ( n22089 & ~n21870 ) | ( n22089 & n22091 ) | ( ~n21870 & n22091 ) ;
  assign n22093 = ( n21870 & ~n3634 ) | ( n21870 & n22092 ) | ( ~n3634 & n22092 ) ;
  assign n22094 = n3634 | n22093 ;
  assign n22101 = n3388 &  n21650 ;
  assign n22102 = n22094 &  n22101 ;
  assign n22095 = ~n21869 |  n3388 ;
  assign n22096 = n22094 &  n22095 ;
  assign n22100 = n21870 | n22091 ;
  assign n22104 = ( n22089 & n22096 ) | ( n22089 & n22100 ) | ( n22096 & n22100 ) ;
  assign n22103 = n22089 | n22100 ;
  assign n22105 = ( n22102 & ~n22104 ) | ( n22102 & n22103 ) | ( ~n22104 & n22103 ) ;
  assign n22109 = n21878 &  n22095 ;
  assign n22110 = n22094 &  n22109 ;
  assign n22097 = x89 | n21878 ;
  assign n22098 = x89 &  n21878 ;
  assign n22099 = ( n22097 & ~n22098 ) | ( n22097 & 1'b0 ) | ( ~n22098 & 1'b0 ) ;
  assign n22112 = ( n22088 & n22096 ) | ( n22088 & n22099 ) | ( n22096 & n22099 ) ;
  assign n22111 = n22088 | n22099 ;
  assign n22113 = ( n22110 & ~n22112 ) | ( n22110 & n22111 ) | ( ~n22112 & n22111 ) ;
  assign n22117 = n21886 &  n22095 ;
  assign n22118 = n22094 &  n22117 ;
  assign n22106 = x88 | n21886 ;
  assign n22107 = x88 &  n21886 ;
  assign n22108 = ( n22106 & ~n22107 ) | ( n22106 & 1'b0 ) | ( ~n22107 & 1'b0 ) ;
  assign n22120 = ( n22087 & n22096 ) | ( n22087 & n22108 ) | ( n22096 & n22108 ) ;
  assign n22119 = n22087 | n22108 ;
  assign n22121 = ( n22118 & ~n22120 ) | ( n22118 & n22119 ) | ( ~n22120 & n22119 ) ;
  assign n22125 = n21894 &  n22095 ;
  assign n22126 = n22094 &  n22125 ;
  assign n22114 = x87 | n21894 ;
  assign n22115 = x87 &  n21894 ;
  assign n22116 = ( n22114 & ~n22115 ) | ( n22114 & 1'b0 ) | ( ~n22115 & 1'b0 ) ;
  assign n22128 = ( n22086 & n22096 ) | ( n22086 & n22116 ) | ( n22096 & n22116 ) ;
  assign n22127 = n22086 | n22116 ;
  assign n22129 = ( n22126 & ~n22128 ) | ( n22126 & n22127 ) | ( ~n22128 & n22127 ) ;
  assign n22133 = n21902 &  n22095 ;
  assign n22134 = n22094 &  n22133 ;
  assign n22122 = x86 | n21902 ;
  assign n22123 = x86 &  n21902 ;
  assign n22124 = ( n22122 & ~n22123 ) | ( n22122 & 1'b0 ) | ( ~n22123 & 1'b0 ) ;
  assign n22136 = ( n22085 & n22096 ) | ( n22085 & n22124 ) | ( n22096 & n22124 ) ;
  assign n22135 = n22085 | n22124 ;
  assign n22137 = ( n22134 & ~n22136 ) | ( n22134 & n22135 ) | ( ~n22136 & n22135 ) ;
  assign n22141 = n21910 &  n22095 ;
  assign n22142 = n22094 &  n22141 ;
  assign n22130 = x85 | n21910 ;
  assign n22131 = x85 &  n21910 ;
  assign n22132 = ( n22130 & ~n22131 ) | ( n22130 & 1'b0 ) | ( ~n22131 & 1'b0 ) ;
  assign n22144 = ( n22084 & n22096 ) | ( n22084 & n22132 ) | ( n22096 & n22132 ) ;
  assign n22143 = n22084 | n22132 ;
  assign n22145 = ( n22142 & ~n22144 ) | ( n22142 & n22143 ) | ( ~n22144 & n22143 ) ;
  assign n22149 = n21918 &  n22095 ;
  assign n22150 = n22094 &  n22149 ;
  assign n22138 = x84 | n21918 ;
  assign n22139 = x84 &  n21918 ;
  assign n22140 = ( n22138 & ~n22139 ) | ( n22138 & 1'b0 ) | ( ~n22139 & 1'b0 ) ;
  assign n22152 = ( n22083 & n22096 ) | ( n22083 & n22140 ) | ( n22096 & n22140 ) ;
  assign n22151 = n22083 | n22140 ;
  assign n22153 = ( n22150 & ~n22152 ) | ( n22150 & n22151 ) | ( ~n22152 & n22151 ) ;
  assign n22157 = n21926 &  n22095 ;
  assign n22158 = n22094 &  n22157 ;
  assign n22146 = x83 | n21926 ;
  assign n22147 = x83 &  n21926 ;
  assign n22148 = ( n22146 & ~n22147 ) | ( n22146 & 1'b0 ) | ( ~n22147 & 1'b0 ) ;
  assign n22160 = ( n22082 & n22096 ) | ( n22082 & n22148 ) | ( n22096 & n22148 ) ;
  assign n22159 = n22082 | n22148 ;
  assign n22161 = ( n22158 & ~n22160 ) | ( n22158 & n22159 ) | ( ~n22160 & n22159 ) ;
  assign n22165 = n21934 &  n22095 ;
  assign n22166 = n22094 &  n22165 ;
  assign n22154 = x82 | n21934 ;
  assign n22155 = x82 &  n21934 ;
  assign n22156 = ( n22154 & ~n22155 ) | ( n22154 & 1'b0 ) | ( ~n22155 & 1'b0 ) ;
  assign n22168 = ( n22081 & n22096 ) | ( n22081 & n22156 ) | ( n22096 & n22156 ) ;
  assign n22167 = n22081 | n22156 ;
  assign n22169 = ( n22166 & ~n22168 ) | ( n22166 & n22167 ) | ( ~n22168 & n22167 ) ;
  assign n22173 = n21942 &  n22095 ;
  assign n22174 = n22094 &  n22173 ;
  assign n22162 = x81 | n21942 ;
  assign n22163 = x81 &  n21942 ;
  assign n22164 = ( n22162 & ~n22163 ) | ( n22162 & 1'b0 ) | ( ~n22163 & 1'b0 ) ;
  assign n22176 = ( n22080 & n22096 ) | ( n22080 & n22164 ) | ( n22096 & n22164 ) ;
  assign n22175 = n22080 | n22164 ;
  assign n22177 = ( n22174 & ~n22176 ) | ( n22174 & n22175 ) | ( ~n22176 & n22175 ) ;
  assign n22181 = n21950 &  n22095 ;
  assign n22182 = n22094 &  n22181 ;
  assign n22170 = x80 | n21950 ;
  assign n22171 = x80 &  n21950 ;
  assign n22172 = ( n22170 & ~n22171 ) | ( n22170 & 1'b0 ) | ( ~n22171 & 1'b0 ) ;
  assign n22184 = ( n22079 & n22096 ) | ( n22079 & n22172 ) | ( n22096 & n22172 ) ;
  assign n22183 = n22079 | n22172 ;
  assign n22185 = ( n22182 & ~n22184 ) | ( n22182 & n22183 ) | ( ~n22184 & n22183 ) ;
  assign n22189 = n21958 &  n22095 ;
  assign n22190 = n22094 &  n22189 ;
  assign n22178 = x79 | n21958 ;
  assign n22179 = x79 &  n21958 ;
  assign n22180 = ( n22178 & ~n22179 ) | ( n22178 & 1'b0 ) | ( ~n22179 & 1'b0 ) ;
  assign n22192 = ( n22078 & n22096 ) | ( n22078 & n22180 ) | ( n22096 & n22180 ) ;
  assign n22191 = n22078 | n22180 ;
  assign n22193 = ( n22190 & ~n22192 ) | ( n22190 & n22191 ) | ( ~n22192 & n22191 ) ;
  assign n22197 = n21966 &  n22095 ;
  assign n22198 = n22094 &  n22197 ;
  assign n22186 = x78 | n21966 ;
  assign n22187 = x78 &  n21966 ;
  assign n22188 = ( n22186 & ~n22187 ) | ( n22186 & 1'b0 ) | ( ~n22187 & 1'b0 ) ;
  assign n22200 = ( n22077 & n22096 ) | ( n22077 & n22188 ) | ( n22096 & n22188 ) ;
  assign n22199 = n22077 | n22188 ;
  assign n22201 = ( n22198 & ~n22200 ) | ( n22198 & n22199 ) | ( ~n22200 & n22199 ) ;
  assign n22205 = n21974 &  n22095 ;
  assign n22206 = n22094 &  n22205 ;
  assign n22194 = x77 | n21974 ;
  assign n22195 = x77 &  n21974 ;
  assign n22196 = ( n22194 & ~n22195 ) | ( n22194 & 1'b0 ) | ( ~n22195 & 1'b0 ) ;
  assign n22208 = ( n22076 & n22096 ) | ( n22076 & n22196 ) | ( n22096 & n22196 ) ;
  assign n22207 = n22076 | n22196 ;
  assign n22209 = ( n22206 & ~n22208 ) | ( n22206 & n22207 ) | ( ~n22208 & n22207 ) ;
  assign n22213 = n21982 &  n22095 ;
  assign n22214 = n22094 &  n22213 ;
  assign n22202 = x76 | n21982 ;
  assign n22203 = x76 &  n21982 ;
  assign n22204 = ( n22202 & ~n22203 ) | ( n22202 & 1'b0 ) | ( ~n22203 & 1'b0 ) ;
  assign n22216 = ( n22075 & n22096 ) | ( n22075 & n22204 ) | ( n22096 & n22204 ) ;
  assign n22215 = n22075 | n22204 ;
  assign n22217 = ( n22214 & ~n22216 ) | ( n22214 & n22215 ) | ( ~n22216 & n22215 ) ;
  assign n22221 = n21990 &  n22095 ;
  assign n22222 = n22094 &  n22221 ;
  assign n22210 = x75 | n21990 ;
  assign n22211 = x75 &  n21990 ;
  assign n22212 = ( n22210 & ~n22211 ) | ( n22210 & 1'b0 ) | ( ~n22211 & 1'b0 ) ;
  assign n22224 = ( n22074 & n22096 ) | ( n22074 & n22212 ) | ( n22096 & n22212 ) ;
  assign n22223 = n22074 | n22212 ;
  assign n22225 = ( n22222 & ~n22224 ) | ( n22222 & n22223 ) | ( ~n22224 & n22223 ) ;
  assign n22229 = n21998 &  n22095 ;
  assign n22230 = n22094 &  n22229 ;
  assign n22218 = x74 | n21998 ;
  assign n22219 = x74 &  n21998 ;
  assign n22220 = ( n22218 & ~n22219 ) | ( n22218 & 1'b0 ) | ( ~n22219 & 1'b0 ) ;
  assign n22232 = ( n22073 & n22096 ) | ( n22073 & n22220 ) | ( n22096 & n22220 ) ;
  assign n22231 = n22073 | n22220 ;
  assign n22233 = ( n22230 & ~n22232 ) | ( n22230 & n22231 ) | ( ~n22232 & n22231 ) ;
  assign n22237 = n22006 &  n22095 ;
  assign n22238 = n22094 &  n22237 ;
  assign n22226 = x73 | n22006 ;
  assign n22227 = x73 &  n22006 ;
  assign n22228 = ( n22226 & ~n22227 ) | ( n22226 & 1'b0 ) | ( ~n22227 & 1'b0 ) ;
  assign n22240 = ( n22072 & n22096 ) | ( n22072 & n22228 ) | ( n22096 & n22228 ) ;
  assign n22239 = n22072 | n22228 ;
  assign n22241 = ( n22238 & ~n22240 ) | ( n22238 & n22239 ) | ( ~n22240 & n22239 ) ;
  assign n22245 = n22014 &  n22095 ;
  assign n22246 = n22094 &  n22245 ;
  assign n22234 = x72 | n22014 ;
  assign n22235 = x72 &  n22014 ;
  assign n22236 = ( n22234 & ~n22235 ) | ( n22234 & 1'b0 ) | ( ~n22235 & 1'b0 ) ;
  assign n22248 = ( n22071 & n22096 ) | ( n22071 & n22236 ) | ( n22096 & n22236 ) ;
  assign n22247 = n22071 | n22236 ;
  assign n22249 = ( n22246 & ~n22248 ) | ( n22246 & n22247 ) | ( ~n22248 & n22247 ) ;
  assign n22253 = n22022 &  n22095 ;
  assign n22254 = n22094 &  n22253 ;
  assign n22242 = x71 | n22022 ;
  assign n22243 = x71 &  n22022 ;
  assign n22244 = ( n22242 & ~n22243 ) | ( n22242 & 1'b0 ) | ( ~n22243 & 1'b0 ) ;
  assign n22256 = ( n22070 & n22096 ) | ( n22070 & n22244 ) | ( n22096 & n22244 ) ;
  assign n22255 = n22070 | n22244 ;
  assign n22257 = ( n22254 & ~n22256 ) | ( n22254 & n22255 ) | ( ~n22256 & n22255 ) ;
  assign n22261 = n22030 &  n22095 ;
  assign n22262 = n22094 &  n22261 ;
  assign n22250 = x70 | n22030 ;
  assign n22251 = x70 &  n22030 ;
  assign n22252 = ( n22250 & ~n22251 ) | ( n22250 & 1'b0 ) | ( ~n22251 & 1'b0 ) ;
  assign n22264 = ( n22069 & n22096 ) | ( n22069 & n22252 ) | ( n22096 & n22252 ) ;
  assign n22263 = n22069 | n22252 ;
  assign n22265 = ( n22262 & ~n22264 ) | ( n22262 & n22263 ) | ( ~n22264 & n22263 ) ;
  assign n22269 = n22038 &  n22095 ;
  assign n22270 = n22094 &  n22269 ;
  assign n22258 = x69 | n22038 ;
  assign n22259 = x69 &  n22038 ;
  assign n22260 = ( n22258 & ~n22259 ) | ( n22258 & 1'b0 ) | ( ~n22259 & 1'b0 ) ;
  assign n22272 = ( n22068 & n22096 ) | ( n22068 & n22260 ) | ( n22096 & n22260 ) ;
  assign n22271 = n22068 | n22260 ;
  assign n22273 = ( n22270 & ~n22272 ) | ( n22270 & n22271 ) | ( ~n22272 & n22271 ) ;
  assign n22277 = n22046 &  n22095 ;
  assign n22278 = n22094 &  n22277 ;
  assign n22266 = x68 | n22046 ;
  assign n22267 = x68 &  n22046 ;
  assign n22268 = ( n22266 & ~n22267 ) | ( n22266 & 1'b0 ) | ( ~n22267 & 1'b0 ) ;
  assign n22280 = ( n22067 & n22096 ) | ( n22067 & n22268 ) | ( n22096 & n22268 ) ;
  assign n22279 = n22067 | n22268 ;
  assign n22281 = ( n22278 & ~n22280 ) | ( n22278 & n22279 ) | ( ~n22280 & n22279 ) ;
  assign n22285 = n22054 &  n22095 ;
  assign n22286 = n22094 &  n22285 ;
  assign n22274 = x67 | n22054 ;
  assign n22275 = x67 &  n22054 ;
  assign n22276 = ( n22274 & ~n22275 ) | ( n22274 & 1'b0 ) | ( ~n22275 & 1'b0 ) ;
  assign n22288 = ( n22066 & n22096 ) | ( n22066 & n22276 ) | ( n22096 & n22276 ) ;
  assign n22287 = n22066 | n22276 ;
  assign n22289 = ( n22286 & ~n22288 ) | ( n22286 & n22287 ) | ( ~n22288 & n22287 ) ;
  assign n22290 = n22060 &  n22095 ;
  assign n22291 = n22094 &  n22290 ;
  assign n22282 = x66 | n22060 ;
  assign n22283 = x66 &  n22060 ;
  assign n22284 = ( n22282 & ~n22283 ) | ( n22282 & 1'b0 ) | ( ~n22283 & 1'b0 ) ;
  assign n22293 = ( n22065 & n22096 ) | ( n22065 & n22284 ) | ( n22096 & n22284 ) ;
  assign n22292 = n22065 | n22284 ;
  assign n22294 = ( n22291 & ~n22293 ) | ( n22291 & n22292 ) | ( ~n22293 & n22292 ) ;
  assign n22295 = ( x65 & ~n3437 ) | ( x65 & n22064 ) | ( ~n3437 & n22064 ) ;
  assign n22296 = ( n22065 & ~x65 ) | ( n22065 & n22295 ) | ( ~x65 & n22295 ) ;
  assign n22297 = ~n22096 & n22296 ;
  assign n22298 = n22064 &  n22095 ;
  assign n22299 = n22094 &  n22298 ;
  assign n22300 = n22297 | n22299 ;
  assign n22301 = ( x64 & ~n22096 ) | ( x64 & 1'b0 ) | ( ~n22096 & 1'b0 ) ;
  assign n22302 = ( x37 & ~n22301 ) | ( x37 & 1'b0 ) | ( ~n22301 & 1'b0 ) ;
  assign n22303 = ( n3437 & ~n22096 ) | ( n3437 & 1'b0 ) | ( ~n22096 & 1'b0 ) ;
  assign n22304 = n22302 | n22303 ;
  assign n22305 = ( x65 & ~n22304 ) | ( x65 & n3844 ) | ( ~n22304 & n3844 ) ;
  assign n22306 = ( x66 & ~n22300 ) | ( x66 & n22305 ) | ( ~n22300 & n22305 ) ;
  assign n22307 = ( x67 & ~n22294 ) | ( x67 & n22306 ) | ( ~n22294 & n22306 ) ;
  assign n22308 = ( x68 & ~n22289 ) | ( x68 & n22307 ) | ( ~n22289 & n22307 ) ;
  assign n22309 = ( x69 & ~n22281 ) | ( x69 & n22308 ) | ( ~n22281 & n22308 ) ;
  assign n22310 = ( x70 & ~n22273 ) | ( x70 & n22309 ) | ( ~n22273 & n22309 ) ;
  assign n22311 = ( x71 & ~n22265 ) | ( x71 & n22310 ) | ( ~n22265 & n22310 ) ;
  assign n22312 = ( x72 & ~n22257 ) | ( x72 & n22311 ) | ( ~n22257 & n22311 ) ;
  assign n22313 = ( x73 & ~n22249 ) | ( x73 & n22312 ) | ( ~n22249 & n22312 ) ;
  assign n22314 = ( x74 & ~n22241 ) | ( x74 & n22313 ) | ( ~n22241 & n22313 ) ;
  assign n22315 = ( x75 & ~n22233 ) | ( x75 & n22314 ) | ( ~n22233 & n22314 ) ;
  assign n22316 = ( x76 & ~n22225 ) | ( x76 & n22315 ) | ( ~n22225 & n22315 ) ;
  assign n22317 = ( x77 & ~n22217 ) | ( x77 & n22316 ) | ( ~n22217 & n22316 ) ;
  assign n22318 = ( x78 & ~n22209 ) | ( x78 & n22317 ) | ( ~n22209 & n22317 ) ;
  assign n22319 = ( x79 & ~n22201 ) | ( x79 & n22318 ) | ( ~n22201 & n22318 ) ;
  assign n22320 = ( x80 & ~n22193 ) | ( x80 & n22319 ) | ( ~n22193 & n22319 ) ;
  assign n22321 = ( x81 & ~n22185 ) | ( x81 & n22320 ) | ( ~n22185 & n22320 ) ;
  assign n22322 = ( x82 & ~n22177 ) | ( x82 & n22321 ) | ( ~n22177 & n22321 ) ;
  assign n22323 = ( x83 & ~n22169 ) | ( x83 & n22322 ) | ( ~n22169 & n22322 ) ;
  assign n22324 = ( x84 & ~n22161 ) | ( x84 & n22323 ) | ( ~n22161 & n22323 ) ;
  assign n22325 = ( x85 & ~n22153 ) | ( x85 & n22324 ) | ( ~n22153 & n22324 ) ;
  assign n22326 = ( x86 & ~n22145 ) | ( x86 & n22325 ) | ( ~n22145 & n22325 ) ;
  assign n22327 = ( x87 & ~n22137 ) | ( x87 & n22326 ) | ( ~n22137 & n22326 ) ;
  assign n22328 = ( x88 & ~n22129 ) | ( x88 & n22327 ) | ( ~n22129 & n22327 ) ;
  assign n22329 = ( x89 & ~n22121 ) | ( x89 & n22328 ) | ( ~n22121 & n22328 ) ;
  assign n22330 = ( x90 & ~n22113 ) | ( x90 & n22329 ) | ( ~n22113 & n22329 ) ;
  assign n22337 = ( x91 & ~n3873 ) | ( x91 & n22330 ) | ( ~n3873 & n22330 ) ;
  assign n22336 = x91 &  n22330 ;
  assign n22338 = ( n22105 & ~n22337 ) | ( n22105 & n22336 ) | ( ~n22337 & n22336 ) ;
  assign n22331 = ( x91 & ~n22105 ) | ( x91 & n22330 ) | ( ~n22105 & n22330 ) ;
  assign n22332 = n3873 | n22331 ;
  assign n22339 = n22113 &  n22332 ;
  assign n22333 = x90 | n22113 ;
  assign n22334 = x90 &  n22113 ;
  assign n22335 = ( n22333 & ~n22334 ) | ( n22333 & 1'b0 ) | ( ~n22334 & 1'b0 ) ;
  assign n22343 = ( n3873 & n22329 ) | ( n3873 & n22335 ) | ( n22329 & n22335 ) ;
  assign n22344 = ( n22329 & ~n22331 ) | ( n22329 & n22335 ) | ( ~n22331 & n22335 ) ;
  assign n22345 = ~n22343 & n22344 ;
  assign n22346 = n22339 | n22345 ;
  assign n22347 = n22121 &  n22332 ;
  assign n22340 = x89 | n22121 ;
  assign n22341 = x89 &  n22121 ;
  assign n22342 = ( n22340 & ~n22341 ) | ( n22340 & 1'b0 ) | ( ~n22341 & 1'b0 ) ;
  assign n22351 = ( n3873 & n22328 ) | ( n3873 & n22342 ) | ( n22328 & n22342 ) ;
  assign n22352 = ( n22328 & ~n22331 ) | ( n22328 & n22342 ) | ( ~n22331 & n22342 ) ;
  assign n22353 = ~n22351 & n22352 ;
  assign n22354 = n22347 | n22353 ;
  assign n22355 = n22129 &  n22332 ;
  assign n22348 = x88 | n22129 ;
  assign n22349 = x88 &  n22129 ;
  assign n22350 = ( n22348 & ~n22349 ) | ( n22348 & 1'b0 ) | ( ~n22349 & 1'b0 ) ;
  assign n22359 = ( n3873 & n22327 ) | ( n3873 & n22350 ) | ( n22327 & n22350 ) ;
  assign n22360 = ( n22327 & ~n22331 ) | ( n22327 & n22350 ) | ( ~n22331 & n22350 ) ;
  assign n22361 = ~n22359 & n22360 ;
  assign n22362 = n22355 | n22361 ;
  assign n22363 = n22137 &  n22332 ;
  assign n22356 = x87 | n22137 ;
  assign n22357 = x87 &  n22137 ;
  assign n22358 = ( n22356 & ~n22357 ) | ( n22356 & 1'b0 ) | ( ~n22357 & 1'b0 ) ;
  assign n22367 = ( n3873 & n22326 ) | ( n3873 & n22358 ) | ( n22326 & n22358 ) ;
  assign n22368 = ( n22326 & ~n22331 ) | ( n22326 & n22358 ) | ( ~n22331 & n22358 ) ;
  assign n22369 = ~n22367 & n22368 ;
  assign n22370 = n22363 | n22369 ;
  assign n22371 = n22145 &  n22332 ;
  assign n22364 = x86 | n22145 ;
  assign n22365 = x86 &  n22145 ;
  assign n22366 = ( n22364 & ~n22365 ) | ( n22364 & 1'b0 ) | ( ~n22365 & 1'b0 ) ;
  assign n22375 = ( n3873 & n22325 ) | ( n3873 & n22366 ) | ( n22325 & n22366 ) ;
  assign n22376 = ( n22325 & ~n22331 ) | ( n22325 & n22366 ) | ( ~n22331 & n22366 ) ;
  assign n22377 = ~n22375 & n22376 ;
  assign n22378 = n22371 | n22377 ;
  assign n22379 = n22153 &  n22332 ;
  assign n22372 = x85 | n22153 ;
  assign n22373 = x85 &  n22153 ;
  assign n22374 = ( n22372 & ~n22373 ) | ( n22372 & 1'b0 ) | ( ~n22373 & 1'b0 ) ;
  assign n22383 = ( n3873 & n22324 ) | ( n3873 & n22374 ) | ( n22324 & n22374 ) ;
  assign n22384 = ( n22324 & ~n22331 ) | ( n22324 & n22374 ) | ( ~n22331 & n22374 ) ;
  assign n22385 = ~n22383 & n22384 ;
  assign n22386 = n22379 | n22385 ;
  assign n22387 = n22161 &  n22332 ;
  assign n22380 = x84 | n22161 ;
  assign n22381 = x84 &  n22161 ;
  assign n22382 = ( n22380 & ~n22381 ) | ( n22380 & 1'b0 ) | ( ~n22381 & 1'b0 ) ;
  assign n22391 = ( n3873 & n22323 ) | ( n3873 & n22382 ) | ( n22323 & n22382 ) ;
  assign n22392 = ( n22323 & ~n22331 ) | ( n22323 & n22382 ) | ( ~n22331 & n22382 ) ;
  assign n22393 = ~n22391 & n22392 ;
  assign n22394 = n22387 | n22393 ;
  assign n22395 = n22169 &  n22332 ;
  assign n22388 = x83 | n22169 ;
  assign n22389 = x83 &  n22169 ;
  assign n22390 = ( n22388 & ~n22389 ) | ( n22388 & 1'b0 ) | ( ~n22389 & 1'b0 ) ;
  assign n22399 = ( n3873 & n22322 ) | ( n3873 & n22390 ) | ( n22322 & n22390 ) ;
  assign n22400 = ( n22322 & ~n22331 ) | ( n22322 & n22390 ) | ( ~n22331 & n22390 ) ;
  assign n22401 = ~n22399 & n22400 ;
  assign n22402 = n22395 | n22401 ;
  assign n22403 = n22177 &  n22332 ;
  assign n22396 = x82 | n22177 ;
  assign n22397 = x82 &  n22177 ;
  assign n22398 = ( n22396 & ~n22397 ) | ( n22396 & 1'b0 ) | ( ~n22397 & 1'b0 ) ;
  assign n22407 = ( n3873 & n22321 ) | ( n3873 & n22398 ) | ( n22321 & n22398 ) ;
  assign n22408 = ( n22321 & ~n22331 ) | ( n22321 & n22398 ) | ( ~n22331 & n22398 ) ;
  assign n22409 = ~n22407 & n22408 ;
  assign n22410 = n22403 | n22409 ;
  assign n22411 = n22185 &  n22332 ;
  assign n22404 = x81 | n22185 ;
  assign n22405 = x81 &  n22185 ;
  assign n22406 = ( n22404 & ~n22405 ) | ( n22404 & 1'b0 ) | ( ~n22405 & 1'b0 ) ;
  assign n22415 = ( n3873 & n22320 ) | ( n3873 & n22406 ) | ( n22320 & n22406 ) ;
  assign n22416 = ( n22320 & ~n22331 ) | ( n22320 & n22406 ) | ( ~n22331 & n22406 ) ;
  assign n22417 = ~n22415 & n22416 ;
  assign n22418 = n22411 | n22417 ;
  assign n22419 = n22193 &  n22332 ;
  assign n22412 = x80 | n22193 ;
  assign n22413 = x80 &  n22193 ;
  assign n22414 = ( n22412 & ~n22413 ) | ( n22412 & 1'b0 ) | ( ~n22413 & 1'b0 ) ;
  assign n22423 = ( n3873 & n22319 ) | ( n3873 & n22414 ) | ( n22319 & n22414 ) ;
  assign n22424 = ( n22319 & ~n22331 ) | ( n22319 & n22414 ) | ( ~n22331 & n22414 ) ;
  assign n22425 = ~n22423 & n22424 ;
  assign n22426 = n22419 | n22425 ;
  assign n22427 = n22201 &  n22332 ;
  assign n22420 = x79 | n22201 ;
  assign n22421 = x79 &  n22201 ;
  assign n22422 = ( n22420 & ~n22421 ) | ( n22420 & 1'b0 ) | ( ~n22421 & 1'b0 ) ;
  assign n22431 = ( n3873 & n22318 ) | ( n3873 & n22422 ) | ( n22318 & n22422 ) ;
  assign n22432 = ( n22318 & ~n22331 ) | ( n22318 & n22422 ) | ( ~n22331 & n22422 ) ;
  assign n22433 = ~n22431 & n22432 ;
  assign n22434 = n22427 | n22433 ;
  assign n22435 = n22209 &  n22332 ;
  assign n22428 = x78 | n22209 ;
  assign n22429 = x78 &  n22209 ;
  assign n22430 = ( n22428 & ~n22429 ) | ( n22428 & 1'b0 ) | ( ~n22429 & 1'b0 ) ;
  assign n22439 = ( n3873 & n22317 ) | ( n3873 & n22430 ) | ( n22317 & n22430 ) ;
  assign n22440 = ( n22317 & ~n22331 ) | ( n22317 & n22430 ) | ( ~n22331 & n22430 ) ;
  assign n22441 = ~n22439 & n22440 ;
  assign n22442 = n22435 | n22441 ;
  assign n22443 = n22217 &  n22332 ;
  assign n22436 = x77 | n22217 ;
  assign n22437 = x77 &  n22217 ;
  assign n22438 = ( n22436 & ~n22437 ) | ( n22436 & 1'b0 ) | ( ~n22437 & 1'b0 ) ;
  assign n22447 = ( n3873 & n22316 ) | ( n3873 & n22438 ) | ( n22316 & n22438 ) ;
  assign n22448 = ( n22316 & ~n22331 ) | ( n22316 & n22438 ) | ( ~n22331 & n22438 ) ;
  assign n22449 = ~n22447 & n22448 ;
  assign n22450 = n22443 | n22449 ;
  assign n22451 = n22225 &  n22332 ;
  assign n22444 = x76 | n22225 ;
  assign n22445 = x76 &  n22225 ;
  assign n22446 = ( n22444 & ~n22445 ) | ( n22444 & 1'b0 ) | ( ~n22445 & 1'b0 ) ;
  assign n22455 = ( n3873 & n22315 ) | ( n3873 & n22446 ) | ( n22315 & n22446 ) ;
  assign n22456 = ( n22315 & ~n22331 ) | ( n22315 & n22446 ) | ( ~n22331 & n22446 ) ;
  assign n22457 = ~n22455 & n22456 ;
  assign n22458 = n22451 | n22457 ;
  assign n22459 = n22233 &  n22332 ;
  assign n22452 = x75 | n22233 ;
  assign n22453 = x75 &  n22233 ;
  assign n22454 = ( n22452 & ~n22453 ) | ( n22452 & 1'b0 ) | ( ~n22453 & 1'b0 ) ;
  assign n22463 = ( n3873 & n22314 ) | ( n3873 & n22454 ) | ( n22314 & n22454 ) ;
  assign n22464 = ( n22314 & ~n22331 ) | ( n22314 & n22454 ) | ( ~n22331 & n22454 ) ;
  assign n22465 = ~n22463 & n22464 ;
  assign n22466 = n22459 | n22465 ;
  assign n22467 = n22241 &  n22332 ;
  assign n22460 = x74 | n22241 ;
  assign n22461 = x74 &  n22241 ;
  assign n22462 = ( n22460 & ~n22461 ) | ( n22460 & 1'b0 ) | ( ~n22461 & 1'b0 ) ;
  assign n22471 = ( n3873 & n22313 ) | ( n3873 & n22462 ) | ( n22313 & n22462 ) ;
  assign n22472 = ( n22313 & ~n22331 ) | ( n22313 & n22462 ) | ( ~n22331 & n22462 ) ;
  assign n22473 = ~n22471 & n22472 ;
  assign n22474 = n22467 | n22473 ;
  assign n22475 = n22249 &  n22332 ;
  assign n22468 = x73 | n22249 ;
  assign n22469 = x73 &  n22249 ;
  assign n22470 = ( n22468 & ~n22469 ) | ( n22468 & 1'b0 ) | ( ~n22469 & 1'b0 ) ;
  assign n22479 = ( n3873 & n22312 ) | ( n3873 & n22470 ) | ( n22312 & n22470 ) ;
  assign n22480 = ( n22312 & ~n22331 ) | ( n22312 & n22470 ) | ( ~n22331 & n22470 ) ;
  assign n22481 = ~n22479 & n22480 ;
  assign n22482 = n22475 | n22481 ;
  assign n22483 = n22257 &  n22332 ;
  assign n22476 = x72 | n22257 ;
  assign n22477 = x72 &  n22257 ;
  assign n22478 = ( n22476 & ~n22477 ) | ( n22476 & 1'b0 ) | ( ~n22477 & 1'b0 ) ;
  assign n22487 = ( n3873 & n22311 ) | ( n3873 & n22478 ) | ( n22311 & n22478 ) ;
  assign n22488 = ( n22311 & ~n22331 ) | ( n22311 & n22478 ) | ( ~n22331 & n22478 ) ;
  assign n22489 = ~n22487 & n22488 ;
  assign n22490 = n22483 | n22489 ;
  assign n22491 = n22265 &  n22332 ;
  assign n22484 = x71 | n22265 ;
  assign n22485 = x71 &  n22265 ;
  assign n22486 = ( n22484 & ~n22485 ) | ( n22484 & 1'b0 ) | ( ~n22485 & 1'b0 ) ;
  assign n22495 = ( n3873 & n22310 ) | ( n3873 & n22486 ) | ( n22310 & n22486 ) ;
  assign n22496 = ( n22310 & ~n22331 ) | ( n22310 & n22486 ) | ( ~n22331 & n22486 ) ;
  assign n22497 = ~n22495 & n22496 ;
  assign n22498 = n22491 | n22497 ;
  assign n22499 = n22273 &  n22332 ;
  assign n22492 = x70 | n22273 ;
  assign n22493 = x70 &  n22273 ;
  assign n22494 = ( n22492 & ~n22493 ) | ( n22492 & 1'b0 ) | ( ~n22493 & 1'b0 ) ;
  assign n22503 = ( n3873 & n22309 ) | ( n3873 & n22494 ) | ( n22309 & n22494 ) ;
  assign n22504 = ( n22309 & ~n22331 ) | ( n22309 & n22494 ) | ( ~n22331 & n22494 ) ;
  assign n22505 = ~n22503 & n22504 ;
  assign n22506 = n22499 | n22505 ;
  assign n22507 = n22281 &  n22332 ;
  assign n22500 = x69 | n22281 ;
  assign n22501 = x69 &  n22281 ;
  assign n22502 = ( n22500 & ~n22501 ) | ( n22500 & 1'b0 ) | ( ~n22501 & 1'b0 ) ;
  assign n22511 = ( n3873 & n22308 ) | ( n3873 & n22502 ) | ( n22308 & n22502 ) ;
  assign n22512 = ( n22308 & ~n22331 ) | ( n22308 & n22502 ) | ( ~n22331 & n22502 ) ;
  assign n22513 = ~n22511 & n22512 ;
  assign n22514 = n22507 | n22513 ;
  assign n22515 = n22289 &  n22332 ;
  assign n22508 = x68 | n22289 ;
  assign n22509 = x68 &  n22289 ;
  assign n22510 = ( n22508 & ~n22509 ) | ( n22508 & 1'b0 ) | ( ~n22509 & 1'b0 ) ;
  assign n22519 = ( n3873 & n22307 ) | ( n3873 & n22510 ) | ( n22307 & n22510 ) ;
  assign n22520 = ( n22307 & ~n22331 ) | ( n22307 & n22510 ) | ( ~n22331 & n22510 ) ;
  assign n22521 = ~n22519 & n22520 ;
  assign n22522 = n22515 | n22521 ;
  assign n22523 = n22294 &  n22332 ;
  assign n22516 = x67 | n22294 ;
  assign n22517 = x67 &  n22294 ;
  assign n22518 = ( n22516 & ~n22517 ) | ( n22516 & 1'b0 ) | ( ~n22517 & 1'b0 ) ;
  assign n22527 = ( n3873 & n22306 ) | ( n3873 & n22518 ) | ( n22306 & n22518 ) ;
  assign n22528 = ( n22306 & ~n22331 ) | ( n22306 & n22518 ) | ( ~n22331 & n22518 ) ;
  assign n22529 = ~n22527 & n22528 ;
  assign n22530 = n22523 | n22529 ;
  assign n22531 = n22300 &  n22332 ;
  assign n22524 = x66 | n22300 ;
  assign n22525 = x66 &  n22300 ;
  assign n22526 = ( n22524 & ~n22525 ) | ( n22524 & 1'b0 ) | ( ~n22525 & 1'b0 ) ;
  assign n22532 = ( n3873 & n22305 ) | ( n3873 & n22526 ) | ( n22305 & n22526 ) ;
  assign n22533 = ( n22305 & ~n22331 ) | ( n22305 & n22526 ) | ( ~n22331 & n22526 ) ;
  assign n22534 = ~n22532 & n22533 ;
  assign n22535 = n22531 | n22534 ;
  assign n22536 = n22304 &  n22332 ;
  assign n22537 = ( x65 & ~x37 ) | ( x65 & n22301 ) | ( ~x37 & n22301 ) ;
  assign n22538 = ( x37 & ~n22301 ) | ( x37 & x65 ) | ( ~n22301 & x65 ) ;
  assign n22539 = ( n22537 & ~x65 ) | ( n22537 & n22538 ) | ( ~x65 & n22538 ) ;
  assign n22540 = ( n3844 & ~n3873 ) | ( n3844 & n22539 ) | ( ~n3873 & n22539 ) ;
  assign n22541 = ( n3844 & n22331 ) | ( n3844 & n22539 ) | ( n22331 & n22539 ) ;
  assign n22542 = ( n22540 & ~n22541 ) | ( n22540 & 1'b0 ) | ( ~n22541 & 1'b0 ) ;
  assign n22543 = n22536 | n22542 ;
  assign n22544 = ( n4091 & ~n22331 ) | ( n4091 & 1'b0 ) | ( ~n22331 & 1'b0 ) ;
  assign n22545 = ( x36 & ~n22544 ) | ( x36 & 1'b0 ) | ( ~n22544 & 1'b0 ) ;
  assign n22546 = ( n4096 & ~n22331 ) | ( n4096 & 1'b0 ) | ( ~n22331 & 1'b0 ) ;
  assign n22547 = n22545 | n22546 ;
  assign n22548 = ( x65 & ~n22547 ) | ( x65 & n4099 ) | ( ~n22547 & n4099 ) ;
  assign n22549 = ( x66 & ~n22543 ) | ( x66 & n22548 ) | ( ~n22543 & n22548 ) ;
  assign n22550 = ( x67 & ~n22535 ) | ( x67 & n22549 ) | ( ~n22535 & n22549 ) ;
  assign n22551 = ( x68 & ~n22530 ) | ( x68 & n22550 ) | ( ~n22530 & n22550 ) ;
  assign n22552 = ( x69 & ~n22522 ) | ( x69 & n22551 ) | ( ~n22522 & n22551 ) ;
  assign n22553 = ( x70 & ~n22514 ) | ( x70 & n22552 ) | ( ~n22514 & n22552 ) ;
  assign n22554 = ( x71 & ~n22506 ) | ( x71 & n22553 ) | ( ~n22506 & n22553 ) ;
  assign n22555 = ( x72 & ~n22498 ) | ( x72 & n22554 ) | ( ~n22498 & n22554 ) ;
  assign n22556 = ( x73 & ~n22490 ) | ( x73 & n22555 ) | ( ~n22490 & n22555 ) ;
  assign n22557 = ( x74 & ~n22482 ) | ( x74 & n22556 ) | ( ~n22482 & n22556 ) ;
  assign n22558 = ( x75 & ~n22474 ) | ( x75 & n22557 ) | ( ~n22474 & n22557 ) ;
  assign n22559 = ( x76 & ~n22466 ) | ( x76 & n22558 ) | ( ~n22466 & n22558 ) ;
  assign n22560 = ( x77 & ~n22458 ) | ( x77 & n22559 ) | ( ~n22458 & n22559 ) ;
  assign n22561 = ( x78 & ~n22450 ) | ( x78 & n22560 ) | ( ~n22450 & n22560 ) ;
  assign n22562 = ( x79 & ~n22442 ) | ( x79 & n22561 ) | ( ~n22442 & n22561 ) ;
  assign n22563 = ( x80 & ~n22434 ) | ( x80 & n22562 ) | ( ~n22434 & n22562 ) ;
  assign n22564 = ( x81 & ~n22426 ) | ( x81 & n22563 ) | ( ~n22426 & n22563 ) ;
  assign n22565 = ( x82 & ~n22418 ) | ( x82 & n22564 ) | ( ~n22418 & n22564 ) ;
  assign n22566 = ( x83 & ~n22410 ) | ( x83 & n22565 ) | ( ~n22410 & n22565 ) ;
  assign n22567 = ( x84 & ~n22402 ) | ( x84 & n22566 ) | ( ~n22402 & n22566 ) ;
  assign n22568 = ( x85 & ~n22394 ) | ( x85 & n22567 ) | ( ~n22394 & n22567 ) ;
  assign n22569 = ( x86 & ~n22386 ) | ( x86 & n22568 ) | ( ~n22386 & n22568 ) ;
  assign n22570 = ( x87 & ~n22378 ) | ( x87 & n22569 ) | ( ~n22378 & n22569 ) ;
  assign n22571 = ( x88 & ~n22370 ) | ( x88 & n22570 ) | ( ~n22370 & n22570 ) ;
  assign n22572 = ( x89 & ~n22362 ) | ( x89 & n22571 ) | ( ~n22362 & n22571 ) ;
  assign n22573 = ( x90 & ~n22354 ) | ( x90 & n22572 ) | ( ~n22354 & n22572 ) ;
  assign n22574 = ( x91 & ~n22346 ) | ( x91 & n22573 ) | ( ~n22346 & n22573 ) ;
  assign n22575 = ( x92 & ~n22338 ) | ( x92 & n22574 ) | ( ~n22338 & n22574 ) ;
  assign n22576 = n4129 | n22575 ;
  assign n22577 = n22338 &  n22576 ;
  assign n22581 = ( n4129 & n22338 ) | ( n4129 & n22574 ) | ( n22338 & n22574 ) ;
  assign n22582 = ( x92 & ~n22581 ) | ( x92 & n22338 ) | ( ~n22581 & n22338 ) ;
  assign n22583 = ~x92 & n22582 ;
  assign n22584 = n22577 | n22583 ;
  assign n22585 = ~x93 & n22584 ;
  assign n22586 = n22346 &  n22576 ;
  assign n22578 = x91 | n22346 ;
  assign n22579 = x91 &  n22346 ;
  assign n22580 = ( n22578 & ~n22579 ) | ( n22578 & 1'b0 ) | ( ~n22579 & 1'b0 ) ;
  assign n22590 = ( n4129 & n22573 ) | ( n4129 & n22580 ) | ( n22573 & n22580 ) ;
  assign n22591 = ( n22573 & ~n22575 ) | ( n22573 & n22580 ) | ( ~n22575 & n22580 ) ;
  assign n22592 = ~n22590 & n22591 ;
  assign n22593 = n22586 | n22592 ;
  assign n22594 = n22354 &  n22576 ;
  assign n22587 = x90 | n22354 ;
  assign n22588 = x90 &  n22354 ;
  assign n22589 = ( n22587 & ~n22588 ) | ( n22587 & 1'b0 ) | ( ~n22588 & 1'b0 ) ;
  assign n22598 = ( n4129 & n22572 ) | ( n4129 & n22589 ) | ( n22572 & n22589 ) ;
  assign n22599 = ( n22572 & ~n22575 ) | ( n22572 & n22589 ) | ( ~n22575 & n22589 ) ;
  assign n22600 = ~n22598 & n22599 ;
  assign n22601 = n22594 | n22600 ;
  assign n22602 = n22362 &  n22576 ;
  assign n22595 = x89 | n22362 ;
  assign n22596 = x89 &  n22362 ;
  assign n22597 = ( n22595 & ~n22596 ) | ( n22595 & 1'b0 ) | ( ~n22596 & 1'b0 ) ;
  assign n22606 = ( n4129 & n22571 ) | ( n4129 & n22597 ) | ( n22571 & n22597 ) ;
  assign n22607 = ( n22571 & ~n22575 ) | ( n22571 & n22597 ) | ( ~n22575 & n22597 ) ;
  assign n22608 = ~n22606 & n22607 ;
  assign n22609 = n22602 | n22608 ;
  assign n22610 = n22370 &  n22576 ;
  assign n22603 = x88 | n22370 ;
  assign n22604 = x88 &  n22370 ;
  assign n22605 = ( n22603 & ~n22604 ) | ( n22603 & 1'b0 ) | ( ~n22604 & 1'b0 ) ;
  assign n22614 = ( n4129 & n22570 ) | ( n4129 & n22605 ) | ( n22570 & n22605 ) ;
  assign n22615 = ( n22570 & ~n22575 ) | ( n22570 & n22605 ) | ( ~n22575 & n22605 ) ;
  assign n22616 = ~n22614 & n22615 ;
  assign n22617 = n22610 | n22616 ;
  assign n22618 = n22378 &  n22576 ;
  assign n22611 = x87 | n22378 ;
  assign n22612 = x87 &  n22378 ;
  assign n22613 = ( n22611 & ~n22612 ) | ( n22611 & 1'b0 ) | ( ~n22612 & 1'b0 ) ;
  assign n22622 = ( n4129 & n22569 ) | ( n4129 & n22613 ) | ( n22569 & n22613 ) ;
  assign n22623 = ( n22569 & ~n22575 ) | ( n22569 & n22613 ) | ( ~n22575 & n22613 ) ;
  assign n22624 = ~n22622 & n22623 ;
  assign n22625 = n22618 | n22624 ;
  assign n22626 = n22386 &  n22576 ;
  assign n22619 = x86 | n22386 ;
  assign n22620 = x86 &  n22386 ;
  assign n22621 = ( n22619 & ~n22620 ) | ( n22619 & 1'b0 ) | ( ~n22620 & 1'b0 ) ;
  assign n22630 = ( n4129 & n22568 ) | ( n4129 & n22621 ) | ( n22568 & n22621 ) ;
  assign n22631 = ( n22568 & ~n22575 ) | ( n22568 & n22621 ) | ( ~n22575 & n22621 ) ;
  assign n22632 = ~n22630 & n22631 ;
  assign n22633 = n22626 | n22632 ;
  assign n22634 = n22394 &  n22576 ;
  assign n22627 = x85 | n22394 ;
  assign n22628 = x85 &  n22394 ;
  assign n22629 = ( n22627 & ~n22628 ) | ( n22627 & 1'b0 ) | ( ~n22628 & 1'b0 ) ;
  assign n22638 = ( n4129 & n22567 ) | ( n4129 & n22629 ) | ( n22567 & n22629 ) ;
  assign n22639 = ( n22567 & ~n22575 ) | ( n22567 & n22629 ) | ( ~n22575 & n22629 ) ;
  assign n22640 = ~n22638 & n22639 ;
  assign n22641 = n22634 | n22640 ;
  assign n22642 = n22402 &  n22576 ;
  assign n22635 = x84 | n22402 ;
  assign n22636 = x84 &  n22402 ;
  assign n22637 = ( n22635 & ~n22636 ) | ( n22635 & 1'b0 ) | ( ~n22636 & 1'b0 ) ;
  assign n22646 = ( n4129 & n22566 ) | ( n4129 & n22637 ) | ( n22566 & n22637 ) ;
  assign n22647 = ( n22566 & ~n22575 ) | ( n22566 & n22637 ) | ( ~n22575 & n22637 ) ;
  assign n22648 = ~n22646 & n22647 ;
  assign n22649 = n22642 | n22648 ;
  assign n22650 = n22410 &  n22576 ;
  assign n22643 = x83 | n22410 ;
  assign n22644 = x83 &  n22410 ;
  assign n22645 = ( n22643 & ~n22644 ) | ( n22643 & 1'b0 ) | ( ~n22644 & 1'b0 ) ;
  assign n22654 = ( n4129 & n22565 ) | ( n4129 & n22645 ) | ( n22565 & n22645 ) ;
  assign n22655 = ( n22565 & ~n22575 ) | ( n22565 & n22645 ) | ( ~n22575 & n22645 ) ;
  assign n22656 = ~n22654 & n22655 ;
  assign n22657 = n22650 | n22656 ;
  assign n22658 = n22418 &  n22576 ;
  assign n22651 = x82 | n22418 ;
  assign n22652 = x82 &  n22418 ;
  assign n22653 = ( n22651 & ~n22652 ) | ( n22651 & 1'b0 ) | ( ~n22652 & 1'b0 ) ;
  assign n22662 = ( n4129 & n22564 ) | ( n4129 & n22653 ) | ( n22564 & n22653 ) ;
  assign n22663 = ( n22564 & ~n22575 ) | ( n22564 & n22653 ) | ( ~n22575 & n22653 ) ;
  assign n22664 = ~n22662 & n22663 ;
  assign n22665 = n22658 | n22664 ;
  assign n22666 = n22426 &  n22576 ;
  assign n22659 = x81 | n22426 ;
  assign n22660 = x81 &  n22426 ;
  assign n22661 = ( n22659 & ~n22660 ) | ( n22659 & 1'b0 ) | ( ~n22660 & 1'b0 ) ;
  assign n22670 = ( n4129 & n22563 ) | ( n4129 & n22661 ) | ( n22563 & n22661 ) ;
  assign n22671 = ( n22563 & ~n22575 ) | ( n22563 & n22661 ) | ( ~n22575 & n22661 ) ;
  assign n22672 = ~n22670 & n22671 ;
  assign n22673 = n22666 | n22672 ;
  assign n22674 = n22434 &  n22576 ;
  assign n22667 = x80 | n22434 ;
  assign n22668 = x80 &  n22434 ;
  assign n22669 = ( n22667 & ~n22668 ) | ( n22667 & 1'b0 ) | ( ~n22668 & 1'b0 ) ;
  assign n22678 = ( n4129 & n22562 ) | ( n4129 & n22669 ) | ( n22562 & n22669 ) ;
  assign n22679 = ( n22562 & ~n22575 ) | ( n22562 & n22669 ) | ( ~n22575 & n22669 ) ;
  assign n22680 = ~n22678 & n22679 ;
  assign n22681 = n22674 | n22680 ;
  assign n22682 = n22442 &  n22576 ;
  assign n22675 = x79 | n22442 ;
  assign n22676 = x79 &  n22442 ;
  assign n22677 = ( n22675 & ~n22676 ) | ( n22675 & 1'b0 ) | ( ~n22676 & 1'b0 ) ;
  assign n22686 = ( n4129 & n22561 ) | ( n4129 & n22677 ) | ( n22561 & n22677 ) ;
  assign n22687 = ( n22561 & ~n22575 ) | ( n22561 & n22677 ) | ( ~n22575 & n22677 ) ;
  assign n22688 = ~n22686 & n22687 ;
  assign n22689 = n22682 | n22688 ;
  assign n22690 = n22450 &  n22576 ;
  assign n22683 = x78 | n22450 ;
  assign n22684 = x78 &  n22450 ;
  assign n22685 = ( n22683 & ~n22684 ) | ( n22683 & 1'b0 ) | ( ~n22684 & 1'b0 ) ;
  assign n22694 = ( n4129 & n22560 ) | ( n4129 & n22685 ) | ( n22560 & n22685 ) ;
  assign n22695 = ( n22560 & ~n22575 ) | ( n22560 & n22685 ) | ( ~n22575 & n22685 ) ;
  assign n22696 = ~n22694 & n22695 ;
  assign n22697 = n22690 | n22696 ;
  assign n22698 = n22458 &  n22576 ;
  assign n22691 = x77 | n22458 ;
  assign n22692 = x77 &  n22458 ;
  assign n22693 = ( n22691 & ~n22692 ) | ( n22691 & 1'b0 ) | ( ~n22692 & 1'b0 ) ;
  assign n22702 = ( n4129 & n22559 ) | ( n4129 & n22693 ) | ( n22559 & n22693 ) ;
  assign n22703 = ( n22559 & ~n22575 ) | ( n22559 & n22693 ) | ( ~n22575 & n22693 ) ;
  assign n22704 = ~n22702 & n22703 ;
  assign n22705 = n22698 | n22704 ;
  assign n22706 = n22466 &  n22576 ;
  assign n22699 = x76 | n22466 ;
  assign n22700 = x76 &  n22466 ;
  assign n22701 = ( n22699 & ~n22700 ) | ( n22699 & 1'b0 ) | ( ~n22700 & 1'b0 ) ;
  assign n22710 = ( n4129 & n22558 ) | ( n4129 & n22701 ) | ( n22558 & n22701 ) ;
  assign n22711 = ( n22558 & ~n22575 ) | ( n22558 & n22701 ) | ( ~n22575 & n22701 ) ;
  assign n22712 = ~n22710 & n22711 ;
  assign n22713 = n22706 | n22712 ;
  assign n22714 = n22474 &  n22576 ;
  assign n22707 = x75 | n22474 ;
  assign n22708 = x75 &  n22474 ;
  assign n22709 = ( n22707 & ~n22708 ) | ( n22707 & 1'b0 ) | ( ~n22708 & 1'b0 ) ;
  assign n22718 = ( n4129 & n22557 ) | ( n4129 & n22709 ) | ( n22557 & n22709 ) ;
  assign n22719 = ( n22557 & ~n22575 ) | ( n22557 & n22709 ) | ( ~n22575 & n22709 ) ;
  assign n22720 = ~n22718 & n22719 ;
  assign n22721 = n22714 | n22720 ;
  assign n22722 = n22482 &  n22576 ;
  assign n22715 = x74 | n22482 ;
  assign n22716 = x74 &  n22482 ;
  assign n22717 = ( n22715 & ~n22716 ) | ( n22715 & 1'b0 ) | ( ~n22716 & 1'b0 ) ;
  assign n22726 = ( n4129 & n22556 ) | ( n4129 & n22717 ) | ( n22556 & n22717 ) ;
  assign n22727 = ( n22556 & ~n22575 ) | ( n22556 & n22717 ) | ( ~n22575 & n22717 ) ;
  assign n22728 = ~n22726 & n22727 ;
  assign n22729 = n22722 | n22728 ;
  assign n22730 = n22490 &  n22576 ;
  assign n22723 = x73 | n22490 ;
  assign n22724 = x73 &  n22490 ;
  assign n22725 = ( n22723 & ~n22724 ) | ( n22723 & 1'b0 ) | ( ~n22724 & 1'b0 ) ;
  assign n22734 = ( n4129 & n22555 ) | ( n4129 & n22725 ) | ( n22555 & n22725 ) ;
  assign n22735 = ( n22555 & ~n22575 ) | ( n22555 & n22725 ) | ( ~n22575 & n22725 ) ;
  assign n22736 = ~n22734 & n22735 ;
  assign n22737 = n22730 | n22736 ;
  assign n22738 = n22498 &  n22576 ;
  assign n22731 = x72 | n22498 ;
  assign n22732 = x72 &  n22498 ;
  assign n22733 = ( n22731 & ~n22732 ) | ( n22731 & 1'b0 ) | ( ~n22732 & 1'b0 ) ;
  assign n22742 = ( n4129 & n22554 ) | ( n4129 & n22733 ) | ( n22554 & n22733 ) ;
  assign n22743 = ( n22554 & ~n22575 ) | ( n22554 & n22733 ) | ( ~n22575 & n22733 ) ;
  assign n22744 = ~n22742 & n22743 ;
  assign n22745 = n22738 | n22744 ;
  assign n22746 = n22506 &  n22576 ;
  assign n22739 = x71 | n22506 ;
  assign n22740 = x71 &  n22506 ;
  assign n22741 = ( n22739 & ~n22740 ) | ( n22739 & 1'b0 ) | ( ~n22740 & 1'b0 ) ;
  assign n22750 = ( n4129 & n22553 ) | ( n4129 & n22741 ) | ( n22553 & n22741 ) ;
  assign n22751 = ( n22553 & ~n22575 ) | ( n22553 & n22741 ) | ( ~n22575 & n22741 ) ;
  assign n22752 = ~n22750 & n22751 ;
  assign n22753 = n22746 | n22752 ;
  assign n22754 = n22514 &  n22576 ;
  assign n22747 = x70 | n22514 ;
  assign n22748 = x70 &  n22514 ;
  assign n22749 = ( n22747 & ~n22748 ) | ( n22747 & 1'b0 ) | ( ~n22748 & 1'b0 ) ;
  assign n22758 = ( n4129 & n22552 ) | ( n4129 & n22749 ) | ( n22552 & n22749 ) ;
  assign n22759 = ( n22552 & ~n22575 ) | ( n22552 & n22749 ) | ( ~n22575 & n22749 ) ;
  assign n22760 = ~n22758 & n22759 ;
  assign n22761 = n22754 | n22760 ;
  assign n22762 = n22522 &  n22576 ;
  assign n22755 = x69 | n22522 ;
  assign n22756 = x69 &  n22522 ;
  assign n22757 = ( n22755 & ~n22756 ) | ( n22755 & 1'b0 ) | ( ~n22756 & 1'b0 ) ;
  assign n22766 = ( n4129 & n22551 ) | ( n4129 & n22757 ) | ( n22551 & n22757 ) ;
  assign n22767 = ( n22551 & ~n22575 ) | ( n22551 & n22757 ) | ( ~n22575 & n22757 ) ;
  assign n22768 = ~n22766 & n22767 ;
  assign n22769 = n22762 | n22768 ;
  assign n22770 = n22530 &  n22576 ;
  assign n22763 = x68 | n22530 ;
  assign n22764 = x68 &  n22530 ;
  assign n22765 = ( n22763 & ~n22764 ) | ( n22763 & 1'b0 ) | ( ~n22764 & 1'b0 ) ;
  assign n22774 = ( n4129 & n22550 ) | ( n4129 & n22765 ) | ( n22550 & n22765 ) ;
  assign n22775 = ( n22550 & ~n22575 ) | ( n22550 & n22765 ) | ( ~n22575 & n22765 ) ;
  assign n22776 = ~n22774 & n22775 ;
  assign n22777 = n22770 | n22776 ;
  assign n22778 = n22535 &  n22576 ;
  assign n22771 = x67 | n22535 ;
  assign n22772 = x67 &  n22535 ;
  assign n22773 = ( n22771 & ~n22772 ) | ( n22771 & 1'b0 ) | ( ~n22772 & 1'b0 ) ;
  assign n22782 = ( n4129 & n22549 ) | ( n4129 & n22773 ) | ( n22549 & n22773 ) ;
  assign n22783 = ( n22549 & ~n22575 ) | ( n22549 & n22773 ) | ( ~n22575 & n22773 ) ;
  assign n22784 = ~n22782 & n22783 ;
  assign n22785 = n22778 | n22784 ;
  assign n22786 = n22543 &  n22576 ;
  assign n22779 = x66 | n22543 ;
  assign n22780 = x66 &  n22543 ;
  assign n22781 = ( n22779 & ~n22780 ) | ( n22779 & 1'b0 ) | ( ~n22780 & 1'b0 ) ;
  assign n22790 = ( n4129 & n22548 ) | ( n4129 & n22781 ) | ( n22548 & n22781 ) ;
  assign n22791 = ( n22548 & ~n22575 ) | ( n22548 & n22781 ) | ( ~n22575 & n22781 ) ;
  assign n22792 = ~n22790 & n22791 ;
  assign n22793 = n22786 | n22792 ;
  assign n22794 = n22547 &  n22576 ;
  assign n22787 = x65 &  n22547 ;
  assign n22788 = x65 | n22546 ;
  assign n22789 = n22545 | n22788 ;
  assign n22795 = ~n22787 & n22789 ;
  assign n22796 = ( n4099 & ~n4129 ) | ( n4099 & n22795 ) | ( ~n4129 & n22795 ) ;
  assign n22797 = ( n4099 & n22575 ) | ( n4099 & n22795 ) | ( n22575 & n22795 ) ;
  assign n22798 = ( n22796 & ~n22797 ) | ( n22796 & 1'b0 ) | ( ~n22797 & 1'b0 ) ;
  assign n22799 = n22794 | n22798 ;
  assign n22800 = ( n4201 & ~n22575 ) | ( n4201 & 1'b0 ) | ( ~n22575 & 1'b0 ) ;
  assign n22801 = ( x35 & ~n22800 ) | ( x35 & 1'b0 ) | ( ~n22800 & 1'b0 ) ;
  assign n22802 = ( n4206 & ~n22575 ) | ( n4206 & 1'b0 ) | ( ~n22575 & 1'b0 ) ;
  assign n22803 = n22801 | n22802 ;
  assign n22804 = ( x65 & ~n22803 ) | ( x65 & n4209 ) | ( ~n22803 & n4209 ) ;
  assign n22805 = ( x66 & ~n22799 ) | ( x66 & n22804 ) | ( ~n22799 & n22804 ) ;
  assign n22806 = ( x67 & ~n22793 ) | ( x67 & n22805 ) | ( ~n22793 & n22805 ) ;
  assign n22807 = ( x68 & ~n22785 ) | ( x68 & n22806 ) | ( ~n22785 & n22806 ) ;
  assign n22808 = ( x69 & ~n22777 ) | ( x69 & n22807 ) | ( ~n22777 & n22807 ) ;
  assign n22809 = ( x70 & ~n22769 ) | ( x70 & n22808 ) | ( ~n22769 & n22808 ) ;
  assign n22810 = ( x71 & ~n22761 ) | ( x71 & n22809 ) | ( ~n22761 & n22809 ) ;
  assign n22811 = ( x72 & ~n22753 ) | ( x72 & n22810 ) | ( ~n22753 & n22810 ) ;
  assign n22812 = ( x73 & ~n22745 ) | ( x73 & n22811 ) | ( ~n22745 & n22811 ) ;
  assign n22813 = ( x74 & ~n22737 ) | ( x74 & n22812 ) | ( ~n22737 & n22812 ) ;
  assign n22814 = ( x75 & ~n22729 ) | ( x75 & n22813 ) | ( ~n22729 & n22813 ) ;
  assign n22815 = ( x76 & ~n22721 ) | ( x76 & n22814 ) | ( ~n22721 & n22814 ) ;
  assign n22816 = ( x77 & ~n22713 ) | ( x77 & n22815 ) | ( ~n22713 & n22815 ) ;
  assign n22817 = ( x78 & ~n22705 ) | ( x78 & n22816 ) | ( ~n22705 & n22816 ) ;
  assign n22818 = ( x79 & ~n22697 ) | ( x79 & n22817 ) | ( ~n22697 & n22817 ) ;
  assign n22819 = ( x80 & ~n22689 ) | ( x80 & n22818 ) | ( ~n22689 & n22818 ) ;
  assign n22820 = ( x81 & ~n22681 ) | ( x81 & n22819 ) | ( ~n22681 & n22819 ) ;
  assign n22821 = ( x82 & ~n22673 ) | ( x82 & n22820 ) | ( ~n22673 & n22820 ) ;
  assign n22822 = ( x83 & ~n22665 ) | ( x83 & n22821 ) | ( ~n22665 & n22821 ) ;
  assign n22823 = ( x84 & ~n22657 ) | ( x84 & n22822 ) | ( ~n22657 & n22822 ) ;
  assign n22824 = ( x85 & ~n22649 ) | ( x85 & n22823 ) | ( ~n22649 & n22823 ) ;
  assign n22825 = ( x86 & ~n22641 ) | ( x86 & n22824 ) | ( ~n22641 & n22824 ) ;
  assign n22826 = ( x87 & ~n22633 ) | ( x87 & n22825 ) | ( ~n22633 & n22825 ) ;
  assign n22827 = ( x88 & ~n22625 ) | ( x88 & n22826 ) | ( ~n22625 & n22826 ) ;
  assign n22828 = ( x89 & ~n22617 ) | ( x89 & n22827 ) | ( ~n22617 & n22827 ) ;
  assign n22829 = ( x90 & ~n22609 ) | ( x90 & n22828 ) | ( ~n22609 & n22828 ) ;
  assign n22830 = ( x91 & ~n22601 ) | ( x91 & n22829 ) | ( ~n22601 & n22829 ) ;
  assign n22831 = ( x92 & ~n22593 ) | ( x92 & n22830 ) | ( ~n22593 & n22830 ) ;
  assign n22832 = ( x93 & ~n22577 ) | ( x93 & 1'b0 ) | ( ~n22577 & 1'b0 ) ;
  assign n22833 = ~n22583 & n22832 ;
  assign n22834 = ( n22831 & ~n22585 ) | ( n22831 & n22833 ) | ( ~n22585 & n22833 ) ;
  assign n22835 = ( n22585 & ~n4401 ) | ( n22585 & n22834 ) | ( ~n4401 & n22834 ) ;
  assign n22836 = n4401 | n22835 ;
  assign n22843 = n4129 &  n22338 ;
  assign n22844 = n22836 &  n22843 ;
  assign n22837 = ~n22584 |  n4129 ;
  assign n22838 = n22836 &  n22837 ;
  assign n22842 = n22585 | n22833 ;
  assign n22846 = ( n22831 & n22838 ) | ( n22831 & n22842 ) | ( n22838 & n22842 ) ;
  assign n22845 = n22831 | n22842 ;
  assign n22847 = ( n22844 & ~n22846 ) | ( n22844 & n22845 ) | ( ~n22846 & n22845 ) ;
  assign n22851 = n22593 &  n22837 ;
  assign n22852 = n22836 &  n22851 ;
  assign n22839 = x92 | n22593 ;
  assign n22840 = x92 &  n22593 ;
  assign n22841 = ( n22839 & ~n22840 ) | ( n22839 & 1'b0 ) | ( ~n22840 & 1'b0 ) ;
  assign n22854 = ( n22830 & n22838 ) | ( n22830 & n22841 ) | ( n22838 & n22841 ) ;
  assign n22853 = n22830 | n22841 ;
  assign n22855 = ( n22852 & ~n22854 ) | ( n22852 & n22853 ) | ( ~n22854 & n22853 ) ;
  assign n22859 = n22601 &  n22837 ;
  assign n22860 = n22836 &  n22859 ;
  assign n22848 = x91 | n22601 ;
  assign n22849 = x91 &  n22601 ;
  assign n22850 = ( n22848 & ~n22849 ) | ( n22848 & 1'b0 ) | ( ~n22849 & 1'b0 ) ;
  assign n22862 = ( n22829 & n22838 ) | ( n22829 & n22850 ) | ( n22838 & n22850 ) ;
  assign n22861 = n22829 | n22850 ;
  assign n22863 = ( n22860 & ~n22862 ) | ( n22860 & n22861 ) | ( ~n22862 & n22861 ) ;
  assign n22867 = n22609 &  n22837 ;
  assign n22868 = n22836 &  n22867 ;
  assign n22856 = x90 | n22609 ;
  assign n22857 = x90 &  n22609 ;
  assign n22858 = ( n22856 & ~n22857 ) | ( n22856 & 1'b0 ) | ( ~n22857 & 1'b0 ) ;
  assign n22870 = ( n22828 & n22838 ) | ( n22828 & n22858 ) | ( n22838 & n22858 ) ;
  assign n22869 = n22828 | n22858 ;
  assign n22871 = ( n22868 & ~n22870 ) | ( n22868 & n22869 ) | ( ~n22870 & n22869 ) ;
  assign n22875 = n22617 &  n22837 ;
  assign n22876 = n22836 &  n22875 ;
  assign n22864 = x89 | n22617 ;
  assign n22865 = x89 &  n22617 ;
  assign n22866 = ( n22864 & ~n22865 ) | ( n22864 & 1'b0 ) | ( ~n22865 & 1'b0 ) ;
  assign n22878 = ( n22827 & n22838 ) | ( n22827 & n22866 ) | ( n22838 & n22866 ) ;
  assign n22877 = n22827 | n22866 ;
  assign n22879 = ( n22876 & ~n22878 ) | ( n22876 & n22877 ) | ( ~n22878 & n22877 ) ;
  assign n22883 = n22625 &  n22837 ;
  assign n22884 = n22836 &  n22883 ;
  assign n22872 = x88 | n22625 ;
  assign n22873 = x88 &  n22625 ;
  assign n22874 = ( n22872 & ~n22873 ) | ( n22872 & 1'b0 ) | ( ~n22873 & 1'b0 ) ;
  assign n22886 = ( n22826 & n22838 ) | ( n22826 & n22874 ) | ( n22838 & n22874 ) ;
  assign n22885 = n22826 | n22874 ;
  assign n22887 = ( n22884 & ~n22886 ) | ( n22884 & n22885 ) | ( ~n22886 & n22885 ) ;
  assign n22891 = n22633 &  n22837 ;
  assign n22892 = n22836 &  n22891 ;
  assign n22880 = x87 | n22633 ;
  assign n22881 = x87 &  n22633 ;
  assign n22882 = ( n22880 & ~n22881 ) | ( n22880 & 1'b0 ) | ( ~n22881 & 1'b0 ) ;
  assign n22894 = ( n22825 & n22838 ) | ( n22825 & n22882 ) | ( n22838 & n22882 ) ;
  assign n22893 = n22825 | n22882 ;
  assign n22895 = ( n22892 & ~n22894 ) | ( n22892 & n22893 ) | ( ~n22894 & n22893 ) ;
  assign n22899 = n22641 &  n22837 ;
  assign n22900 = n22836 &  n22899 ;
  assign n22888 = x86 | n22641 ;
  assign n22889 = x86 &  n22641 ;
  assign n22890 = ( n22888 & ~n22889 ) | ( n22888 & 1'b0 ) | ( ~n22889 & 1'b0 ) ;
  assign n22902 = ( n22824 & n22838 ) | ( n22824 & n22890 ) | ( n22838 & n22890 ) ;
  assign n22901 = n22824 | n22890 ;
  assign n22903 = ( n22900 & ~n22902 ) | ( n22900 & n22901 ) | ( ~n22902 & n22901 ) ;
  assign n22907 = n22649 &  n22837 ;
  assign n22908 = n22836 &  n22907 ;
  assign n22896 = x85 | n22649 ;
  assign n22897 = x85 &  n22649 ;
  assign n22898 = ( n22896 & ~n22897 ) | ( n22896 & 1'b0 ) | ( ~n22897 & 1'b0 ) ;
  assign n22910 = ( n22823 & n22838 ) | ( n22823 & n22898 ) | ( n22838 & n22898 ) ;
  assign n22909 = n22823 | n22898 ;
  assign n22911 = ( n22908 & ~n22910 ) | ( n22908 & n22909 ) | ( ~n22910 & n22909 ) ;
  assign n22915 = n22657 &  n22837 ;
  assign n22916 = n22836 &  n22915 ;
  assign n22904 = x84 | n22657 ;
  assign n22905 = x84 &  n22657 ;
  assign n22906 = ( n22904 & ~n22905 ) | ( n22904 & 1'b0 ) | ( ~n22905 & 1'b0 ) ;
  assign n22918 = ( n22822 & n22838 ) | ( n22822 & n22906 ) | ( n22838 & n22906 ) ;
  assign n22917 = n22822 | n22906 ;
  assign n22919 = ( n22916 & ~n22918 ) | ( n22916 & n22917 ) | ( ~n22918 & n22917 ) ;
  assign n22923 = n22665 &  n22837 ;
  assign n22924 = n22836 &  n22923 ;
  assign n22912 = x83 | n22665 ;
  assign n22913 = x83 &  n22665 ;
  assign n22914 = ( n22912 & ~n22913 ) | ( n22912 & 1'b0 ) | ( ~n22913 & 1'b0 ) ;
  assign n22926 = ( n22821 & n22838 ) | ( n22821 & n22914 ) | ( n22838 & n22914 ) ;
  assign n22925 = n22821 | n22914 ;
  assign n22927 = ( n22924 & ~n22926 ) | ( n22924 & n22925 ) | ( ~n22926 & n22925 ) ;
  assign n22931 = n22673 &  n22837 ;
  assign n22932 = n22836 &  n22931 ;
  assign n22920 = x82 | n22673 ;
  assign n22921 = x82 &  n22673 ;
  assign n22922 = ( n22920 & ~n22921 ) | ( n22920 & 1'b0 ) | ( ~n22921 & 1'b0 ) ;
  assign n22934 = ( n22820 & n22838 ) | ( n22820 & n22922 ) | ( n22838 & n22922 ) ;
  assign n22933 = n22820 | n22922 ;
  assign n22935 = ( n22932 & ~n22934 ) | ( n22932 & n22933 ) | ( ~n22934 & n22933 ) ;
  assign n22939 = n22681 &  n22837 ;
  assign n22940 = n22836 &  n22939 ;
  assign n22928 = x81 | n22681 ;
  assign n22929 = x81 &  n22681 ;
  assign n22930 = ( n22928 & ~n22929 ) | ( n22928 & 1'b0 ) | ( ~n22929 & 1'b0 ) ;
  assign n22942 = ( n22819 & n22838 ) | ( n22819 & n22930 ) | ( n22838 & n22930 ) ;
  assign n22941 = n22819 | n22930 ;
  assign n22943 = ( n22940 & ~n22942 ) | ( n22940 & n22941 ) | ( ~n22942 & n22941 ) ;
  assign n22947 = n22689 &  n22837 ;
  assign n22948 = n22836 &  n22947 ;
  assign n22936 = x80 | n22689 ;
  assign n22937 = x80 &  n22689 ;
  assign n22938 = ( n22936 & ~n22937 ) | ( n22936 & 1'b0 ) | ( ~n22937 & 1'b0 ) ;
  assign n22950 = ( n22818 & n22838 ) | ( n22818 & n22938 ) | ( n22838 & n22938 ) ;
  assign n22949 = n22818 | n22938 ;
  assign n22951 = ( n22948 & ~n22950 ) | ( n22948 & n22949 ) | ( ~n22950 & n22949 ) ;
  assign n22955 = n22697 &  n22837 ;
  assign n22956 = n22836 &  n22955 ;
  assign n22944 = x79 | n22697 ;
  assign n22945 = x79 &  n22697 ;
  assign n22946 = ( n22944 & ~n22945 ) | ( n22944 & 1'b0 ) | ( ~n22945 & 1'b0 ) ;
  assign n22958 = ( n22817 & n22838 ) | ( n22817 & n22946 ) | ( n22838 & n22946 ) ;
  assign n22957 = n22817 | n22946 ;
  assign n22959 = ( n22956 & ~n22958 ) | ( n22956 & n22957 ) | ( ~n22958 & n22957 ) ;
  assign n22963 = n22705 &  n22837 ;
  assign n22964 = n22836 &  n22963 ;
  assign n22952 = x78 | n22705 ;
  assign n22953 = x78 &  n22705 ;
  assign n22954 = ( n22952 & ~n22953 ) | ( n22952 & 1'b0 ) | ( ~n22953 & 1'b0 ) ;
  assign n22966 = ( n22816 & n22838 ) | ( n22816 & n22954 ) | ( n22838 & n22954 ) ;
  assign n22965 = n22816 | n22954 ;
  assign n22967 = ( n22964 & ~n22966 ) | ( n22964 & n22965 ) | ( ~n22966 & n22965 ) ;
  assign n22971 = n22713 &  n22837 ;
  assign n22972 = n22836 &  n22971 ;
  assign n22960 = x77 | n22713 ;
  assign n22961 = x77 &  n22713 ;
  assign n22962 = ( n22960 & ~n22961 ) | ( n22960 & 1'b0 ) | ( ~n22961 & 1'b0 ) ;
  assign n22974 = ( n22815 & n22838 ) | ( n22815 & n22962 ) | ( n22838 & n22962 ) ;
  assign n22973 = n22815 | n22962 ;
  assign n22975 = ( n22972 & ~n22974 ) | ( n22972 & n22973 ) | ( ~n22974 & n22973 ) ;
  assign n22979 = n22721 &  n22837 ;
  assign n22980 = n22836 &  n22979 ;
  assign n22968 = x76 | n22721 ;
  assign n22969 = x76 &  n22721 ;
  assign n22970 = ( n22968 & ~n22969 ) | ( n22968 & 1'b0 ) | ( ~n22969 & 1'b0 ) ;
  assign n22982 = ( n22814 & n22838 ) | ( n22814 & n22970 ) | ( n22838 & n22970 ) ;
  assign n22981 = n22814 | n22970 ;
  assign n22983 = ( n22980 & ~n22982 ) | ( n22980 & n22981 ) | ( ~n22982 & n22981 ) ;
  assign n22987 = n22729 &  n22837 ;
  assign n22988 = n22836 &  n22987 ;
  assign n22976 = x75 | n22729 ;
  assign n22977 = x75 &  n22729 ;
  assign n22978 = ( n22976 & ~n22977 ) | ( n22976 & 1'b0 ) | ( ~n22977 & 1'b0 ) ;
  assign n22990 = ( n22813 & n22838 ) | ( n22813 & n22978 ) | ( n22838 & n22978 ) ;
  assign n22989 = n22813 | n22978 ;
  assign n22991 = ( n22988 & ~n22990 ) | ( n22988 & n22989 ) | ( ~n22990 & n22989 ) ;
  assign n22995 = n22737 &  n22837 ;
  assign n22996 = n22836 &  n22995 ;
  assign n22984 = x74 | n22737 ;
  assign n22985 = x74 &  n22737 ;
  assign n22986 = ( n22984 & ~n22985 ) | ( n22984 & 1'b0 ) | ( ~n22985 & 1'b0 ) ;
  assign n22998 = ( n22812 & n22838 ) | ( n22812 & n22986 ) | ( n22838 & n22986 ) ;
  assign n22997 = n22812 | n22986 ;
  assign n22999 = ( n22996 & ~n22998 ) | ( n22996 & n22997 ) | ( ~n22998 & n22997 ) ;
  assign n23003 = n22745 &  n22837 ;
  assign n23004 = n22836 &  n23003 ;
  assign n22992 = x73 | n22745 ;
  assign n22993 = x73 &  n22745 ;
  assign n22994 = ( n22992 & ~n22993 ) | ( n22992 & 1'b0 ) | ( ~n22993 & 1'b0 ) ;
  assign n23006 = ( n22811 & n22838 ) | ( n22811 & n22994 ) | ( n22838 & n22994 ) ;
  assign n23005 = n22811 | n22994 ;
  assign n23007 = ( n23004 & ~n23006 ) | ( n23004 & n23005 ) | ( ~n23006 & n23005 ) ;
  assign n23011 = n22753 &  n22837 ;
  assign n23012 = n22836 &  n23011 ;
  assign n23000 = x72 | n22753 ;
  assign n23001 = x72 &  n22753 ;
  assign n23002 = ( n23000 & ~n23001 ) | ( n23000 & 1'b0 ) | ( ~n23001 & 1'b0 ) ;
  assign n23014 = ( n22810 & n22838 ) | ( n22810 & n23002 ) | ( n22838 & n23002 ) ;
  assign n23013 = n22810 | n23002 ;
  assign n23015 = ( n23012 & ~n23014 ) | ( n23012 & n23013 ) | ( ~n23014 & n23013 ) ;
  assign n23019 = n22761 &  n22837 ;
  assign n23020 = n22836 &  n23019 ;
  assign n23008 = x71 | n22761 ;
  assign n23009 = x71 &  n22761 ;
  assign n23010 = ( n23008 & ~n23009 ) | ( n23008 & 1'b0 ) | ( ~n23009 & 1'b0 ) ;
  assign n23022 = ( n22809 & n22838 ) | ( n22809 & n23010 ) | ( n22838 & n23010 ) ;
  assign n23021 = n22809 | n23010 ;
  assign n23023 = ( n23020 & ~n23022 ) | ( n23020 & n23021 ) | ( ~n23022 & n23021 ) ;
  assign n23027 = n22769 &  n22837 ;
  assign n23028 = n22836 &  n23027 ;
  assign n23016 = x70 | n22769 ;
  assign n23017 = x70 &  n22769 ;
  assign n23018 = ( n23016 & ~n23017 ) | ( n23016 & 1'b0 ) | ( ~n23017 & 1'b0 ) ;
  assign n23030 = ( n22808 & n22838 ) | ( n22808 & n23018 ) | ( n22838 & n23018 ) ;
  assign n23029 = n22808 | n23018 ;
  assign n23031 = ( n23028 & ~n23030 ) | ( n23028 & n23029 ) | ( ~n23030 & n23029 ) ;
  assign n23035 = n22777 &  n22837 ;
  assign n23036 = n22836 &  n23035 ;
  assign n23024 = x69 | n22777 ;
  assign n23025 = x69 &  n22777 ;
  assign n23026 = ( n23024 & ~n23025 ) | ( n23024 & 1'b0 ) | ( ~n23025 & 1'b0 ) ;
  assign n23038 = ( n22807 & n22838 ) | ( n22807 & n23026 ) | ( n22838 & n23026 ) ;
  assign n23037 = n22807 | n23026 ;
  assign n23039 = ( n23036 & ~n23038 ) | ( n23036 & n23037 ) | ( ~n23038 & n23037 ) ;
  assign n23043 = n22785 &  n22837 ;
  assign n23044 = n22836 &  n23043 ;
  assign n23032 = x68 | n22785 ;
  assign n23033 = x68 &  n22785 ;
  assign n23034 = ( n23032 & ~n23033 ) | ( n23032 & 1'b0 ) | ( ~n23033 & 1'b0 ) ;
  assign n23046 = ( n22806 & n22838 ) | ( n22806 & n23034 ) | ( n22838 & n23034 ) ;
  assign n23045 = n22806 | n23034 ;
  assign n23047 = ( n23044 & ~n23046 ) | ( n23044 & n23045 ) | ( ~n23046 & n23045 ) ;
  assign n23051 = n22793 &  n22837 ;
  assign n23052 = n22836 &  n23051 ;
  assign n23040 = x67 | n22793 ;
  assign n23041 = x67 &  n22793 ;
  assign n23042 = ( n23040 & ~n23041 ) | ( n23040 & 1'b0 ) | ( ~n23041 & 1'b0 ) ;
  assign n23054 = ( n22805 & n22838 ) | ( n22805 & n23042 ) | ( n22838 & n23042 ) ;
  assign n23053 = n22805 | n23042 ;
  assign n23055 = ( n23052 & ~n23054 ) | ( n23052 & n23053 ) | ( ~n23054 & n23053 ) ;
  assign n23056 = n22799 &  n22837 ;
  assign n23057 = n22836 &  n23056 ;
  assign n23048 = x66 | n22799 ;
  assign n23049 = x66 &  n22799 ;
  assign n23050 = ( n23048 & ~n23049 ) | ( n23048 & 1'b0 ) | ( ~n23049 & 1'b0 ) ;
  assign n23059 = ( n22804 & n22838 ) | ( n22804 & n23050 ) | ( n22838 & n23050 ) ;
  assign n23058 = n22804 | n23050 ;
  assign n23060 = ( n23057 & ~n23059 ) | ( n23057 & n23058 ) | ( ~n23059 & n23058 ) ;
  assign n23061 = ( x65 & ~n4209 ) | ( x65 & n22803 ) | ( ~n4209 & n22803 ) ;
  assign n23062 = ( n22804 & ~x65 ) | ( n22804 & n23061 ) | ( ~x65 & n23061 ) ;
  assign n23063 = ~n22838 & n23062 ;
  assign n23064 = n22803 &  n22837 ;
  assign n23065 = n22836 &  n23064 ;
  assign n23066 = n23063 | n23065 ;
  assign n23067 = ( x64 & ~n22838 ) | ( x64 & 1'b0 ) | ( ~n22838 & 1'b0 ) ;
  assign n23068 = ( x34 & ~n23067 ) | ( x34 & 1'b0 ) | ( ~n23067 & 1'b0 ) ;
  assign n23069 = ( n4209 & ~n22838 ) | ( n4209 & 1'b0 ) | ( ~n22838 & 1'b0 ) ;
  assign n23070 = n23068 | n23069 ;
  assign n23071 = ( x65 & ~n23070 ) | ( x65 & n4635 ) | ( ~n23070 & n4635 ) ;
  assign n23072 = ( x66 & ~n23066 ) | ( x66 & n23071 ) | ( ~n23066 & n23071 ) ;
  assign n23073 = ( x67 & ~n23060 ) | ( x67 & n23072 ) | ( ~n23060 & n23072 ) ;
  assign n23074 = ( x68 & ~n23055 ) | ( x68 & n23073 ) | ( ~n23055 & n23073 ) ;
  assign n23075 = ( x69 & ~n23047 ) | ( x69 & n23074 ) | ( ~n23047 & n23074 ) ;
  assign n23076 = ( x70 & ~n23039 ) | ( x70 & n23075 ) | ( ~n23039 & n23075 ) ;
  assign n23077 = ( x71 & ~n23031 ) | ( x71 & n23076 ) | ( ~n23031 & n23076 ) ;
  assign n23078 = ( x72 & ~n23023 ) | ( x72 & n23077 ) | ( ~n23023 & n23077 ) ;
  assign n23079 = ( x73 & ~n23015 ) | ( x73 & n23078 ) | ( ~n23015 & n23078 ) ;
  assign n23080 = ( x74 & ~n23007 ) | ( x74 & n23079 ) | ( ~n23007 & n23079 ) ;
  assign n23081 = ( x75 & ~n22999 ) | ( x75 & n23080 ) | ( ~n22999 & n23080 ) ;
  assign n23082 = ( x76 & ~n22991 ) | ( x76 & n23081 ) | ( ~n22991 & n23081 ) ;
  assign n23083 = ( x77 & ~n22983 ) | ( x77 & n23082 ) | ( ~n22983 & n23082 ) ;
  assign n23084 = ( x78 & ~n22975 ) | ( x78 & n23083 ) | ( ~n22975 & n23083 ) ;
  assign n23085 = ( x79 & ~n22967 ) | ( x79 & n23084 ) | ( ~n22967 & n23084 ) ;
  assign n23086 = ( x80 & ~n22959 ) | ( x80 & n23085 ) | ( ~n22959 & n23085 ) ;
  assign n23087 = ( x81 & ~n22951 ) | ( x81 & n23086 ) | ( ~n22951 & n23086 ) ;
  assign n23088 = ( x82 & ~n22943 ) | ( x82 & n23087 ) | ( ~n22943 & n23087 ) ;
  assign n23089 = ( x83 & ~n22935 ) | ( x83 & n23088 ) | ( ~n22935 & n23088 ) ;
  assign n23090 = ( x84 & ~n22927 ) | ( x84 & n23089 ) | ( ~n22927 & n23089 ) ;
  assign n23091 = ( x85 & ~n22919 ) | ( x85 & n23090 ) | ( ~n22919 & n23090 ) ;
  assign n23092 = ( x86 & ~n22911 ) | ( x86 & n23091 ) | ( ~n22911 & n23091 ) ;
  assign n23093 = ( x87 & ~n22903 ) | ( x87 & n23092 ) | ( ~n22903 & n23092 ) ;
  assign n23094 = ( x88 & ~n22895 ) | ( x88 & n23093 ) | ( ~n22895 & n23093 ) ;
  assign n23095 = ( x89 & ~n22887 ) | ( x89 & n23094 ) | ( ~n22887 & n23094 ) ;
  assign n23096 = ( x90 & ~n22879 ) | ( x90 & n23095 ) | ( ~n22879 & n23095 ) ;
  assign n23097 = ( x91 & ~n22871 ) | ( x91 & n23096 ) | ( ~n22871 & n23096 ) ;
  assign n23098 = ( x92 & ~n22863 ) | ( x92 & n23097 ) | ( ~n22863 & n23097 ) ;
  assign n23099 = ( x93 & ~n22855 ) | ( x93 & n23098 ) | ( ~n22855 & n23098 ) ;
  assign n23106 = ( x94 & ~n4668 ) | ( x94 & n23099 ) | ( ~n4668 & n23099 ) ;
  assign n23105 = x94 &  n23099 ;
  assign n23107 = ( n22847 & ~n23106 ) | ( n22847 & n23105 ) | ( ~n23106 & n23105 ) ;
  assign n23100 = ( x94 & ~n22847 ) | ( x94 & n23099 ) | ( ~n22847 & n23099 ) ;
  assign n23101 = n4668 | n23100 ;
  assign n23108 = n22855 &  n23101 ;
  assign n23102 = x93 | n22855 ;
  assign n23103 = x93 &  n22855 ;
  assign n23104 = ( n23102 & ~n23103 ) | ( n23102 & 1'b0 ) | ( ~n23103 & 1'b0 ) ;
  assign n23112 = ( n4668 & n23098 ) | ( n4668 & n23104 ) | ( n23098 & n23104 ) ;
  assign n23113 = ( n23098 & ~n23100 ) | ( n23098 & n23104 ) | ( ~n23100 & n23104 ) ;
  assign n23114 = ~n23112 & n23113 ;
  assign n23115 = n23108 | n23114 ;
  assign n23116 = n22863 &  n23101 ;
  assign n23109 = x92 | n22863 ;
  assign n23110 = x92 &  n22863 ;
  assign n23111 = ( n23109 & ~n23110 ) | ( n23109 & 1'b0 ) | ( ~n23110 & 1'b0 ) ;
  assign n23120 = ( n4668 & n23097 ) | ( n4668 & n23111 ) | ( n23097 & n23111 ) ;
  assign n23121 = ( n23097 & ~n23100 ) | ( n23097 & n23111 ) | ( ~n23100 & n23111 ) ;
  assign n23122 = ~n23120 & n23121 ;
  assign n23123 = n23116 | n23122 ;
  assign n23124 = n22871 &  n23101 ;
  assign n23117 = x91 | n22871 ;
  assign n23118 = x91 &  n22871 ;
  assign n23119 = ( n23117 & ~n23118 ) | ( n23117 & 1'b0 ) | ( ~n23118 & 1'b0 ) ;
  assign n23128 = ( n4668 & n23096 ) | ( n4668 & n23119 ) | ( n23096 & n23119 ) ;
  assign n23129 = ( n23096 & ~n23100 ) | ( n23096 & n23119 ) | ( ~n23100 & n23119 ) ;
  assign n23130 = ~n23128 & n23129 ;
  assign n23131 = n23124 | n23130 ;
  assign n23132 = n22879 &  n23101 ;
  assign n23125 = x90 | n22879 ;
  assign n23126 = x90 &  n22879 ;
  assign n23127 = ( n23125 & ~n23126 ) | ( n23125 & 1'b0 ) | ( ~n23126 & 1'b0 ) ;
  assign n23136 = ( n4668 & n23095 ) | ( n4668 & n23127 ) | ( n23095 & n23127 ) ;
  assign n23137 = ( n23095 & ~n23100 ) | ( n23095 & n23127 ) | ( ~n23100 & n23127 ) ;
  assign n23138 = ~n23136 & n23137 ;
  assign n23139 = n23132 | n23138 ;
  assign n23140 = n22887 &  n23101 ;
  assign n23133 = x89 | n22887 ;
  assign n23134 = x89 &  n22887 ;
  assign n23135 = ( n23133 & ~n23134 ) | ( n23133 & 1'b0 ) | ( ~n23134 & 1'b0 ) ;
  assign n23144 = ( n4668 & n23094 ) | ( n4668 & n23135 ) | ( n23094 & n23135 ) ;
  assign n23145 = ( n23094 & ~n23100 ) | ( n23094 & n23135 ) | ( ~n23100 & n23135 ) ;
  assign n23146 = ~n23144 & n23145 ;
  assign n23147 = n23140 | n23146 ;
  assign n23148 = n22895 &  n23101 ;
  assign n23141 = x88 | n22895 ;
  assign n23142 = x88 &  n22895 ;
  assign n23143 = ( n23141 & ~n23142 ) | ( n23141 & 1'b0 ) | ( ~n23142 & 1'b0 ) ;
  assign n23152 = ( n4668 & n23093 ) | ( n4668 & n23143 ) | ( n23093 & n23143 ) ;
  assign n23153 = ( n23093 & ~n23100 ) | ( n23093 & n23143 ) | ( ~n23100 & n23143 ) ;
  assign n23154 = ~n23152 & n23153 ;
  assign n23155 = n23148 | n23154 ;
  assign n23156 = n22903 &  n23101 ;
  assign n23149 = x87 | n22903 ;
  assign n23150 = x87 &  n22903 ;
  assign n23151 = ( n23149 & ~n23150 ) | ( n23149 & 1'b0 ) | ( ~n23150 & 1'b0 ) ;
  assign n23160 = ( n4668 & n23092 ) | ( n4668 & n23151 ) | ( n23092 & n23151 ) ;
  assign n23161 = ( n23092 & ~n23100 ) | ( n23092 & n23151 ) | ( ~n23100 & n23151 ) ;
  assign n23162 = ~n23160 & n23161 ;
  assign n23163 = n23156 | n23162 ;
  assign n23164 = n22911 &  n23101 ;
  assign n23157 = x86 | n22911 ;
  assign n23158 = x86 &  n22911 ;
  assign n23159 = ( n23157 & ~n23158 ) | ( n23157 & 1'b0 ) | ( ~n23158 & 1'b0 ) ;
  assign n23168 = ( n4668 & n23091 ) | ( n4668 & n23159 ) | ( n23091 & n23159 ) ;
  assign n23169 = ( n23091 & ~n23100 ) | ( n23091 & n23159 ) | ( ~n23100 & n23159 ) ;
  assign n23170 = ~n23168 & n23169 ;
  assign n23171 = n23164 | n23170 ;
  assign n23172 = n22919 &  n23101 ;
  assign n23165 = x85 | n22919 ;
  assign n23166 = x85 &  n22919 ;
  assign n23167 = ( n23165 & ~n23166 ) | ( n23165 & 1'b0 ) | ( ~n23166 & 1'b0 ) ;
  assign n23176 = ( n4668 & n23090 ) | ( n4668 & n23167 ) | ( n23090 & n23167 ) ;
  assign n23177 = ( n23090 & ~n23100 ) | ( n23090 & n23167 ) | ( ~n23100 & n23167 ) ;
  assign n23178 = ~n23176 & n23177 ;
  assign n23179 = n23172 | n23178 ;
  assign n23180 = n22927 &  n23101 ;
  assign n23173 = x84 | n22927 ;
  assign n23174 = x84 &  n22927 ;
  assign n23175 = ( n23173 & ~n23174 ) | ( n23173 & 1'b0 ) | ( ~n23174 & 1'b0 ) ;
  assign n23184 = ( n4668 & n23089 ) | ( n4668 & n23175 ) | ( n23089 & n23175 ) ;
  assign n23185 = ( n23089 & ~n23100 ) | ( n23089 & n23175 ) | ( ~n23100 & n23175 ) ;
  assign n23186 = ~n23184 & n23185 ;
  assign n23187 = n23180 | n23186 ;
  assign n23188 = n22935 &  n23101 ;
  assign n23181 = x83 | n22935 ;
  assign n23182 = x83 &  n22935 ;
  assign n23183 = ( n23181 & ~n23182 ) | ( n23181 & 1'b0 ) | ( ~n23182 & 1'b0 ) ;
  assign n23192 = ( n4668 & n23088 ) | ( n4668 & n23183 ) | ( n23088 & n23183 ) ;
  assign n23193 = ( n23088 & ~n23100 ) | ( n23088 & n23183 ) | ( ~n23100 & n23183 ) ;
  assign n23194 = ~n23192 & n23193 ;
  assign n23195 = n23188 | n23194 ;
  assign n23196 = n22943 &  n23101 ;
  assign n23189 = x82 | n22943 ;
  assign n23190 = x82 &  n22943 ;
  assign n23191 = ( n23189 & ~n23190 ) | ( n23189 & 1'b0 ) | ( ~n23190 & 1'b0 ) ;
  assign n23200 = ( n4668 & n23087 ) | ( n4668 & n23191 ) | ( n23087 & n23191 ) ;
  assign n23201 = ( n23087 & ~n23100 ) | ( n23087 & n23191 ) | ( ~n23100 & n23191 ) ;
  assign n23202 = ~n23200 & n23201 ;
  assign n23203 = n23196 | n23202 ;
  assign n23204 = n22951 &  n23101 ;
  assign n23197 = x81 | n22951 ;
  assign n23198 = x81 &  n22951 ;
  assign n23199 = ( n23197 & ~n23198 ) | ( n23197 & 1'b0 ) | ( ~n23198 & 1'b0 ) ;
  assign n23208 = ( n4668 & n23086 ) | ( n4668 & n23199 ) | ( n23086 & n23199 ) ;
  assign n23209 = ( n23086 & ~n23100 ) | ( n23086 & n23199 ) | ( ~n23100 & n23199 ) ;
  assign n23210 = ~n23208 & n23209 ;
  assign n23211 = n23204 | n23210 ;
  assign n23212 = n22959 &  n23101 ;
  assign n23205 = x80 | n22959 ;
  assign n23206 = x80 &  n22959 ;
  assign n23207 = ( n23205 & ~n23206 ) | ( n23205 & 1'b0 ) | ( ~n23206 & 1'b0 ) ;
  assign n23216 = ( n4668 & n23085 ) | ( n4668 & n23207 ) | ( n23085 & n23207 ) ;
  assign n23217 = ( n23085 & ~n23100 ) | ( n23085 & n23207 ) | ( ~n23100 & n23207 ) ;
  assign n23218 = ~n23216 & n23217 ;
  assign n23219 = n23212 | n23218 ;
  assign n23220 = n22967 &  n23101 ;
  assign n23213 = x79 | n22967 ;
  assign n23214 = x79 &  n22967 ;
  assign n23215 = ( n23213 & ~n23214 ) | ( n23213 & 1'b0 ) | ( ~n23214 & 1'b0 ) ;
  assign n23224 = ( n4668 & n23084 ) | ( n4668 & n23215 ) | ( n23084 & n23215 ) ;
  assign n23225 = ( n23084 & ~n23100 ) | ( n23084 & n23215 ) | ( ~n23100 & n23215 ) ;
  assign n23226 = ~n23224 & n23225 ;
  assign n23227 = n23220 | n23226 ;
  assign n23228 = n22975 &  n23101 ;
  assign n23221 = x78 | n22975 ;
  assign n23222 = x78 &  n22975 ;
  assign n23223 = ( n23221 & ~n23222 ) | ( n23221 & 1'b0 ) | ( ~n23222 & 1'b0 ) ;
  assign n23232 = ( n4668 & n23083 ) | ( n4668 & n23223 ) | ( n23083 & n23223 ) ;
  assign n23233 = ( n23083 & ~n23100 ) | ( n23083 & n23223 ) | ( ~n23100 & n23223 ) ;
  assign n23234 = ~n23232 & n23233 ;
  assign n23235 = n23228 | n23234 ;
  assign n23236 = n22983 &  n23101 ;
  assign n23229 = x77 | n22983 ;
  assign n23230 = x77 &  n22983 ;
  assign n23231 = ( n23229 & ~n23230 ) | ( n23229 & 1'b0 ) | ( ~n23230 & 1'b0 ) ;
  assign n23240 = ( n4668 & n23082 ) | ( n4668 & n23231 ) | ( n23082 & n23231 ) ;
  assign n23241 = ( n23082 & ~n23100 ) | ( n23082 & n23231 ) | ( ~n23100 & n23231 ) ;
  assign n23242 = ~n23240 & n23241 ;
  assign n23243 = n23236 | n23242 ;
  assign n23244 = n22991 &  n23101 ;
  assign n23237 = x76 | n22991 ;
  assign n23238 = x76 &  n22991 ;
  assign n23239 = ( n23237 & ~n23238 ) | ( n23237 & 1'b0 ) | ( ~n23238 & 1'b0 ) ;
  assign n23248 = ( n4668 & n23081 ) | ( n4668 & n23239 ) | ( n23081 & n23239 ) ;
  assign n23249 = ( n23081 & ~n23100 ) | ( n23081 & n23239 ) | ( ~n23100 & n23239 ) ;
  assign n23250 = ~n23248 & n23249 ;
  assign n23251 = n23244 | n23250 ;
  assign n23252 = n22999 &  n23101 ;
  assign n23245 = x75 | n22999 ;
  assign n23246 = x75 &  n22999 ;
  assign n23247 = ( n23245 & ~n23246 ) | ( n23245 & 1'b0 ) | ( ~n23246 & 1'b0 ) ;
  assign n23256 = ( n4668 & n23080 ) | ( n4668 & n23247 ) | ( n23080 & n23247 ) ;
  assign n23257 = ( n23080 & ~n23100 ) | ( n23080 & n23247 ) | ( ~n23100 & n23247 ) ;
  assign n23258 = ~n23256 & n23257 ;
  assign n23259 = n23252 | n23258 ;
  assign n23260 = n23007 &  n23101 ;
  assign n23253 = x74 | n23007 ;
  assign n23254 = x74 &  n23007 ;
  assign n23255 = ( n23253 & ~n23254 ) | ( n23253 & 1'b0 ) | ( ~n23254 & 1'b0 ) ;
  assign n23264 = ( n4668 & n23079 ) | ( n4668 & n23255 ) | ( n23079 & n23255 ) ;
  assign n23265 = ( n23079 & ~n23100 ) | ( n23079 & n23255 ) | ( ~n23100 & n23255 ) ;
  assign n23266 = ~n23264 & n23265 ;
  assign n23267 = n23260 | n23266 ;
  assign n23268 = n23015 &  n23101 ;
  assign n23261 = x73 | n23015 ;
  assign n23262 = x73 &  n23015 ;
  assign n23263 = ( n23261 & ~n23262 ) | ( n23261 & 1'b0 ) | ( ~n23262 & 1'b0 ) ;
  assign n23272 = ( n4668 & n23078 ) | ( n4668 & n23263 ) | ( n23078 & n23263 ) ;
  assign n23273 = ( n23078 & ~n23100 ) | ( n23078 & n23263 ) | ( ~n23100 & n23263 ) ;
  assign n23274 = ~n23272 & n23273 ;
  assign n23275 = n23268 | n23274 ;
  assign n23276 = n23023 &  n23101 ;
  assign n23269 = x72 | n23023 ;
  assign n23270 = x72 &  n23023 ;
  assign n23271 = ( n23269 & ~n23270 ) | ( n23269 & 1'b0 ) | ( ~n23270 & 1'b0 ) ;
  assign n23280 = ( n4668 & n23077 ) | ( n4668 & n23271 ) | ( n23077 & n23271 ) ;
  assign n23281 = ( n23077 & ~n23100 ) | ( n23077 & n23271 ) | ( ~n23100 & n23271 ) ;
  assign n23282 = ~n23280 & n23281 ;
  assign n23283 = n23276 | n23282 ;
  assign n23284 = n23031 &  n23101 ;
  assign n23277 = x71 | n23031 ;
  assign n23278 = x71 &  n23031 ;
  assign n23279 = ( n23277 & ~n23278 ) | ( n23277 & 1'b0 ) | ( ~n23278 & 1'b0 ) ;
  assign n23288 = ( n4668 & n23076 ) | ( n4668 & n23279 ) | ( n23076 & n23279 ) ;
  assign n23289 = ( n23076 & ~n23100 ) | ( n23076 & n23279 ) | ( ~n23100 & n23279 ) ;
  assign n23290 = ~n23288 & n23289 ;
  assign n23291 = n23284 | n23290 ;
  assign n23292 = n23039 &  n23101 ;
  assign n23285 = x70 | n23039 ;
  assign n23286 = x70 &  n23039 ;
  assign n23287 = ( n23285 & ~n23286 ) | ( n23285 & 1'b0 ) | ( ~n23286 & 1'b0 ) ;
  assign n23296 = ( n4668 & n23075 ) | ( n4668 & n23287 ) | ( n23075 & n23287 ) ;
  assign n23297 = ( n23075 & ~n23100 ) | ( n23075 & n23287 ) | ( ~n23100 & n23287 ) ;
  assign n23298 = ~n23296 & n23297 ;
  assign n23299 = n23292 | n23298 ;
  assign n23300 = n23047 &  n23101 ;
  assign n23293 = x69 | n23047 ;
  assign n23294 = x69 &  n23047 ;
  assign n23295 = ( n23293 & ~n23294 ) | ( n23293 & 1'b0 ) | ( ~n23294 & 1'b0 ) ;
  assign n23304 = ( n4668 & n23074 ) | ( n4668 & n23295 ) | ( n23074 & n23295 ) ;
  assign n23305 = ( n23074 & ~n23100 ) | ( n23074 & n23295 ) | ( ~n23100 & n23295 ) ;
  assign n23306 = ~n23304 & n23305 ;
  assign n23307 = n23300 | n23306 ;
  assign n23308 = n23055 &  n23101 ;
  assign n23301 = x68 | n23055 ;
  assign n23302 = x68 &  n23055 ;
  assign n23303 = ( n23301 & ~n23302 ) | ( n23301 & 1'b0 ) | ( ~n23302 & 1'b0 ) ;
  assign n23312 = ( n4668 & n23073 ) | ( n4668 & n23303 ) | ( n23073 & n23303 ) ;
  assign n23313 = ( n23073 & ~n23100 ) | ( n23073 & n23303 ) | ( ~n23100 & n23303 ) ;
  assign n23314 = ~n23312 & n23313 ;
  assign n23315 = n23308 | n23314 ;
  assign n23316 = n23060 &  n23101 ;
  assign n23309 = x67 | n23060 ;
  assign n23310 = x67 &  n23060 ;
  assign n23311 = ( n23309 & ~n23310 ) | ( n23309 & 1'b0 ) | ( ~n23310 & 1'b0 ) ;
  assign n23320 = ( n4668 & n23072 ) | ( n4668 & n23311 ) | ( n23072 & n23311 ) ;
  assign n23321 = ( n23072 & ~n23100 ) | ( n23072 & n23311 ) | ( ~n23100 & n23311 ) ;
  assign n23322 = ~n23320 & n23321 ;
  assign n23323 = n23316 | n23322 ;
  assign n23324 = n23066 &  n23101 ;
  assign n23317 = x66 | n23066 ;
  assign n23318 = x66 &  n23066 ;
  assign n23319 = ( n23317 & ~n23318 ) | ( n23317 & 1'b0 ) | ( ~n23318 & 1'b0 ) ;
  assign n23325 = ( n4668 & n23071 ) | ( n4668 & n23319 ) | ( n23071 & n23319 ) ;
  assign n23326 = ( n23071 & ~n23100 ) | ( n23071 & n23319 ) | ( ~n23100 & n23319 ) ;
  assign n23327 = ~n23325 & n23326 ;
  assign n23328 = n23324 | n23327 ;
  assign n23329 = n23070 &  n23101 ;
  assign n23330 = ( x65 & ~x34 ) | ( x65 & n23067 ) | ( ~x34 & n23067 ) ;
  assign n23331 = ( x34 & ~n23067 ) | ( x34 & x65 ) | ( ~n23067 & x65 ) ;
  assign n23332 = ( n23330 & ~x65 ) | ( n23330 & n23331 ) | ( ~x65 & n23331 ) ;
  assign n23333 = ( n4635 & ~n4668 ) | ( n4635 & n23332 ) | ( ~n4668 & n23332 ) ;
  assign n23334 = ( n4635 & n23100 ) | ( n4635 & n23332 ) | ( n23100 & n23332 ) ;
  assign n23335 = ( n23333 & ~n23334 ) | ( n23333 & 1'b0 ) | ( ~n23334 & 1'b0 ) ;
  assign n23336 = n23329 | n23335 ;
  assign n23337 = ( n4910 & ~n23100 ) | ( n4910 & 1'b0 ) | ( ~n23100 & 1'b0 ) ;
  assign n23338 = ( x33 & ~n23337 ) | ( x33 & 1'b0 ) | ( ~n23337 & 1'b0 ) ;
  assign n23339 = ( n4916 & ~n23100 ) | ( n4916 & 1'b0 ) | ( ~n23100 & 1'b0 ) ;
  assign n23340 = n23338 | n23339 ;
  assign n23341 = ( x65 & ~n23340 ) | ( x65 & n4919 ) | ( ~n23340 & n4919 ) ;
  assign n23342 = ( x66 & ~n23336 ) | ( x66 & n23341 ) | ( ~n23336 & n23341 ) ;
  assign n23343 = ( x67 & ~n23328 ) | ( x67 & n23342 ) | ( ~n23328 & n23342 ) ;
  assign n23344 = ( x68 & ~n23323 ) | ( x68 & n23343 ) | ( ~n23323 & n23343 ) ;
  assign n23345 = ( x69 & ~n23315 ) | ( x69 & n23344 ) | ( ~n23315 & n23344 ) ;
  assign n23346 = ( x70 & ~n23307 ) | ( x70 & n23345 ) | ( ~n23307 & n23345 ) ;
  assign n23347 = ( x71 & ~n23299 ) | ( x71 & n23346 ) | ( ~n23299 & n23346 ) ;
  assign n23348 = ( x72 & ~n23291 ) | ( x72 & n23347 ) | ( ~n23291 & n23347 ) ;
  assign n23349 = ( x73 & ~n23283 ) | ( x73 & n23348 ) | ( ~n23283 & n23348 ) ;
  assign n23350 = ( x74 & ~n23275 ) | ( x74 & n23349 ) | ( ~n23275 & n23349 ) ;
  assign n23351 = ( x75 & ~n23267 ) | ( x75 & n23350 ) | ( ~n23267 & n23350 ) ;
  assign n23352 = ( x76 & ~n23259 ) | ( x76 & n23351 ) | ( ~n23259 & n23351 ) ;
  assign n23353 = ( x77 & ~n23251 ) | ( x77 & n23352 ) | ( ~n23251 & n23352 ) ;
  assign n23354 = ( x78 & ~n23243 ) | ( x78 & n23353 ) | ( ~n23243 & n23353 ) ;
  assign n23355 = ( x79 & ~n23235 ) | ( x79 & n23354 ) | ( ~n23235 & n23354 ) ;
  assign n23356 = ( x80 & ~n23227 ) | ( x80 & n23355 ) | ( ~n23227 & n23355 ) ;
  assign n23357 = ( x81 & ~n23219 ) | ( x81 & n23356 ) | ( ~n23219 & n23356 ) ;
  assign n23358 = ( x82 & ~n23211 ) | ( x82 & n23357 ) | ( ~n23211 & n23357 ) ;
  assign n23359 = ( x83 & ~n23203 ) | ( x83 & n23358 ) | ( ~n23203 & n23358 ) ;
  assign n23360 = ( x84 & ~n23195 ) | ( x84 & n23359 ) | ( ~n23195 & n23359 ) ;
  assign n23361 = ( x85 & ~n23187 ) | ( x85 & n23360 ) | ( ~n23187 & n23360 ) ;
  assign n23362 = ( x86 & ~n23179 ) | ( x86 & n23361 ) | ( ~n23179 & n23361 ) ;
  assign n23363 = ( x87 & ~n23171 ) | ( x87 & n23362 ) | ( ~n23171 & n23362 ) ;
  assign n23364 = ( x88 & ~n23163 ) | ( x88 & n23363 ) | ( ~n23163 & n23363 ) ;
  assign n23365 = ( x89 & ~n23155 ) | ( x89 & n23364 ) | ( ~n23155 & n23364 ) ;
  assign n23366 = ( x90 & ~n23147 ) | ( x90 & n23365 ) | ( ~n23147 & n23365 ) ;
  assign n23367 = ( x91 & ~n23139 ) | ( x91 & n23366 ) | ( ~n23139 & n23366 ) ;
  assign n23368 = ( x92 & ~n23131 ) | ( x92 & n23367 ) | ( ~n23131 & n23367 ) ;
  assign n23369 = ( x93 & ~n23123 ) | ( x93 & n23368 ) | ( ~n23123 & n23368 ) ;
  assign n23370 = ( x94 & ~n23115 ) | ( x94 & n23369 ) | ( ~n23115 & n23369 ) ;
  assign n23371 = ( x95 & ~n23107 ) | ( x95 & n23370 ) | ( ~n23107 & n23370 ) ;
  assign n23372 = n274 | n23371 ;
  assign n23373 = n23107 &  n23372 ;
  assign n23377 = ( n274 & n23107 ) | ( n274 & n23370 ) | ( n23107 & n23370 ) ;
  assign n23378 = ( x95 & ~n23377 ) | ( x95 & n23107 ) | ( ~n23377 & n23107 ) ;
  assign n23379 = ~x95 & n23378 ;
  assign n23380 = n23373 | n23379 ;
  assign n23381 = ~x96 & n23380 ;
  assign n23382 = n23115 &  n23372 ;
  assign n23374 = x94 | n23115 ;
  assign n23375 = x94 &  n23115 ;
  assign n23376 = ( n23374 & ~n23375 ) | ( n23374 & 1'b0 ) | ( ~n23375 & 1'b0 ) ;
  assign n23386 = ( n274 & n23369 ) | ( n274 & n23376 ) | ( n23369 & n23376 ) ;
  assign n23387 = ( n23369 & ~n23371 ) | ( n23369 & n23376 ) | ( ~n23371 & n23376 ) ;
  assign n23388 = ~n23386 & n23387 ;
  assign n23389 = n23382 | n23388 ;
  assign n23390 = n23123 &  n23372 ;
  assign n23383 = x93 | n23123 ;
  assign n23384 = x93 &  n23123 ;
  assign n23385 = ( n23383 & ~n23384 ) | ( n23383 & 1'b0 ) | ( ~n23384 & 1'b0 ) ;
  assign n23394 = ( n274 & n23368 ) | ( n274 & n23385 ) | ( n23368 & n23385 ) ;
  assign n23395 = ( n23368 & ~n23371 ) | ( n23368 & n23385 ) | ( ~n23371 & n23385 ) ;
  assign n23396 = ~n23394 & n23395 ;
  assign n23397 = n23390 | n23396 ;
  assign n23398 = n23131 &  n23372 ;
  assign n23391 = x92 | n23131 ;
  assign n23392 = x92 &  n23131 ;
  assign n23393 = ( n23391 & ~n23392 ) | ( n23391 & 1'b0 ) | ( ~n23392 & 1'b0 ) ;
  assign n23402 = ( n274 & n23367 ) | ( n274 & n23393 ) | ( n23367 & n23393 ) ;
  assign n23403 = ( n23367 & ~n23371 ) | ( n23367 & n23393 ) | ( ~n23371 & n23393 ) ;
  assign n23404 = ~n23402 & n23403 ;
  assign n23405 = n23398 | n23404 ;
  assign n23406 = n23139 &  n23372 ;
  assign n23399 = x91 | n23139 ;
  assign n23400 = x91 &  n23139 ;
  assign n23401 = ( n23399 & ~n23400 ) | ( n23399 & 1'b0 ) | ( ~n23400 & 1'b0 ) ;
  assign n23410 = ( n274 & n23366 ) | ( n274 & n23401 ) | ( n23366 & n23401 ) ;
  assign n23411 = ( n23366 & ~n23371 ) | ( n23366 & n23401 ) | ( ~n23371 & n23401 ) ;
  assign n23412 = ~n23410 & n23411 ;
  assign n23413 = n23406 | n23412 ;
  assign n23414 = n23147 &  n23372 ;
  assign n23407 = x90 | n23147 ;
  assign n23408 = x90 &  n23147 ;
  assign n23409 = ( n23407 & ~n23408 ) | ( n23407 & 1'b0 ) | ( ~n23408 & 1'b0 ) ;
  assign n23418 = ( n274 & n23365 ) | ( n274 & n23409 ) | ( n23365 & n23409 ) ;
  assign n23419 = ( n23365 & ~n23371 ) | ( n23365 & n23409 ) | ( ~n23371 & n23409 ) ;
  assign n23420 = ~n23418 & n23419 ;
  assign n23421 = n23414 | n23420 ;
  assign n23422 = n23155 &  n23372 ;
  assign n23415 = x89 | n23155 ;
  assign n23416 = x89 &  n23155 ;
  assign n23417 = ( n23415 & ~n23416 ) | ( n23415 & 1'b0 ) | ( ~n23416 & 1'b0 ) ;
  assign n23426 = ( n274 & n23364 ) | ( n274 & n23417 ) | ( n23364 & n23417 ) ;
  assign n23427 = ( n23364 & ~n23371 ) | ( n23364 & n23417 ) | ( ~n23371 & n23417 ) ;
  assign n23428 = ~n23426 & n23427 ;
  assign n23429 = n23422 | n23428 ;
  assign n23430 = n23163 &  n23372 ;
  assign n23423 = x88 | n23163 ;
  assign n23424 = x88 &  n23163 ;
  assign n23425 = ( n23423 & ~n23424 ) | ( n23423 & 1'b0 ) | ( ~n23424 & 1'b0 ) ;
  assign n23434 = ( n274 & n23363 ) | ( n274 & n23425 ) | ( n23363 & n23425 ) ;
  assign n23435 = ( n23363 & ~n23371 ) | ( n23363 & n23425 ) | ( ~n23371 & n23425 ) ;
  assign n23436 = ~n23434 & n23435 ;
  assign n23437 = n23430 | n23436 ;
  assign n23438 = n23171 &  n23372 ;
  assign n23431 = x87 | n23171 ;
  assign n23432 = x87 &  n23171 ;
  assign n23433 = ( n23431 & ~n23432 ) | ( n23431 & 1'b0 ) | ( ~n23432 & 1'b0 ) ;
  assign n23442 = ( n274 & n23362 ) | ( n274 & n23433 ) | ( n23362 & n23433 ) ;
  assign n23443 = ( n23362 & ~n23371 ) | ( n23362 & n23433 ) | ( ~n23371 & n23433 ) ;
  assign n23444 = ~n23442 & n23443 ;
  assign n23445 = n23438 | n23444 ;
  assign n23446 = n23179 &  n23372 ;
  assign n23439 = x86 | n23179 ;
  assign n23440 = x86 &  n23179 ;
  assign n23441 = ( n23439 & ~n23440 ) | ( n23439 & 1'b0 ) | ( ~n23440 & 1'b0 ) ;
  assign n23450 = ( n274 & n23361 ) | ( n274 & n23441 ) | ( n23361 & n23441 ) ;
  assign n23451 = ( n23361 & ~n23371 ) | ( n23361 & n23441 ) | ( ~n23371 & n23441 ) ;
  assign n23452 = ~n23450 & n23451 ;
  assign n23453 = n23446 | n23452 ;
  assign n23454 = n23187 &  n23372 ;
  assign n23447 = x85 | n23187 ;
  assign n23448 = x85 &  n23187 ;
  assign n23449 = ( n23447 & ~n23448 ) | ( n23447 & 1'b0 ) | ( ~n23448 & 1'b0 ) ;
  assign n23458 = ( n274 & n23360 ) | ( n274 & n23449 ) | ( n23360 & n23449 ) ;
  assign n23459 = ( n23360 & ~n23371 ) | ( n23360 & n23449 ) | ( ~n23371 & n23449 ) ;
  assign n23460 = ~n23458 & n23459 ;
  assign n23461 = n23454 | n23460 ;
  assign n23462 = n23195 &  n23372 ;
  assign n23455 = x84 | n23195 ;
  assign n23456 = x84 &  n23195 ;
  assign n23457 = ( n23455 & ~n23456 ) | ( n23455 & 1'b0 ) | ( ~n23456 & 1'b0 ) ;
  assign n23466 = ( n274 & n23359 ) | ( n274 & n23457 ) | ( n23359 & n23457 ) ;
  assign n23467 = ( n23359 & ~n23371 ) | ( n23359 & n23457 ) | ( ~n23371 & n23457 ) ;
  assign n23468 = ~n23466 & n23467 ;
  assign n23469 = n23462 | n23468 ;
  assign n23470 = n23203 &  n23372 ;
  assign n23463 = x83 | n23203 ;
  assign n23464 = x83 &  n23203 ;
  assign n23465 = ( n23463 & ~n23464 ) | ( n23463 & 1'b0 ) | ( ~n23464 & 1'b0 ) ;
  assign n23474 = ( n274 & n23358 ) | ( n274 & n23465 ) | ( n23358 & n23465 ) ;
  assign n23475 = ( n23358 & ~n23371 ) | ( n23358 & n23465 ) | ( ~n23371 & n23465 ) ;
  assign n23476 = ~n23474 & n23475 ;
  assign n23477 = n23470 | n23476 ;
  assign n23478 = n23211 &  n23372 ;
  assign n23471 = x82 | n23211 ;
  assign n23472 = x82 &  n23211 ;
  assign n23473 = ( n23471 & ~n23472 ) | ( n23471 & 1'b0 ) | ( ~n23472 & 1'b0 ) ;
  assign n23482 = ( n274 & n23357 ) | ( n274 & n23473 ) | ( n23357 & n23473 ) ;
  assign n23483 = ( n23357 & ~n23371 ) | ( n23357 & n23473 ) | ( ~n23371 & n23473 ) ;
  assign n23484 = ~n23482 & n23483 ;
  assign n23485 = n23478 | n23484 ;
  assign n23486 = n23219 &  n23372 ;
  assign n23479 = x81 | n23219 ;
  assign n23480 = x81 &  n23219 ;
  assign n23481 = ( n23479 & ~n23480 ) | ( n23479 & 1'b0 ) | ( ~n23480 & 1'b0 ) ;
  assign n23490 = ( n274 & n23356 ) | ( n274 & n23481 ) | ( n23356 & n23481 ) ;
  assign n23491 = ( n23356 & ~n23371 ) | ( n23356 & n23481 ) | ( ~n23371 & n23481 ) ;
  assign n23492 = ~n23490 & n23491 ;
  assign n23493 = n23486 | n23492 ;
  assign n23494 = n23227 &  n23372 ;
  assign n23487 = x80 | n23227 ;
  assign n23488 = x80 &  n23227 ;
  assign n23489 = ( n23487 & ~n23488 ) | ( n23487 & 1'b0 ) | ( ~n23488 & 1'b0 ) ;
  assign n23498 = ( n274 & n23355 ) | ( n274 & n23489 ) | ( n23355 & n23489 ) ;
  assign n23499 = ( n23355 & ~n23371 ) | ( n23355 & n23489 ) | ( ~n23371 & n23489 ) ;
  assign n23500 = ~n23498 & n23499 ;
  assign n23501 = n23494 | n23500 ;
  assign n23502 = n23235 &  n23372 ;
  assign n23495 = x79 | n23235 ;
  assign n23496 = x79 &  n23235 ;
  assign n23497 = ( n23495 & ~n23496 ) | ( n23495 & 1'b0 ) | ( ~n23496 & 1'b0 ) ;
  assign n23506 = ( n274 & n23354 ) | ( n274 & n23497 ) | ( n23354 & n23497 ) ;
  assign n23507 = ( n23354 & ~n23371 ) | ( n23354 & n23497 ) | ( ~n23371 & n23497 ) ;
  assign n23508 = ~n23506 & n23507 ;
  assign n23509 = n23502 | n23508 ;
  assign n23510 = n23243 &  n23372 ;
  assign n23503 = x78 | n23243 ;
  assign n23504 = x78 &  n23243 ;
  assign n23505 = ( n23503 & ~n23504 ) | ( n23503 & 1'b0 ) | ( ~n23504 & 1'b0 ) ;
  assign n23514 = ( n274 & n23353 ) | ( n274 & n23505 ) | ( n23353 & n23505 ) ;
  assign n23515 = ( n23353 & ~n23371 ) | ( n23353 & n23505 ) | ( ~n23371 & n23505 ) ;
  assign n23516 = ~n23514 & n23515 ;
  assign n23517 = n23510 | n23516 ;
  assign n23518 = n23251 &  n23372 ;
  assign n23511 = x77 | n23251 ;
  assign n23512 = x77 &  n23251 ;
  assign n23513 = ( n23511 & ~n23512 ) | ( n23511 & 1'b0 ) | ( ~n23512 & 1'b0 ) ;
  assign n23522 = ( n274 & n23352 ) | ( n274 & n23513 ) | ( n23352 & n23513 ) ;
  assign n23523 = ( n23352 & ~n23371 ) | ( n23352 & n23513 ) | ( ~n23371 & n23513 ) ;
  assign n23524 = ~n23522 & n23523 ;
  assign n23525 = n23518 | n23524 ;
  assign n23526 = n23259 &  n23372 ;
  assign n23519 = x76 | n23259 ;
  assign n23520 = x76 &  n23259 ;
  assign n23521 = ( n23519 & ~n23520 ) | ( n23519 & 1'b0 ) | ( ~n23520 & 1'b0 ) ;
  assign n23530 = ( n274 & n23351 ) | ( n274 & n23521 ) | ( n23351 & n23521 ) ;
  assign n23531 = ( n23351 & ~n23371 ) | ( n23351 & n23521 ) | ( ~n23371 & n23521 ) ;
  assign n23532 = ~n23530 & n23531 ;
  assign n23533 = n23526 | n23532 ;
  assign n23534 = n23267 &  n23372 ;
  assign n23527 = x75 | n23267 ;
  assign n23528 = x75 &  n23267 ;
  assign n23529 = ( n23527 & ~n23528 ) | ( n23527 & 1'b0 ) | ( ~n23528 & 1'b0 ) ;
  assign n23538 = ( n274 & n23350 ) | ( n274 & n23529 ) | ( n23350 & n23529 ) ;
  assign n23539 = ( n23350 & ~n23371 ) | ( n23350 & n23529 ) | ( ~n23371 & n23529 ) ;
  assign n23540 = ~n23538 & n23539 ;
  assign n23541 = n23534 | n23540 ;
  assign n23542 = n23275 &  n23372 ;
  assign n23535 = x74 | n23275 ;
  assign n23536 = x74 &  n23275 ;
  assign n23537 = ( n23535 & ~n23536 ) | ( n23535 & 1'b0 ) | ( ~n23536 & 1'b0 ) ;
  assign n23546 = ( n274 & n23349 ) | ( n274 & n23537 ) | ( n23349 & n23537 ) ;
  assign n23547 = ( n23349 & ~n23371 ) | ( n23349 & n23537 ) | ( ~n23371 & n23537 ) ;
  assign n23548 = ~n23546 & n23547 ;
  assign n23549 = n23542 | n23548 ;
  assign n23550 = n23283 &  n23372 ;
  assign n23543 = x73 | n23283 ;
  assign n23544 = x73 &  n23283 ;
  assign n23545 = ( n23543 & ~n23544 ) | ( n23543 & 1'b0 ) | ( ~n23544 & 1'b0 ) ;
  assign n23554 = ( n274 & n23348 ) | ( n274 & n23545 ) | ( n23348 & n23545 ) ;
  assign n23555 = ( n23348 & ~n23371 ) | ( n23348 & n23545 ) | ( ~n23371 & n23545 ) ;
  assign n23556 = ~n23554 & n23555 ;
  assign n23557 = n23550 | n23556 ;
  assign n23558 = n23291 &  n23372 ;
  assign n23551 = x72 | n23291 ;
  assign n23552 = x72 &  n23291 ;
  assign n23553 = ( n23551 & ~n23552 ) | ( n23551 & 1'b0 ) | ( ~n23552 & 1'b0 ) ;
  assign n23562 = ( n274 & n23347 ) | ( n274 & n23553 ) | ( n23347 & n23553 ) ;
  assign n23563 = ( n23347 & ~n23371 ) | ( n23347 & n23553 ) | ( ~n23371 & n23553 ) ;
  assign n23564 = ~n23562 & n23563 ;
  assign n23565 = n23558 | n23564 ;
  assign n23566 = n23299 &  n23372 ;
  assign n23559 = x71 | n23299 ;
  assign n23560 = x71 &  n23299 ;
  assign n23561 = ( n23559 & ~n23560 ) | ( n23559 & 1'b0 ) | ( ~n23560 & 1'b0 ) ;
  assign n23570 = ( n274 & n23346 ) | ( n274 & n23561 ) | ( n23346 & n23561 ) ;
  assign n23571 = ( n23346 & ~n23371 ) | ( n23346 & n23561 ) | ( ~n23371 & n23561 ) ;
  assign n23572 = ~n23570 & n23571 ;
  assign n23573 = n23566 | n23572 ;
  assign n23574 = n23307 &  n23372 ;
  assign n23567 = x70 | n23307 ;
  assign n23568 = x70 &  n23307 ;
  assign n23569 = ( n23567 & ~n23568 ) | ( n23567 & 1'b0 ) | ( ~n23568 & 1'b0 ) ;
  assign n23578 = ( n274 & n23345 ) | ( n274 & n23569 ) | ( n23345 & n23569 ) ;
  assign n23579 = ( n23345 & ~n23371 ) | ( n23345 & n23569 ) | ( ~n23371 & n23569 ) ;
  assign n23580 = ~n23578 & n23579 ;
  assign n23581 = n23574 | n23580 ;
  assign n23582 = n23315 &  n23372 ;
  assign n23575 = x69 | n23315 ;
  assign n23576 = x69 &  n23315 ;
  assign n23577 = ( n23575 & ~n23576 ) | ( n23575 & 1'b0 ) | ( ~n23576 & 1'b0 ) ;
  assign n23586 = ( n274 & n23344 ) | ( n274 & n23577 ) | ( n23344 & n23577 ) ;
  assign n23587 = ( n23344 & ~n23371 ) | ( n23344 & n23577 ) | ( ~n23371 & n23577 ) ;
  assign n23588 = ~n23586 & n23587 ;
  assign n23589 = n23582 | n23588 ;
  assign n23590 = n23323 &  n23372 ;
  assign n23583 = x68 | n23323 ;
  assign n23584 = x68 &  n23323 ;
  assign n23585 = ( n23583 & ~n23584 ) | ( n23583 & 1'b0 ) | ( ~n23584 & 1'b0 ) ;
  assign n23594 = ( n274 & n23343 ) | ( n274 & n23585 ) | ( n23343 & n23585 ) ;
  assign n23595 = ( n23343 & ~n23371 ) | ( n23343 & n23585 ) | ( ~n23371 & n23585 ) ;
  assign n23596 = ~n23594 & n23595 ;
  assign n23597 = n23590 | n23596 ;
  assign n23598 = n23328 &  n23372 ;
  assign n23591 = x67 | n23328 ;
  assign n23592 = x67 &  n23328 ;
  assign n23593 = ( n23591 & ~n23592 ) | ( n23591 & 1'b0 ) | ( ~n23592 & 1'b0 ) ;
  assign n23602 = ( n274 & n23342 ) | ( n274 & n23593 ) | ( n23342 & n23593 ) ;
  assign n23603 = ( n23342 & ~n23371 ) | ( n23342 & n23593 ) | ( ~n23371 & n23593 ) ;
  assign n23604 = ~n23602 & n23603 ;
  assign n23605 = n23598 | n23604 ;
  assign n23606 = n23336 &  n23372 ;
  assign n23599 = x66 | n23336 ;
  assign n23600 = x66 &  n23336 ;
  assign n23601 = ( n23599 & ~n23600 ) | ( n23599 & 1'b0 ) | ( ~n23600 & 1'b0 ) ;
  assign n23610 = ( n274 & n23341 ) | ( n274 & n23601 ) | ( n23341 & n23601 ) ;
  assign n23611 = ( n23341 & ~n23371 ) | ( n23341 & n23601 ) | ( ~n23371 & n23601 ) ;
  assign n23612 = ~n23610 & n23611 ;
  assign n23613 = n23606 | n23612 ;
  assign n23614 = n23340 &  n23372 ;
  assign n23607 = x65 &  n23340 ;
  assign n23608 = x65 | n23339 ;
  assign n23609 = n23338 | n23608 ;
  assign n23615 = ~n23607 & n23609 ;
  assign n23616 = ( n4919 & ~n23371 ) | ( n4919 & n23615 ) | ( ~n23371 & n23615 ) ;
  assign n23617 = ( n274 & n4919 ) | ( n274 & n23615 ) | ( n4919 & n23615 ) ;
  assign n23618 = ( n23616 & ~n23617 ) | ( n23616 & 1'b0 ) | ( ~n23617 & 1'b0 ) ;
  assign n23619 = n23614 | n23618 ;
  assign n23620 = ( n5052 & ~n23371 ) | ( n5052 & 1'b0 ) | ( ~n23371 & 1'b0 ) ;
  assign n23621 = ( x32 & ~n23620 ) | ( x32 & 1'b0 ) | ( ~n23620 & 1'b0 ) ;
  assign n23622 = ( n5057 & ~n23371 ) | ( n5057 & 1'b0 ) | ( ~n23371 & 1'b0 ) ;
  assign n23623 = n23621 | n23622 ;
  assign n23624 = ( x65 & ~n23623 ) | ( x65 & n5060 ) | ( ~n23623 & n5060 ) ;
  assign n23625 = ( x66 & ~n23619 ) | ( x66 & n23624 ) | ( ~n23619 & n23624 ) ;
  assign n23626 = ( x67 & ~n23613 ) | ( x67 & n23625 ) | ( ~n23613 & n23625 ) ;
  assign n23627 = ( x68 & ~n23605 ) | ( x68 & n23626 ) | ( ~n23605 & n23626 ) ;
  assign n23628 = ( x69 & ~n23597 ) | ( x69 & n23627 ) | ( ~n23597 & n23627 ) ;
  assign n23629 = ( x70 & ~n23589 ) | ( x70 & n23628 ) | ( ~n23589 & n23628 ) ;
  assign n23630 = ( x71 & ~n23581 ) | ( x71 & n23629 ) | ( ~n23581 & n23629 ) ;
  assign n23631 = ( x72 & ~n23573 ) | ( x72 & n23630 ) | ( ~n23573 & n23630 ) ;
  assign n23632 = ( x73 & ~n23565 ) | ( x73 & n23631 ) | ( ~n23565 & n23631 ) ;
  assign n23633 = ( x74 & ~n23557 ) | ( x74 & n23632 ) | ( ~n23557 & n23632 ) ;
  assign n23634 = ( x75 & ~n23549 ) | ( x75 & n23633 ) | ( ~n23549 & n23633 ) ;
  assign n23635 = ( x76 & ~n23541 ) | ( x76 & n23634 ) | ( ~n23541 & n23634 ) ;
  assign n23636 = ( x77 & ~n23533 ) | ( x77 & n23635 ) | ( ~n23533 & n23635 ) ;
  assign n23637 = ( x78 & ~n23525 ) | ( x78 & n23636 ) | ( ~n23525 & n23636 ) ;
  assign n23638 = ( x79 & ~n23517 ) | ( x79 & n23637 ) | ( ~n23517 & n23637 ) ;
  assign n23639 = ( x80 & ~n23509 ) | ( x80 & n23638 ) | ( ~n23509 & n23638 ) ;
  assign n23640 = ( x81 & ~n23501 ) | ( x81 & n23639 ) | ( ~n23501 & n23639 ) ;
  assign n23641 = ( x82 & ~n23493 ) | ( x82 & n23640 ) | ( ~n23493 & n23640 ) ;
  assign n23642 = ( x83 & ~n23485 ) | ( x83 & n23641 ) | ( ~n23485 & n23641 ) ;
  assign n23643 = ( x84 & ~n23477 ) | ( x84 & n23642 ) | ( ~n23477 & n23642 ) ;
  assign n23644 = ( x85 & ~n23469 ) | ( x85 & n23643 ) | ( ~n23469 & n23643 ) ;
  assign n23645 = ( x86 & ~n23461 ) | ( x86 & n23644 ) | ( ~n23461 & n23644 ) ;
  assign n23646 = ( x87 & ~n23453 ) | ( x87 & n23645 ) | ( ~n23453 & n23645 ) ;
  assign n23647 = ( x88 & ~n23445 ) | ( x88 & n23646 ) | ( ~n23445 & n23646 ) ;
  assign n23648 = ( x89 & ~n23437 ) | ( x89 & n23647 ) | ( ~n23437 & n23647 ) ;
  assign n23649 = ( x90 & ~n23429 ) | ( x90 & n23648 ) | ( ~n23429 & n23648 ) ;
  assign n23650 = ( x91 & ~n23421 ) | ( x91 & n23649 ) | ( ~n23421 & n23649 ) ;
  assign n23651 = ( x92 & ~n23413 ) | ( x92 & n23650 ) | ( ~n23413 & n23650 ) ;
  assign n23652 = ( x93 & ~n23405 ) | ( x93 & n23651 ) | ( ~n23405 & n23651 ) ;
  assign n23653 = ( x94 & ~n23397 ) | ( x94 & n23652 ) | ( ~n23397 & n23652 ) ;
  assign n23654 = ( x95 & ~n23389 ) | ( x95 & n23653 ) | ( ~n23389 & n23653 ) ;
  assign n23655 = ( x96 & ~n23373 ) | ( x96 & 1'b0 ) | ( ~n23373 & 1'b0 ) ;
  assign n23656 = ~n23379 & n23655 ;
  assign n23657 = ( n23654 & ~n23381 ) | ( n23654 & n23656 ) | ( ~n23381 & n23656 ) ;
  assign n23658 = ( n23381 & ~n256 ) | ( n23381 & n23657 ) | ( ~n256 & n23657 ) ;
  assign n23659 = n256 | n23658 ;
  assign n23666 = n274 &  n23107 ;
  assign n23667 = n23659 &  n23666 ;
  assign n23660 = ~n23380 |  n274 ;
  assign n23661 = n23659 &  n23660 ;
  assign n23665 = n23381 | n23656 ;
  assign n23669 = ( n23654 & n23661 ) | ( n23654 & n23665 ) | ( n23661 & n23665 ) ;
  assign n23668 = n23654 | n23665 ;
  assign n23670 = ( n23667 & ~n23669 ) | ( n23667 & n23668 ) | ( ~n23669 & n23668 ) ;
  assign n23674 = n23389 &  n23660 ;
  assign n23675 = n23659 &  n23674 ;
  assign n23662 = x95 | n23389 ;
  assign n23663 = x95 &  n23389 ;
  assign n23664 = ( n23662 & ~n23663 ) | ( n23662 & 1'b0 ) | ( ~n23663 & 1'b0 ) ;
  assign n23677 = ( n23653 & n23661 ) | ( n23653 & n23664 ) | ( n23661 & n23664 ) ;
  assign n23676 = n23653 | n23664 ;
  assign n23678 = ( n23675 & ~n23677 ) | ( n23675 & n23676 ) | ( ~n23677 & n23676 ) ;
  assign n23682 = n23397 &  n23660 ;
  assign n23683 = n23659 &  n23682 ;
  assign n23671 = x94 | n23397 ;
  assign n23672 = x94 &  n23397 ;
  assign n23673 = ( n23671 & ~n23672 ) | ( n23671 & 1'b0 ) | ( ~n23672 & 1'b0 ) ;
  assign n23685 = ( n23652 & n23661 ) | ( n23652 & n23673 ) | ( n23661 & n23673 ) ;
  assign n23684 = n23652 | n23673 ;
  assign n23686 = ( n23683 & ~n23685 ) | ( n23683 & n23684 ) | ( ~n23685 & n23684 ) ;
  assign n23690 = n23405 &  n23660 ;
  assign n23691 = n23659 &  n23690 ;
  assign n23679 = x93 | n23405 ;
  assign n23680 = x93 &  n23405 ;
  assign n23681 = ( n23679 & ~n23680 ) | ( n23679 & 1'b0 ) | ( ~n23680 & 1'b0 ) ;
  assign n23693 = ( n23651 & n23661 ) | ( n23651 & n23681 ) | ( n23661 & n23681 ) ;
  assign n23692 = n23651 | n23681 ;
  assign n23694 = ( n23691 & ~n23693 ) | ( n23691 & n23692 ) | ( ~n23693 & n23692 ) ;
  assign n23698 = n23413 &  n23660 ;
  assign n23699 = n23659 &  n23698 ;
  assign n23687 = x92 | n23413 ;
  assign n23688 = x92 &  n23413 ;
  assign n23689 = ( n23687 & ~n23688 ) | ( n23687 & 1'b0 ) | ( ~n23688 & 1'b0 ) ;
  assign n23701 = ( n23650 & n23661 ) | ( n23650 & n23689 ) | ( n23661 & n23689 ) ;
  assign n23700 = n23650 | n23689 ;
  assign n23702 = ( n23699 & ~n23701 ) | ( n23699 & n23700 ) | ( ~n23701 & n23700 ) ;
  assign n23706 = n23421 &  n23660 ;
  assign n23707 = n23659 &  n23706 ;
  assign n23695 = x91 | n23421 ;
  assign n23696 = x91 &  n23421 ;
  assign n23697 = ( n23695 & ~n23696 ) | ( n23695 & 1'b0 ) | ( ~n23696 & 1'b0 ) ;
  assign n23709 = ( n23649 & n23661 ) | ( n23649 & n23697 ) | ( n23661 & n23697 ) ;
  assign n23708 = n23649 | n23697 ;
  assign n23710 = ( n23707 & ~n23709 ) | ( n23707 & n23708 ) | ( ~n23709 & n23708 ) ;
  assign n23714 = n23429 &  n23660 ;
  assign n23715 = n23659 &  n23714 ;
  assign n23703 = x90 | n23429 ;
  assign n23704 = x90 &  n23429 ;
  assign n23705 = ( n23703 & ~n23704 ) | ( n23703 & 1'b0 ) | ( ~n23704 & 1'b0 ) ;
  assign n23717 = ( n23648 & n23661 ) | ( n23648 & n23705 ) | ( n23661 & n23705 ) ;
  assign n23716 = n23648 | n23705 ;
  assign n23718 = ( n23715 & ~n23717 ) | ( n23715 & n23716 ) | ( ~n23717 & n23716 ) ;
  assign n23722 = n23437 &  n23660 ;
  assign n23723 = n23659 &  n23722 ;
  assign n23711 = x89 | n23437 ;
  assign n23712 = x89 &  n23437 ;
  assign n23713 = ( n23711 & ~n23712 ) | ( n23711 & 1'b0 ) | ( ~n23712 & 1'b0 ) ;
  assign n23725 = ( n23647 & n23661 ) | ( n23647 & n23713 ) | ( n23661 & n23713 ) ;
  assign n23724 = n23647 | n23713 ;
  assign n23726 = ( n23723 & ~n23725 ) | ( n23723 & n23724 ) | ( ~n23725 & n23724 ) ;
  assign n23730 = n23445 &  n23660 ;
  assign n23731 = n23659 &  n23730 ;
  assign n23719 = x88 | n23445 ;
  assign n23720 = x88 &  n23445 ;
  assign n23721 = ( n23719 & ~n23720 ) | ( n23719 & 1'b0 ) | ( ~n23720 & 1'b0 ) ;
  assign n23733 = ( n23646 & n23661 ) | ( n23646 & n23721 ) | ( n23661 & n23721 ) ;
  assign n23732 = n23646 | n23721 ;
  assign n23734 = ( n23731 & ~n23733 ) | ( n23731 & n23732 ) | ( ~n23733 & n23732 ) ;
  assign n23738 = n23453 &  n23660 ;
  assign n23739 = n23659 &  n23738 ;
  assign n23727 = x87 | n23453 ;
  assign n23728 = x87 &  n23453 ;
  assign n23729 = ( n23727 & ~n23728 ) | ( n23727 & 1'b0 ) | ( ~n23728 & 1'b0 ) ;
  assign n23741 = ( n23645 & n23661 ) | ( n23645 & n23729 ) | ( n23661 & n23729 ) ;
  assign n23740 = n23645 | n23729 ;
  assign n23742 = ( n23739 & ~n23741 ) | ( n23739 & n23740 ) | ( ~n23741 & n23740 ) ;
  assign n23746 = n23461 &  n23660 ;
  assign n23747 = n23659 &  n23746 ;
  assign n23735 = x86 | n23461 ;
  assign n23736 = x86 &  n23461 ;
  assign n23737 = ( n23735 & ~n23736 ) | ( n23735 & 1'b0 ) | ( ~n23736 & 1'b0 ) ;
  assign n23749 = ( n23644 & n23661 ) | ( n23644 & n23737 ) | ( n23661 & n23737 ) ;
  assign n23748 = n23644 | n23737 ;
  assign n23750 = ( n23747 & ~n23749 ) | ( n23747 & n23748 ) | ( ~n23749 & n23748 ) ;
  assign n23754 = n23469 &  n23660 ;
  assign n23755 = n23659 &  n23754 ;
  assign n23743 = x85 | n23469 ;
  assign n23744 = x85 &  n23469 ;
  assign n23745 = ( n23743 & ~n23744 ) | ( n23743 & 1'b0 ) | ( ~n23744 & 1'b0 ) ;
  assign n23757 = ( n23643 & n23661 ) | ( n23643 & n23745 ) | ( n23661 & n23745 ) ;
  assign n23756 = n23643 | n23745 ;
  assign n23758 = ( n23755 & ~n23757 ) | ( n23755 & n23756 ) | ( ~n23757 & n23756 ) ;
  assign n23762 = n23477 &  n23660 ;
  assign n23763 = n23659 &  n23762 ;
  assign n23751 = x84 | n23477 ;
  assign n23752 = x84 &  n23477 ;
  assign n23753 = ( n23751 & ~n23752 ) | ( n23751 & 1'b0 ) | ( ~n23752 & 1'b0 ) ;
  assign n23765 = ( n23642 & n23661 ) | ( n23642 & n23753 ) | ( n23661 & n23753 ) ;
  assign n23764 = n23642 | n23753 ;
  assign n23766 = ( n23763 & ~n23765 ) | ( n23763 & n23764 ) | ( ~n23765 & n23764 ) ;
  assign n23770 = n23485 &  n23660 ;
  assign n23771 = n23659 &  n23770 ;
  assign n23759 = x83 | n23485 ;
  assign n23760 = x83 &  n23485 ;
  assign n23761 = ( n23759 & ~n23760 ) | ( n23759 & 1'b0 ) | ( ~n23760 & 1'b0 ) ;
  assign n23773 = ( n23641 & n23661 ) | ( n23641 & n23761 ) | ( n23661 & n23761 ) ;
  assign n23772 = n23641 | n23761 ;
  assign n23774 = ( n23771 & ~n23773 ) | ( n23771 & n23772 ) | ( ~n23773 & n23772 ) ;
  assign n23778 = n23493 &  n23660 ;
  assign n23779 = n23659 &  n23778 ;
  assign n23767 = x82 | n23493 ;
  assign n23768 = x82 &  n23493 ;
  assign n23769 = ( n23767 & ~n23768 ) | ( n23767 & 1'b0 ) | ( ~n23768 & 1'b0 ) ;
  assign n23781 = ( n23640 & n23661 ) | ( n23640 & n23769 ) | ( n23661 & n23769 ) ;
  assign n23780 = n23640 | n23769 ;
  assign n23782 = ( n23779 & ~n23781 ) | ( n23779 & n23780 ) | ( ~n23781 & n23780 ) ;
  assign n23786 = n23501 &  n23660 ;
  assign n23787 = n23659 &  n23786 ;
  assign n23775 = x81 | n23501 ;
  assign n23776 = x81 &  n23501 ;
  assign n23777 = ( n23775 & ~n23776 ) | ( n23775 & 1'b0 ) | ( ~n23776 & 1'b0 ) ;
  assign n23789 = ( n23639 & n23661 ) | ( n23639 & n23777 ) | ( n23661 & n23777 ) ;
  assign n23788 = n23639 | n23777 ;
  assign n23790 = ( n23787 & ~n23789 ) | ( n23787 & n23788 ) | ( ~n23789 & n23788 ) ;
  assign n23794 = n23509 &  n23660 ;
  assign n23795 = n23659 &  n23794 ;
  assign n23783 = x80 | n23509 ;
  assign n23784 = x80 &  n23509 ;
  assign n23785 = ( n23783 & ~n23784 ) | ( n23783 & 1'b0 ) | ( ~n23784 & 1'b0 ) ;
  assign n23797 = ( n23638 & n23661 ) | ( n23638 & n23785 ) | ( n23661 & n23785 ) ;
  assign n23796 = n23638 | n23785 ;
  assign n23798 = ( n23795 & ~n23797 ) | ( n23795 & n23796 ) | ( ~n23797 & n23796 ) ;
  assign n23802 = n23517 &  n23660 ;
  assign n23803 = n23659 &  n23802 ;
  assign n23791 = x79 | n23517 ;
  assign n23792 = x79 &  n23517 ;
  assign n23793 = ( n23791 & ~n23792 ) | ( n23791 & 1'b0 ) | ( ~n23792 & 1'b0 ) ;
  assign n23805 = ( n23637 & n23661 ) | ( n23637 & n23793 ) | ( n23661 & n23793 ) ;
  assign n23804 = n23637 | n23793 ;
  assign n23806 = ( n23803 & ~n23805 ) | ( n23803 & n23804 ) | ( ~n23805 & n23804 ) ;
  assign n23810 = n23525 &  n23660 ;
  assign n23811 = n23659 &  n23810 ;
  assign n23799 = x78 | n23525 ;
  assign n23800 = x78 &  n23525 ;
  assign n23801 = ( n23799 & ~n23800 ) | ( n23799 & 1'b0 ) | ( ~n23800 & 1'b0 ) ;
  assign n23813 = ( n23636 & n23661 ) | ( n23636 & n23801 ) | ( n23661 & n23801 ) ;
  assign n23812 = n23636 | n23801 ;
  assign n23814 = ( n23811 & ~n23813 ) | ( n23811 & n23812 ) | ( ~n23813 & n23812 ) ;
  assign n23818 = n23533 &  n23660 ;
  assign n23819 = n23659 &  n23818 ;
  assign n23807 = x77 | n23533 ;
  assign n23808 = x77 &  n23533 ;
  assign n23809 = ( n23807 & ~n23808 ) | ( n23807 & 1'b0 ) | ( ~n23808 & 1'b0 ) ;
  assign n23821 = ( n23635 & n23661 ) | ( n23635 & n23809 ) | ( n23661 & n23809 ) ;
  assign n23820 = n23635 | n23809 ;
  assign n23822 = ( n23819 & ~n23821 ) | ( n23819 & n23820 ) | ( ~n23821 & n23820 ) ;
  assign n23826 = n23541 &  n23660 ;
  assign n23827 = n23659 &  n23826 ;
  assign n23815 = x76 | n23541 ;
  assign n23816 = x76 &  n23541 ;
  assign n23817 = ( n23815 & ~n23816 ) | ( n23815 & 1'b0 ) | ( ~n23816 & 1'b0 ) ;
  assign n23829 = ( n23634 & n23661 ) | ( n23634 & n23817 ) | ( n23661 & n23817 ) ;
  assign n23828 = n23634 | n23817 ;
  assign n23830 = ( n23827 & ~n23829 ) | ( n23827 & n23828 ) | ( ~n23829 & n23828 ) ;
  assign n23834 = n23549 &  n23660 ;
  assign n23835 = n23659 &  n23834 ;
  assign n23823 = x75 | n23549 ;
  assign n23824 = x75 &  n23549 ;
  assign n23825 = ( n23823 & ~n23824 ) | ( n23823 & 1'b0 ) | ( ~n23824 & 1'b0 ) ;
  assign n23837 = ( n23633 & n23661 ) | ( n23633 & n23825 ) | ( n23661 & n23825 ) ;
  assign n23836 = n23633 | n23825 ;
  assign n23838 = ( n23835 & ~n23837 ) | ( n23835 & n23836 ) | ( ~n23837 & n23836 ) ;
  assign n23842 = n23557 &  n23660 ;
  assign n23843 = n23659 &  n23842 ;
  assign n23831 = x74 | n23557 ;
  assign n23832 = x74 &  n23557 ;
  assign n23833 = ( n23831 & ~n23832 ) | ( n23831 & 1'b0 ) | ( ~n23832 & 1'b0 ) ;
  assign n23845 = ( n23632 & n23661 ) | ( n23632 & n23833 ) | ( n23661 & n23833 ) ;
  assign n23844 = n23632 | n23833 ;
  assign n23846 = ( n23843 & ~n23845 ) | ( n23843 & n23844 ) | ( ~n23845 & n23844 ) ;
  assign n23850 = n23565 &  n23660 ;
  assign n23851 = n23659 &  n23850 ;
  assign n23839 = x73 | n23565 ;
  assign n23840 = x73 &  n23565 ;
  assign n23841 = ( n23839 & ~n23840 ) | ( n23839 & 1'b0 ) | ( ~n23840 & 1'b0 ) ;
  assign n23853 = ( n23631 & n23661 ) | ( n23631 & n23841 ) | ( n23661 & n23841 ) ;
  assign n23852 = n23631 | n23841 ;
  assign n23854 = ( n23851 & ~n23853 ) | ( n23851 & n23852 ) | ( ~n23853 & n23852 ) ;
  assign n23858 = n23573 &  n23660 ;
  assign n23859 = n23659 &  n23858 ;
  assign n23847 = x72 | n23573 ;
  assign n23848 = x72 &  n23573 ;
  assign n23849 = ( n23847 & ~n23848 ) | ( n23847 & 1'b0 ) | ( ~n23848 & 1'b0 ) ;
  assign n23861 = ( n23630 & n23661 ) | ( n23630 & n23849 ) | ( n23661 & n23849 ) ;
  assign n23860 = n23630 | n23849 ;
  assign n23862 = ( n23859 & ~n23861 ) | ( n23859 & n23860 ) | ( ~n23861 & n23860 ) ;
  assign n23866 = n23581 &  n23660 ;
  assign n23867 = n23659 &  n23866 ;
  assign n23855 = x71 | n23581 ;
  assign n23856 = x71 &  n23581 ;
  assign n23857 = ( n23855 & ~n23856 ) | ( n23855 & 1'b0 ) | ( ~n23856 & 1'b0 ) ;
  assign n23869 = ( n23629 & n23661 ) | ( n23629 & n23857 ) | ( n23661 & n23857 ) ;
  assign n23868 = n23629 | n23857 ;
  assign n23870 = ( n23867 & ~n23869 ) | ( n23867 & n23868 ) | ( ~n23869 & n23868 ) ;
  assign n23874 = n23589 &  n23660 ;
  assign n23875 = n23659 &  n23874 ;
  assign n23863 = x70 | n23589 ;
  assign n23864 = x70 &  n23589 ;
  assign n23865 = ( n23863 & ~n23864 ) | ( n23863 & 1'b0 ) | ( ~n23864 & 1'b0 ) ;
  assign n23877 = ( n23628 & n23661 ) | ( n23628 & n23865 ) | ( n23661 & n23865 ) ;
  assign n23876 = n23628 | n23865 ;
  assign n23878 = ( n23875 & ~n23877 ) | ( n23875 & n23876 ) | ( ~n23877 & n23876 ) ;
  assign n23882 = n23597 &  n23660 ;
  assign n23883 = n23659 &  n23882 ;
  assign n23871 = x69 | n23597 ;
  assign n23872 = x69 &  n23597 ;
  assign n23873 = ( n23871 & ~n23872 ) | ( n23871 & 1'b0 ) | ( ~n23872 & 1'b0 ) ;
  assign n23885 = ( n23627 & n23661 ) | ( n23627 & n23873 ) | ( n23661 & n23873 ) ;
  assign n23884 = n23627 | n23873 ;
  assign n23886 = ( n23883 & ~n23885 ) | ( n23883 & n23884 ) | ( ~n23885 & n23884 ) ;
  assign n23890 = n23605 &  n23660 ;
  assign n23891 = n23659 &  n23890 ;
  assign n23879 = x68 | n23605 ;
  assign n23880 = x68 &  n23605 ;
  assign n23881 = ( n23879 & ~n23880 ) | ( n23879 & 1'b0 ) | ( ~n23880 & 1'b0 ) ;
  assign n23893 = ( n23626 & n23661 ) | ( n23626 & n23881 ) | ( n23661 & n23881 ) ;
  assign n23892 = n23626 | n23881 ;
  assign n23894 = ( n23891 & ~n23893 ) | ( n23891 & n23892 ) | ( ~n23893 & n23892 ) ;
  assign n23898 = n23613 &  n23660 ;
  assign n23899 = n23659 &  n23898 ;
  assign n23887 = x67 | n23613 ;
  assign n23888 = x67 &  n23613 ;
  assign n23889 = ( n23887 & ~n23888 ) | ( n23887 & 1'b0 ) | ( ~n23888 & 1'b0 ) ;
  assign n23901 = ( n23625 & n23661 ) | ( n23625 & n23889 ) | ( n23661 & n23889 ) ;
  assign n23900 = n23625 | n23889 ;
  assign n23902 = ( n23899 & ~n23901 ) | ( n23899 & n23900 ) | ( ~n23901 & n23900 ) ;
  assign n23903 = n23619 &  n23660 ;
  assign n23904 = n23659 &  n23903 ;
  assign n23895 = x66 | n23619 ;
  assign n23896 = x66 &  n23619 ;
  assign n23897 = ( n23895 & ~n23896 ) | ( n23895 & 1'b0 ) | ( ~n23896 & 1'b0 ) ;
  assign n23906 = ( n23624 & n23661 ) | ( n23624 & n23897 ) | ( n23661 & n23897 ) ;
  assign n23905 = n23624 | n23897 ;
  assign n23907 = ( n23904 & ~n23906 ) | ( n23904 & n23905 ) | ( ~n23906 & n23905 ) ;
  assign n23908 = ( x65 & ~n5060 ) | ( x65 & n23623 ) | ( ~n5060 & n23623 ) ;
  assign n23909 = ( n23624 & ~x65 ) | ( n23624 & n23908 ) | ( ~x65 & n23908 ) ;
  assign n23910 = ~n23661 & n23909 ;
  assign n23911 = n23623 &  n23660 ;
  assign n23912 = n23659 &  n23911 ;
  assign n23913 = n23910 | n23912 ;
  assign n23914 = ( x64 & ~n23661 ) | ( x64 & 1'b0 ) | ( ~n23661 & 1'b0 ) ;
  assign n23915 = ( x31 & ~n23914 ) | ( x31 & 1'b0 ) | ( ~n23914 & 1'b0 ) ;
  assign n23916 = ( n5060 & ~n23661 ) | ( n5060 & 1'b0 ) | ( ~n23661 & 1'b0 ) ;
  assign n23917 = n23915 | n23916 ;
  assign n23918 = ( x65 & ~n23917 ) | ( x65 & n5505 ) | ( ~n23917 & n5505 ) ;
  assign n23919 = ( x66 & ~n23913 ) | ( x66 & n23918 ) | ( ~n23913 & n23918 ) ;
  assign n23920 = ( x67 & ~n23907 ) | ( x67 & n23919 ) | ( ~n23907 & n23919 ) ;
  assign n23921 = ( x68 & ~n23902 ) | ( x68 & n23920 ) | ( ~n23902 & n23920 ) ;
  assign n23922 = ( x69 & ~n23894 ) | ( x69 & n23921 ) | ( ~n23894 & n23921 ) ;
  assign n23923 = ( x70 & ~n23886 ) | ( x70 & n23922 ) | ( ~n23886 & n23922 ) ;
  assign n23924 = ( x71 & ~n23878 ) | ( x71 & n23923 ) | ( ~n23878 & n23923 ) ;
  assign n23925 = ( x72 & ~n23870 ) | ( x72 & n23924 ) | ( ~n23870 & n23924 ) ;
  assign n23926 = ( x73 & ~n23862 ) | ( x73 & n23925 ) | ( ~n23862 & n23925 ) ;
  assign n23927 = ( x74 & ~n23854 ) | ( x74 & n23926 ) | ( ~n23854 & n23926 ) ;
  assign n23928 = ( x75 & ~n23846 ) | ( x75 & n23927 ) | ( ~n23846 & n23927 ) ;
  assign n23929 = ( x76 & ~n23838 ) | ( x76 & n23928 ) | ( ~n23838 & n23928 ) ;
  assign n23930 = ( x77 & ~n23830 ) | ( x77 & n23929 ) | ( ~n23830 & n23929 ) ;
  assign n23931 = ( x78 & ~n23822 ) | ( x78 & n23930 ) | ( ~n23822 & n23930 ) ;
  assign n23932 = ( x79 & ~n23814 ) | ( x79 & n23931 ) | ( ~n23814 & n23931 ) ;
  assign n23933 = ( x80 & ~n23806 ) | ( x80 & n23932 ) | ( ~n23806 & n23932 ) ;
  assign n23934 = ( x81 & ~n23798 ) | ( x81 & n23933 ) | ( ~n23798 & n23933 ) ;
  assign n23935 = ( x82 & ~n23790 ) | ( x82 & n23934 ) | ( ~n23790 & n23934 ) ;
  assign n23936 = ( x83 & ~n23782 ) | ( x83 & n23935 ) | ( ~n23782 & n23935 ) ;
  assign n23937 = ( x84 & ~n23774 ) | ( x84 & n23936 ) | ( ~n23774 & n23936 ) ;
  assign n23938 = ( x85 & ~n23766 ) | ( x85 & n23937 ) | ( ~n23766 & n23937 ) ;
  assign n23939 = ( x86 & ~n23758 ) | ( x86 & n23938 ) | ( ~n23758 & n23938 ) ;
  assign n23940 = ( x87 & ~n23750 ) | ( x87 & n23939 ) | ( ~n23750 & n23939 ) ;
  assign n23941 = ( x88 & ~n23742 ) | ( x88 & n23940 ) | ( ~n23742 & n23940 ) ;
  assign n23942 = ( x89 & ~n23734 ) | ( x89 & n23941 ) | ( ~n23734 & n23941 ) ;
  assign n23943 = ( x90 & ~n23726 ) | ( x90 & n23942 ) | ( ~n23726 & n23942 ) ;
  assign n23944 = ( x91 & ~n23718 ) | ( x91 & n23943 ) | ( ~n23718 & n23943 ) ;
  assign n23945 = ( x92 & ~n23710 ) | ( x92 & n23944 ) | ( ~n23710 & n23944 ) ;
  assign n23946 = ( x93 & ~n23702 ) | ( x93 & n23945 ) | ( ~n23702 & n23945 ) ;
  assign n23947 = ( x94 & ~n23694 ) | ( x94 & n23946 ) | ( ~n23694 & n23946 ) ;
  assign n23948 = ( x95 & ~n23686 ) | ( x95 & n23947 ) | ( ~n23686 & n23947 ) ;
  assign n23949 = ( x96 & ~n23678 ) | ( x96 & n23948 ) | ( ~n23678 & n23948 ) ;
  assign n23956 = ( x97 & ~n5541 ) | ( x97 & n23949 ) | ( ~n5541 & n23949 ) ;
  assign n23955 = x97 &  n23949 ;
  assign n23957 = ( n23670 & ~n23956 ) | ( n23670 & n23955 ) | ( ~n23956 & n23955 ) ;
  assign n23950 = ( x97 & ~n23670 ) | ( x97 & n23949 ) | ( ~n23670 & n23949 ) ;
  assign n23951 = n5541 | n23950 ;
  assign n23958 = n23678 &  n23951 ;
  assign n23952 = x96 | n23678 ;
  assign n23953 = x96 &  n23678 ;
  assign n23954 = ( n23952 & ~n23953 ) | ( n23952 & 1'b0 ) | ( ~n23953 & 1'b0 ) ;
  assign n23962 = ( n5541 & n23948 ) | ( n5541 & n23954 ) | ( n23948 & n23954 ) ;
  assign n23963 = ( n23948 & ~n23950 ) | ( n23948 & n23954 ) | ( ~n23950 & n23954 ) ;
  assign n23964 = ~n23962 & n23963 ;
  assign n23965 = n23958 | n23964 ;
  assign n23966 = n23686 &  n23951 ;
  assign n23959 = x95 | n23686 ;
  assign n23960 = x95 &  n23686 ;
  assign n23961 = ( n23959 & ~n23960 ) | ( n23959 & 1'b0 ) | ( ~n23960 & 1'b0 ) ;
  assign n23970 = ( n5541 & n23947 ) | ( n5541 & n23961 ) | ( n23947 & n23961 ) ;
  assign n23971 = ( n23947 & ~n23950 ) | ( n23947 & n23961 ) | ( ~n23950 & n23961 ) ;
  assign n23972 = ~n23970 & n23971 ;
  assign n23973 = n23966 | n23972 ;
  assign n23974 = n23694 &  n23951 ;
  assign n23967 = x94 | n23694 ;
  assign n23968 = x94 &  n23694 ;
  assign n23969 = ( n23967 & ~n23968 ) | ( n23967 & 1'b0 ) | ( ~n23968 & 1'b0 ) ;
  assign n23978 = ( n5541 & n23946 ) | ( n5541 & n23969 ) | ( n23946 & n23969 ) ;
  assign n23979 = ( n23946 & ~n23950 ) | ( n23946 & n23969 ) | ( ~n23950 & n23969 ) ;
  assign n23980 = ~n23978 & n23979 ;
  assign n23981 = n23974 | n23980 ;
  assign n23982 = n23702 &  n23951 ;
  assign n23975 = x93 | n23702 ;
  assign n23976 = x93 &  n23702 ;
  assign n23977 = ( n23975 & ~n23976 ) | ( n23975 & 1'b0 ) | ( ~n23976 & 1'b0 ) ;
  assign n23986 = ( n5541 & n23945 ) | ( n5541 & n23977 ) | ( n23945 & n23977 ) ;
  assign n23987 = ( n23945 & ~n23950 ) | ( n23945 & n23977 ) | ( ~n23950 & n23977 ) ;
  assign n23988 = ~n23986 & n23987 ;
  assign n23989 = n23982 | n23988 ;
  assign n23990 = n23710 &  n23951 ;
  assign n23983 = x92 | n23710 ;
  assign n23984 = x92 &  n23710 ;
  assign n23985 = ( n23983 & ~n23984 ) | ( n23983 & 1'b0 ) | ( ~n23984 & 1'b0 ) ;
  assign n23994 = ( n5541 & n23944 ) | ( n5541 & n23985 ) | ( n23944 & n23985 ) ;
  assign n23995 = ( n23944 & ~n23950 ) | ( n23944 & n23985 ) | ( ~n23950 & n23985 ) ;
  assign n23996 = ~n23994 & n23995 ;
  assign n23997 = n23990 | n23996 ;
  assign n23998 = n23718 &  n23951 ;
  assign n23991 = x91 | n23718 ;
  assign n23992 = x91 &  n23718 ;
  assign n23993 = ( n23991 & ~n23992 ) | ( n23991 & 1'b0 ) | ( ~n23992 & 1'b0 ) ;
  assign n24002 = ( n5541 & n23943 ) | ( n5541 & n23993 ) | ( n23943 & n23993 ) ;
  assign n24003 = ( n23943 & ~n23950 ) | ( n23943 & n23993 ) | ( ~n23950 & n23993 ) ;
  assign n24004 = ~n24002 & n24003 ;
  assign n24005 = n23998 | n24004 ;
  assign n24006 = n23726 &  n23951 ;
  assign n23999 = x90 | n23726 ;
  assign n24000 = x90 &  n23726 ;
  assign n24001 = ( n23999 & ~n24000 ) | ( n23999 & 1'b0 ) | ( ~n24000 & 1'b0 ) ;
  assign n24010 = ( n5541 & n23942 ) | ( n5541 & n24001 ) | ( n23942 & n24001 ) ;
  assign n24011 = ( n23942 & ~n23950 ) | ( n23942 & n24001 ) | ( ~n23950 & n24001 ) ;
  assign n24012 = ~n24010 & n24011 ;
  assign n24013 = n24006 | n24012 ;
  assign n24014 = n23734 &  n23951 ;
  assign n24007 = x89 | n23734 ;
  assign n24008 = x89 &  n23734 ;
  assign n24009 = ( n24007 & ~n24008 ) | ( n24007 & 1'b0 ) | ( ~n24008 & 1'b0 ) ;
  assign n24018 = ( n5541 & n23941 ) | ( n5541 & n24009 ) | ( n23941 & n24009 ) ;
  assign n24019 = ( n23941 & ~n23950 ) | ( n23941 & n24009 ) | ( ~n23950 & n24009 ) ;
  assign n24020 = ~n24018 & n24019 ;
  assign n24021 = n24014 | n24020 ;
  assign n24022 = n23742 &  n23951 ;
  assign n24015 = x88 | n23742 ;
  assign n24016 = x88 &  n23742 ;
  assign n24017 = ( n24015 & ~n24016 ) | ( n24015 & 1'b0 ) | ( ~n24016 & 1'b0 ) ;
  assign n24026 = ( n5541 & n23940 ) | ( n5541 & n24017 ) | ( n23940 & n24017 ) ;
  assign n24027 = ( n23940 & ~n23950 ) | ( n23940 & n24017 ) | ( ~n23950 & n24017 ) ;
  assign n24028 = ~n24026 & n24027 ;
  assign n24029 = n24022 | n24028 ;
  assign n24030 = n23750 &  n23951 ;
  assign n24023 = x87 | n23750 ;
  assign n24024 = x87 &  n23750 ;
  assign n24025 = ( n24023 & ~n24024 ) | ( n24023 & 1'b0 ) | ( ~n24024 & 1'b0 ) ;
  assign n24034 = ( n5541 & n23939 ) | ( n5541 & n24025 ) | ( n23939 & n24025 ) ;
  assign n24035 = ( n23939 & ~n23950 ) | ( n23939 & n24025 ) | ( ~n23950 & n24025 ) ;
  assign n24036 = ~n24034 & n24035 ;
  assign n24037 = n24030 | n24036 ;
  assign n24038 = n23758 &  n23951 ;
  assign n24031 = x86 | n23758 ;
  assign n24032 = x86 &  n23758 ;
  assign n24033 = ( n24031 & ~n24032 ) | ( n24031 & 1'b0 ) | ( ~n24032 & 1'b0 ) ;
  assign n24042 = ( n5541 & n23938 ) | ( n5541 & n24033 ) | ( n23938 & n24033 ) ;
  assign n24043 = ( n23938 & ~n23950 ) | ( n23938 & n24033 ) | ( ~n23950 & n24033 ) ;
  assign n24044 = ~n24042 & n24043 ;
  assign n24045 = n24038 | n24044 ;
  assign n24046 = n23766 &  n23951 ;
  assign n24039 = x85 | n23766 ;
  assign n24040 = x85 &  n23766 ;
  assign n24041 = ( n24039 & ~n24040 ) | ( n24039 & 1'b0 ) | ( ~n24040 & 1'b0 ) ;
  assign n24050 = ( n5541 & n23937 ) | ( n5541 & n24041 ) | ( n23937 & n24041 ) ;
  assign n24051 = ( n23937 & ~n23950 ) | ( n23937 & n24041 ) | ( ~n23950 & n24041 ) ;
  assign n24052 = ~n24050 & n24051 ;
  assign n24053 = n24046 | n24052 ;
  assign n24054 = n23774 &  n23951 ;
  assign n24047 = x84 | n23774 ;
  assign n24048 = x84 &  n23774 ;
  assign n24049 = ( n24047 & ~n24048 ) | ( n24047 & 1'b0 ) | ( ~n24048 & 1'b0 ) ;
  assign n24058 = ( n5541 & n23936 ) | ( n5541 & n24049 ) | ( n23936 & n24049 ) ;
  assign n24059 = ( n23936 & ~n23950 ) | ( n23936 & n24049 ) | ( ~n23950 & n24049 ) ;
  assign n24060 = ~n24058 & n24059 ;
  assign n24061 = n24054 | n24060 ;
  assign n24062 = n23782 &  n23951 ;
  assign n24055 = x83 | n23782 ;
  assign n24056 = x83 &  n23782 ;
  assign n24057 = ( n24055 & ~n24056 ) | ( n24055 & 1'b0 ) | ( ~n24056 & 1'b0 ) ;
  assign n24066 = ( n5541 & n23935 ) | ( n5541 & n24057 ) | ( n23935 & n24057 ) ;
  assign n24067 = ( n23935 & ~n23950 ) | ( n23935 & n24057 ) | ( ~n23950 & n24057 ) ;
  assign n24068 = ~n24066 & n24067 ;
  assign n24069 = n24062 | n24068 ;
  assign n24070 = n23790 &  n23951 ;
  assign n24063 = x82 | n23790 ;
  assign n24064 = x82 &  n23790 ;
  assign n24065 = ( n24063 & ~n24064 ) | ( n24063 & 1'b0 ) | ( ~n24064 & 1'b0 ) ;
  assign n24074 = ( n5541 & n23934 ) | ( n5541 & n24065 ) | ( n23934 & n24065 ) ;
  assign n24075 = ( n23934 & ~n23950 ) | ( n23934 & n24065 ) | ( ~n23950 & n24065 ) ;
  assign n24076 = ~n24074 & n24075 ;
  assign n24077 = n24070 | n24076 ;
  assign n24078 = n23798 &  n23951 ;
  assign n24071 = x81 | n23798 ;
  assign n24072 = x81 &  n23798 ;
  assign n24073 = ( n24071 & ~n24072 ) | ( n24071 & 1'b0 ) | ( ~n24072 & 1'b0 ) ;
  assign n24082 = ( n5541 & n23933 ) | ( n5541 & n24073 ) | ( n23933 & n24073 ) ;
  assign n24083 = ( n23933 & ~n23950 ) | ( n23933 & n24073 ) | ( ~n23950 & n24073 ) ;
  assign n24084 = ~n24082 & n24083 ;
  assign n24085 = n24078 | n24084 ;
  assign n24086 = n23806 &  n23951 ;
  assign n24079 = x80 | n23806 ;
  assign n24080 = x80 &  n23806 ;
  assign n24081 = ( n24079 & ~n24080 ) | ( n24079 & 1'b0 ) | ( ~n24080 & 1'b0 ) ;
  assign n24090 = ( n5541 & n23932 ) | ( n5541 & n24081 ) | ( n23932 & n24081 ) ;
  assign n24091 = ( n23932 & ~n23950 ) | ( n23932 & n24081 ) | ( ~n23950 & n24081 ) ;
  assign n24092 = ~n24090 & n24091 ;
  assign n24093 = n24086 | n24092 ;
  assign n24094 = n23814 &  n23951 ;
  assign n24087 = x79 | n23814 ;
  assign n24088 = x79 &  n23814 ;
  assign n24089 = ( n24087 & ~n24088 ) | ( n24087 & 1'b0 ) | ( ~n24088 & 1'b0 ) ;
  assign n24098 = ( n5541 & n23931 ) | ( n5541 & n24089 ) | ( n23931 & n24089 ) ;
  assign n24099 = ( n23931 & ~n23950 ) | ( n23931 & n24089 ) | ( ~n23950 & n24089 ) ;
  assign n24100 = ~n24098 & n24099 ;
  assign n24101 = n24094 | n24100 ;
  assign n24102 = n23822 &  n23951 ;
  assign n24095 = x78 | n23822 ;
  assign n24096 = x78 &  n23822 ;
  assign n24097 = ( n24095 & ~n24096 ) | ( n24095 & 1'b0 ) | ( ~n24096 & 1'b0 ) ;
  assign n24106 = ( n5541 & n23930 ) | ( n5541 & n24097 ) | ( n23930 & n24097 ) ;
  assign n24107 = ( n23930 & ~n23950 ) | ( n23930 & n24097 ) | ( ~n23950 & n24097 ) ;
  assign n24108 = ~n24106 & n24107 ;
  assign n24109 = n24102 | n24108 ;
  assign n24110 = n23830 &  n23951 ;
  assign n24103 = x77 | n23830 ;
  assign n24104 = x77 &  n23830 ;
  assign n24105 = ( n24103 & ~n24104 ) | ( n24103 & 1'b0 ) | ( ~n24104 & 1'b0 ) ;
  assign n24114 = ( n5541 & n23929 ) | ( n5541 & n24105 ) | ( n23929 & n24105 ) ;
  assign n24115 = ( n23929 & ~n23950 ) | ( n23929 & n24105 ) | ( ~n23950 & n24105 ) ;
  assign n24116 = ~n24114 & n24115 ;
  assign n24117 = n24110 | n24116 ;
  assign n24118 = n23838 &  n23951 ;
  assign n24111 = x76 | n23838 ;
  assign n24112 = x76 &  n23838 ;
  assign n24113 = ( n24111 & ~n24112 ) | ( n24111 & 1'b0 ) | ( ~n24112 & 1'b0 ) ;
  assign n24122 = ( n5541 & n23928 ) | ( n5541 & n24113 ) | ( n23928 & n24113 ) ;
  assign n24123 = ( n23928 & ~n23950 ) | ( n23928 & n24113 ) | ( ~n23950 & n24113 ) ;
  assign n24124 = ~n24122 & n24123 ;
  assign n24125 = n24118 | n24124 ;
  assign n24126 = n23846 &  n23951 ;
  assign n24119 = x75 | n23846 ;
  assign n24120 = x75 &  n23846 ;
  assign n24121 = ( n24119 & ~n24120 ) | ( n24119 & 1'b0 ) | ( ~n24120 & 1'b0 ) ;
  assign n24130 = ( n5541 & n23927 ) | ( n5541 & n24121 ) | ( n23927 & n24121 ) ;
  assign n24131 = ( n23927 & ~n23950 ) | ( n23927 & n24121 ) | ( ~n23950 & n24121 ) ;
  assign n24132 = ~n24130 & n24131 ;
  assign n24133 = n24126 | n24132 ;
  assign n24134 = n23854 &  n23951 ;
  assign n24127 = x74 | n23854 ;
  assign n24128 = x74 &  n23854 ;
  assign n24129 = ( n24127 & ~n24128 ) | ( n24127 & 1'b0 ) | ( ~n24128 & 1'b0 ) ;
  assign n24138 = ( n5541 & n23926 ) | ( n5541 & n24129 ) | ( n23926 & n24129 ) ;
  assign n24139 = ( n23926 & ~n23950 ) | ( n23926 & n24129 ) | ( ~n23950 & n24129 ) ;
  assign n24140 = ~n24138 & n24139 ;
  assign n24141 = n24134 | n24140 ;
  assign n24142 = n23862 &  n23951 ;
  assign n24135 = x73 | n23862 ;
  assign n24136 = x73 &  n23862 ;
  assign n24137 = ( n24135 & ~n24136 ) | ( n24135 & 1'b0 ) | ( ~n24136 & 1'b0 ) ;
  assign n24146 = ( n5541 & n23925 ) | ( n5541 & n24137 ) | ( n23925 & n24137 ) ;
  assign n24147 = ( n23925 & ~n23950 ) | ( n23925 & n24137 ) | ( ~n23950 & n24137 ) ;
  assign n24148 = ~n24146 & n24147 ;
  assign n24149 = n24142 | n24148 ;
  assign n24150 = n23870 &  n23951 ;
  assign n24143 = x72 | n23870 ;
  assign n24144 = x72 &  n23870 ;
  assign n24145 = ( n24143 & ~n24144 ) | ( n24143 & 1'b0 ) | ( ~n24144 & 1'b0 ) ;
  assign n24154 = ( n5541 & n23924 ) | ( n5541 & n24145 ) | ( n23924 & n24145 ) ;
  assign n24155 = ( n23924 & ~n23950 ) | ( n23924 & n24145 ) | ( ~n23950 & n24145 ) ;
  assign n24156 = ~n24154 & n24155 ;
  assign n24157 = n24150 | n24156 ;
  assign n24158 = n23878 &  n23951 ;
  assign n24151 = x71 | n23878 ;
  assign n24152 = x71 &  n23878 ;
  assign n24153 = ( n24151 & ~n24152 ) | ( n24151 & 1'b0 ) | ( ~n24152 & 1'b0 ) ;
  assign n24162 = ( n5541 & n23923 ) | ( n5541 & n24153 ) | ( n23923 & n24153 ) ;
  assign n24163 = ( n23923 & ~n23950 ) | ( n23923 & n24153 ) | ( ~n23950 & n24153 ) ;
  assign n24164 = ~n24162 & n24163 ;
  assign n24165 = n24158 | n24164 ;
  assign n24166 = n23886 &  n23951 ;
  assign n24159 = x70 | n23886 ;
  assign n24160 = x70 &  n23886 ;
  assign n24161 = ( n24159 & ~n24160 ) | ( n24159 & 1'b0 ) | ( ~n24160 & 1'b0 ) ;
  assign n24170 = ( n5541 & n23922 ) | ( n5541 & n24161 ) | ( n23922 & n24161 ) ;
  assign n24171 = ( n23922 & ~n23950 ) | ( n23922 & n24161 ) | ( ~n23950 & n24161 ) ;
  assign n24172 = ~n24170 & n24171 ;
  assign n24173 = n24166 | n24172 ;
  assign n24174 = n23894 &  n23951 ;
  assign n24167 = x69 | n23894 ;
  assign n24168 = x69 &  n23894 ;
  assign n24169 = ( n24167 & ~n24168 ) | ( n24167 & 1'b0 ) | ( ~n24168 & 1'b0 ) ;
  assign n24178 = ( n5541 & n23921 ) | ( n5541 & n24169 ) | ( n23921 & n24169 ) ;
  assign n24179 = ( n23921 & ~n23950 ) | ( n23921 & n24169 ) | ( ~n23950 & n24169 ) ;
  assign n24180 = ~n24178 & n24179 ;
  assign n24181 = n24174 | n24180 ;
  assign n24182 = n23902 &  n23951 ;
  assign n24175 = x68 | n23902 ;
  assign n24176 = x68 &  n23902 ;
  assign n24177 = ( n24175 & ~n24176 ) | ( n24175 & 1'b0 ) | ( ~n24176 & 1'b0 ) ;
  assign n24186 = ( n5541 & n23920 ) | ( n5541 & n24177 ) | ( n23920 & n24177 ) ;
  assign n24187 = ( n23920 & ~n23950 ) | ( n23920 & n24177 ) | ( ~n23950 & n24177 ) ;
  assign n24188 = ~n24186 & n24187 ;
  assign n24189 = n24182 | n24188 ;
  assign n24190 = n23907 &  n23951 ;
  assign n24183 = x67 | n23907 ;
  assign n24184 = x67 &  n23907 ;
  assign n24185 = ( n24183 & ~n24184 ) | ( n24183 & 1'b0 ) | ( ~n24184 & 1'b0 ) ;
  assign n24194 = ( n5541 & n23919 ) | ( n5541 & n24185 ) | ( n23919 & n24185 ) ;
  assign n24195 = ( n23919 & ~n23950 ) | ( n23919 & n24185 ) | ( ~n23950 & n24185 ) ;
  assign n24196 = ~n24194 & n24195 ;
  assign n24197 = n24190 | n24196 ;
  assign n24198 = n23913 &  n23951 ;
  assign n24191 = x66 | n23913 ;
  assign n24192 = x66 &  n23913 ;
  assign n24193 = ( n24191 & ~n24192 ) | ( n24191 & 1'b0 ) | ( ~n24192 & 1'b0 ) ;
  assign n24199 = ( n5541 & n23918 ) | ( n5541 & n24193 ) | ( n23918 & n24193 ) ;
  assign n24200 = ( n23918 & ~n23950 ) | ( n23918 & n24193 ) | ( ~n23950 & n24193 ) ;
  assign n24201 = ~n24199 & n24200 ;
  assign n24202 = n24198 | n24201 ;
  assign n24203 = n23917 &  n23951 ;
  assign n24204 = ( x65 & ~x31 ) | ( x65 & n23914 ) | ( ~x31 & n23914 ) ;
  assign n24205 = ( x31 & ~n23914 ) | ( x31 & x65 ) | ( ~n23914 & x65 ) ;
  assign n24206 = ( n24204 & ~x65 ) | ( n24204 & n24205 ) | ( ~x65 & n24205 ) ;
  assign n24207 = ( n5505 & ~n5541 ) | ( n5505 & n24206 ) | ( ~n5541 & n24206 ) ;
  assign n24208 = ( n5505 & n23950 ) | ( n5505 & n24206 ) | ( n23950 & n24206 ) ;
  assign n24209 = ( n24207 & ~n24208 ) | ( n24207 & 1'b0 ) | ( ~n24208 & 1'b0 ) ;
  assign n24210 = n24203 | n24209 ;
  assign n24211 = ( n5808 & ~n23950 ) | ( n5808 & 1'b0 ) | ( ~n23950 & 1'b0 ) ;
  assign n24212 = ( x30 & ~n24211 ) | ( x30 & 1'b0 ) | ( ~n24211 & 1'b0 ) ;
  assign n24213 = ( n5814 & ~n23950 ) | ( n5814 & 1'b0 ) | ( ~n23950 & 1'b0 ) ;
  assign n24214 = n24212 | n24213 ;
  assign n24215 = ( x65 & ~n24214 ) | ( x65 & n5817 ) | ( ~n24214 & n5817 ) ;
  assign n24216 = ( x66 & ~n24210 ) | ( x66 & n24215 ) | ( ~n24210 & n24215 ) ;
  assign n24217 = ( x67 & ~n24202 ) | ( x67 & n24216 ) | ( ~n24202 & n24216 ) ;
  assign n24218 = ( x68 & ~n24197 ) | ( x68 & n24217 ) | ( ~n24197 & n24217 ) ;
  assign n24219 = ( x69 & ~n24189 ) | ( x69 & n24218 ) | ( ~n24189 & n24218 ) ;
  assign n24220 = ( x70 & ~n24181 ) | ( x70 & n24219 ) | ( ~n24181 & n24219 ) ;
  assign n24221 = ( x71 & ~n24173 ) | ( x71 & n24220 ) | ( ~n24173 & n24220 ) ;
  assign n24222 = ( x72 & ~n24165 ) | ( x72 & n24221 ) | ( ~n24165 & n24221 ) ;
  assign n24223 = ( x73 & ~n24157 ) | ( x73 & n24222 ) | ( ~n24157 & n24222 ) ;
  assign n24224 = ( x74 & ~n24149 ) | ( x74 & n24223 ) | ( ~n24149 & n24223 ) ;
  assign n24225 = ( x75 & ~n24141 ) | ( x75 & n24224 ) | ( ~n24141 & n24224 ) ;
  assign n24226 = ( x76 & ~n24133 ) | ( x76 & n24225 ) | ( ~n24133 & n24225 ) ;
  assign n24227 = ( x77 & ~n24125 ) | ( x77 & n24226 ) | ( ~n24125 & n24226 ) ;
  assign n24228 = ( x78 & ~n24117 ) | ( x78 & n24227 ) | ( ~n24117 & n24227 ) ;
  assign n24229 = ( x79 & ~n24109 ) | ( x79 & n24228 ) | ( ~n24109 & n24228 ) ;
  assign n24230 = ( x80 & ~n24101 ) | ( x80 & n24229 ) | ( ~n24101 & n24229 ) ;
  assign n24231 = ( x81 & ~n24093 ) | ( x81 & n24230 ) | ( ~n24093 & n24230 ) ;
  assign n24232 = ( x82 & ~n24085 ) | ( x82 & n24231 ) | ( ~n24085 & n24231 ) ;
  assign n24233 = ( x83 & ~n24077 ) | ( x83 & n24232 ) | ( ~n24077 & n24232 ) ;
  assign n24234 = ( x84 & ~n24069 ) | ( x84 & n24233 ) | ( ~n24069 & n24233 ) ;
  assign n24235 = ( x85 & ~n24061 ) | ( x85 & n24234 ) | ( ~n24061 & n24234 ) ;
  assign n24236 = ( x86 & ~n24053 ) | ( x86 & n24235 ) | ( ~n24053 & n24235 ) ;
  assign n24237 = ( x87 & ~n24045 ) | ( x87 & n24236 ) | ( ~n24045 & n24236 ) ;
  assign n24238 = ( x88 & ~n24037 ) | ( x88 & n24237 ) | ( ~n24037 & n24237 ) ;
  assign n24239 = ( x89 & ~n24029 ) | ( x89 & n24238 ) | ( ~n24029 & n24238 ) ;
  assign n24240 = ( x90 & ~n24021 ) | ( x90 & n24239 ) | ( ~n24021 & n24239 ) ;
  assign n24241 = ( x91 & ~n24013 ) | ( x91 & n24240 ) | ( ~n24013 & n24240 ) ;
  assign n24242 = ( x92 & ~n24005 ) | ( x92 & n24241 ) | ( ~n24005 & n24241 ) ;
  assign n24243 = ( x93 & ~n23997 ) | ( x93 & n24242 ) | ( ~n23997 & n24242 ) ;
  assign n24244 = ( x94 & ~n23989 ) | ( x94 & n24243 ) | ( ~n23989 & n24243 ) ;
  assign n24245 = ( x95 & ~n23981 ) | ( x95 & n24244 ) | ( ~n23981 & n24244 ) ;
  assign n24246 = ( x96 & ~n23973 ) | ( x96 & n24245 ) | ( ~n23973 & n24245 ) ;
  assign n24247 = ( x97 & ~n23965 ) | ( x97 & n24246 ) | ( ~n23965 & n24246 ) ;
  assign n24248 = ( x98 & ~n23957 ) | ( x98 & n24247 ) | ( ~n23957 & n24247 ) ;
  assign n24249 = n5854 | n24248 ;
  assign n24250 = n23957 &  n24249 ;
  assign n24254 = ( n5854 & n23957 ) | ( n5854 & n24247 ) | ( n23957 & n24247 ) ;
  assign n24255 = ( x98 & ~n24254 ) | ( x98 & n23957 ) | ( ~n24254 & n23957 ) ;
  assign n24256 = ~x98 & n24255 ;
  assign n24257 = n24250 | n24256 ;
  assign n24258 = ~x99 & n24257 ;
  assign n24259 = n23965 &  n24249 ;
  assign n24251 = x97 | n23965 ;
  assign n24252 = x97 &  n23965 ;
  assign n24253 = ( n24251 & ~n24252 ) | ( n24251 & 1'b0 ) | ( ~n24252 & 1'b0 ) ;
  assign n24263 = ( n5854 & n24246 ) | ( n5854 & n24253 ) | ( n24246 & n24253 ) ;
  assign n24264 = ( n24246 & ~n24248 ) | ( n24246 & n24253 ) | ( ~n24248 & n24253 ) ;
  assign n24265 = ~n24263 & n24264 ;
  assign n24266 = n24259 | n24265 ;
  assign n24267 = n23973 &  n24249 ;
  assign n24260 = x96 | n23973 ;
  assign n24261 = x96 &  n23973 ;
  assign n24262 = ( n24260 & ~n24261 ) | ( n24260 & 1'b0 ) | ( ~n24261 & 1'b0 ) ;
  assign n24271 = ( n5854 & n24245 ) | ( n5854 & n24262 ) | ( n24245 & n24262 ) ;
  assign n24272 = ( n24245 & ~n24248 ) | ( n24245 & n24262 ) | ( ~n24248 & n24262 ) ;
  assign n24273 = ~n24271 & n24272 ;
  assign n24274 = n24267 | n24273 ;
  assign n24275 = n23981 &  n24249 ;
  assign n24268 = x95 | n23981 ;
  assign n24269 = x95 &  n23981 ;
  assign n24270 = ( n24268 & ~n24269 ) | ( n24268 & 1'b0 ) | ( ~n24269 & 1'b0 ) ;
  assign n24279 = ( n5854 & n24244 ) | ( n5854 & n24270 ) | ( n24244 & n24270 ) ;
  assign n24280 = ( n24244 & ~n24248 ) | ( n24244 & n24270 ) | ( ~n24248 & n24270 ) ;
  assign n24281 = ~n24279 & n24280 ;
  assign n24282 = n24275 | n24281 ;
  assign n24283 = n23989 &  n24249 ;
  assign n24276 = x94 | n23989 ;
  assign n24277 = x94 &  n23989 ;
  assign n24278 = ( n24276 & ~n24277 ) | ( n24276 & 1'b0 ) | ( ~n24277 & 1'b0 ) ;
  assign n24287 = ( n5854 & n24243 ) | ( n5854 & n24278 ) | ( n24243 & n24278 ) ;
  assign n24288 = ( n24243 & ~n24248 ) | ( n24243 & n24278 ) | ( ~n24248 & n24278 ) ;
  assign n24289 = ~n24287 & n24288 ;
  assign n24290 = n24283 | n24289 ;
  assign n24291 = n23997 &  n24249 ;
  assign n24284 = x93 | n23997 ;
  assign n24285 = x93 &  n23997 ;
  assign n24286 = ( n24284 & ~n24285 ) | ( n24284 & 1'b0 ) | ( ~n24285 & 1'b0 ) ;
  assign n24295 = ( n5854 & n24242 ) | ( n5854 & n24286 ) | ( n24242 & n24286 ) ;
  assign n24296 = ( n24242 & ~n24248 ) | ( n24242 & n24286 ) | ( ~n24248 & n24286 ) ;
  assign n24297 = ~n24295 & n24296 ;
  assign n24298 = n24291 | n24297 ;
  assign n24299 = n24005 &  n24249 ;
  assign n24292 = x92 | n24005 ;
  assign n24293 = x92 &  n24005 ;
  assign n24294 = ( n24292 & ~n24293 ) | ( n24292 & 1'b0 ) | ( ~n24293 & 1'b0 ) ;
  assign n24303 = ( n5854 & n24241 ) | ( n5854 & n24294 ) | ( n24241 & n24294 ) ;
  assign n24304 = ( n24241 & ~n24248 ) | ( n24241 & n24294 ) | ( ~n24248 & n24294 ) ;
  assign n24305 = ~n24303 & n24304 ;
  assign n24306 = n24299 | n24305 ;
  assign n24307 = n24013 &  n24249 ;
  assign n24300 = x91 | n24013 ;
  assign n24301 = x91 &  n24013 ;
  assign n24302 = ( n24300 & ~n24301 ) | ( n24300 & 1'b0 ) | ( ~n24301 & 1'b0 ) ;
  assign n24311 = ( n5854 & n24240 ) | ( n5854 & n24302 ) | ( n24240 & n24302 ) ;
  assign n24312 = ( n24240 & ~n24248 ) | ( n24240 & n24302 ) | ( ~n24248 & n24302 ) ;
  assign n24313 = ~n24311 & n24312 ;
  assign n24314 = n24307 | n24313 ;
  assign n24315 = n24021 &  n24249 ;
  assign n24308 = x90 | n24021 ;
  assign n24309 = x90 &  n24021 ;
  assign n24310 = ( n24308 & ~n24309 ) | ( n24308 & 1'b0 ) | ( ~n24309 & 1'b0 ) ;
  assign n24319 = ( n5854 & n24239 ) | ( n5854 & n24310 ) | ( n24239 & n24310 ) ;
  assign n24320 = ( n24239 & ~n24248 ) | ( n24239 & n24310 ) | ( ~n24248 & n24310 ) ;
  assign n24321 = ~n24319 & n24320 ;
  assign n24322 = n24315 | n24321 ;
  assign n24323 = n24029 &  n24249 ;
  assign n24316 = x89 | n24029 ;
  assign n24317 = x89 &  n24029 ;
  assign n24318 = ( n24316 & ~n24317 ) | ( n24316 & 1'b0 ) | ( ~n24317 & 1'b0 ) ;
  assign n24327 = ( n5854 & n24238 ) | ( n5854 & n24318 ) | ( n24238 & n24318 ) ;
  assign n24328 = ( n24238 & ~n24248 ) | ( n24238 & n24318 ) | ( ~n24248 & n24318 ) ;
  assign n24329 = ~n24327 & n24328 ;
  assign n24330 = n24323 | n24329 ;
  assign n24331 = n24037 &  n24249 ;
  assign n24324 = x88 | n24037 ;
  assign n24325 = x88 &  n24037 ;
  assign n24326 = ( n24324 & ~n24325 ) | ( n24324 & 1'b0 ) | ( ~n24325 & 1'b0 ) ;
  assign n24335 = ( n5854 & n24237 ) | ( n5854 & n24326 ) | ( n24237 & n24326 ) ;
  assign n24336 = ( n24237 & ~n24248 ) | ( n24237 & n24326 ) | ( ~n24248 & n24326 ) ;
  assign n24337 = ~n24335 & n24336 ;
  assign n24338 = n24331 | n24337 ;
  assign n24339 = n24045 &  n24249 ;
  assign n24332 = x87 | n24045 ;
  assign n24333 = x87 &  n24045 ;
  assign n24334 = ( n24332 & ~n24333 ) | ( n24332 & 1'b0 ) | ( ~n24333 & 1'b0 ) ;
  assign n24343 = ( n5854 & n24236 ) | ( n5854 & n24334 ) | ( n24236 & n24334 ) ;
  assign n24344 = ( n24236 & ~n24248 ) | ( n24236 & n24334 ) | ( ~n24248 & n24334 ) ;
  assign n24345 = ~n24343 & n24344 ;
  assign n24346 = n24339 | n24345 ;
  assign n24347 = n24053 &  n24249 ;
  assign n24340 = x86 | n24053 ;
  assign n24341 = x86 &  n24053 ;
  assign n24342 = ( n24340 & ~n24341 ) | ( n24340 & 1'b0 ) | ( ~n24341 & 1'b0 ) ;
  assign n24351 = ( n5854 & n24235 ) | ( n5854 & n24342 ) | ( n24235 & n24342 ) ;
  assign n24352 = ( n24235 & ~n24248 ) | ( n24235 & n24342 ) | ( ~n24248 & n24342 ) ;
  assign n24353 = ~n24351 & n24352 ;
  assign n24354 = n24347 | n24353 ;
  assign n24355 = n24061 &  n24249 ;
  assign n24348 = x85 | n24061 ;
  assign n24349 = x85 &  n24061 ;
  assign n24350 = ( n24348 & ~n24349 ) | ( n24348 & 1'b0 ) | ( ~n24349 & 1'b0 ) ;
  assign n24359 = ( n5854 & n24234 ) | ( n5854 & n24350 ) | ( n24234 & n24350 ) ;
  assign n24360 = ( n24234 & ~n24248 ) | ( n24234 & n24350 ) | ( ~n24248 & n24350 ) ;
  assign n24361 = ~n24359 & n24360 ;
  assign n24362 = n24355 | n24361 ;
  assign n24363 = n24069 &  n24249 ;
  assign n24356 = x84 | n24069 ;
  assign n24357 = x84 &  n24069 ;
  assign n24358 = ( n24356 & ~n24357 ) | ( n24356 & 1'b0 ) | ( ~n24357 & 1'b0 ) ;
  assign n24367 = ( n5854 & n24233 ) | ( n5854 & n24358 ) | ( n24233 & n24358 ) ;
  assign n24368 = ( n24233 & ~n24248 ) | ( n24233 & n24358 ) | ( ~n24248 & n24358 ) ;
  assign n24369 = ~n24367 & n24368 ;
  assign n24370 = n24363 | n24369 ;
  assign n24371 = n24077 &  n24249 ;
  assign n24364 = x83 | n24077 ;
  assign n24365 = x83 &  n24077 ;
  assign n24366 = ( n24364 & ~n24365 ) | ( n24364 & 1'b0 ) | ( ~n24365 & 1'b0 ) ;
  assign n24375 = ( n5854 & n24232 ) | ( n5854 & n24366 ) | ( n24232 & n24366 ) ;
  assign n24376 = ( n24232 & ~n24248 ) | ( n24232 & n24366 ) | ( ~n24248 & n24366 ) ;
  assign n24377 = ~n24375 & n24376 ;
  assign n24378 = n24371 | n24377 ;
  assign n24379 = n24085 &  n24249 ;
  assign n24372 = x82 | n24085 ;
  assign n24373 = x82 &  n24085 ;
  assign n24374 = ( n24372 & ~n24373 ) | ( n24372 & 1'b0 ) | ( ~n24373 & 1'b0 ) ;
  assign n24383 = ( n5854 & n24231 ) | ( n5854 & n24374 ) | ( n24231 & n24374 ) ;
  assign n24384 = ( n24231 & ~n24248 ) | ( n24231 & n24374 ) | ( ~n24248 & n24374 ) ;
  assign n24385 = ~n24383 & n24384 ;
  assign n24386 = n24379 | n24385 ;
  assign n24387 = n24093 &  n24249 ;
  assign n24380 = x81 | n24093 ;
  assign n24381 = x81 &  n24093 ;
  assign n24382 = ( n24380 & ~n24381 ) | ( n24380 & 1'b0 ) | ( ~n24381 & 1'b0 ) ;
  assign n24391 = ( n5854 & n24230 ) | ( n5854 & n24382 ) | ( n24230 & n24382 ) ;
  assign n24392 = ( n24230 & ~n24248 ) | ( n24230 & n24382 ) | ( ~n24248 & n24382 ) ;
  assign n24393 = ~n24391 & n24392 ;
  assign n24394 = n24387 | n24393 ;
  assign n24395 = n24101 &  n24249 ;
  assign n24388 = x80 | n24101 ;
  assign n24389 = x80 &  n24101 ;
  assign n24390 = ( n24388 & ~n24389 ) | ( n24388 & 1'b0 ) | ( ~n24389 & 1'b0 ) ;
  assign n24399 = ( n5854 & n24229 ) | ( n5854 & n24390 ) | ( n24229 & n24390 ) ;
  assign n24400 = ( n24229 & ~n24248 ) | ( n24229 & n24390 ) | ( ~n24248 & n24390 ) ;
  assign n24401 = ~n24399 & n24400 ;
  assign n24402 = n24395 | n24401 ;
  assign n24403 = n24109 &  n24249 ;
  assign n24396 = x79 | n24109 ;
  assign n24397 = x79 &  n24109 ;
  assign n24398 = ( n24396 & ~n24397 ) | ( n24396 & 1'b0 ) | ( ~n24397 & 1'b0 ) ;
  assign n24407 = ( n5854 & n24228 ) | ( n5854 & n24398 ) | ( n24228 & n24398 ) ;
  assign n24408 = ( n24228 & ~n24248 ) | ( n24228 & n24398 ) | ( ~n24248 & n24398 ) ;
  assign n24409 = ~n24407 & n24408 ;
  assign n24410 = n24403 | n24409 ;
  assign n24411 = n24117 &  n24249 ;
  assign n24404 = x78 | n24117 ;
  assign n24405 = x78 &  n24117 ;
  assign n24406 = ( n24404 & ~n24405 ) | ( n24404 & 1'b0 ) | ( ~n24405 & 1'b0 ) ;
  assign n24415 = ( n5854 & n24227 ) | ( n5854 & n24406 ) | ( n24227 & n24406 ) ;
  assign n24416 = ( n24227 & ~n24248 ) | ( n24227 & n24406 ) | ( ~n24248 & n24406 ) ;
  assign n24417 = ~n24415 & n24416 ;
  assign n24418 = n24411 | n24417 ;
  assign n24419 = n24125 &  n24249 ;
  assign n24412 = x77 | n24125 ;
  assign n24413 = x77 &  n24125 ;
  assign n24414 = ( n24412 & ~n24413 ) | ( n24412 & 1'b0 ) | ( ~n24413 & 1'b0 ) ;
  assign n24423 = ( n5854 & n24226 ) | ( n5854 & n24414 ) | ( n24226 & n24414 ) ;
  assign n24424 = ( n24226 & ~n24248 ) | ( n24226 & n24414 ) | ( ~n24248 & n24414 ) ;
  assign n24425 = ~n24423 & n24424 ;
  assign n24426 = n24419 | n24425 ;
  assign n24427 = n24133 &  n24249 ;
  assign n24420 = x76 | n24133 ;
  assign n24421 = x76 &  n24133 ;
  assign n24422 = ( n24420 & ~n24421 ) | ( n24420 & 1'b0 ) | ( ~n24421 & 1'b0 ) ;
  assign n24431 = ( n5854 & n24225 ) | ( n5854 & n24422 ) | ( n24225 & n24422 ) ;
  assign n24432 = ( n24225 & ~n24248 ) | ( n24225 & n24422 ) | ( ~n24248 & n24422 ) ;
  assign n24433 = ~n24431 & n24432 ;
  assign n24434 = n24427 | n24433 ;
  assign n24435 = n24141 &  n24249 ;
  assign n24428 = x75 | n24141 ;
  assign n24429 = x75 &  n24141 ;
  assign n24430 = ( n24428 & ~n24429 ) | ( n24428 & 1'b0 ) | ( ~n24429 & 1'b0 ) ;
  assign n24439 = ( n5854 & n24224 ) | ( n5854 & n24430 ) | ( n24224 & n24430 ) ;
  assign n24440 = ( n24224 & ~n24248 ) | ( n24224 & n24430 ) | ( ~n24248 & n24430 ) ;
  assign n24441 = ~n24439 & n24440 ;
  assign n24442 = n24435 | n24441 ;
  assign n24443 = n24149 &  n24249 ;
  assign n24436 = x74 | n24149 ;
  assign n24437 = x74 &  n24149 ;
  assign n24438 = ( n24436 & ~n24437 ) | ( n24436 & 1'b0 ) | ( ~n24437 & 1'b0 ) ;
  assign n24447 = ( n5854 & n24223 ) | ( n5854 & n24438 ) | ( n24223 & n24438 ) ;
  assign n24448 = ( n24223 & ~n24248 ) | ( n24223 & n24438 ) | ( ~n24248 & n24438 ) ;
  assign n24449 = ~n24447 & n24448 ;
  assign n24450 = n24443 | n24449 ;
  assign n24451 = n24157 &  n24249 ;
  assign n24444 = x73 | n24157 ;
  assign n24445 = x73 &  n24157 ;
  assign n24446 = ( n24444 & ~n24445 ) | ( n24444 & 1'b0 ) | ( ~n24445 & 1'b0 ) ;
  assign n24455 = ( n5854 & n24222 ) | ( n5854 & n24446 ) | ( n24222 & n24446 ) ;
  assign n24456 = ( n24222 & ~n24248 ) | ( n24222 & n24446 ) | ( ~n24248 & n24446 ) ;
  assign n24457 = ~n24455 & n24456 ;
  assign n24458 = n24451 | n24457 ;
  assign n24459 = n24165 &  n24249 ;
  assign n24452 = x72 | n24165 ;
  assign n24453 = x72 &  n24165 ;
  assign n24454 = ( n24452 & ~n24453 ) | ( n24452 & 1'b0 ) | ( ~n24453 & 1'b0 ) ;
  assign n24463 = ( n5854 & n24221 ) | ( n5854 & n24454 ) | ( n24221 & n24454 ) ;
  assign n24464 = ( n24221 & ~n24248 ) | ( n24221 & n24454 ) | ( ~n24248 & n24454 ) ;
  assign n24465 = ~n24463 & n24464 ;
  assign n24466 = n24459 | n24465 ;
  assign n24467 = n24173 &  n24249 ;
  assign n24460 = x71 | n24173 ;
  assign n24461 = x71 &  n24173 ;
  assign n24462 = ( n24460 & ~n24461 ) | ( n24460 & 1'b0 ) | ( ~n24461 & 1'b0 ) ;
  assign n24471 = ( n5854 & n24220 ) | ( n5854 & n24462 ) | ( n24220 & n24462 ) ;
  assign n24472 = ( n24220 & ~n24248 ) | ( n24220 & n24462 ) | ( ~n24248 & n24462 ) ;
  assign n24473 = ~n24471 & n24472 ;
  assign n24474 = n24467 | n24473 ;
  assign n24475 = n24181 &  n24249 ;
  assign n24468 = x70 | n24181 ;
  assign n24469 = x70 &  n24181 ;
  assign n24470 = ( n24468 & ~n24469 ) | ( n24468 & 1'b0 ) | ( ~n24469 & 1'b0 ) ;
  assign n24479 = ( n5854 & n24219 ) | ( n5854 & n24470 ) | ( n24219 & n24470 ) ;
  assign n24480 = ( n24219 & ~n24248 ) | ( n24219 & n24470 ) | ( ~n24248 & n24470 ) ;
  assign n24481 = ~n24479 & n24480 ;
  assign n24482 = n24475 | n24481 ;
  assign n24483 = n24189 &  n24249 ;
  assign n24476 = x69 | n24189 ;
  assign n24477 = x69 &  n24189 ;
  assign n24478 = ( n24476 & ~n24477 ) | ( n24476 & 1'b0 ) | ( ~n24477 & 1'b0 ) ;
  assign n24487 = ( n5854 & n24218 ) | ( n5854 & n24478 ) | ( n24218 & n24478 ) ;
  assign n24488 = ( n24218 & ~n24248 ) | ( n24218 & n24478 ) | ( ~n24248 & n24478 ) ;
  assign n24489 = ~n24487 & n24488 ;
  assign n24490 = n24483 | n24489 ;
  assign n24491 = n24197 &  n24249 ;
  assign n24484 = x68 | n24197 ;
  assign n24485 = x68 &  n24197 ;
  assign n24486 = ( n24484 & ~n24485 ) | ( n24484 & 1'b0 ) | ( ~n24485 & 1'b0 ) ;
  assign n24495 = ( n5854 & n24217 ) | ( n5854 & n24486 ) | ( n24217 & n24486 ) ;
  assign n24496 = ( n24217 & ~n24248 ) | ( n24217 & n24486 ) | ( ~n24248 & n24486 ) ;
  assign n24497 = ~n24495 & n24496 ;
  assign n24498 = n24491 | n24497 ;
  assign n24499 = n24202 &  n24249 ;
  assign n24492 = x67 | n24202 ;
  assign n24493 = x67 &  n24202 ;
  assign n24494 = ( n24492 & ~n24493 ) | ( n24492 & 1'b0 ) | ( ~n24493 & 1'b0 ) ;
  assign n24503 = ( n5854 & n24216 ) | ( n5854 & n24494 ) | ( n24216 & n24494 ) ;
  assign n24504 = ( n24216 & ~n24248 ) | ( n24216 & n24494 ) | ( ~n24248 & n24494 ) ;
  assign n24505 = ~n24503 & n24504 ;
  assign n24506 = n24499 | n24505 ;
  assign n24507 = n24210 &  n24249 ;
  assign n24500 = x66 | n24210 ;
  assign n24501 = x66 &  n24210 ;
  assign n24502 = ( n24500 & ~n24501 ) | ( n24500 & 1'b0 ) | ( ~n24501 & 1'b0 ) ;
  assign n24511 = ( n5854 & n24215 ) | ( n5854 & n24502 ) | ( n24215 & n24502 ) ;
  assign n24512 = ( n24215 & ~n24248 ) | ( n24215 & n24502 ) | ( ~n24248 & n24502 ) ;
  assign n24513 = ~n24511 & n24512 ;
  assign n24514 = n24507 | n24513 ;
  assign n24515 = n24214 &  n24249 ;
  assign n24508 = x65 &  n24214 ;
  assign n24509 = x65 | n24213 ;
  assign n24510 = n24212 | n24509 ;
  assign n24516 = ~n24508 & n24510 ;
  assign n24517 = ( n5817 & ~n5854 ) | ( n5817 & n24516 ) | ( ~n5854 & n24516 ) ;
  assign n24518 = ( n5817 & n24248 ) | ( n5817 & n24516 ) | ( n24248 & n24516 ) ;
  assign n24519 = ( n24517 & ~n24518 ) | ( n24517 & 1'b0 ) | ( ~n24518 & 1'b0 ) ;
  assign n24520 = n24515 | n24519 ;
  assign n24521 = ( n5989 & ~n24248 ) | ( n5989 & 1'b0 ) | ( ~n24248 & 1'b0 ) ;
  assign n24522 = ( x29 & ~n24521 ) | ( x29 & 1'b0 ) | ( ~n24521 & 1'b0 ) ;
  assign n24523 = ( n5995 & ~n24248 ) | ( n5995 & 1'b0 ) | ( ~n24248 & 1'b0 ) ;
  assign n24524 = n24522 | n24523 ;
  assign n24525 = ( x65 & ~n24524 ) | ( x65 & n5998 ) | ( ~n24524 & n5998 ) ;
  assign n24526 = ( x66 & ~n24520 ) | ( x66 & n24525 ) | ( ~n24520 & n24525 ) ;
  assign n24527 = ( x67 & ~n24514 ) | ( x67 & n24526 ) | ( ~n24514 & n24526 ) ;
  assign n24528 = ( x68 & ~n24506 ) | ( x68 & n24527 ) | ( ~n24506 & n24527 ) ;
  assign n24529 = ( x69 & ~n24498 ) | ( x69 & n24528 ) | ( ~n24498 & n24528 ) ;
  assign n24530 = ( x70 & ~n24490 ) | ( x70 & n24529 ) | ( ~n24490 & n24529 ) ;
  assign n24531 = ( x71 & ~n24482 ) | ( x71 & n24530 ) | ( ~n24482 & n24530 ) ;
  assign n24532 = ( x72 & ~n24474 ) | ( x72 & n24531 ) | ( ~n24474 & n24531 ) ;
  assign n24533 = ( x73 & ~n24466 ) | ( x73 & n24532 ) | ( ~n24466 & n24532 ) ;
  assign n24534 = ( x74 & ~n24458 ) | ( x74 & n24533 ) | ( ~n24458 & n24533 ) ;
  assign n24535 = ( x75 & ~n24450 ) | ( x75 & n24534 ) | ( ~n24450 & n24534 ) ;
  assign n24536 = ( x76 & ~n24442 ) | ( x76 & n24535 ) | ( ~n24442 & n24535 ) ;
  assign n24537 = ( x77 & ~n24434 ) | ( x77 & n24536 ) | ( ~n24434 & n24536 ) ;
  assign n24538 = ( x78 & ~n24426 ) | ( x78 & n24537 ) | ( ~n24426 & n24537 ) ;
  assign n24539 = ( x79 & ~n24418 ) | ( x79 & n24538 ) | ( ~n24418 & n24538 ) ;
  assign n24540 = ( x80 & ~n24410 ) | ( x80 & n24539 ) | ( ~n24410 & n24539 ) ;
  assign n24541 = ( x81 & ~n24402 ) | ( x81 & n24540 ) | ( ~n24402 & n24540 ) ;
  assign n24542 = ( x82 & ~n24394 ) | ( x82 & n24541 ) | ( ~n24394 & n24541 ) ;
  assign n24543 = ( x83 & ~n24386 ) | ( x83 & n24542 ) | ( ~n24386 & n24542 ) ;
  assign n24544 = ( x84 & ~n24378 ) | ( x84 & n24543 ) | ( ~n24378 & n24543 ) ;
  assign n24545 = ( x85 & ~n24370 ) | ( x85 & n24544 ) | ( ~n24370 & n24544 ) ;
  assign n24546 = ( x86 & ~n24362 ) | ( x86 & n24545 ) | ( ~n24362 & n24545 ) ;
  assign n24547 = ( x87 & ~n24354 ) | ( x87 & n24546 ) | ( ~n24354 & n24546 ) ;
  assign n24548 = ( x88 & ~n24346 ) | ( x88 & n24547 ) | ( ~n24346 & n24547 ) ;
  assign n24549 = ( x89 & ~n24338 ) | ( x89 & n24548 ) | ( ~n24338 & n24548 ) ;
  assign n24550 = ( x90 & ~n24330 ) | ( x90 & n24549 ) | ( ~n24330 & n24549 ) ;
  assign n24551 = ( x91 & ~n24322 ) | ( x91 & n24550 ) | ( ~n24322 & n24550 ) ;
  assign n24552 = ( x92 & ~n24314 ) | ( x92 & n24551 ) | ( ~n24314 & n24551 ) ;
  assign n24553 = ( x93 & ~n24306 ) | ( x93 & n24552 ) | ( ~n24306 & n24552 ) ;
  assign n24554 = ( x94 & ~n24298 ) | ( x94 & n24553 ) | ( ~n24298 & n24553 ) ;
  assign n24555 = ( x95 & ~n24290 ) | ( x95 & n24554 ) | ( ~n24290 & n24554 ) ;
  assign n24556 = ( x96 & ~n24282 ) | ( x96 & n24555 ) | ( ~n24282 & n24555 ) ;
  assign n24557 = ( x97 & ~n24274 ) | ( x97 & n24556 ) | ( ~n24274 & n24556 ) ;
  assign n24558 = ( x98 & ~n24266 ) | ( x98 & n24557 ) | ( ~n24266 & n24557 ) ;
  assign n24559 = ( x99 & ~n24250 ) | ( x99 & 1'b0 ) | ( ~n24250 & 1'b0 ) ;
  assign n24560 = ~n24256 & n24559 ;
  assign n24561 = ( n24558 & ~n24258 ) | ( n24558 & n24560 ) | ( ~n24258 & n24560 ) ;
  assign n24562 = ( n24258 & ~n356 ) | ( n24258 & n24561 ) | ( ~n356 & n24561 ) ;
  assign n24563 = n356 | n24562 ;
  assign n24570 = n5854 &  n23957 ;
  assign n24571 = n24563 &  n24570 ;
  assign n24564 = ~n24257 |  n5854 ;
  assign n24565 = n24563 &  n24564 ;
  assign n24569 = n24258 | n24560 ;
  assign n24573 = ( n24558 & n24565 ) | ( n24558 & n24569 ) | ( n24565 & n24569 ) ;
  assign n24572 = n24558 | n24569 ;
  assign n24574 = ( n24571 & ~n24573 ) | ( n24571 & n24572 ) | ( ~n24573 & n24572 ) ;
  assign n24578 = n24266 &  n24564 ;
  assign n24579 = n24563 &  n24578 ;
  assign n24566 = x98 | n24266 ;
  assign n24567 = x98 &  n24266 ;
  assign n24568 = ( n24566 & ~n24567 ) | ( n24566 & 1'b0 ) | ( ~n24567 & 1'b0 ) ;
  assign n24581 = ( n24557 & n24565 ) | ( n24557 & n24568 ) | ( n24565 & n24568 ) ;
  assign n24580 = n24557 | n24568 ;
  assign n24582 = ( n24579 & ~n24581 ) | ( n24579 & n24580 ) | ( ~n24581 & n24580 ) ;
  assign n24586 = n24274 &  n24564 ;
  assign n24587 = n24563 &  n24586 ;
  assign n24575 = x97 | n24274 ;
  assign n24576 = x97 &  n24274 ;
  assign n24577 = ( n24575 & ~n24576 ) | ( n24575 & 1'b0 ) | ( ~n24576 & 1'b0 ) ;
  assign n24589 = ( n24556 & n24565 ) | ( n24556 & n24577 ) | ( n24565 & n24577 ) ;
  assign n24588 = n24556 | n24577 ;
  assign n24590 = ( n24587 & ~n24589 ) | ( n24587 & n24588 ) | ( ~n24589 & n24588 ) ;
  assign n24594 = n24282 &  n24564 ;
  assign n24595 = n24563 &  n24594 ;
  assign n24583 = x96 | n24282 ;
  assign n24584 = x96 &  n24282 ;
  assign n24585 = ( n24583 & ~n24584 ) | ( n24583 & 1'b0 ) | ( ~n24584 & 1'b0 ) ;
  assign n24597 = ( n24555 & n24565 ) | ( n24555 & n24585 ) | ( n24565 & n24585 ) ;
  assign n24596 = n24555 | n24585 ;
  assign n24598 = ( n24595 & ~n24597 ) | ( n24595 & n24596 ) | ( ~n24597 & n24596 ) ;
  assign n24602 = n24290 &  n24564 ;
  assign n24603 = n24563 &  n24602 ;
  assign n24591 = x95 | n24290 ;
  assign n24592 = x95 &  n24290 ;
  assign n24593 = ( n24591 & ~n24592 ) | ( n24591 & 1'b0 ) | ( ~n24592 & 1'b0 ) ;
  assign n24605 = ( n24554 & n24565 ) | ( n24554 & n24593 ) | ( n24565 & n24593 ) ;
  assign n24604 = n24554 | n24593 ;
  assign n24606 = ( n24603 & ~n24605 ) | ( n24603 & n24604 ) | ( ~n24605 & n24604 ) ;
  assign n24610 = n24298 &  n24564 ;
  assign n24611 = n24563 &  n24610 ;
  assign n24599 = x94 | n24298 ;
  assign n24600 = x94 &  n24298 ;
  assign n24601 = ( n24599 & ~n24600 ) | ( n24599 & 1'b0 ) | ( ~n24600 & 1'b0 ) ;
  assign n24613 = ( n24553 & n24565 ) | ( n24553 & n24601 ) | ( n24565 & n24601 ) ;
  assign n24612 = n24553 | n24601 ;
  assign n24614 = ( n24611 & ~n24613 ) | ( n24611 & n24612 ) | ( ~n24613 & n24612 ) ;
  assign n24618 = n24306 &  n24564 ;
  assign n24619 = n24563 &  n24618 ;
  assign n24607 = x93 | n24306 ;
  assign n24608 = x93 &  n24306 ;
  assign n24609 = ( n24607 & ~n24608 ) | ( n24607 & 1'b0 ) | ( ~n24608 & 1'b0 ) ;
  assign n24621 = ( n24552 & n24565 ) | ( n24552 & n24609 ) | ( n24565 & n24609 ) ;
  assign n24620 = n24552 | n24609 ;
  assign n24622 = ( n24619 & ~n24621 ) | ( n24619 & n24620 ) | ( ~n24621 & n24620 ) ;
  assign n24626 = n24314 &  n24564 ;
  assign n24627 = n24563 &  n24626 ;
  assign n24615 = x92 | n24314 ;
  assign n24616 = x92 &  n24314 ;
  assign n24617 = ( n24615 & ~n24616 ) | ( n24615 & 1'b0 ) | ( ~n24616 & 1'b0 ) ;
  assign n24629 = ( n24551 & n24565 ) | ( n24551 & n24617 ) | ( n24565 & n24617 ) ;
  assign n24628 = n24551 | n24617 ;
  assign n24630 = ( n24627 & ~n24629 ) | ( n24627 & n24628 ) | ( ~n24629 & n24628 ) ;
  assign n24634 = n24322 &  n24564 ;
  assign n24635 = n24563 &  n24634 ;
  assign n24623 = x91 | n24322 ;
  assign n24624 = x91 &  n24322 ;
  assign n24625 = ( n24623 & ~n24624 ) | ( n24623 & 1'b0 ) | ( ~n24624 & 1'b0 ) ;
  assign n24637 = ( n24550 & n24565 ) | ( n24550 & n24625 ) | ( n24565 & n24625 ) ;
  assign n24636 = n24550 | n24625 ;
  assign n24638 = ( n24635 & ~n24637 ) | ( n24635 & n24636 ) | ( ~n24637 & n24636 ) ;
  assign n24642 = n24330 &  n24564 ;
  assign n24643 = n24563 &  n24642 ;
  assign n24631 = x90 | n24330 ;
  assign n24632 = x90 &  n24330 ;
  assign n24633 = ( n24631 & ~n24632 ) | ( n24631 & 1'b0 ) | ( ~n24632 & 1'b0 ) ;
  assign n24645 = ( n24549 & n24565 ) | ( n24549 & n24633 ) | ( n24565 & n24633 ) ;
  assign n24644 = n24549 | n24633 ;
  assign n24646 = ( n24643 & ~n24645 ) | ( n24643 & n24644 ) | ( ~n24645 & n24644 ) ;
  assign n24650 = n24338 &  n24564 ;
  assign n24651 = n24563 &  n24650 ;
  assign n24639 = x89 | n24338 ;
  assign n24640 = x89 &  n24338 ;
  assign n24641 = ( n24639 & ~n24640 ) | ( n24639 & 1'b0 ) | ( ~n24640 & 1'b0 ) ;
  assign n24653 = ( n24548 & n24565 ) | ( n24548 & n24641 ) | ( n24565 & n24641 ) ;
  assign n24652 = n24548 | n24641 ;
  assign n24654 = ( n24651 & ~n24653 ) | ( n24651 & n24652 ) | ( ~n24653 & n24652 ) ;
  assign n24658 = n24346 &  n24564 ;
  assign n24659 = n24563 &  n24658 ;
  assign n24647 = x88 | n24346 ;
  assign n24648 = x88 &  n24346 ;
  assign n24649 = ( n24647 & ~n24648 ) | ( n24647 & 1'b0 ) | ( ~n24648 & 1'b0 ) ;
  assign n24661 = ( n24547 & n24565 ) | ( n24547 & n24649 ) | ( n24565 & n24649 ) ;
  assign n24660 = n24547 | n24649 ;
  assign n24662 = ( n24659 & ~n24661 ) | ( n24659 & n24660 ) | ( ~n24661 & n24660 ) ;
  assign n24666 = n24354 &  n24564 ;
  assign n24667 = n24563 &  n24666 ;
  assign n24655 = x87 | n24354 ;
  assign n24656 = x87 &  n24354 ;
  assign n24657 = ( n24655 & ~n24656 ) | ( n24655 & 1'b0 ) | ( ~n24656 & 1'b0 ) ;
  assign n24669 = ( n24546 & n24565 ) | ( n24546 & n24657 ) | ( n24565 & n24657 ) ;
  assign n24668 = n24546 | n24657 ;
  assign n24670 = ( n24667 & ~n24669 ) | ( n24667 & n24668 ) | ( ~n24669 & n24668 ) ;
  assign n24674 = n24362 &  n24564 ;
  assign n24675 = n24563 &  n24674 ;
  assign n24663 = x86 | n24362 ;
  assign n24664 = x86 &  n24362 ;
  assign n24665 = ( n24663 & ~n24664 ) | ( n24663 & 1'b0 ) | ( ~n24664 & 1'b0 ) ;
  assign n24677 = ( n24545 & n24565 ) | ( n24545 & n24665 ) | ( n24565 & n24665 ) ;
  assign n24676 = n24545 | n24665 ;
  assign n24678 = ( n24675 & ~n24677 ) | ( n24675 & n24676 ) | ( ~n24677 & n24676 ) ;
  assign n24682 = n24370 &  n24564 ;
  assign n24683 = n24563 &  n24682 ;
  assign n24671 = x85 | n24370 ;
  assign n24672 = x85 &  n24370 ;
  assign n24673 = ( n24671 & ~n24672 ) | ( n24671 & 1'b0 ) | ( ~n24672 & 1'b0 ) ;
  assign n24685 = ( n24544 & n24565 ) | ( n24544 & n24673 ) | ( n24565 & n24673 ) ;
  assign n24684 = n24544 | n24673 ;
  assign n24686 = ( n24683 & ~n24685 ) | ( n24683 & n24684 ) | ( ~n24685 & n24684 ) ;
  assign n24690 = n24378 &  n24564 ;
  assign n24691 = n24563 &  n24690 ;
  assign n24679 = x84 | n24378 ;
  assign n24680 = x84 &  n24378 ;
  assign n24681 = ( n24679 & ~n24680 ) | ( n24679 & 1'b0 ) | ( ~n24680 & 1'b0 ) ;
  assign n24693 = ( n24543 & n24565 ) | ( n24543 & n24681 ) | ( n24565 & n24681 ) ;
  assign n24692 = n24543 | n24681 ;
  assign n24694 = ( n24691 & ~n24693 ) | ( n24691 & n24692 ) | ( ~n24693 & n24692 ) ;
  assign n24698 = n24386 &  n24564 ;
  assign n24699 = n24563 &  n24698 ;
  assign n24687 = x83 | n24386 ;
  assign n24688 = x83 &  n24386 ;
  assign n24689 = ( n24687 & ~n24688 ) | ( n24687 & 1'b0 ) | ( ~n24688 & 1'b0 ) ;
  assign n24701 = ( n24542 & n24565 ) | ( n24542 & n24689 ) | ( n24565 & n24689 ) ;
  assign n24700 = n24542 | n24689 ;
  assign n24702 = ( n24699 & ~n24701 ) | ( n24699 & n24700 ) | ( ~n24701 & n24700 ) ;
  assign n24706 = n24394 &  n24564 ;
  assign n24707 = n24563 &  n24706 ;
  assign n24695 = x82 | n24394 ;
  assign n24696 = x82 &  n24394 ;
  assign n24697 = ( n24695 & ~n24696 ) | ( n24695 & 1'b0 ) | ( ~n24696 & 1'b0 ) ;
  assign n24709 = ( n24541 & n24565 ) | ( n24541 & n24697 ) | ( n24565 & n24697 ) ;
  assign n24708 = n24541 | n24697 ;
  assign n24710 = ( n24707 & ~n24709 ) | ( n24707 & n24708 ) | ( ~n24709 & n24708 ) ;
  assign n24714 = n24402 &  n24564 ;
  assign n24715 = n24563 &  n24714 ;
  assign n24703 = x81 | n24402 ;
  assign n24704 = x81 &  n24402 ;
  assign n24705 = ( n24703 & ~n24704 ) | ( n24703 & 1'b0 ) | ( ~n24704 & 1'b0 ) ;
  assign n24717 = ( n24540 & n24565 ) | ( n24540 & n24705 ) | ( n24565 & n24705 ) ;
  assign n24716 = n24540 | n24705 ;
  assign n24718 = ( n24715 & ~n24717 ) | ( n24715 & n24716 ) | ( ~n24717 & n24716 ) ;
  assign n24722 = n24410 &  n24564 ;
  assign n24723 = n24563 &  n24722 ;
  assign n24711 = x80 | n24410 ;
  assign n24712 = x80 &  n24410 ;
  assign n24713 = ( n24711 & ~n24712 ) | ( n24711 & 1'b0 ) | ( ~n24712 & 1'b0 ) ;
  assign n24725 = ( n24539 & n24565 ) | ( n24539 & n24713 ) | ( n24565 & n24713 ) ;
  assign n24724 = n24539 | n24713 ;
  assign n24726 = ( n24723 & ~n24725 ) | ( n24723 & n24724 ) | ( ~n24725 & n24724 ) ;
  assign n24730 = n24418 &  n24564 ;
  assign n24731 = n24563 &  n24730 ;
  assign n24719 = x79 | n24418 ;
  assign n24720 = x79 &  n24418 ;
  assign n24721 = ( n24719 & ~n24720 ) | ( n24719 & 1'b0 ) | ( ~n24720 & 1'b0 ) ;
  assign n24733 = ( n24538 & n24565 ) | ( n24538 & n24721 ) | ( n24565 & n24721 ) ;
  assign n24732 = n24538 | n24721 ;
  assign n24734 = ( n24731 & ~n24733 ) | ( n24731 & n24732 ) | ( ~n24733 & n24732 ) ;
  assign n24738 = n24426 &  n24564 ;
  assign n24739 = n24563 &  n24738 ;
  assign n24727 = x78 | n24426 ;
  assign n24728 = x78 &  n24426 ;
  assign n24729 = ( n24727 & ~n24728 ) | ( n24727 & 1'b0 ) | ( ~n24728 & 1'b0 ) ;
  assign n24741 = ( n24537 & n24565 ) | ( n24537 & n24729 ) | ( n24565 & n24729 ) ;
  assign n24740 = n24537 | n24729 ;
  assign n24742 = ( n24739 & ~n24741 ) | ( n24739 & n24740 ) | ( ~n24741 & n24740 ) ;
  assign n24746 = n24434 &  n24564 ;
  assign n24747 = n24563 &  n24746 ;
  assign n24735 = x77 | n24434 ;
  assign n24736 = x77 &  n24434 ;
  assign n24737 = ( n24735 & ~n24736 ) | ( n24735 & 1'b0 ) | ( ~n24736 & 1'b0 ) ;
  assign n24749 = ( n24536 & n24565 ) | ( n24536 & n24737 ) | ( n24565 & n24737 ) ;
  assign n24748 = n24536 | n24737 ;
  assign n24750 = ( n24747 & ~n24749 ) | ( n24747 & n24748 ) | ( ~n24749 & n24748 ) ;
  assign n24754 = n24442 &  n24564 ;
  assign n24755 = n24563 &  n24754 ;
  assign n24743 = x76 | n24442 ;
  assign n24744 = x76 &  n24442 ;
  assign n24745 = ( n24743 & ~n24744 ) | ( n24743 & 1'b0 ) | ( ~n24744 & 1'b0 ) ;
  assign n24757 = ( n24535 & n24565 ) | ( n24535 & n24745 ) | ( n24565 & n24745 ) ;
  assign n24756 = n24535 | n24745 ;
  assign n24758 = ( n24755 & ~n24757 ) | ( n24755 & n24756 ) | ( ~n24757 & n24756 ) ;
  assign n24762 = n24450 &  n24564 ;
  assign n24763 = n24563 &  n24762 ;
  assign n24751 = x75 | n24450 ;
  assign n24752 = x75 &  n24450 ;
  assign n24753 = ( n24751 & ~n24752 ) | ( n24751 & 1'b0 ) | ( ~n24752 & 1'b0 ) ;
  assign n24765 = ( n24534 & n24565 ) | ( n24534 & n24753 ) | ( n24565 & n24753 ) ;
  assign n24764 = n24534 | n24753 ;
  assign n24766 = ( n24763 & ~n24765 ) | ( n24763 & n24764 ) | ( ~n24765 & n24764 ) ;
  assign n24770 = n24458 &  n24564 ;
  assign n24771 = n24563 &  n24770 ;
  assign n24759 = x74 | n24458 ;
  assign n24760 = x74 &  n24458 ;
  assign n24761 = ( n24759 & ~n24760 ) | ( n24759 & 1'b0 ) | ( ~n24760 & 1'b0 ) ;
  assign n24773 = ( n24533 & n24565 ) | ( n24533 & n24761 ) | ( n24565 & n24761 ) ;
  assign n24772 = n24533 | n24761 ;
  assign n24774 = ( n24771 & ~n24773 ) | ( n24771 & n24772 ) | ( ~n24773 & n24772 ) ;
  assign n24778 = n24466 &  n24564 ;
  assign n24779 = n24563 &  n24778 ;
  assign n24767 = x73 | n24466 ;
  assign n24768 = x73 &  n24466 ;
  assign n24769 = ( n24767 & ~n24768 ) | ( n24767 & 1'b0 ) | ( ~n24768 & 1'b0 ) ;
  assign n24781 = ( n24532 & n24565 ) | ( n24532 & n24769 ) | ( n24565 & n24769 ) ;
  assign n24780 = n24532 | n24769 ;
  assign n24782 = ( n24779 & ~n24781 ) | ( n24779 & n24780 ) | ( ~n24781 & n24780 ) ;
  assign n24786 = n24474 &  n24564 ;
  assign n24787 = n24563 &  n24786 ;
  assign n24775 = x72 | n24474 ;
  assign n24776 = x72 &  n24474 ;
  assign n24777 = ( n24775 & ~n24776 ) | ( n24775 & 1'b0 ) | ( ~n24776 & 1'b0 ) ;
  assign n24789 = ( n24531 & n24565 ) | ( n24531 & n24777 ) | ( n24565 & n24777 ) ;
  assign n24788 = n24531 | n24777 ;
  assign n24790 = ( n24787 & ~n24789 ) | ( n24787 & n24788 ) | ( ~n24789 & n24788 ) ;
  assign n24794 = n24482 &  n24564 ;
  assign n24795 = n24563 &  n24794 ;
  assign n24783 = x71 | n24482 ;
  assign n24784 = x71 &  n24482 ;
  assign n24785 = ( n24783 & ~n24784 ) | ( n24783 & 1'b0 ) | ( ~n24784 & 1'b0 ) ;
  assign n24797 = ( n24530 & n24565 ) | ( n24530 & n24785 ) | ( n24565 & n24785 ) ;
  assign n24796 = n24530 | n24785 ;
  assign n24798 = ( n24795 & ~n24797 ) | ( n24795 & n24796 ) | ( ~n24797 & n24796 ) ;
  assign n24802 = n24490 &  n24564 ;
  assign n24803 = n24563 &  n24802 ;
  assign n24791 = x70 | n24490 ;
  assign n24792 = x70 &  n24490 ;
  assign n24793 = ( n24791 & ~n24792 ) | ( n24791 & 1'b0 ) | ( ~n24792 & 1'b0 ) ;
  assign n24805 = ( n24529 & n24565 ) | ( n24529 & n24793 ) | ( n24565 & n24793 ) ;
  assign n24804 = n24529 | n24793 ;
  assign n24806 = ( n24803 & ~n24805 ) | ( n24803 & n24804 ) | ( ~n24805 & n24804 ) ;
  assign n24810 = n24498 &  n24564 ;
  assign n24811 = n24563 &  n24810 ;
  assign n24799 = x69 | n24498 ;
  assign n24800 = x69 &  n24498 ;
  assign n24801 = ( n24799 & ~n24800 ) | ( n24799 & 1'b0 ) | ( ~n24800 & 1'b0 ) ;
  assign n24813 = ( n24528 & n24565 ) | ( n24528 & n24801 ) | ( n24565 & n24801 ) ;
  assign n24812 = n24528 | n24801 ;
  assign n24814 = ( n24811 & ~n24813 ) | ( n24811 & n24812 ) | ( ~n24813 & n24812 ) ;
  assign n24818 = n24506 &  n24564 ;
  assign n24819 = n24563 &  n24818 ;
  assign n24807 = x68 | n24506 ;
  assign n24808 = x68 &  n24506 ;
  assign n24809 = ( n24807 & ~n24808 ) | ( n24807 & 1'b0 ) | ( ~n24808 & 1'b0 ) ;
  assign n24821 = ( n24527 & n24565 ) | ( n24527 & n24809 ) | ( n24565 & n24809 ) ;
  assign n24820 = n24527 | n24809 ;
  assign n24822 = ( n24819 & ~n24821 ) | ( n24819 & n24820 ) | ( ~n24821 & n24820 ) ;
  assign n24826 = n24514 &  n24564 ;
  assign n24827 = n24563 &  n24826 ;
  assign n24815 = x67 | n24514 ;
  assign n24816 = x67 &  n24514 ;
  assign n24817 = ( n24815 & ~n24816 ) | ( n24815 & 1'b0 ) | ( ~n24816 & 1'b0 ) ;
  assign n24829 = ( n24526 & n24565 ) | ( n24526 & n24817 ) | ( n24565 & n24817 ) ;
  assign n24828 = n24526 | n24817 ;
  assign n24830 = ( n24827 & ~n24829 ) | ( n24827 & n24828 ) | ( ~n24829 & n24828 ) ;
  assign n24831 = n24520 &  n24564 ;
  assign n24832 = n24563 &  n24831 ;
  assign n24823 = x66 | n24520 ;
  assign n24824 = x66 &  n24520 ;
  assign n24825 = ( n24823 & ~n24824 ) | ( n24823 & 1'b0 ) | ( ~n24824 & 1'b0 ) ;
  assign n24834 = ( n24525 & n24565 ) | ( n24525 & n24825 ) | ( n24565 & n24825 ) ;
  assign n24833 = n24525 | n24825 ;
  assign n24835 = ( n24832 & ~n24834 ) | ( n24832 & n24833 ) | ( ~n24834 & n24833 ) ;
  assign n24836 = ( x65 & ~n5998 ) | ( x65 & n24524 ) | ( ~n5998 & n24524 ) ;
  assign n24837 = ( n24525 & ~x65 ) | ( n24525 & n24836 ) | ( ~x65 & n24836 ) ;
  assign n24838 = ~n24565 & n24837 ;
  assign n24839 = n24524 &  n24564 ;
  assign n24840 = n24563 &  n24839 ;
  assign n24841 = n24838 | n24840 ;
  assign n24842 = ( x64 & ~n24565 ) | ( x64 & 1'b0 ) | ( ~n24565 & 1'b0 ) ;
  assign n24843 = ( x28 & ~n24842 ) | ( x28 & 1'b0 ) | ( ~n24842 & 1'b0 ) ;
  assign n24844 = ( n5998 & ~n24565 ) | ( n5998 & 1'b0 ) | ( ~n24565 & 1'b0 ) ;
  assign n24845 = n24843 | n24844 ;
  assign n24846 = ( x65 & ~n24845 ) | ( x65 & n6462 ) | ( ~n24845 & n6462 ) ;
  assign n24847 = ( x66 & ~n24841 ) | ( x66 & n24846 ) | ( ~n24841 & n24846 ) ;
  assign n24848 = ( x67 & ~n24835 ) | ( x67 & n24847 ) | ( ~n24835 & n24847 ) ;
  assign n24849 = ( x68 & ~n24830 ) | ( x68 & n24848 ) | ( ~n24830 & n24848 ) ;
  assign n24850 = ( x69 & ~n24822 ) | ( x69 & n24849 ) | ( ~n24822 & n24849 ) ;
  assign n24851 = ( x70 & ~n24814 ) | ( x70 & n24850 ) | ( ~n24814 & n24850 ) ;
  assign n24852 = ( x71 & ~n24806 ) | ( x71 & n24851 ) | ( ~n24806 & n24851 ) ;
  assign n24853 = ( x72 & ~n24798 ) | ( x72 & n24852 ) | ( ~n24798 & n24852 ) ;
  assign n24854 = ( x73 & ~n24790 ) | ( x73 & n24853 ) | ( ~n24790 & n24853 ) ;
  assign n24855 = ( x74 & ~n24782 ) | ( x74 & n24854 ) | ( ~n24782 & n24854 ) ;
  assign n24856 = ( x75 & ~n24774 ) | ( x75 & n24855 ) | ( ~n24774 & n24855 ) ;
  assign n24857 = ( x76 & ~n24766 ) | ( x76 & n24856 ) | ( ~n24766 & n24856 ) ;
  assign n24858 = ( x77 & ~n24758 ) | ( x77 & n24857 ) | ( ~n24758 & n24857 ) ;
  assign n24859 = ( x78 & ~n24750 ) | ( x78 & n24858 ) | ( ~n24750 & n24858 ) ;
  assign n24860 = ( x79 & ~n24742 ) | ( x79 & n24859 ) | ( ~n24742 & n24859 ) ;
  assign n24861 = ( x80 & ~n24734 ) | ( x80 & n24860 ) | ( ~n24734 & n24860 ) ;
  assign n24862 = ( x81 & ~n24726 ) | ( x81 & n24861 ) | ( ~n24726 & n24861 ) ;
  assign n24863 = ( x82 & ~n24718 ) | ( x82 & n24862 ) | ( ~n24718 & n24862 ) ;
  assign n24864 = ( x83 & ~n24710 ) | ( x83 & n24863 ) | ( ~n24710 & n24863 ) ;
  assign n24865 = ( x84 & ~n24702 ) | ( x84 & n24864 ) | ( ~n24702 & n24864 ) ;
  assign n24866 = ( x85 & ~n24694 ) | ( x85 & n24865 ) | ( ~n24694 & n24865 ) ;
  assign n24867 = ( x86 & ~n24686 ) | ( x86 & n24866 ) | ( ~n24686 & n24866 ) ;
  assign n24868 = ( x87 & ~n24678 ) | ( x87 & n24867 ) | ( ~n24678 & n24867 ) ;
  assign n24869 = ( x88 & ~n24670 ) | ( x88 & n24868 ) | ( ~n24670 & n24868 ) ;
  assign n24870 = ( x89 & ~n24662 ) | ( x89 & n24869 ) | ( ~n24662 & n24869 ) ;
  assign n24871 = ( x90 & ~n24654 ) | ( x90 & n24870 ) | ( ~n24654 & n24870 ) ;
  assign n24872 = ( x91 & ~n24646 ) | ( x91 & n24871 ) | ( ~n24646 & n24871 ) ;
  assign n24873 = ( x92 & ~n24638 ) | ( x92 & n24872 ) | ( ~n24638 & n24872 ) ;
  assign n24874 = ( x93 & ~n24630 ) | ( x93 & n24873 ) | ( ~n24630 & n24873 ) ;
  assign n24875 = ( x94 & ~n24622 ) | ( x94 & n24874 ) | ( ~n24622 & n24874 ) ;
  assign n24876 = ( x95 & ~n24614 ) | ( x95 & n24875 ) | ( ~n24614 & n24875 ) ;
  assign n24877 = ( x96 & ~n24606 ) | ( x96 & n24876 ) | ( ~n24606 & n24876 ) ;
  assign n24878 = ( x97 & ~n24598 ) | ( x97 & n24877 ) | ( ~n24598 & n24877 ) ;
  assign n24879 = ( x98 & ~n24590 ) | ( x98 & n24878 ) | ( ~n24590 & n24878 ) ;
  assign n24880 = ( x99 & ~n24582 ) | ( x99 & n24879 ) | ( ~n24582 & n24879 ) ;
  assign n24887 = ( x100 & ~n429 ) | ( x100 & n24880 ) | ( ~n429 & n24880 ) ;
  assign n24886 = x100 &  n24880 ;
  assign n24888 = ( n24574 & ~n24887 ) | ( n24574 & n24886 ) | ( ~n24887 & n24886 ) ;
  assign n24881 = ( x100 & ~n24574 ) | ( x100 & n24880 ) | ( ~n24574 & n24880 ) ;
  assign n24882 = n429 | n24881 ;
  assign n24889 = n24582 &  n24882 ;
  assign n24883 = x99 | n24582 ;
  assign n24884 = x99 &  n24582 ;
  assign n24885 = ( n24883 & ~n24884 ) | ( n24883 & 1'b0 ) | ( ~n24884 & 1'b0 ) ;
  assign n24893 = ( n429 & n24879 ) | ( n429 & n24885 ) | ( n24879 & n24885 ) ;
  assign n24894 = ( n24879 & ~n24881 ) | ( n24879 & n24885 ) | ( ~n24881 & n24885 ) ;
  assign n24895 = ~n24893 & n24894 ;
  assign n24896 = n24889 | n24895 ;
  assign n24897 = n24590 &  n24882 ;
  assign n24890 = x98 | n24590 ;
  assign n24891 = x98 &  n24590 ;
  assign n24892 = ( n24890 & ~n24891 ) | ( n24890 & 1'b0 ) | ( ~n24891 & 1'b0 ) ;
  assign n24901 = ( n429 & n24878 ) | ( n429 & n24892 ) | ( n24878 & n24892 ) ;
  assign n24902 = ( n24878 & ~n24881 ) | ( n24878 & n24892 ) | ( ~n24881 & n24892 ) ;
  assign n24903 = ~n24901 & n24902 ;
  assign n24904 = n24897 | n24903 ;
  assign n24905 = n24598 &  n24882 ;
  assign n24898 = x97 | n24598 ;
  assign n24899 = x97 &  n24598 ;
  assign n24900 = ( n24898 & ~n24899 ) | ( n24898 & 1'b0 ) | ( ~n24899 & 1'b0 ) ;
  assign n24909 = ( n429 & n24877 ) | ( n429 & n24900 ) | ( n24877 & n24900 ) ;
  assign n24910 = ( n24877 & ~n24881 ) | ( n24877 & n24900 ) | ( ~n24881 & n24900 ) ;
  assign n24911 = ~n24909 & n24910 ;
  assign n24912 = n24905 | n24911 ;
  assign n24913 = n24606 &  n24882 ;
  assign n24906 = x96 | n24606 ;
  assign n24907 = x96 &  n24606 ;
  assign n24908 = ( n24906 & ~n24907 ) | ( n24906 & 1'b0 ) | ( ~n24907 & 1'b0 ) ;
  assign n24917 = ( n429 & n24876 ) | ( n429 & n24908 ) | ( n24876 & n24908 ) ;
  assign n24918 = ( n24876 & ~n24881 ) | ( n24876 & n24908 ) | ( ~n24881 & n24908 ) ;
  assign n24919 = ~n24917 & n24918 ;
  assign n24920 = n24913 | n24919 ;
  assign n24921 = n24614 &  n24882 ;
  assign n24914 = x95 | n24614 ;
  assign n24915 = x95 &  n24614 ;
  assign n24916 = ( n24914 & ~n24915 ) | ( n24914 & 1'b0 ) | ( ~n24915 & 1'b0 ) ;
  assign n24925 = ( n429 & n24875 ) | ( n429 & n24916 ) | ( n24875 & n24916 ) ;
  assign n24926 = ( n24875 & ~n24881 ) | ( n24875 & n24916 ) | ( ~n24881 & n24916 ) ;
  assign n24927 = ~n24925 & n24926 ;
  assign n24928 = n24921 | n24927 ;
  assign n24929 = n24622 &  n24882 ;
  assign n24922 = x94 | n24622 ;
  assign n24923 = x94 &  n24622 ;
  assign n24924 = ( n24922 & ~n24923 ) | ( n24922 & 1'b0 ) | ( ~n24923 & 1'b0 ) ;
  assign n24933 = ( n429 & n24874 ) | ( n429 & n24924 ) | ( n24874 & n24924 ) ;
  assign n24934 = ( n24874 & ~n24881 ) | ( n24874 & n24924 ) | ( ~n24881 & n24924 ) ;
  assign n24935 = ~n24933 & n24934 ;
  assign n24936 = n24929 | n24935 ;
  assign n24937 = n24630 &  n24882 ;
  assign n24930 = x93 | n24630 ;
  assign n24931 = x93 &  n24630 ;
  assign n24932 = ( n24930 & ~n24931 ) | ( n24930 & 1'b0 ) | ( ~n24931 & 1'b0 ) ;
  assign n24941 = ( n429 & n24873 ) | ( n429 & n24932 ) | ( n24873 & n24932 ) ;
  assign n24942 = ( n24873 & ~n24881 ) | ( n24873 & n24932 ) | ( ~n24881 & n24932 ) ;
  assign n24943 = ~n24941 & n24942 ;
  assign n24944 = n24937 | n24943 ;
  assign n24945 = n24638 &  n24882 ;
  assign n24938 = x92 | n24638 ;
  assign n24939 = x92 &  n24638 ;
  assign n24940 = ( n24938 & ~n24939 ) | ( n24938 & 1'b0 ) | ( ~n24939 & 1'b0 ) ;
  assign n24949 = ( n429 & n24872 ) | ( n429 & n24940 ) | ( n24872 & n24940 ) ;
  assign n24950 = ( n24872 & ~n24881 ) | ( n24872 & n24940 ) | ( ~n24881 & n24940 ) ;
  assign n24951 = ~n24949 & n24950 ;
  assign n24952 = n24945 | n24951 ;
  assign n24953 = n24646 &  n24882 ;
  assign n24946 = x91 | n24646 ;
  assign n24947 = x91 &  n24646 ;
  assign n24948 = ( n24946 & ~n24947 ) | ( n24946 & 1'b0 ) | ( ~n24947 & 1'b0 ) ;
  assign n24957 = ( n429 & n24871 ) | ( n429 & n24948 ) | ( n24871 & n24948 ) ;
  assign n24958 = ( n24871 & ~n24881 ) | ( n24871 & n24948 ) | ( ~n24881 & n24948 ) ;
  assign n24959 = ~n24957 & n24958 ;
  assign n24960 = n24953 | n24959 ;
  assign n24961 = n24654 &  n24882 ;
  assign n24954 = x90 | n24654 ;
  assign n24955 = x90 &  n24654 ;
  assign n24956 = ( n24954 & ~n24955 ) | ( n24954 & 1'b0 ) | ( ~n24955 & 1'b0 ) ;
  assign n24965 = ( n429 & n24870 ) | ( n429 & n24956 ) | ( n24870 & n24956 ) ;
  assign n24966 = ( n24870 & ~n24881 ) | ( n24870 & n24956 ) | ( ~n24881 & n24956 ) ;
  assign n24967 = ~n24965 & n24966 ;
  assign n24968 = n24961 | n24967 ;
  assign n24969 = n24662 &  n24882 ;
  assign n24962 = x89 | n24662 ;
  assign n24963 = x89 &  n24662 ;
  assign n24964 = ( n24962 & ~n24963 ) | ( n24962 & 1'b0 ) | ( ~n24963 & 1'b0 ) ;
  assign n24973 = ( n429 & n24869 ) | ( n429 & n24964 ) | ( n24869 & n24964 ) ;
  assign n24974 = ( n24869 & ~n24881 ) | ( n24869 & n24964 ) | ( ~n24881 & n24964 ) ;
  assign n24975 = ~n24973 & n24974 ;
  assign n24976 = n24969 | n24975 ;
  assign n24977 = n24670 &  n24882 ;
  assign n24970 = x88 | n24670 ;
  assign n24971 = x88 &  n24670 ;
  assign n24972 = ( n24970 & ~n24971 ) | ( n24970 & 1'b0 ) | ( ~n24971 & 1'b0 ) ;
  assign n24981 = ( n429 & n24868 ) | ( n429 & n24972 ) | ( n24868 & n24972 ) ;
  assign n24982 = ( n24868 & ~n24881 ) | ( n24868 & n24972 ) | ( ~n24881 & n24972 ) ;
  assign n24983 = ~n24981 & n24982 ;
  assign n24984 = n24977 | n24983 ;
  assign n24985 = n24678 &  n24882 ;
  assign n24978 = x87 | n24678 ;
  assign n24979 = x87 &  n24678 ;
  assign n24980 = ( n24978 & ~n24979 ) | ( n24978 & 1'b0 ) | ( ~n24979 & 1'b0 ) ;
  assign n24989 = ( n429 & n24867 ) | ( n429 & n24980 ) | ( n24867 & n24980 ) ;
  assign n24990 = ( n24867 & ~n24881 ) | ( n24867 & n24980 ) | ( ~n24881 & n24980 ) ;
  assign n24991 = ~n24989 & n24990 ;
  assign n24992 = n24985 | n24991 ;
  assign n24993 = n24686 &  n24882 ;
  assign n24986 = x86 | n24686 ;
  assign n24987 = x86 &  n24686 ;
  assign n24988 = ( n24986 & ~n24987 ) | ( n24986 & 1'b0 ) | ( ~n24987 & 1'b0 ) ;
  assign n24997 = ( n429 & n24866 ) | ( n429 & n24988 ) | ( n24866 & n24988 ) ;
  assign n24998 = ( n24866 & ~n24881 ) | ( n24866 & n24988 ) | ( ~n24881 & n24988 ) ;
  assign n24999 = ~n24997 & n24998 ;
  assign n25000 = n24993 | n24999 ;
  assign n25001 = n24694 &  n24882 ;
  assign n24994 = x85 | n24694 ;
  assign n24995 = x85 &  n24694 ;
  assign n24996 = ( n24994 & ~n24995 ) | ( n24994 & 1'b0 ) | ( ~n24995 & 1'b0 ) ;
  assign n25005 = ( n429 & n24865 ) | ( n429 & n24996 ) | ( n24865 & n24996 ) ;
  assign n25006 = ( n24865 & ~n24881 ) | ( n24865 & n24996 ) | ( ~n24881 & n24996 ) ;
  assign n25007 = ~n25005 & n25006 ;
  assign n25008 = n25001 | n25007 ;
  assign n25009 = n24702 &  n24882 ;
  assign n25002 = x84 | n24702 ;
  assign n25003 = x84 &  n24702 ;
  assign n25004 = ( n25002 & ~n25003 ) | ( n25002 & 1'b0 ) | ( ~n25003 & 1'b0 ) ;
  assign n25013 = ( n429 & n24864 ) | ( n429 & n25004 ) | ( n24864 & n25004 ) ;
  assign n25014 = ( n24864 & ~n24881 ) | ( n24864 & n25004 ) | ( ~n24881 & n25004 ) ;
  assign n25015 = ~n25013 & n25014 ;
  assign n25016 = n25009 | n25015 ;
  assign n25017 = n24710 &  n24882 ;
  assign n25010 = x83 | n24710 ;
  assign n25011 = x83 &  n24710 ;
  assign n25012 = ( n25010 & ~n25011 ) | ( n25010 & 1'b0 ) | ( ~n25011 & 1'b0 ) ;
  assign n25021 = ( n429 & n24863 ) | ( n429 & n25012 ) | ( n24863 & n25012 ) ;
  assign n25022 = ( n24863 & ~n24881 ) | ( n24863 & n25012 ) | ( ~n24881 & n25012 ) ;
  assign n25023 = ~n25021 & n25022 ;
  assign n25024 = n25017 | n25023 ;
  assign n25025 = n24718 &  n24882 ;
  assign n25018 = x82 | n24718 ;
  assign n25019 = x82 &  n24718 ;
  assign n25020 = ( n25018 & ~n25019 ) | ( n25018 & 1'b0 ) | ( ~n25019 & 1'b0 ) ;
  assign n25029 = ( n429 & n24862 ) | ( n429 & n25020 ) | ( n24862 & n25020 ) ;
  assign n25030 = ( n24862 & ~n24881 ) | ( n24862 & n25020 ) | ( ~n24881 & n25020 ) ;
  assign n25031 = ~n25029 & n25030 ;
  assign n25032 = n25025 | n25031 ;
  assign n25033 = n24726 &  n24882 ;
  assign n25026 = x81 | n24726 ;
  assign n25027 = x81 &  n24726 ;
  assign n25028 = ( n25026 & ~n25027 ) | ( n25026 & 1'b0 ) | ( ~n25027 & 1'b0 ) ;
  assign n25037 = ( n429 & n24861 ) | ( n429 & n25028 ) | ( n24861 & n25028 ) ;
  assign n25038 = ( n24861 & ~n24881 ) | ( n24861 & n25028 ) | ( ~n24881 & n25028 ) ;
  assign n25039 = ~n25037 & n25038 ;
  assign n25040 = n25033 | n25039 ;
  assign n25041 = n24734 &  n24882 ;
  assign n25034 = x80 | n24734 ;
  assign n25035 = x80 &  n24734 ;
  assign n25036 = ( n25034 & ~n25035 ) | ( n25034 & 1'b0 ) | ( ~n25035 & 1'b0 ) ;
  assign n25045 = ( n429 & n24860 ) | ( n429 & n25036 ) | ( n24860 & n25036 ) ;
  assign n25046 = ( n24860 & ~n24881 ) | ( n24860 & n25036 ) | ( ~n24881 & n25036 ) ;
  assign n25047 = ~n25045 & n25046 ;
  assign n25048 = n25041 | n25047 ;
  assign n25049 = n24742 &  n24882 ;
  assign n25042 = x79 | n24742 ;
  assign n25043 = x79 &  n24742 ;
  assign n25044 = ( n25042 & ~n25043 ) | ( n25042 & 1'b0 ) | ( ~n25043 & 1'b0 ) ;
  assign n25053 = ( n429 & n24859 ) | ( n429 & n25044 ) | ( n24859 & n25044 ) ;
  assign n25054 = ( n24859 & ~n24881 ) | ( n24859 & n25044 ) | ( ~n24881 & n25044 ) ;
  assign n25055 = ~n25053 & n25054 ;
  assign n25056 = n25049 | n25055 ;
  assign n25057 = n24750 &  n24882 ;
  assign n25050 = x78 | n24750 ;
  assign n25051 = x78 &  n24750 ;
  assign n25052 = ( n25050 & ~n25051 ) | ( n25050 & 1'b0 ) | ( ~n25051 & 1'b0 ) ;
  assign n25061 = ( n429 & n24858 ) | ( n429 & n25052 ) | ( n24858 & n25052 ) ;
  assign n25062 = ( n24858 & ~n24881 ) | ( n24858 & n25052 ) | ( ~n24881 & n25052 ) ;
  assign n25063 = ~n25061 & n25062 ;
  assign n25064 = n25057 | n25063 ;
  assign n25065 = n24758 &  n24882 ;
  assign n25058 = x77 | n24758 ;
  assign n25059 = x77 &  n24758 ;
  assign n25060 = ( n25058 & ~n25059 ) | ( n25058 & 1'b0 ) | ( ~n25059 & 1'b0 ) ;
  assign n25069 = ( n429 & n24857 ) | ( n429 & n25060 ) | ( n24857 & n25060 ) ;
  assign n25070 = ( n24857 & ~n24881 ) | ( n24857 & n25060 ) | ( ~n24881 & n25060 ) ;
  assign n25071 = ~n25069 & n25070 ;
  assign n25072 = n25065 | n25071 ;
  assign n25073 = n24766 &  n24882 ;
  assign n25066 = x76 | n24766 ;
  assign n25067 = x76 &  n24766 ;
  assign n25068 = ( n25066 & ~n25067 ) | ( n25066 & 1'b0 ) | ( ~n25067 & 1'b0 ) ;
  assign n25077 = ( n429 & n24856 ) | ( n429 & n25068 ) | ( n24856 & n25068 ) ;
  assign n25078 = ( n24856 & ~n24881 ) | ( n24856 & n25068 ) | ( ~n24881 & n25068 ) ;
  assign n25079 = ~n25077 & n25078 ;
  assign n25080 = n25073 | n25079 ;
  assign n25081 = n24774 &  n24882 ;
  assign n25074 = x75 | n24774 ;
  assign n25075 = x75 &  n24774 ;
  assign n25076 = ( n25074 & ~n25075 ) | ( n25074 & 1'b0 ) | ( ~n25075 & 1'b0 ) ;
  assign n25085 = ( n429 & n24855 ) | ( n429 & n25076 ) | ( n24855 & n25076 ) ;
  assign n25086 = ( n24855 & ~n24881 ) | ( n24855 & n25076 ) | ( ~n24881 & n25076 ) ;
  assign n25087 = ~n25085 & n25086 ;
  assign n25088 = n25081 | n25087 ;
  assign n25089 = n24782 &  n24882 ;
  assign n25082 = x74 | n24782 ;
  assign n25083 = x74 &  n24782 ;
  assign n25084 = ( n25082 & ~n25083 ) | ( n25082 & 1'b0 ) | ( ~n25083 & 1'b0 ) ;
  assign n25093 = ( n429 & n24854 ) | ( n429 & n25084 ) | ( n24854 & n25084 ) ;
  assign n25094 = ( n24854 & ~n24881 ) | ( n24854 & n25084 ) | ( ~n24881 & n25084 ) ;
  assign n25095 = ~n25093 & n25094 ;
  assign n25096 = n25089 | n25095 ;
  assign n25097 = n24790 &  n24882 ;
  assign n25090 = x73 | n24790 ;
  assign n25091 = x73 &  n24790 ;
  assign n25092 = ( n25090 & ~n25091 ) | ( n25090 & 1'b0 ) | ( ~n25091 & 1'b0 ) ;
  assign n25101 = ( n429 & n24853 ) | ( n429 & n25092 ) | ( n24853 & n25092 ) ;
  assign n25102 = ( n24853 & ~n24881 ) | ( n24853 & n25092 ) | ( ~n24881 & n25092 ) ;
  assign n25103 = ~n25101 & n25102 ;
  assign n25104 = n25097 | n25103 ;
  assign n25105 = n24798 &  n24882 ;
  assign n25098 = x72 | n24798 ;
  assign n25099 = x72 &  n24798 ;
  assign n25100 = ( n25098 & ~n25099 ) | ( n25098 & 1'b0 ) | ( ~n25099 & 1'b0 ) ;
  assign n25109 = ( n429 & n24852 ) | ( n429 & n25100 ) | ( n24852 & n25100 ) ;
  assign n25110 = ( n24852 & ~n24881 ) | ( n24852 & n25100 ) | ( ~n24881 & n25100 ) ;
  assign n25111 = ~n25109 & n25110 ;
  assign n25112 = n25105 | n25111 ;
  assign n25113 = n24806 &  n24882 ;
  assign n25106 = x71 | n24806 ;
  assign n25107 = x71 &  n24806 ;
  assign n25108 = ( n25106 & ~n25107 ) | ( n25106 & 1'b0 ) | ( ~n25107 & 1'b0 ) ;
  assign n25117 = ( n429 & n24851 ) | ( n429 & n25108 ) | ( n24851 & n25108 ) ;
  assign n25118 = ( n24851 & ~n24881 ) | ( n24851 & n25108 ) | ( ~n24881 & n25108 ) ;
  assign n25119 = ~n25117 & n25118 ;
  assign n25120 = n25113 | n25119 ;
  assign n25121 = n24814 &  n24882 ;
  assign n25114 = x70 | n24814 ;
  assign n25115 = x70 &  n24814 ;
  assign n25116 = ( n25114 & ~n25115 ) | ( n25114 & 1'b0 ) | ( ~n25115 & 1'b0 ) ;
  assign n25125 = ( n429 & n24850 ) | ( n429 & n25116 ) | ( n24850 & n25116 ) ;
  assign n25126 = ( n24850 & ~n24881 ) | ( n24850 & n25116 ) | ( ~n24881 & n25116 ) ;
  assign n25127 = ~n25125 & n25126 ;
  assign n25128 = n25121 | n25127 ;
  assign n25129 = n24822 &  n24882 ;
  assign n25122 = x69 | n24822 ;
  assign n25123 = x69 &  n24822 ;
  assign n25124 = ( n25122 & ~n25123 ) | ( n25122 & 1'b0 ) | ( ~n25123 & 1'b0 ) ;
  assign n25133 = ( n429 & n24849 ) | ( n429 & n25124 ) | ( n24849 & n25124 ) ;
  assign n25134 = ( n24849 & ~n24881 ) | ( n24849 & n25124 ) | ( ~n24881 & n25124 ) ;
  assign n25135 = ~n25133 & n25134 ;
  assign n25136 = n25129 | n25135 ;
  assign n25137 = n24830 &  n24882 ;
  assign n25130 = x68 | n24830 ;
  assign n25131 = x68 &  n24830 ;
  assign n25132 = ( n25130 & ~n25131 ) | ( n25130 & 1'b0 ) | ( ~n25131 & 1'b0 ) ;
  assign n25141 = ( n429 & n24848 ) | ( n429 & n25132 ) | ( n24848 & n25132 ) ;
  assign n25142 = ( n24848 & ~n24881 ) | ( n24848 & n25132 ) | ( ~n24881 & n25132 ) ;
  assign n25143 = ~n25141 & n25142 ;
  assign n25144 = n25137 | n25143 ;
  assign n25145 = n24835 &  n24882 ;
  assign n25138 = x67 | n24835 ;
  assign n25139 = x67 &  n24835 ;
  assign n25140 = ( n25138 & ~n25139 ) | ( n25138 & 1'b0 ) | ( ~n25139 & 1'b0 ) ;
  assign n25149 = ( n429 & n24847 ) | ( n429 & n25140 ) | ( n24847 & n25140 ) ;
  assign n25150 = ( n24847 & ~n24881 ) | ( n24847 & n25140 ) | ( ~n24881 & n25140 ) ;
  assign n25151 = ~n25149 & n25150 ;
  assign n25152 = n25145 | n25151 ;
  assign n25153 = n24841 &  n24882 ;
  assign n25146 = x66 | n24841 ;
  assign n25147 = x66 &  n24841 ;
  assign n25148 = ( n25146 & ~n25147 ) | ( n25146 & 1'b0 ) | ( ~n25147 & 1'b0 ) ;
  assign n25154 = ( n429 & n24846 ) | ( n429 & n25148 ) | ( n24846 & n25148 ) ;
  assign n25155 = ( n24846 & ~n24881 ) | ( n24846 & n25148 ) | ( ~n24881 & n25148 ) ;
  assign n25156 = ~n25154 & n25155 ;
  assign n25157 = n25153 | n25156 ;
  assign n25158 = n24845 &  n24882 ;
  assign n25159 = ( x65 & ~x28 ) | ( x65 & n24842 ) | ( ~x28 & n24842 ) ;
  assign n25160 = ( x28 & ~n24842 ) | ( x28 & x65 ) | ( ~n24842 & x65 ) ;
  assign n25161 = ( n25159 & ~x65 ) | ( n25159 & n25160 ) | ( ~x65 & n25160 ) ;
  assign n25162 = ( n6462 & ~n24881 ) | ( n6462 & n25161 ) | ( ~n24881 & n25161 ) ;
  assign n25163 = ( n429 & n6462 ) | ( n429 & n25161 ) | ( n6462 & n25161 ) ;
  assign n25164 = ( n25162 & ~n25163 ) | ( n25162 & 1'b0 ) | ( ~n25163 & 1'b0 ) ;
  assign n25165 = n25158 | n25164 ;
  assign n25166 = ( n6787 & ~n24881 ) | ( n6787 & 1'b0 ) | ( ~n24881 & 1'b0 ) ;
  assign n25167 = ( x27 & ~n25166 ) | ( x27 & 1'b0 ) | ( ~n25166 & 1'b0 ) ;
  assign n25168 = ( n6792 & ~n24881 ) | ( n6792 & 1'b0 ) | ( ~n24881 & 1'b0 ) ;
  assign n25169 = n25167 | n25168 ;
  assign n25170 = ( x65 & ~n25169 ) | ( x65 & n6795 ) | ( ~n25169 & n6795 ) ;
  assign n25171 = ( x66 & ~n25165 ) | ( x66 & n25170 ) | ( ~n25165 & n25170 ) ;
  assign n25172 = ( x67 & ~n25157 ) | ( x67 & n25171 ) | ( ~n25157 & n25171 ) ;
  assign n25173 = ( x68 & ~n25152 ) | ( x68 & n25172 ) | ( ~n25152 & n25172 ) ;
  assign n25174 = ( x69 & ~n25144 ) | ( x69 & n25173 ) | ( ~n25144 & n25173 ) ;
  assign n25175 = ( x70 & ~n25136 ) | ( x70 & n25174 ) | ( ~n25136 & n25174 ) ;
  assign n25176 = ( x71 & ~n25128 ) | ( x71 & n25175 ) | ( ~n25128 & n25175 ) ;
  assign n25177 = ( x72 & ~n25120 ) | ( x72 & n25176 ) | ( ~n25120 & n25176 ) ;
  assign n25178 = ( x73 & ~n25112 ) | ( x73 & n25177 ) | ( ~n25112 & n25177 ) ;
  assign n25179 = ( x74 & ~n25104 ) | ( x74 & n25178 ) | ( ~n25104 & n25178 ) ;
  assign n25180 = ( x75 & ~n25096 ) | ( x75 & n25179 ) | ( ~n25096 & n25179 ) ;
  assign n25181 = ( x76 & ~n25088 ) | ( x76 & n25180 ) | ( ~n25088 & n25180 ) ;
  assign n25182 = ( x77 & ~n25080 ) | ( x77 & n25181 ) | ( ~n25080 & n25181 ) ;
  assign n25183 = ( x78 & ~n25072 ) | ( x78 & n25182 ) | ( ~n25072 & n25182 ) ;
  assign n25184 = ( x79 & ~n25064 ) | ( x79 & n25183 ) | ( ~n25064 & n25183 ) ;
  assign n25185 = ( x80 & ~n25056 ) | ( x80 & n25184 ) | ( ~n25056 & n25184 ) ;
  assign n25186 = ( x81 & ~n25048 ) | ( x81 & n25185 ) | ( ~n25048 & n25185 ) ;
  assign n25187 = ( x82 & ~n25040 ) | ( x82 & n25186 ) | ( ~n25040 & n25186 ) ;
  assign n25188 = ( x83 & ~n25032 ) | ( x83 & n25187 ) | ( ~n25032 & n25187 ) ;
  assign n25189 = ( x84 & ~n25024 ) | ( x84 & n25188 ) | ( ~n25024 & n25188 ) ;
  assign n25190 = ( x85 & ~n25016 ) | ( x85 & n25189 ) | ( ~n25016 & n25189 ) ;
  assign n25191 = ( x86 & ~n25008 ) | ( x86 & n25190 ) | ( ~n25008 & n25190 ) ;
  assign n25192 = ( x87 & ~n25000 ) | ( x87 & n25191 ) | ( ~n25000 & n25191 ) ;
  assign n25193 = ( x88 & ~n24992 ) | ( x88 & n25192 ) | ( ~n24992 & n25192 ) ;
  assign n25194 = ( x89 & ~n24984 ) | ( x89 & n25193 ) | ( ~n24984 & n25193 ) ;
  assign n25195 = ( x90 & ~n24976 ) | ( x90 & n25194 ) | ( ~n24976 & n25194 ) ;
  assign n25196 = ( x91 & ~n24968 ) | ( x91 & n25195 ) | ( ~n24968 & n25195 ) ;
  assign n25197 = ( x92 & ~n24960 ) | ( x92 & n25196 ) | ( ~n24960 & n25196 ) ;
  assign n25198 = ( x93 & ~n24952 ) | ( x93 & n25197 ) | ( ~n24952 & n25197 ) ;
  assign n25199 = ( x94 & ~n24944 ) | ( x94 & n25198 ) | ( ~n24944 & n25198 ) ;
  assign n25200 = ( x95 & ~n24936 ) | ( x95 & n25199 ) | ( ~n24936 & n25199 ) ;
  assign n25201 = ( x96 & ~n24928 ) | ( x96 & n25200 ) | ( ~n24928 & n25200 ) ;
  assign n25202 = ( x97 & ~n24920 ) | ( x97 & n25201 ) | ( ~n24920 & n25201 ) ;
  assign n25203 = ( x98 & ~n24912 ) | ( x98 & n25202 ) | ( ~n24912 & n25202 ) ;
  assign n25204 = ( x99 & ~n24904 ) | ( x99 & n25203 ) | ( ~n24904 & n25203 ) ;
  assign n25205 = ( x100 & ~n24896 ) | ( x100 & n25204 ) | ( ~n24896 & n25204 ) ;
  assign n25206 = ( x101 & ~n24888 ) | ( x101 & n25205 ) | ( ~n24888 & n25205 ) ;
  assign n25207 = n6835 | n25206 ;
  assign n25208 = n24888 &  n25207 ;
  assign n25212 = ( n6835 & n24888 ) | ( n6835 & n25205 ) | ( n24888 & n25205 ) ;
  assign n25213 = ( x101 & ~n25212 ) | ( x101 & n24888 ) | ( ~n25212 & n24888 ) ;
  assign n25214 = ~x101 & n25213 ;
  assign n25215 = n25208 | n25214 ;
  assign n25216 = ~x102 & n25215 ;
  assign n25217 = n24896 &  n25207 ;
  assign n25209 = x100 | n24896 ;
  assign n25210 = x100 &  n24896 ;
  assign n25211 = ( n25209 & ~n25210 ) | ( n25209 & 1'b0 ) | ( ~n25210 & 1'b0 ) ;
  assign n25221 = ( n6835 & n25204 ) | ( n6835 & n25211 ) | ( n25204 & n25211 ) ;
  assign n25222 = ( n25204 & ~n25206 ) | ( n25204 & n25211 ) | ( ~n25206 & n25211 ) ;
  assign n25223 = ~n25221 & n25222 ;
  assign n25224 = n25217 | n25223 ;
  assign n25225 = n24904 &  n25207 ;
  assign n25218 = x99 | n24904 ;
  assign n25219 = x99 &  n24904 ;
  assign n25220 = ( n25218 & ~n25219 ) | ( n25218 & 1'b0 ) | ( ~n25219 & 1'b0 ) ;
  assign n25229 = ( n6835 & n25203 ) | ( n6835 & n25220 ) | ( n25203 & n25220 ) ;
  assign n25230 = ( n25203 & ~n25206 ) | ( n25203 & n25220 ) | ( ~n25206 & n25220 ) ;
  assign n25231 = ~n25229 & n25230 ;
  assign n25232 = n25225 | n25231 ;
  assign n25233 = n24912 &  n25207 ;
  assign n25226 = x98 | n24912 ;
  assign n25227 = x98 &  n24912 ;
  assign n25228 = ( n25226 & ~n25227 ) | ( n25226 & 1'b0 ) | ( ~n25227 & 1'b0 ) ;
  assign n25237 = ( n6835 & n25202 ) | ( n6835 & n25228 ) | ( n25202 & n25228 ) ;
  assign n25238 = ( n25202 & ~n25206 ) | ( n25202 & n25228 ) | ( ~n25206 & n25228 ) ;
  assign n25239 = ~n25237 & n25238 ;
  assign n25240 = n25233 | n25239 ;
  assign n25241 = n24920 &  n25207 ;
  assign n25234 = x97 | n24920 ;
  assign n25235 = x97 &  n24920 ;
  assign n25236 = ( n25234 & ~n25235 ) | ( n25234 & 1'b0 ) | ( ~n25235 & 1'b0 ) ;
  assign n25245 = ( n6835 & n25201 ) | ( n6835 & n25236 ) | ( n25201 & n25236 ) ;
  assign n25246 = ( n25201 & ~n25206 ) | ( n25201 & n25236 ) | ( ~n25206 & n25236 ) ;
  assign n25247 = ~n25245 & n25246 ;
  assign n25248 = n25241 | n25247 ;
  assign n25249 = n24928 &  n25207 ;
  assign n25242 = x96 | n24928 ;
  assign n25243 = x96 &  n24928 ;
  assign n25244 = ( n25242 & ~n25243 ) | ( n25242 & 1'b0 ) | ( ~n25243 & 1'b0 ) ;
  assign n25253 = ( n6835 & n25200 ) | ( n6835 & n25244 ) | ( n25200 & n25244 ) ;
  assign n25254 = ( n25200 & ~n25206 ) | ( n25200 & n25244 ) | ( ~n25206 & n25244 ) ;
  assign n25255 = ~n25253 & n25254 ;
  assign n25256 = n25249 | n25255 ;
  assign n25257 = n24936 &  n25207 ;
  assign n25250 = x95 | n24936 ;
  assign n25251 = x95 &  n24936 ;
  assign n25252 = ( n25250 & ~n25251 ) | ( n25250 & 1'b0 ) | ( ~n25251 & 1'b0 ) ;
  assign n25261 = ( n6835 & n25199 ) | ( n6835 & n25252 ) | ( n25199 & n25252 ) ;
  assign n25262 = ( n25199 & ~n25206 ) | ( n25199 & n25252 ) | ( ~n25206 & n25252 ) ;
  assign n25263 = ~n25261 & n25262 ;
  assign n25264 = n25257 | n25263 ;
  assign n25265 = n24944 &  n25207 ;
  assign n25258 = x94 | n24944 ;
  assign n25259 = x94 &  n24944 ;
  assign n25260 = ( n25258 & ~n25259 ) | ( n25258 & 1'b0 ) | ( ~n25259 & 1'b0 ) ;
  assign n25269 = ( n6835 & n25198 ) | ( n6835 & n25260 ) | ( n25198 & n25260 ) ;
  assign n25270 = ( n25198 & ~n25206 ) | ( n25198 & n25260 ) | ( ~n25206 & n25260 ) ;
  assign n25271 = ~n25269 & n25270 ;
  assign n25272 = n25265 | n25271 ;
  assign n25273 = n24952 &  n25207 ;
  assign n25266 = x93 | n24952 ;
  assign n25267 = x93 &  n24952 ;
  assign n25268 = ( n25266 & ~n25267 ) | ( n25266 & 1'b0 ) | ( ~n25267 & 1'b0 ) ;
  assign n25277 = ( n6835 & n25197 ) | ( n6835 & n25268 ) | ( n25197 & n25268 ) ;
  assign n25278 = ( n25197 & ~n25206 ) | ( n25197 & n25268 ) | ( ~n25206 & n25268 ) ;
  assign n25279 = ~n25277 & n25278 ;
  assign n25280 = n25273 | n25279 ;
  assign n25281 = n24960 &  n25207 ;
  assign n25274 = x92 | n24960 ;
  assign n25275 = x92 &  n24960 ;
  assign n25276 = ( n25274 & ~n25275 ) | ( n25274 & 1'b0 ) | ( ~n25275 & 1'b0 ) ;
  assign n25285 = ( n6835 & n25196 ) | ( n6835 & n25276 ) | ( n25196 & n25276 ) ;
  assign n25286 = ( n25196 & ~n25206 ) | ( n25196 & n25276 ) | ( ~n25206 & n25276 ) ;
  assign n25287 = ~n25285 & n25286 ;
  assign n25288 = n25281 | n25287 ;
  assign n25289 = n24968 &  n25207 ;
  assign n25282 = x91 | n24968 ;
  assign n25283 = x91 &  n24968 ;
  assign n25284 = ( n25282 & ~n25283 ) | ( n25282 & 1'b0 ) | ( ~n25283 & 1'b0 ) ;
  assign n25293 = ( n6835 & n25195 ) | ( n6835 & n25284 ) | ( n25195 & n25284 ) ;
  assign n25294 = ( n25195 & ~n25206 ) | ( n25195 & n25284 ) | ( ~n25206 & n25284 ) ;
  assign n25295 = ~n25293 & n25294 ;
  assign n25296 = n25289 | n25295 ;
  assign n25297 = n24976 &  n25207 ;
  assign n25290 = x90 | n24976 ;
  assign n25291 = x90 &  n24976 ;
  assign n25292 = ( n25290 & ~n25291 ) | ( n25290 & 1'b0 ) | ( ~n25291 & 1'b0 ) ;
  assign n25301 = ( n6835 & n25194 ) | ( n6835 & n25292 ) | ( n25194 & n25292 ) ;
  assign n25302 = ( n25194 & ~n25206 ) | ( n25194 & n25292 ) | ( ~n25206 & n25292 ) ;
  assign n25303 = ~n25301 & n25302 ;
  assign n25304 = n25297 | n25303 ;
  assign n25305 = n24984 &  n25207 ;
  assign n25298 = x89 | n24984 ;
  assign n25299 = x89 &  n24984 ;
  assign n25300 = ( n25298 & ~n25299 ) | ( n25298 & 1'b0 ) | ( ~n25299 & 1'b0 ) ;
  assign n25309 = ( n6835 & n25193 ) | ( n6835 & n25300 ) | ( n25193 & n25300 ) ;
  assign n25310 = ( n25193 & ~n25206 ) | ( n25193 & n25300 ) | ( ~n25206 & n25300 ) ;
  assign n25311 = ~n25309 & n25310 ;
  assign n25312 = n25305 | n25311 ;
  assign n25313 = n24992 &  n25207 ;
  assign n25306 = x88 | n24992 ;
  assign n25307 = x88 &  n24992 ;
  assign n25308 = ( n25306 & ~n25307 ) | ( n25306 & 1'b0 ) | ( ~n25307 & 1'b0 ) ;
  assign n25317 = ( n6835 & n25192 ) | ( n6835 & n25308 ) | ( n25192 & n25308 ) ;
  assign n25318 = ( n25192 & ~n25206 ) | ( n25192 & n25308 ) | ( ~n25206 & n25308 ) ;
  assign n25319 = ~n25317 & n25318 ;
  assign n25320 = n25313 | n25319 ;
  assign n25321 = n25000 &  n25207 ;
  assign n25314 = x87 | n25000 ;
  assign n25315 = x87 &  n25000 ;
  assign n25316 = ( n25314 & ~n25315 ) | ( n25314 & 1'b0 ) | ( ~n25315 & 1'b0 ) ;
  assign n25325 = ( n6835 & n25191 ) | ( n6835 & n25316 ) | ( n25191 & n25316 ) ;
  assign n25326 = ( n25191 & ~n25206 ) | ( n25191 & n25316 ) | ( ~n25206 & n25316 ) ;
  assign n25327 = ~n25325 & n25326 ;
  assign n25328 = n25321 | n25327 ;
  assign n25329 = n25008 &  n25207 ;
  assign n25322 = x86 | n25008 ;
  assign n25323 = x86 &  n25008 ;
  assign n25324 = ( n25322 & ~n25323 ) | ( n25322 & 1'b0 ) | ( ~n25323 & 1'b0 ) ;
  assign n25333 = ( n6835 & n25190 ) | ( n6835 & n25324 ) | ( n25190 & n25324 ) ;
  assign n25334 = ( n25190 & ~n25206 ) | ( n25190 & n25324 ) | ( ~n25206 & n25324 ) ;
  assign n25335 = ~n25333 & n25334 ;
  assign n25336 = n25329 | n25335 ;
  assign n25337 = n25016 &  n25207 ;
  assign n25330 = x85 | n25016 ;
  assign n25331 = x85 &  n25016 ;
  assign n25332 = ( n25330 & ~n25331 ) | ( n25330 & 1'b0 ) | ( ~n25331 & 1'b0 ) ;
  assign n25341 = ( n6835 & n25189 ) | ( n6835 & n25332 ) | ( n25189 & n25332 ) ;
  assign n25342 = ( n25189 & ~n25206 ) | ( n25189 & n25332 ) | ( ~n25206 & n25332 ) ;
  assign n25343 = ~n25341 & n25342 ;
  assign n25344 = n25337 | n25343 ;
  assign n25345 = n25024 &  n25207 ;
  assign n25338 = x84 | n25024 ;
  assign n25339 = x84 &  n25024 ;
  assign n25340 = ( n25338 & ~n25339 ) | ( n25338 & 1'b0 ) | ( ~n25339 & 1'b0 ) ;
  assign n25349 = ( n6835 & n25188 ) | ( n6835 & n25340 ) | ( n25188 & n25340 ) ;
  assign n25350 = ( n25188 & ~n25206 ) | ( n25188 & n25340 ) | ( ~n25206 & n25340 ) ;
  assign n25351 = ~n25349 & n25350 ;
  assign n25352 = n25345 | n25351 ;
  assign n25353 = n25032 &  n25207 ;
  assign n25346 = x83 | n25032 ;
  assign n25347 = x83 &  n25032 ;
  assign n25348 = ( n25346 & ~n25347 ) | ( n25346 & 1'b0 ) | ( ~n25347 & 1'b0 ) ;
  assign n25357 = ( n6835 & n25187 ) | ( n6835 & n25348 ) | ( n25187 & n25348 ) ;
  assign n25358 = ( n25187 & ~n25206 ) | ( n25187 & n25348 ) | ( ~n25206 & n25348 ) ;
  assign n25359 = ~n25357 & n25358 ;
  assign n25360 = n25353 | n25359 ;
  assign n25361 = n25040 &  n25207 ;
  assign n25354 = x82 | n25040 ;
  assign n25355 = x82 &  n25040 ;
  assign n25356 = ( n25354 & ~n25355 ) | ( n25354 & 1'b0 ) | ( ~n25355 & 1'b0 ) ;
  assign n25365 = ( n6835 & n25186 ) | ( n6835 & n25356 ) | ( n25186 & n25356 ) ;
  assign n25366 = ( n25186 & ~n25206 ) | ( n25186 & n25356 ) | ( ~n25206 & n25356 ) ;
  assign n25367 = ~n25365 & n25366 ;
  assign n25368 = n25361 | n25367 ;
  assign n25369 = n25048 &  n25207 ;
  assign n25362 = x81 | n25048 ;
  assign n25363 = x81 &  n25048 ;
  assign n25364 = ( n25362 & ~n25363 ) | ( n25362 & 1'b0 ) | ( ~n25363 & 1'b0 ) ;
  assign n25373 = ( n6835 & n25185 ) | ( n6835 & n25364 ) | ( n25185 & n25364 ) ;
  assign n25374 = ( n25185 & ~n25206 ) | ( n25185 & n25364 ) | ( ~n25206 & n25364 ) ;
  assign n25375 = ~n25373 & n25374 ;
  assign n25376 = n25369 | n25375 ;
  assign n25377 = n25056 &  n25207 ;
  assign n25370 = x80 | n25056 ;
  assign n25371 = x80 &  n25056 ;
  assign n25372 = ( n25370 & ~n25371 ) | ( n25370 & 1'b0 ) | ( ~n25371 & 1'b0 ) ;
  assign n25381 = ( n6835 & n25184 ) | ( n6835 & n25372 ) | ( n25184 & n25372 ) ;
  assign n25382 = ( n25184 & ~n25206 ) | ( n25184 & n25372 ) | ( ~n25206 & n25372 ) ;
  assign n25383 = ~n25381 & n25382 ;
  assign n25384 = n25377 | n25383 ;
  assign n25385 = n25064 &  n25207 ;
  assign n25378 = x79 | n25064 ;
  assign n25379 = x79 &  n25064 ;
  assign n25380 = ( n25378 & ~n25379 ) | ( n25378 & 1'b0 ) | ( ~n25379 & 1'b0 ) ;
  assign n25389 = ( n6835 & n25183 ) | ( n6835 & n25380 ) | ( n25183 & n25380 ) ;
  assign n25390 = ( n25183 & ~n25206 ) | ( n25183 & n25380 ) | ( ~n25206 & n25380 ) ;
  assign n25391 = ~n25389 & n25390 ;
  assign n25392 = n25385 | n25391 ;
  assign n25393 = n25072 &  n25207 ;
  assign n25386 = x78 | n25072 ;
  assign n25387 = x78 &  n25072 ;
  assign n25388 = ( n25386 & ~n25387 ) | ( n25386 & 1'b0 ) | ( ~n25387 & 1'b0 ) ;
  assign n25397 = ( n6835 & n25182 ) | ( n6835 & n25388 ) | ( n25182 & n25388 ) ;
  assign n25398 = ( n25182 & ~n25206 ) | ( n25182 & n25388 ) | ( ~n25206 & n25388 ) ;
  assign n25399 = ~n25397 & n25398 ;
  assign n25400 = n25393 | n25399 ;
  assign n25401 = n25080 &  n25207 ;
  assign n25394 = x77 | n25080 ;
  assign n25395 = x77 &  n25080 ;
  assign n25396 = ( n25394 & ~n25395 ) | ( n25394 & 1'b0 ) | ( ~n25395 & 1'b0 ) ;
  assign n25405 = ( n6835 & n25181 ) | ( n6835 & n25396 ) | ( n25181 & n25396 ) ;
  assign n25406 = ( n25181 & ~n25206 ) | ( n25181 & n25396 ) | ( ~n25206 & n25396 ) ;
  assign n25407 = ~n25405 & n25406 ;
  assign n25408 = n25401 | n25407 ;
  assign n25409 = n25088 &  n25207 ;
  assign n25402 = x76 | n25088 ;
  assign n25403 = x76 &  n25088 ;
  assign n25404 = ( n25402 & ~n25403 ) | ( n25402 & 1'b0 ) | ( ~n25403 & 1'b0 ) ;
  assign n25413 = ( n6835 & n25180 ) | ( n6835 & n25404 ) | ( n25180 & n25404 ) ;
  assign n25414 = ( n25180 & ~n25206 ) | ( n25180 & n25404 ) | ( ~n25206 & n25404 ) ;
  assign n25415 = ~n25413 & n25414 ;
  assign n25416 = n25409 | n25415 ;
  assign n25417 = n25096 &  n25207 ;
  assign n25410 = x75 | n25096 ;
  assign n25411 = x75 &  n25096 ;
  assign n25412 = ( n25410 & ~n25411 ) | ( n25410 & 1'b0 ) | ( ~n25411 & 1'b0 ) ;
  assign n25421 = ( n6835 & n25179 ) | ( n6835 & n25412 ) | ( n25179 & n25412 ) ;
  assign n25422 = ( n25179 & ~n25206 ) | ( n25179 & n25412 ) | ( ~n25206 & n25412 ) ;
  assign n25423 = ~n25421 & n25422 ;
  assign n25424 = n25417 | n25423 ;
  assign n25425 = n25104 &  n25207 ;
  assign n25418 = x74 | n25104 ;
  assign n25419 = x74 &  n25104 ;
  assign n25420 = ( n25418 & ~n25419 ) | ( n25418 & 1'b0 ) | ( ~n25419 & 1'b0 ) ;
  assign n25429 = ( n6835 & n25178 ) | ( n6835 & n25420 ) | ( n25178 & n25420 ) ;
  assign n25430 = ( n25178 & ~n25206 ) | ( n25178 & n25420 ) | ( ~n25206 & n25420 ) ;
  assign n25431 = ~n25429 & n25430 ;
  assign n25432 = n25425 | n25431 ;
  assign n25433 = n25112 &  n25207 ;
  assign n25426 = x73 | n25112 ;
  assign n25427 = x73 &  n25112 ;
  assign n25428 = ( n25426 & ~n25427 ) | ( n25426 & 1'b0 ) | ( ~n25427 & 1'b0 ) ;
  assign n25437 = ( n6835 & n25177 ) | ( n6835 & n25428 ) | ( n25177 & n25428 ) ;
  assign n25438 = ( n25177 & ~n25206 ) | ( n25177 & n25428 ) | ( ~n25206 & n25428 ) ;
  assign n25439 = ~n25437 & n25438 ;
  assign n25440 = n25433 | n25439 ;
  assign n25441 = n25120 &  n25207 ;
  assign n25434 = x72 | n25120 ;
  assign n25435 = x72 &  n25120 ;
  assign n25436 = ( n25434 & ~n25435 ) | ( n25434 & 1'b0 ) | ( ~n25435 & 1'b0 ) ;
  assign n25445 = ( n6835 & n25176 ) | ( n6835 & n25436 ) | ( n25176 & n25436 ) ;
  assign n25446 = ( n25176 & ~n25206 ) | ( n25176 & n25436 ) | ( ~n25206 & n25436 ) ;
  assign n25447 = ~n25445 & n25446 ;
  assign n25448 = n25441 | n25447 ;
  assign n25449 = n25128 &  n25207 ;
  assign n25442 = x71 | n25128 ;
  assign n25443 = x71 &  n25128 ;
  assign n25444 = ( n25442 & ~n25443 ) | ( n25442 & 1'b0 ) | ( ~n25443 & 1'b0 ) ;
  assign n25453 = ( n6835 & n25175 ) | ( n6835 & n25444 ) | ( n25175 & n25444 ) ;
  assign n25454 = ( n25175 & ~n25206 ) | ( n25175 & n25444 ) | ( ~n25206 & n25444 ) ;
  assign n25455 = ~n25453 & n25454 ;
  assign n25456 = n25449 | n25455 ;
  assign n25457 = n25136 &  n25207 ;
  assign n25450 = x70 | n25136 ;
  assign n25451 = x70 &  n25136 ;
  assign n25452 = ( n25450 & ~n25451 ) | ( n25450 & 1'b0 ) | ( ~n25451 & 1'b0 ) ;
  assign n25461 = ( n6835 & n25174 ) | ( n6835 & n25452 ) | ( n25174 & n25452 ) ;
  assign n25462 = ( n25174 & ~n25206 ) | ( n25174 & n25452 ) | ( ~n25206 & n25452 ) ;
  assign n25463 = ~n25461 & n25462 ;
  assign n25464 = n25457 | n25463 ;
  assign n25465 = n25144 &  n25207 ;
  assign n25458 = x69 | n25144 ;
  assign n25459 = x69 &  n25144 ;
  assign n25460 = ( n25458 & ~n25459 ) | ( n25458 & 1'b0 ) | ( ~n25459 & 1'b0 ) ;
  assign n25469 = ( n6835 & n25173 ) | ( n6835 & n25460 ) | ( n25173 & n25460 ) ;
  assign n25470 = ( n25173 & ~n25206 ) | ( n25173 & n25460 ) | ( ~n25206 & n25460 ) ;
  assign n25471 = ~n25469 & n25470 ;
  assign n25472 = n25465 | n25471 ;
  assign n25473 = n25152 &  n25207 ;
  assign n25466 = x68 | n25152 ;
  assign n25467 = x68 &  n25152 ;
  assign n25468 = ( n25466 & ~n25467 ) | ( n25466 & 1'b0 ) | ( ~n25467 & 1'b0 ) ;
  assign n25477 = ( n6835 & n25172 ) | ( n6835 & n25468 ) | ( n25172 & n25468 ) ;
  assign n25478 = ( n25172 & ~n25206 ) | ( n25172 & n25468 ) | ( ~n25206 & n25468 ) ;
  assign n25479 = ~n25477 & n25478 ;
  assign n25480 = n25473 | n25479 ;
  assign n25481 = n25157 &  n25207 ;
  assign n25474 = x67 | n25157 ;
  assign n25475 = x67 &  n25157 ;
  assign n25476 = ( n25474 & ~n25475 ) | ( n25474 & 1'b0 ) | ( ~n25475 & 1'b0 ) ;
  assign n25485 = ( n6835 & n25171 ) | ( n6835 & n25476 ) | ( n25171 & n25476 ) ;
  assign n25486 = ( n25171 & ~n25206 ) | ( n25171 & n25476 ) | ( ~n25206 & n25476 ) ;
  assign n25487 = ~n25485 & n25486 ;
  assign n25488 = n25481 | n25487 ;
  assign n25489 = n25165 &  n25207 ;
  assign n25482 = x66 | n25165 ;
  assign n25483 = x66 &  n25165 ;
  assign n25484 = ( n25482 & ~n25483 ) | ( n25482 & 1'b0 ) | ( ~n25483 & 1'b0 ) ;
  assign n25493 = ( n6835 & n25170 ) | ( n6835 & n25484 ) | ( n25170 & n25484 ) ;
  assign n25494 = ( n25170 & ~n25206 ) | ( n25170 & n25484 ) | ( ~n25206 & n25484 ) ;
  assign n25495 = ~n25493 & n25494 ;
  assign n25496 = n25489 | n25495 ;
  assign n25497 = n25169 &  n25207 ;
  assign n25490 = x65 &  n25169 ;
  assign n25491 = x65 | n25168 ;
  assign n25492 = n25167 | n25491 ;
  assign n25498 = ~n25490 & n25492 ;
  assign n25499 = ( n6795 & ~n6835 ) | ( n6795 & n25498 ) | ( ~n6835 & n25498 ) ;
  assign n25500 = ( n6795 & n25206 ) | ( n6795 & n25498 ) | ( n25206 & n25498 ) ;
  assign n25501 = ( n25499 & ~n25500 ) | ( n25499 & 1'b0 ) | ( ~n25500 & 1'b0 ) ;
  assign n25502 = n25497 | n25501 ;
  assign n25503 = ( n7003 & ~n25206 ) | ( n7003 & 1'b0 ) | ( ~n25206 & 1'b0 ) ;
  assign n25504 = ( x26 & ~n25503 ) | ( x26 & 1'b0 ) | ( ~n25503 & 1'b0 ) ;
  assign n25505 = ( n7009 & ~n25206 ) | ( n7009 & 1'b0 ) | ( ~n25206 & 1'b0 ) ;
  assign n25506 = n25504 | n25505 ;
  assign n25507 = ( x65 & ~n25506 ) | ( x65 & n7012 ) | ( ~n25506 & n7012 ) ;
  assign n25508 = ( x66 & ~n25502 ) | ( x66 & n25507 ) | ( ~n25502 & n25507 ) ;
  assign n25509 = ( x67 & ~n25496 ) | ( x67 & n25508 ) | ( ~n25496 & n25508 ) ;
  assign n25510 = ( x68 & ~n25488 ) | ( x68 & n25509 ) | ( ~n25488 & n25509 ) ;
  assign n25511 = ( x69 & ~n25480 ) | ( x69 & n25510 ) | ( ~n25480 & n25510 ) ;
  assign n25512 = ( x70 & ~n25472 ) | ( x70 & n25511 ) | ( ~n25472 & n25511 ) ;
  assign n25513 = ( x71 & ~n25464 ) | ( x71 & n25512 ) | ( ~n25464 & n25512 ) ;
  assign n25514 = ( x72 & ~n25456 ) | ( x72 & n25513 ) | ( ~n25456 & n25513 ) ;
  assign n25515 = ( x73 & ~n25448 ) | ( x73 & n25514 ) | ( ~n25448 & n25514 ) ;
  assign n25516 = ( x74 & ~n25440 ) | ( x74 & n25515 ) | ( ~n25440 & n25515 ) ;
  assign n25517 = ( x75 & ~n25432 ) | ( x75 & n25516 ) | ( ~n25432 & n25516 ) ;
  assign n25518 = ( x76 & ~n25424 ) | ( x76 & n25517 ) | ( ~n25424 & n25517 ) ;
  assign n25519 = ( x77 & ~n25416 ) | ( x77 & n25518 ) | ( ~n25416 & n25518 ) ;
  assign n25520 = ( x78 & ~n25408 ) | ( x78 & n25519 ) | ( ~n25408 & n25519 ) ;
  assign n25521 = ( x79 & ~n25400 ) | ( x79 & n25520 ) | ( ~n25400 & n25520 ) ;
  assign n25522 = ( x80 & ~n25392 ) | ( x80 & n25521 ) | ( ~n25392 & n25521 ) ;
  assign n25523 = ( x81 & ~n25384 ) | ( x81 & n25522 ) | ( ~n25384 & n25522 ) ;
  assign n25524 = ( x82 & ~n25376 ) | ( x82 & n25523 ) | ( ~n25376 & n25523 ) ;
  assign n25525 = ( x83 & ~n25368 ) | ( x83 & n25524 ) | ( ~n25368 & n25524 ) ;
  assign n25526 = ( x84 & ~n25360 ) | ( x84 & n25525 ) | ( ~n25360 & n25525 ) ;
  assign n25527 = ( x85 & ~n25352 ) | ( x85 & n25526 ) | ( ~n25352 & n25526 ) ;
  assign n25528 = ( x86 & ~n25344 ) | ( x86 & n25527 ) | ( ~n25344 & n25527 ) ;
  assign n25529 = ( x87 & ~n25336 ) | ( x87 & n25528 ) | ( ~n25336 & n25528 ) ;
  assign n25530 = ( x88 & ~n25328 ) | ( x88 & n25529 ) | ( ~n25328 & n25529 ) ;
  assign n25531 = ( x89 & ~n25320 ) | ( x89 & n25530 ) | ( ~n25320 & n25530 ) ;
  assign n25532 = ( x90 & ~n25312 ) | ( x90 & n25531 ) | ( ~n25312 & n25531 ) ;
  assign n25533 = ( x91 & ~n25304 ) | ( x91 & n25532 ) | ( ~n25304 & n25532 ) ;
  assign n25534 = ( x92 & ~n25296 ) | ( x92 & n25533 ) | ( ~n25296 & n25533 ) ;
  assign n25535 = ( x93 & ~n25288 ) | ( x93 & n25534 ) | ( ~n25288 & n25534 ) ;
  assign n25536 = ( x94 & ~n25280 ) | ( x94 & n25535 ) | ( ~n25280 & n25535 ) ;
  assign n25537 = ( x95 & ~n25272 ) | ( x95 & n25536 ) | ( ~n25272 & n25536 ) ;
  assign n25538 = ( x96 & ~n25264 ) | ( x96 & n25537 ) | ( ~n25264 & n25537 ) ;
  assign n25539 = ( x97 & ~n25256 ) | ( x97 & n25538 ) | ( ~n25256 & n25538 ) ;
  assign n25540 = ( x98 & ~n25248 ) | ( x98 & n25539 ) | ( ~n25248 & n25539 ) ;
  assign n25541 = ( x99 & ~n25240 ) | ( x99 & n25540 ) | ( ~n25240 & n25540 ) ;
  assign n25542 = ( x100 & ~n25232 ) | ( x100 & n25541 ) | ( ~n25232 & n25541 ) ;
  assign n25543 = ( x101 & ~n25224 ) | ( x101 & n25542 ) | ( ~n25224 & n25542 ) ;
  assign n25544 = ( x102 & ~n25208 ) | ( x102 & 1'b0 ) | ( ~n25208 & 1'b0 ) ;
  assign n25545 = ~n25214 & n25544 ;
  assign n25546 = ( n25543 & ~n25216 ) | ( n25543 & n25545 ) | ( ~n25216 & n25545 ) ;
  assign n25547 = ( n25216 & ~n7189 ) | ( n25216 & n25546 ) | ( ~n7189 & n25546 ) ;
  assign n25548 = n7189 | n25547 ;
  assign n25555 = n6835 &  n24888 ;
  assign n25556 = n25548 &  n25555 ;
  assign n25549 = ~n25215 |  n6835 ;
  assign n25550 = n25548 &  n25549 ;
  assign n25554 = n25216 | n25545 ;
  assign n25558 = ( n25543 & n25550 ) | ( n25543 & n25554 ) | ( n25550 & n25554 ) ;
  assign n25557 = n25543 | n25554 ;
  assign n25559 = ( n25556 & ~n25558 ) | ( n25556 & n25557 ) | ( ~n25558 & n25557 ) ;
  assign n25563 = n25224 &  n25549 ;
  assign n25564 = n25548 &  n25563 ;
  assign n25551 = x101 | n25224 ;
  assign n25552 = x101 &  n25224 ;
  assign n25553 = ( n25551 & ~n25552 ) | ( n25551 & 1'b0 ) | ( ~n25552 & 1'b0 ) ;
  assign n25566 = ( n25542 & n25550 ) | ( n25542 & n25553 ) | ( n25550 & n25553 ) ;
  assign n25565 = n25542 | n25553 ;
  assign n25567 = ( n25564 & ~n25566 ) | ( n25564 & n25565 ) | ( ~n25566 & n25565 ) ;
  assign n25571 = n25232 &  n25549 ;
  assign n25572 = n25548 &  n25571 ;
  assign n25560 = x100 | n25232 ;
  assign n25561 = x100 &  n25232 ;
  assign n25562 = ( n25560 & ~n25561 ) | ( n25560 & 1'b0 ) | ( ~n25561 & 1'b0 ) ;
  assign n25574 = ( n25541 & n25550 ) | ( n25541 & n25562 ) | ( n25550 & n25562 ) ;
  assign n25573 = n25541 | n25562 ;
  assign n25575 = ( n25572 & ~n25574 ) | ( n25572 & n25573 ) | ( ~n25574 & n25573 ) ;
  assign n25579 = n25240 &  n25549 ;
  assign n25580 = n25548 &  n25579 ;
  assign n25568 = x99 | n25240 ;
  assign n25569 = x99 &  n25240 ;
  assign n25570 = ( n25568 & ~n25569 ) | ( n25568 & 1'b0 ) | ( ~n25569 & 1'b0 ) ;
  assign n25582 = ( n25540 & n25550 ) | ( n25540 & n25570 ) | ( n25550 & n25570 ) ;
  assign n25581 = n25540 | n25570 ;
  assign n25583 = ( n25580 & ~n25582 ) | ( n25580 & n25581 ) | ( ~n25582 & n25581 ) ;
  assign n25587 = n25248 &  n25549 ;
  assign n25588 = n25548 &  n25587 ;
  assign n25576 = x98 | n25248 ;
  assign n25577 = x98 &  n25248 ;
  assign n25578 = ( n25576 & ~n25577 ) | ( n25576 & 1'b0 ) | ( ~n25577 & 1'b0 ) ;
  assign n25590 = ( n25539 & n25550 ) | ( n25539 & n25578 ) | ( n25550 & n25578 ) ;
  assign n25589 = n25539 | n25578 ;
  assign n25591 = ( n25588 & ~n25590 ) | ( n25588 & n25589 ) | ( ~n25590 & n25589 ) ;
  assign n25595 = n25256 &  n25549 ;
  assign n25596 = n25548 &  n25595 ;
  assign n25584 = x97 | n25256 ;
  assign n25585 = x97 &  n25256 ;
  assign n25586 = ( n25584 & ~n25585 ) | ( n25584 & 1'b0 ) | ( ~n25585 & 1'b0 ) ;
  assign n25598 = ( n25538 & n25550 ) | ( n25538 & n25586 ) | ( n25550 & n25586 ) ;
  assign n25597 = n25538 | n25586 ;
  assign n25599 = ( n25596 & ~n25598 ) | ( n25596 & n25597 ) | ( ~n25598 & n25597 ) ;
  assign n25603 = n25264 &  n25549 ;
  assign n25604 = n25548 &  n25603 ;
  assign n25592 = x96 | n25264 ;
  assign n25593 = x96 &  n25264 ;
  assign n25594 = ( n25592 & ~n25593 ) | ( n25592 & 1'b0 ) | ( ~n25593 & 1'b0 ) ;
  assign n25606 = ( n25537 & n25550 ) | ( n25537 & n25594 ) | ( n25550 & n25594 ) ;
  assign n25605 = n25537 | n25594 ;
  assign n25607 = ( n25604 & ~n25606 ) | ( n25604 & n25605 ) | ( ~n25606 & n25605 ) ;
  assign n25611 = n25272 &  n25549 ;
  assign n25612 = n25548 &  n25611 ;
  assign n25600 = x95 | n25272 ;
  assign n25601 = x95 &  n25272 ;
  assign n25602 = ( n25600 & ~n25601 ) | ( n25600 & 1'b0 ) | ( ~n25601 & 1'b0 ) ;
  assign n25614 = ( n25536 & n25550 ) | ( n25536 & n25602 ) | ( n25550 & n25602 ) ;
  assign n25613 = n25536 | n25602 ;
  assign n25615 = ( n25612 & ~n25614 ) | ( n25612 & n25613 ) | ( ~n25614 & n25613 ) ;
  assign n25619 = n25280 &  n25549 ;
  assign n25620 = n25548 &  n25619 ;
  assign n25608 = x94 | n25280 ;
  assign n25609 = x94 &  n25280 ;
  assign n25610 = ( n25608 & ~n25609 ) | ( n25608 & 1'b0 ) | ( ~n25609 & 1'b0 ) ;
  assign n25622 = ( n25535 & n25550 ) | ( n25535 & n25610 ) | ( n25550 & n25610 ) ;
  assign n25621 = n25535 | n25610 ;
  assign n25623 = ( n25620 & ~n25622 ) | ( n25620 & n25621 ) | ( ~n25622 & n25621 ) ;
  assign n25627 = n25288 &  n25549 ;
  assign n25628 = n25548 &  n25627 ;
  assign n25616 = x93 | n25288 ;
  assign n25617 = x93 &  n25288 ;
  assign n25618 = ( n25616 & ~n25617 ) | ( n25616 & 1'b0 ) | ( ~n25617 & 1'b0 ) ;
  assign n25630 = ( n25534 & n25550 ) | ( n25534 & n25618 ) | ( n25550 & n25618 ) ;
  assign n25629 = n25534 | n25618 ;
  assign n25631 = ( n25628 & ~n25630 ) | ( n25628 & n25629 ) | ( ~n25630 & n25629 ) ;
  assign n25635 = n25296 &  n25549 ;
  assign n25636 = n25548 &  n25635 ;
  assign n25624 = x92 | n25296 ;
  assign n25625 = x92 &  n25296 ;
  assign n25626 = ( n25624 & ~n25625 ) | ( n25624 & 1'b0 ) | ( ~n25625 & 1'b0 ) ;
  assign n25638 = ( n25533 & n25550 ) | ( n25533 & n25626 ) | ( n25550 & n25626 ) ;
  assign n25637 = n25533 | n25626 ;
  assign n25639 = ( n25636 & ~n25638 ) | ( n25636 & n25637 ) | ( ~n25638 & n25637 ) ;
  assign n25643 = n25304 &  n25549 ;
  assign n25644 = n25548 &  n25643 ;
  assign n25632 = x91 | n25304 ;
  assign n25633 = x91 &  n25304 ;
  assign n25634 = ( n25632 & ~n25633 ) | ( n25632 & 1'b0 ) | ( ~n25633 & 1'b0 ) ;
  assign n25646 = ( n25532 & n25550 ) | ( n25532 & n25634 ) | ( n25550 & n25634 ) ;
  assign n25645 = n25532 | n25634 ;
  assign n25647 = ( n25644 & ~n25646 ) | ( n25644 & n25645 ) | ( ~n25646 & n25645 ) ;
  assign n25651 = n25312 &  n25549 ;
  assign n25652 = n25548 &  n25651 ;
  assign n25640 = x90 | n25312 ;
  assign n25641 = x90 &  n25312 ;
  assign n25642 = ( n25640 & ~n25641 ) | ( n25640 & 1'b0 ) | ( ~n25641 & 1'b0 ) ;
  assign n25654 = ( n25531 & n25550 ) | ( n25531 & n25642 ) | ( n25550 & n25642 ) ;
  assign n25653 = n25531 | n25642 ;
  assign n25655 = ( n25652 & ~n25654 ) | ( n25652 & n25653 ) | ( ~n25654 & n25653 ) ;
  assign n25659 = n25320 &  n25549 ;
  assign n25660 = n25548 &  n25659 ;
  assign n25648 = x89 | n25320 ;
  assign n25649 = x89 &  n25320 ;
  assign n25650 = ( n25648 & ~n25649 ) | ( n25648 & 1'b0 ) | ( ~n25649 & 1'b0 ) ;
  assign n25662 = ( n25530 & n25550 ) | ( n25530 & n25650 ) | ( n25550 & n25650 ) ;
  assign n25661 = n25530 | n25650 ;
  assign n25663 = ( n25660 & ~n25662 ) | ( n25660 & n25661 ) | ( ~n25662 & n25661 ) ;
  assign n25667 = n25328 &  n25549 ;
  assign n25668 = n25548 &  n25667 ;
  assign n25656 = x88 | n25328 ;
  assign n25657 = x88 &  n25328 ;
  assign n25658 = ( n25656 & ~n25657 ) | ( n25656 & 1'b0 ) | ( ~n25657 & 1'b0 ) ;
  assign n25670 = ( n25529 & n25550 ) | ( n25529 & n25658 ) | ( n25550 & n25658 ) ;
  assign n25669 = n25529 | n25658 ;
  assign n25671 = ( n25668 & ~n25670 ) | ( n25668 & n25669 ) | ( ~n25670 & n25669 ) ;
  assign n25675 = n25336 &  n25549 ;
  assign n25676 = n25548 &  n25675 ;
  assign n25664 = x87 | n25336 ;
  assign n25665 = x87 &  n25336 ;
  assign n25666 = ( n25664 & ~n25665 ) | ( n25664 & 1'b0 ) | ( ~n25665 & 1'b0 ) ;
  assign n25678 = ( n25528 & n25550 ) | ( n25528 & n25666 ) | ( n25550 & n25666 ) ;
  assign n25677 = n25528 | n25666 ;
  assign n25679 = ( n25676 & ~n25678 ) | ( n25676 & n25677 ) | ( ~n25678 & n25677 ) ;
  assign n25683 = n25344 &  n25549 ;
  assign n25684 = n25548 &  n25683 ;
  assign n25672 = x86 | n25344 ;
  assign n25673 = x86 &  n25344 ;
  assign n25674 = ( n25672 & ~n25673 ) | ( n25672 & 1'b0 ) | ( ~n25673 & 1'b0 ) ;
  assign n25686 = ( n25527 & n25550 ) | ( n25527 & n25674 ) | ( n25550 & n25674 ) ;
  assign n25685 = n25527 | n25674 ;
  assign n25687 = ( n25684 & ~n25686 ) | ( n25684 & n25685 ) | ( ~n25686 & n25685 ) ;
  assign n25691 = n25352 &  n25549 ;
  assign n25692 = n25548 &  n25691 ;
  assign n25680 = x85 | n25352 ;
  assign n25681 = x85 &  n25352 ;
  assign n25682 = ( n25680 & ~n25681 ) | ( n25680 & 1'b0 ) | ( ~n25681 & 1'b0 ) ;
  assign n25694 = ( n25526 & n25550 ) | ( n25526 & n25682 ) | ( n25550 & n25682 ) ;
  assign n25693 = n25526 | n25682 ;
  assign n25695 = ( n25692 & ~n25694 ) | ( n25692 & n25693 ) | ( ~n25694 & n25693 ) ;
  assign n25699 = n25360 &  n25549 ;
  assign n25700 = n25548 &  n25699 ;
  assign n25688 = x84 | n25360 ;
  assign n25689 = x84 &  n25360 ;
  assign n25690 = ( n25688 & ~n25689 ) | ( n25688 & 1'b0 ) | ( ~n25689 & 1'b0 ) ;
  assign n25702 = ( n25525 & n25550 ) | ( n25525 & n25690 ) | ( n25550 & n25690 ) ;
  assign n25701 = n25525 | n25690 ;
  assign n25703 = ( n25700 & ~n25702 ) | ( n25700 & n25701 ) | ( ~n25702 & n25701 ) ;
  assign n25707 = n25368 &  n25549 ;
  assign n25708 = n25548 &  n25707 ;
  assign n25696 = x83 | n25368 ;
  assign n25697 = x83 &  n25368 ;
  assign n25698 = ( n25696 & ~n25697 ) | ( n25696 & 1'b0 ) | ( ~n25697 & 1'b0 ) ;
  assign n25710 = ( n25524 & n25550 ) | ( n25524 & n25698 ) | ( n25550 & n25698 ) ;
  assign n25709 = n25524 | n25698 ;
  assign n25711 = ( n25708 & ~n25710 ) | ( n25708 & n25709 ) | ( ~n25710 & n25709 ) ;
  assign n25715 = n25376 &  n25549 ;
  assign n25716 = n25548 &  n25715 ;
  assign n25704 = x82 | n25376 ;
  assign n25705 = x82 &  n25376 ;
  assign n25706 = ( n25704 & ~n25705 ) | ( n25704 & 1'b0 ) | ( ~n25705 & 1'b0 ) ;
  assign n25718 = ( n25523 & n25550 ) | ( n25523 & n25706 ) | ( n25550 & n25706 ) ;
  assign n25717 = n25523 | n25706 ;
  assign n25719 = ( n25716 & ~n25718 ) | ( n25716 & n25717 ) | ( ~n25718 & n25717 ) ;
  assign n25723 = n25384 &  n25549 ;
  assign n25724 = n25548 &  n25723 ;
  assign n25712 = x81 | n25384 ;
  assign n25713 = x81 &  n25384 ;
  assign n25714 = ( n25712 & ~n25713 ) | ( n25712 & 1'b0 ) | ( ~n25713 & 1'b0 ) ;
  assign n25726 = ( n25522 & n25550 ) | ( n25522 & n25714 ) | ( n25550 & n25714 ) ;
  assign n25725 = n25522 | n25714 ;
  assign n25727 = ( n25724 & ~n25726 ) | ( n25724 & n25725 ) | ( ~n25726 & n25725 ) ;
  assign n25731 = n25392 &  n25549 ;
  assign n25732 = n25548 &  n25731 ;
  assign n25720 = x80 | n25392 ;
  assign n25721 = x80 &  n25392 ;
  assign n25722 = ( n25720 & ~n25721 ) | ( n25720 & 1'b0 ) | ( ~n25721 & 1'b0 ) ;
  assign n25734 = ( n25521 & n25550 ) | ( n25521 & n25722 ) | ( n25550 & n25722 ) ;
  assign n25733 = n25521 | n25722 ;
  assign n25735 = ( n25732 & ~n25734 ) | ( n25732 & n25733 ) | ( ~n25734 & n25733 ) ;
  assign n25739 = n25400 &  n25549 ;
  assign n25740 = n25548 &  n25739 ;
  assign n25728 = x79 | n25400 ;
  assign n25729 = x79 &  n25400 ;
  assign n25730 = ( n25728 & ~n25729 ) | ( n25728 & 1'b0 ) | ( ~n25729 & 1'b0 ) ;
  assign n25742 = ( n25520 & n25550 ) | ( n25520 & n25730 ) | ( n25550 & n25730 ) ;
  assign n25741 = n25520 | n25730 ;
  assign n25743 = ( n25740 & ~n25742 ) | ( n25740 & n25741 ) | ( ~n25742 & n25741 ) ;
  assign n25747 = n25408 &  n25549 ;
  assign n25748 = n25548 &  n25747 ;
  assign n25736 = x78 | n25408 ;
  assign n25737 = x78 &  n25408 ;
  assign n25738 = ( n25736 & ~n25737 ) | ( n25736 & 1'b0 ) | ( ~n25737 & 1'b0 ) ;
  assign n25750 = ( n25519 & n25550 ) | ( n25519 & n25738 ) | ( n25550 & n25738 ) ;
  assign n25749 = n25519 | n25738 ;
  assign n25751 = ( n25748 & ~n25750 ) | ( n25748 & n25749 ) | ( ~n25750 & n25749 ) ;
  assign n25755 = n25416 &  n25549 ;
  assign n25756 = n25548 &  n25755 ;
  assign n25744 = x77 | n25416 ;
  assign n25745 = x77 &  n25416 ;
  assign n25746 = ( n25744 & ~n25745 ) | ( n25744 & 1'b0 ) | ( ~n25745 & 1'b0 ) ;
  assign n25758 = ( n25518 & n25550 ) | ( n25518 & n25746 ) | ( n25550 & n25746 ) ;
  assign n25757 = n25518 | n25746 ;
  assign n25759 = ( n25756 & ~n25758 ) | ( n25756 & n25757 ) | ( ~n25758 & n25757 ) ;
  assign n25763 = n25424 &  n25549 ;
  assign n25764 = n25548 &  n25763 ;
  assign n25752 = x76 | n25424 ;
  assign n25753 = x76 &  n25424 ;
  assign n25754 = ( n25752 & ~n25753 ) | ( n25752 & 1'b0 ) | ( ~n25753 & 1'b0 ) ;
  assign n25766 = ( n25517 & n25550 ) | ( n25517 & n25754 ) | ( n25550 & n25754 ) ;
  assign n25765 = n25517 | n25754 ;
  assign n25767 = ( n25764 & ~n25766 ) | ( n25764 & n25765 ) | ( ~n25766 & n25765 ) ;
  assign n25771 = n25432 &  n25549 ;
  assign n25772 = n25548 &  n25771 ;
  assign n25760 = x75 | n25432 ;
  assign n25761 = x75 &  n25432 ;
  assign n25762 = ( n25760 & ~n25761 ) | ( n25760 & 1'b0 ) | ( ~n25761 & 1'b0 ) ;
  assign n25774 = ( n25516 & n25550 ) | ( n25516 & n25762 ) | ( n25550 & n25762 ) ;
  assign n25773 = n25516 | n25762 ;
  assign n25775 = ( n25772 & ~n25774 ) | ( n25772 & n25773 ) | ( ~n25774 & n25773 ) ;
  assign n25779 = n25440 &  n25549 ;
  assign n25780 = n25548 &  n25779 ;
  assign n25768 = x74 | n25440 ;
  assign n25769 = x74 &  n25440 ;
  assign n25770 = ( n25768 & ~n25769 ) | ( n25768 & 1'b0 ) | ( ~n25769 & 1'b0 ) ;
  assign n25782 = ( n25515 & n25550 ) | ( n25515 & n25770 ) | ( n25550 & n25770 ) ;
  assign n25781 = n25515 | n25770 ;
  assign n25783 = ( n25780 & ~n25782 ) | ( n25780 & n25781 ) | ( ~n25782 & n25781 ) ;
  assign n25787 = n25448 &  n25549 ;
  assign n25788 = n25548 &  n25787 ;
  assign n25776 = x73 | n25448 ;
  assign n25777 = x73 &  n25448 ;
  assign n25778 = ( n25776 & ~n25777 ) | ( n25776 & 1'b0 ) | ( ~n25777 & 1'b0 ) ;
  assign n25790 = ( n25514 & n25550 ) | ( n25514 & n25778 ) | ( n25550 & n25778 ) ;
  assign n25789 = n25514 | n25778 ;
  assign n25791 = ( n25788 & ~n25790 ) | ( n25788 & n25789 ) | ( ~n25790 & n25789 ) ;
  assign n25795 = n25456 &  n25549 ;
  assign n25796 = n25548 &  n25795 ;
  assign n25784 = x72 | n25456 ;
  assign n25785 = x72 &  n25456 ;
  assign n25786 = ( n25784 & ~n25785 ) | ( n25784 & 1'b0 ) | ( ~n25785 & 1'b0 ) ;
  assign n25798 = ( n25513 & n25550 ) | ( n25513 & n25786 ) | ( n25550 & n25786 ) ;
  assign n25797 = n25513 | n25786 ;
  assign n25799 = ( n25796 & ~n25798 ) | ( n25796 & n25797 ) | ( ~n25798 & n25797 ) ;
  assign n25803 = n25464 &  n25549 ;
  assign n25804 = n25548 &  n25803 ;
  assign n25792 = x71 | n25464 ;
  assign n25793 = x71 &  n25464 ;
  assign n25794 = ( n25792 & ~n25793 ) | ( n25792 & 1'b0 ) | ( ~n25793 & 1'b0 ) ;
  assign n25806 = ( n25512 & n25550 ) | ( n25512 & n25794 ) | ( n25550 & n25794 ) ;
  assign n25805 = n25512 | n25794 ;
  assign n25807 = ( n25804 & ~n25806 ) | ( n25804 & n25805 ) | ( ~n25806 & n25805 ) ;
  assign n25811 = n25472 &  n25549 ;
  assign n25812 = n25548 &  n25811 ;
  assign n25800 = x70 | n25472 ;
  assign n25801 = x70 &  n25472 ;
  assign n25802 = ( n25800 & ~n25801 ) | ( n25800 & 1'b0 ) | ( ~n25801 & 1'b0 ) ;
  assign n25814 = ( n25511 & n25550 ) | ( n25511 & n25802 ) | ( n25550 & n25802 ) ;
  assign n25813 = n25511 | n25802 ;
  assign n25815 = ( n25812 & ~n25814 ) | ( n25812 & n25813 ) | ( ~n25814 & n25813 ) ;
  assign n25819 = n25480 &  n25549 ;
  assign n25820 = n25548 &  n25819 ;
  assign n25808 = x69 | n25480 ;
  assign n25809 = x69 &  n25480 ;
  assign n25810 = ( n25808 & ~n25809 ) | ( n25808 & 1'b0 ) | ( ~n25809 & 1'b0 ) ;
  assign n25822 = ( n25510 & n25550 ) | ( n25510 & n25810 ) | ( n25550 & n25810 ) ;
  assign n25821 = n25510 | n25810 ;
  assign n25823 = ( n25820 & ~n25822 ) | ( n25820 & n25821 ) | ( ~n25822 & n25821 ) ;
  assign n25827 = n25488 &  n25549 ;
  assign n25828 = n25548 &  n25827 ;
  assign n25816 = x68 | n25488 ;
  assign n25817 = x68 &  n25488 ;
  assign n25818 = ( n25816 & ~n25817 ) | ( n25816 & 1'b0 ) | ( ~n25817 & 1'b0 ) ;
  assign n25830 = ( n25509 & n25550 ) | ( n25509 & n25818 ) | ( n25550 & n25818 ) ;
  assign n25829 = n25509 | n25818 ;
  assign n25831 = ( n25828 & ~n25830 ) | ( n25828 & n25829 ) | ( ~n25830 & n25829 ) ;
  assign n25835 = n25496 &  n25549 ;
  assign n25836 = n25548 &  n25835 ;
  assign n25824 = x67 | n25496 ;
  assign n25825 = x67 &  n25496 ;
  assign n25826 = ( n25824 & ~n25825 ) | ( n25824 & 1'b0 ) | ( ~n25825 & 1'b0 ) ;
  assign n25838 = ( n25508 & n25550 ) | ( n25508 & n25826 ) | ( n25550 & n25826 ) ;
  assign n25837 = n25508 | n25826 ;
  assign n25839 = ( n25836 & ~n25838 ) | ( n25836 & n25837 ) | ( ~n25838 & n25837 ) ;
  assign n25840 = n25502 &  n25549 ;
  assign n25841 = n25548 &  n25840 ;
  assign n25832 = x66 | n25502 ;
  assign n25833 = x66 &  n25502 ;
  assign n25834 = ( n25832 & ~n25833 ) | ( n25832 & 1'b0 ) | ( ~n25833 & 1'b0 ) ;
  assign n25843 = ( n25507 & n25550 ) | ( n25507 & n25834 ) | ( n25550 & n25834 ) ;
  assign n25842 = n25507 | n25834 ;
  assign n25844 = ( n25841 & ~n25843 ) | ( n25841 & n25842 ) | ( ~n25843 & n25842 ) ;
  assign n25845 = ( x65 & ~n7012 ) | ( x65 & n25506 ) | ( ~n7012 & n25506 ) ;
  assign n25846 = ( n25507 & ~x65 ) | ( n25507 & n25845 ) | ( ~x65 & n25845 ) ;
  assign n25847 = ~n25550 & n25846 ;
  assign n25848 = n25506 &  n25549 ;
  assign n25849 = n25548 &  n25848 ;
  assign n25850 = n25847 | n25849 ;
  assign n25851 = ( x64 & ~n25550 ) | ( x64 & 1'b0 ) | ( ~n25550 & 1'b0 ) ;
  assign n25852 = ( x25 & ~n25851 ) | ( x25 & 1'b0 ) | ( ~n25851 & 1'b0 ) ;
  assign n25853 = ( n7012 & ~n25550 ) | ( n7012 & 1'b0 ) | ( ~n25550 & 1'b0 ) ;
  assign n25854 = n25852 | n25853 ;
  assign n25855 = ( x65 & ~n25854 ) | ( x65 & n7495 ) | ( ~n25854 & n7495 ) ;
  assign n25856 = ( x66 & ~n25850 ) | ( x66 & n25855 ) | ( ~n25850 & n25855 ) ;
  assign n25857 = ( x67 & ~n25844 ) | ( x67 & n25856 ) | ( ~n25844 & n25856 ) ;
  assign n25858 = ( x68 & ~n25839 ) | ( x68 & n25857 ) | ( ~n25839 & n25857 ) ;
  assign n25859 = ( x69 & ~n25831 ) | ( x69 & n25858 ) | ( ~n25831 & n25858 ) ;
  assign n25860 = ( x70 & ~n25823 ) | ( x70 & n25859 ) | ( ~n25823 & n25859 ) ;
  assign n25861 = ( x71 & ~n25815 ) | ( x71 & n25860 ) | ( ~n25815 & n25860 ) ;
  assign n25862 = ( x72 & ~n25807 ) | ( x72 & n25861 ) | ( ~n25807 & n25861 ) ;
  assign n25863 = ( x73 & ~n25799 ) | ( x73 & n25862 ) | ( ~n25799 & n25862 ) ;
  assign n25864 = ( x74 & ~n25791 ) | ( x74 & n25863 ) | ( ~n25791 & n25863 ) ;
  assign n25865 = ( x75 & ~n25783 ) | ( x75 & n25864 ) | ( ~n25783 & n25864 ) ;
  assign n25866 = ( x76 & ~n25775 ) | ( x76 & n25865 ) | ( ~n25775 & n25865 ) ;
  assign n25867 = ( x77 & ~n25767 ) | ( x77 & n25866 ) | ( ~n25767 & n25866 ) ;
  assign n25868 = ( x78 & ~n25759 ) | ( x78 & n25867 ) | ( ~n25759 & n25867 ) ;
  assign n25869 = ( x79 & ~n25751 ) | ( x79 & n25868 ) | ( ~n25751 & n25868 ) ;
  assign n25870 = ( x80 & ~n25743 ) | ( x80 & n25869 ) | ( ~n25743 & n25869 ) ;
  assign n25871 = ( x81 & ~n25735 ) | ( x81 & n25870 ) | ( ~n25735 & n25870 ) ;
  assign n25872 = ( x82 & ~n25727 ) | ( x82 & n25871 ) | ( ~n25727 & n25871 ) ;
  assign n25873 = ( x83 & ~n25719 ) | ( x83 & n25872 ) | ( ~n25719 & n25872 ) ;
  assign n25874 = ( x84 & ~n25711 ) | ( x84 & n25873 ) | ( ~n25711 & n25873 ) ;
  assign n25875 = ( x85 & ~n25703 ) | ( x85 & n25874 ) | ( ~n25703 & n25874 ) ;
  assign n25876 = ( x86 & ~n25695 ) | ( x86 & n25875 ) | ( ~n25695 & n25875 ) ;
  assign n25877 = ( x87 & ~n25687 ) | ( x87 & n25876 ) | ( ~n25687 & n25876 ) ;
  assign n25878 = ( x88 & ~n25679 ) | ( x88 & n25877 ) | ( ~n25679 & n25877 ) ;
  assign n25879 = ( x89 & ~n25671 ) | ( x89 & n25878 ) | ( ~n25671 & n25878 ) ;
  assign n25880 = ( x90 & ~n25663 ) | ( x90 & n25879 ) | ( ~n25663 & n25879 ) ;
  assign n25881 = ( x91 & ~n25655 ) | ( x91 & n25880 ) | ( ~n25655 & n25880 ) ;
  assign n25882 = ( x92 & ~n25647 ) | ( x92 & n25881 ) | ( ~n25647 & n25881 ) ;
  assign n25883 = ( x93 & ~n25639 ) | ( x93 & n25882 ) | ( ~n25639 & n25882 ) ;
  assign n25884 = ( x94 & ~n25631 ) | ( x94 & n25883 ) | ( ~n25631 & n25883 ) ;
  assign n25885 = ( x95 & ~n25623 ) | ( x95 & n25884 ) | ( ~n25623 & n25884 ) ;
  assign n25886 = ( x96 & ~n25615 ) | ( x96 & n25885 ) | ( ~n25615 & n25885 ) ;
  assign n25887 = ( x97 & ~n25607 ) | ( x97 & n25886 ) | ( ~n25607 & n25886 ) ;
  assign n25888 = ( x98 & ~n25599 ) | ( x98 & n25887 ) | ( ~n25599 & n25887 ) ;
  assign n25889 = ( x99 & ~n25591 ) | ( x99 & n25888 ) | ( ~n25591 & n25888 ) ;
  assign n25890 = ( x100 & ~n25583 ) | ( x100 & n25889 ) | ( ~n25583 & n25889 ) ;
  assign n25891 = ( x101 & ~n25575 ) | ( x101 & n25890 ) | ( ~n25575 & n25890 ) ;
  assign n25892 = ( x102 & ~n25567 ) | ( x102 & n25891 ) | ( ~n25567 & n25891 ) ;
  assign n25899 = ( x103 & ~n7535 ) | ( x103 & n25892 ) | ( ~n7535 & n25892 ) ;
  assign n25898 = x103 &  n25892 ;
  assign n25900 = ( n25559 & ~n25899 ) | ( n25559 & n25898 ) | ( ~n25899 & n25898 ) ;
  assign n25893 = ( x103 & ~n25559 ) | ( x103 & n25892 ) | ( ~n25559 & n25892 ) ;
  assign n25894 = n7535 | n25893 ;
  assign n25901 = n25567 &  n25894 ;
  assign n25895 = x102 | n25567 ;
  assign n25896 = x102 &  n25567 ;
  assign n25897 = ( n25895 & ~n25896 ) | ( n25895 & 1'b0 ) | ( ~n25896 & 1'b0 ) ;
  assign n25905 = ( n7535 & n25891 ) | ( n7535 & n25897 ) | ( n25891 & n25897 ) ;
  assign n25906 = ( n25891 & ~n25893 ) | ( n25891 & n25897 ) | ( ~n25893 & n25897 ) ;
  assign n25907 = ~n25905 & n25906 ;
  assign n25908 = n25901 | n25907 ;
  assign n25909 = n25575 &  n25894 ;
  assign n25902 = x101 | n25575 ;
  assign n25903 = x101 &  n25575 ;
  assign n25904 = ( n25902 & ~n25903 ) | ( n25902 & 1'b0 ) | ( ~n25903 & 1'b0 ) ;
  assign n25913 = ( n7535 & n25890 ) | ( n7535 & n25904 ) | ( n25890 & n25904 ) ;
  assign n25914 = ( n25890 & ~n25893 ) | ( n25890 & n25904 ) | ( ~n25893 & n25904 ) ;
  assign n25915 = ~n25913 & n25914 ;
  assign n25916 = n25909 | n25915 ;
  assign n25917 = n25583 &  n25894 ;
  assign n25910 = x100 | n25583 ;
  assign n25911 = x100 &  n25583 ;
  assign n25912 = ( n25910 & ~n25911 ) | ( n25910 & 1'b0 ) | ( ~n25911 & 1'b0 ) ;
  assign n25921 = ( n7535 & n25889 ) | ( n7535 & n25912 ) | ( n25889 & n25912 ) ;
  assign n25922 = ( n25889 & ~n25893 ) | ( n25889 & n25912 ) | ( ~n25893 & n25912 ) ;
  assign n25923 = ~n25921 & n25922 ;
  assign n25924 = n25917 | n25923 ;
  assign n25925 = n25591 &  n25894 ;
  assign n25918 = x99 | n25591 ;
  assign n25919 = x99 &  n25591 ;
  assign n25920 = ( n25918 & ~n25919 ) | ( n25918 & 1'b0 ) | ( ~n25919 & 1'b0 ) ;
  assign n25929 = ( n7535 & n25888 ) | ( n7535 & n25920 ) | ( n25888 & n25920 ) ;
  assign n25930 = ( n25888 & ~n25893 ) | ( n25888 & n25920 ) | ( ~n25893 & n25920 ) ;
  assign n25931 = ~n25929 & n25930 ;
  assign n25932 = n25925 | n25931 ;
  assign n25933 = n25599 &  n25894 ;
  assign n25926 = x98 | n25599 ;
  assign n25927 = x98 &  n25599 ;
  assign n25928 = ( n25926 & ~n25927 ) | ( n25926 & 1'b0 ) | ( ~n25927 & 1'b0 ) ;
  assign n25937 = ( n7535 & n25887 ) | ( n7535 & n25928 ) | ( n25887 & n25928 ) ;
  assign n25938 = ( n25887 & ~n25893 ) | ( n25887 & n25928 ) | ( ~n25893 & n25928 ) ;
  assign n25939 = ~n25937 & n25938 ;
  assign n25940 = n25933 | n25939 ;
  assign n25941 = n25607 &  n25894 ;
  assign n25934 = x97 | n25607 ;
  assign n25935 = x97 &  n25607 ;
  assign n25936 = ( n25934 & ~n25935 ) | ( n25934 & 1'b0 ) | ( ~n25935 & 1'b0 ) ;
  assign n25945 = ( n7535 & n25886 ) | ( n7535 & n25936 ) | ( n25886 & n25936 ) ;
  assign n25946 = ( n25886 & ~n25893 ) | ( n25886 & n25936 ) | ( ~n25893 & n25936 ) ;
  assign n25947 = ~n25945 & n25946 ;
  assign n25948 = n25941 | n25947 ;
  assign n25949 = n25615 &  n25894 ;
  assign n25942 = x96 | n25615 ;
  assign n25943 = x96 &  n25615 ;
  assign n25944 = ( n25942 & ~n25943 ) | ( n25942 & 1'b0 ) | ( ~n25943 & 1'b0 ) ;
  assign n25953 = ( n7535 & n25885 ) | ( n7535 & n25944 ) | ( n25885 & n25944 ) ;
  assign n25954 = ( n25885 & ~n25893 ) | ( n25885 & n25944 ) | ( ~n25893 & n25944 ) ;
  assign n25955 = ~n25953 & n25954 ;
  assign n25956 = n25949 | n25955 ;
  assign n25957 = n25623 &  n25894 ;
  assign n25950 = x95 | n25623 ;
  assign n25951 = x95 &  n25623 ;
  assign n25952 = ( n25950 & ~n25951 ) | ( n25950 & 1'b0 ) | ( ~n25951 & 1'b0 ) ;
  assign n25961 = ( n7535 & n25884 ) | ( n7535 & n25952 ) | ( n25884 & n25952 ) ;
  assign n25962 = ( n25884 & ~n25893 ) | ( n25884 & n25952 ) | ( ~n25893 & n25952 ) ;
  assign n25963 = ~n25961 & n25962 ;
  assign n25964 = n25957 | n25963 ;
  assign n25965 = n25631 &  n25894 ;
  assign n25958 = x94 | n25631 ;
  assign n25959 = x94 &  n25631 ;
  assign n25960 = ( n25958 & ~n25959 ) | ( n25958 & 1'b0 ) | ( ~n25959 & 1'b0 ) ;
  assign n25969 = ( n7535 & n25883 ) | ( n7535 & n25960 ) | ( n25883 & n25960 ) ;
  assign n25970 = ( n25883 & ~n25893 ) | ( n25883 & n25960 ) | ( ~n25893 & n25960 ) ;
  assign n25971 = ~n25969 & n25970 ;
  assign n25972 = n25965 | n25971 ;
  assign n25973 = n25639 &  n25894 ;
  assign n25966 = x93 | n25639 ;
  assign n25967 = x93 &  n25639 ;
  assign n25968 = ( n25966 & ~n25967 ) | ( n25966 & 1'b0 ) | ( ~n25967 & 1'b0 ) ;
  assign n25977 = ( n7535 & n25882 ) | ( n7535 & n25968 ) | ( n25882 & n25968 ) ;
  assign n25978 = ( n25882 & ~n25893 ) | ( n25882 & n25968 ) | ( ~n25893 & n25968 ) ;
  assign n25979 = ~n25977 & n25978 ;
  assign n25980 = n25973 | n25979 ;
  assign n25981 = n25647 &  n25894 ;
  assign n25974 = x92 | n25647 ;
  assign n25975 = x92 &  n25647 ;
  assign n25976 = ( n25974 & ~n25975 ) | ( n25974 & 1'b0 ) | ( ~n25975 & 1'b0 ) ;
  assign n25985 = ( n7535 & n25881 ) | ( n7535 & n25976 ) | ( n25881 & n25976 ) ;
  assign n25986 = ( n25881 & ~n25893 ) | ( n25881 & n25976 ) | ( ~n25893 & n25976 ) ;
  assign n25987 = ~n25985 & n25986 ;
  assign n25988 = n25981 | n25987 ;
  assign n25989 = n25655 &  n25894 ;
  assign n25982 = x91 | n25655 ;
  assign n25983 = x91 &  n25655 ;
  assign n25984 = ( n25982 & ~n25983 ) | ( n25982 & 1'b0 ) | ( ~n25983 & 1'b0 ) ;
  assign n25993 = ( n7535 & n25880 ) | ( n7535 & n25984 ) | ( n25880 & n25984 ) ;
  assign n25994 = ( n25880 & ~n25893 ) | ( n25880 & n25984 ) | ( ~n25893 & n25984 ) ;
  assign n25995 = ~n25993 & n25994 ;
  assign n25996 = n25989 | n25995 ;
  assign n25997 = n25663 &  n25894 ;
  assign n25990 = x90 | n25663 ;
  assign n25991 = x90 &  n25663 ;
  assign n25992 = ( n25990 & ~n25991 ) | ( n25990 & 1'b0 ) | ( ~n25991 & 1'b0 ) ;
  assign n26001 = ( n7535 & n25879 ) | ( n7535 & n25992 ) | ( n25879 & n25992 ) ;
  assign n26002 = ( n25879 & ~n25893 ) | ( n25879 & n25992 ) | ( ~n25893 & n25992 ) ;
  assign n26003 = ~n26001 & n26002 ;
  assign n26004 = n25997 | n26003 ;
  assign n26005 = n25671 &  n25894 ;
  assign n25998 = x89 | n25671 ;
  assign n25999 = x89 &  n25671 ;
  assign n26000 = ( n25998 & ~n25999 ) | ( n25998 & 1'b0 ) | ( ~n25999 & 1'b0 ) ;
  assign n26009 = ( n7535 & n25878 ) | ( n7535 & n26000 ) | ( n25878 & n26000 ) ;
  assign n26010 = ( n25878 & ~n25893 ) | ( n25878 & n26000 ) | ( ~n25893 & n26000 ) ;
  assign n26011 = ~n26009 & n26010 ;
  assign n26012 = n26005 | n26011 ;
  assign n26013 = n25679 &  n25894 ;
  assign n26006 = x88 | n25679 ;
  assign n26007 = x88 &  n25679 ;
  assign n26008 = ( n26006 & ~n26007 ) | ( n26006 & 1'b0 ) | ( ~n26007 & 1'b0 ) ;
  assign n26017 = ( n7535 & n25877 ) | ( n7535 & n26008 ) | ( n25877 & n26008 ) ;
  assign n26018 = ( n25877 & ~n25893 ) | ( n25877 & n26008 ) | ( ~n25893 & n26008 ) ;
  assign n26019 = ~n26017 & n26018 ;
  assign n26020 = n26013 | n26019 ;
  assign n26021 = n25687 &  n25894 ;
  assign n26014 = x87 | n25687 ;
  assign n26015 = x87 &  n25687 ;
  assign n26016 = ( n26014 & ~n26015 ) | ( n26014 & 1'b0 ) | ( ~n26015 & 1'b0 ) ;
  assign n26025 = ( n7535 & n25876 ) | ( n7535 & n26016 ) | ( n25876 & n26016 ) ;
  assign n26026 = ( n25876 & ~n25893 ) | ( n25876 & n26016 ) | ( ~n25893 & n26016 ) ;
  assign n26027 = ~n26025 & n26026 ;
  assign n26028 = n26021 | n26027 ;
  assign n26029 = n25695 &  n25894 ;
  assign n26022 = x86 | n25695 ;
  assign n26023 = x86 &  n25695 ;
  assign n26024 = ( n26022 & ~n26023 ) | ( n26022 & 1'b0 ) | ( ~n26023 & 1'b0 ) ;
  assign n26033 = ( n7535 & n25875 ) | ( n7535 & n26024 ) | ( n25875 & n26024 ) ;
  assign n26034 = ( n25875 & ~n25893 ) | ( n25875 & n26024 ) | ( ~n25893 & n26024 ) ;
  assign n26035 = ~n26033 & n26034 ;
  assign n26036 = n26029 | n26035 ;
  assign n26037 = n25703 &  n25894 ;
  assign n26030 = x85 | n25703 ;
  assign n26031 = x85 &  n25703 ;
  assign n26032 = ( n26030 & ~n26031 ) | ( n26030 & 1'b0 ) | ( ~n26031 & 1'b0 ) ;
  assign n26041 = ( n7535 & n25874 ) | ( n7535 & n26032 ) | ( n25874 & n26032 ) ;
  assign n26042 = ( n25874 & ~n25893 ) | ( n25874 & n26032 ) | ( ~n25893 & n26032 ) ;
  assign n26043 = ~n26041 & n26042 ;
  assign n26044 = n26037 | n26043 ;
  assign n26045 = n25711 &  n25894 ;
  assign n26038 = x84 | n25711 ;
  assign n26039 = x84 &  n25711 ;
  assign n26040 = ( n26038 & ~n26039 ) | ( n26038 & 1'b0 ) | ( ~n26039 & 1'b0 ) ;
  assign n26049 = ( n7535 & n25873 ) | ( n7535 & n26040 ) | ( n25873 & n26040 ) ;
  assign n26050 = ( n25873 & ~n25893 ) | ( n25873 & n26040 ) | ( ~n25893 & n26040 ) ;
  assign n26051 = ~n26049 & n26050 ;
  assign n26052 = n26045 | n26051 ;
  assign n26053 = n25719 &  n25894 ;
  assign n26046 = x83 | n25719 ;
  assign n26047 = x83 &  n25719 ;
  assign n26048 = ( n26046 & ~n26047 ) | ( n26046 & 1'b0 ) | ( ~n26047 & 1'b0 ) ;
  assign n26057 = ( n7535 & n25872 ) | ( n7535 & n26048 ) | ( n25872 & n26048 ) ;
  assign n26058 = ( n25872 & ~n25893 ) | ( n25872 & n26048 ) | ( ~n25893 & n26048 ) ;
  assign n26059 = ~n26057 & n26058 ;
  assign n26060 = n26053 | n26059 ;
  assign n26061 = n25727 &  n25894 ;
  assign n26054 = x82 | n25727 ;
  assign n26055 = x82 &  n25727 ;
  assign n26056 = ( n26054 & ~n26055 ) | ( n26054 & 1'b0 ) | ( ~n26055 & 1'b0 ) ;
  assign n26065 = ( n7535 & n25871 ) | ( n7535 & n26056 ) | ( n25871 & n26056 ) ;
  assign n26066 = ( n25871 & ~n25893 ) | ( n25871 & n26056 ) | ( ~n25893 & n26056 ) ;
  assign n26067 = ~n26065 & n26066 ;
  assign n26068 = n26061 | n26067 ;
  assign n26069 = n25735 &  n25894 ;
  assign n26062 = x81 | n25735 ;
  assign n26063 = x81 &  n25735 ;
  assign n26064 = ( n26062 & ~n26063 ) | ( n26062 & 1'b0 ) | ( ~n26063 & 1'b0 ) ;
  assign n26073 = ( n7535 & n25870 ) | ( n7535 & n26064 ) | ( n25870 & n26064 ) ;
  assign n26074 = ( n25870 & ~n25893 ) | ( n25870 & n26064 ) | ( ~n25893 & n26064 ) ;
  assign n26075 = ~n26073 & n26074 ;
  assign n26076 = n26069 | n26075 ;
  assign n26077 = n25743 &  n25894 ;
  assign n26070 = x80 | n25743 ;
  assign n26071 = x80 &  n25743 ;
  assign n26072 = ( n26070 & ~n26071 ) | ( n26070 & 1'b0 ) | ( ~n26071 & 1'b0 ) ;
  assign n26081 = ( n7535 & n25869 ) | ( n7535 & n26072 ) | ( n25869 & n26072 ) ;
  assign n26082 = ( n25869 & ~n25893 ) | ( n25869 & n26072 ) | ( ~n25893 & n26072 ) ;
  assign n26083 = ~n26081 & n26082 ;
  assign n26084 = n26077 | n26083 ;
  assign n26085 = n25751 &  n25894 ;
  assign n26078 = x79 | n25751 ;
  assign n26079 = x79 &  n25751 ;
  assign n26080 = ( n26078 & ~n26079 ) | ( n26078 & 1'b0 ) | ( ~n26079 & 1'b0 ) ;
  assign n26089 = ( n7535 & n25868 ) | ( n7535 & n26080 ) | ( n25868 & n26080 ) ;
  assign n26090 = ( n25868 & ~n25893 ) | ( n25868 & n26080 ) | ( ~n25893 & n26080 ) ;
  assign n26091 = ~n26089 & n26090 ;
  assign n26092 = n26085 | n26091 ;
  assign n26093 = n25759 &  n25894 ;
  assign n26086 = x78 | n25759 ;
  assign n26087 = x78 &  n25759 ;
  assign n26088 = ( n26086 & ~n26087 ) | ( n26086 & 1'b0 ) | ( ~n26087 & 1'b0 ) ;
  assign n26097 = ( n7535 & n25867 ) | ( n7535 & n26088 ) | ( n25867 & n26088 ) ;
  assign n26098 = ( n25867 & ~n25893 ) | ( n25867 & n26088 ) | ( ~n25893 & n26088 ) ;
  assign n26099 = ~n26097 & n26098 ;
  assign n26100 = n26093 | n26099 ;
  assign n26101 = n25767 &  n25894 ;
  assign n26094 = x77 | n25767 ;
  assign n26095 = x77 &  n25767 ;
  assign n26096 = ( n26094 & ~n26095 ) | ( n26094 & 1'b0 ) | ( ~n26095 & 1'b0 ) ;
  assign n26105 = ( n7535 & n25866 ) | ( n7535 & n26096 ) | ( n25866 & n26096 ) ;
  assign n26106 = ( n25866 & ~n25893 ) | ( n25866 & n26096 ) | ( ~n25893 & n26096 ) ;
  assign n26107 = ~n26105 & n26106 ;
  assign n26108 = n26101 | n26107 ;
  assign n26109 = n25775 &  n25894 ;
  assign n26102 = x76 | n25775 ;
  assign n26103 = x76 &  n25775 ;
  assign n26104 = ( n26102 & ~n26103 ) | ( n26102 & 1'b0 ) | ( ~n26103 & 1'b0 ) ;
  assign n26113 = ( n7535 & n25865 ) | ( n7535 & n26104 ) | ( n25865 & n26104 ) ;
  assign n26114 = ( n25865 & ~n25893 ) | ( n25865 & n26104 ) | ( ~n25893 & n26104 ) ;
  assign n26115 = ~n26113 & n26114 ;
  assign n26116 = n26109 | n26115 ;
  assign n26117 = n25783 &  n25894 ;
  assign n26110 = x75 | n25783 ;
  assign n26111 = x75 &  n25783 ;
  assign n26112 = ( n26110 & ~n26111 ) | ( n26110 & 1'b0 ) | ( ~n26111 & 1'b0 ) ;
  assign n26121 = ( n7535 & n25864 ) | ( n7535 & n26112 ) | ( n25864 & n26112 ) ;
  assign n26122 = ( n25864 & ~n25893 ) | ( n25864 & n26112 ) | ( ~n25893 & n26112 ) ;
  assign n26123 = ~n26121 & n26122 ;
  assign n26124 = n26117 | n26123 ;
  assign n26125 = n25791 &  n25894 ;
  assign n26118 = x74 | n25791 ;
  assign n26119 = x74 &  n25791 ;
  assign n26120 = ( n26118 & ~n26119 ) | ( n26118 & 1'b0 ) | ( ~n26119 & 1'b0 ) ;
  assign n26129 = ( n7535 & n25863 ) | ( n7535 & n26120 ) | ( n25863 & n26120 ) ;
  assign n26130 = ( n25863 & ~n25893 ) | ( n25863 & n26120 ) | ( ~n25893 & n26120 ) ;
  assign n26131 = ~n26129 & n26130 ;
  assign n26132 = n26125 | n26131 ;
  assign n26133 = n25799 &  n25894 ;
  assign n26126 = x73 | n25799 ;
  assign n26127 = x73 &  n25799 ;
  assign n26128 = ( n26126 & ~n26127 ) | ( n26126 & 1'b0 ) | ( ~n26127 & 1'b0 ) ;
  assign n26137 = ( n7535 & n25862 ) | ( n7535 & n26128 ) | ( n25862 & n26128 ) ;
  assign n26138 = ( n25862 & ~n25893 ) | ( n25862 & n26128 ) | ( ~n25893 & n26128 ) ;
  assign n26139 = ~n26137 & n26138 ;
  assign n26140 = n26133 | n26139 ;
  assign n26141 = n25807 &  n25894 ;
  assign n26134 = x72 | n25807 ;
  assign n26135 = x72 &  n25807 ;
  assign n26136 = ( n26134 & ~n26135 ) | ( n26134 & 1'b0 ) | ( ~n26135 & 1'b0 ) ;
  assign n26145 = ( n7535 & n25861 ) | ( n7535 & n26136 ) | ( n25861 & n26136 ) ;
  assign n26146 = ( n25861 & ~n25893 ) | ( n25861 & n26136 ) | ( ~n25893 & n26136 ) ;
  assign n26147 = ~n26145 & n26146 ;
  assign n26148 = n26141 | n26147 ;
  assign n26149 = n25815 &  n25894 ;
  assign n26142 = x71 | n25815 ;
  assign n26143 = x71 &  n25815 ;
  assign n26144 = ( n26142 & ~n26143 ) | ( n26142 & 1'b0 ) | ( ~n26143 & 1'b0 ) ;
  assign n26153 = ( n7535 & n25860 ) | ( n7535 & n26144 ) | ( n25860 & n26144 ) ;
  assign n26154 = ( n25860 & ~n25893 ) | ( n25860 & n26144 ) | ( ~n25893 & n26144 ) ;
  assign n26155 = ~n26153 & n26154 ;
  assign n26156 = n26149 | n26155 ;
  assign n26157 = n25823 &  n25894 ;
  assign n26150 = x70 | n25823 ;
  assign n26151 = x70 &  n25823 ;
  assign n26152 = ( n26150 & ~n26151 ) | ( n26150 & 1'b0 ) | ( ~n26151 & 1'b0 ) ;
  assign n26161 = ( n7535 & n25859 ) | ( n7535 & n26152 ) | ( n25859 & n26152 ) ;
  assign n26162 = ( n25859 & ~n25893 ) | ( n25859 & n26152 ) | ( ~n25893 & n26152 ) ;
  assign n26163 = ~n26161 & n26162 ;
  assign n26164 = n26157 | n26163 ;
  assign n26165 = n25831 &  n25894 ;
  assign n26158 = x69 | n25831 ;
  assign n26159 = x69 &  n25831 ;
  assign n26160 = ( n26158 & ~n26159 ) | ( n26158 & 1'b0 ) | ( ~n26159 & 1'b0 ) ;
  assign n26169 = ( n7535 & n25858 ) | ( n7535 & n26160 ) | ( n25858 & n26160 ) ;
  assign n26170 = ( n25858 & ~n25893 ) | ( n25858 & n26160 ) | ( ~n25893 & n26160 ) ;
  assign n26171 = ~n26169 & n26170 ;
  assign n26172 = n26165 | n26171 ;
  assign n26173 = n25839 &  n25894 ;
  assign n26166 = x68 | n25839 ;
  assign n26167 = x68 &  n25839 ;
  assign n26168 = ( n26166 & ~n26167 ) | ( n26166 & 1'b0 ) | ( ~n26167 & 1'b0 ) ;
  assign n26177 = ( n7535 & n25857 ) | ( n7535 & n26168 ) | ( n25857 & n26168 ) ;
  assign n26178 = ( n25857 & ~n25893 ) | ( n25857 & n26168 ) | ( ~n25893 & n26168 ) ;
  assign n26179 = ~n26177 & n26178 ;
  assign n26180 = n26173 | n26179 ;
  assign n26181 = n25844 &  n25894 ;
  assign n26174 = x67 | n25844 ;
  assign n26175 = x67 &  n25844 ;
  assign n26176 = ( n26174 & ~n26175 ) | ( n26174 & 1'b0 ) | ( ~n26175 & 1'b0 ) ;
  assign n26185 = ( n7535 & n25856 ) | ( n7535 & n26176 ) | ( n25856 & n26176 ) ;
  assign n26186 = ( n25856 & ~n25893 ) | ( n25856 & n26176 ) | ( ~n25893 & n26176 ) ;
  assign n26187 = ~n26185 & n26186 ;
  assign n26188 = n26181 | n26187 ;
  assign n26189 = n25850 &  n25894 ;
  assign n26182 = x66 | n25850 ;
  assign n26183 = x66 &  n25850 ;
  assign n26184 = ( n26182 & ~n26183 ) | ( n26182 & 1'b0 ) | ( ~n26183 & 1'b0 ) ;
  assign n26190 = ( n7535 & n25855 ) | ( n7535 & n26184 ) | ( n25855 & n26184 ) ;
  assign n26191 = ( n25855 & ~n25893 ) | ( n25855 & n26184 ) | ( ~n25893 & n26184 ) ;
  assign n26192 = ~n26190 & n26191 ;
  assign n26193 = n26189 | n26192 ;
  assign n26194 = n25854 &  n25894 ;
  assign n26195 = ( x65 & ~x25 ) | ( x65 & n25851 ) | ( ~x25 & n25851 ) ;
  assign n26196 = ( x25 & ~n25851 ) | ( x25 & x65 ) | ( ~n25851 & x65 ) ;
  assign n26197 = ( n26195 & ~x65 ) | ( n26195 & n26196 ) | ( ~x65 & n26196 ) ;
  assign n26198 = ( n7495 & ~n7535 ) | ( n7495 & n26197 ) | ( ~n7535 & n26197 ) ;
  assign n26199 = ( n7495 & n25893 ) | ( n7495 & n26197 ) | ( n25893 & n26197 ) ;
  assign n26200 = ( n26198 & ~n26199 ) | ( n26198 & 1'b0 ) | ( ~n26199 & 1'b0 ) ;
  assign n26201 = n26194 | n26200 ;
  assign n26202 = ( n7849 & ~n25893 ) | ( n7849 & 1'b0 ) | ( ~n25893 & 1'b0 ) ;
  assign n26203 = ( x24 & ~n26202 ) | ( x24 & 1'b0 ) | ( ~n26202 & 1'b0 ) ;
  assign n26204 = ( n7854 & ~n25893 ) | ( n7854 & 1'b0 ) | ( ~n25893 & 1'b0 ) ;
  assign n26205 = n26203 | n26204 ;
  assign n26206 = ( x65 & ~n26205 ) | ( x65 & n7857 ) | ( ~n26205 & n7857 ) ;
  assign n26207 = ( x66 & ~n26201 ) | ( x66 & n26206 ) | ( ~n26201 & n26206 ) ;
  assign n26208 = ( x67 & ~n26193 ) | ( x67 & n26207 ) | ( ~n26193 & n26207 ) ;
  assign n26209 = ( x68 & ~n26188 ) | ( x68 & n26208 ) | ( ~n26188 & n26208 ) ;
  assign n26210 = ( x69 & ~n26180 ) | ( x69 & n26209 ) | ( ~n26180 & n26209 ) ;
  assign n26211 = ( x70 & ~n26172 ) | ( x70 & n26210 ) | ( ~n26172 & n26210 ) ;
  assign n26212 = ( x71 & ~n26164 ) | ( x71 & n26211 ) | ( ~n26164 & n26211 ) ;
  assign n26213 = ( x72 & ~n26156 ) | ( x72 & n26212 ) | ( ~n26156 & n26212 ) ;
  assign n26214 = ( x73 & ~n26148 ) | ( x73 & n26213 ) | ( ~n26148 & n26213 ) ;
  assign n26215 = ( x74 & ~n26140 ) | ( x74 & n26214 ) | ( ~n26140 & n26214 ) ;
  assign n26216 = ( x75 & ~n26132 ) | ( x75 & n26215 ) | ( ~n26132 & n26215 ) ;
  assign n26217 = ( x76 & ~n26124 ) | ( x76 & n26216 ) | ( ~n26124 & n26216 ) ;
  assign n26218 = ( x77 & ~n26116 ) | ( x77 & n26217 ) | ( ~n26116 & n26217 ) ;
  assign n26219 = ( x78 & ~n26108 ) | ( x78 & n26218 ) | ( ~n26108 & n26218 ) ;
  assign n26220 = ( x79 & ~n26100 ) | ( x79 & n26219 ) | ( ~n26100 & n26219 ) ;
  assign n26221 = ( x80 & ~n26092 ) | ( x80 & n26220 ) | ( ~n26092 & n26220 ) ;
  assign n26222 = ( x81 & ~n26084 ) | ( x81 & n26221 ) | ( ~n26084 & n26221 ) ;
  assign n26223 = ( x82 & ~n26076 ) | ( x82 & n26222 ) | ( ~n26076 & n26222 ) ;
  assign n26224 = ( x83 & ~n26068 ) | ( x83 & n26223 ) | ( ~n26068 & n26223 ) ;
  assign n26225 = ( x84 & ~n26060 ) | ( x84 & n26224 ) | ( ~n26060 & n26224 ) ;
  assign n26226 = ( x85 & ~n26052 ) | ( x85 & n26225 ) | ( ~n26052 & n26225 ) ;
  assign n26227 = ( x86 & ~n26044 ) | ( x86 & n26226 ) | ( ~n26044 & n26226 ) ;
  assign n26228 = ( x87 & ~n26036 ) | ( x87 & n26227 ) | ( ~n26036 & n26227 ) ;
  assign n26229 = ( x88 & ~n26028 ) | ( x88 & n26228 ) | ( ~n26028 & n26228 ) ;
  assign n26230 = ( x89 & ~n26020 ) | ( x89 & n26229 ) | ( ~n26020 & n26229 ) ;
  assign n26231 = ( x90 & ~n26012 ) | ( x90 & n26230 ) | ( ~n26012 & n26230 ) ;
  assign n26232 = ( x91 & ~n26004 ) | ( x91 & n26231 ) | ( ~n26004 & n26231 ) ;
  assign n26233 = ( x92 & ~n25996 ) | ( x92 & n26232 ) | ( ~n25996 & n26232 ) ;
  assign n26234 = ( x93 & ~n25988 ) | ( x93 & n26233 ) | ( ~n25988 & n26233 ) ;
  assign n26235 = ( x94 & ~n25980 ) | ( x94 & n26234 ) | ( ~n25980 & n26234 ) ;
  assign n26236 = ( x95 & ~n25972 ) | ( x95 & n26235 ) | ( ~n25972 & n26235 ) ;
  assign n26237 = ( x96 & ~n25964 ) | ( x96 & n26236 ) | ( ~n25964 & n26236 ) ;
  assign n26238 = ( x97 & ~n25956 ) | ( x97 & n26237 ) | ( ~n25956 & n26237 ) ;
  assign n26239 = ( x98 & ~n25948 ) | ( x98 & n26238 ) | ( ~n25948 & n26238 ) ;
  assign n26240 = ( x99 & ~n25940 ) | ( x99 & n26239 ) | ( ~n25940 & n26239 ) ;
  assign n26241 = ( x100 & ~n25932 ) | ( x100 & n26240 ) | ( ~n25932 & n26240 ) ;
  assign n26242 = ( x101 & ~n25924 ) | ( x101 & n26241 ) | ( ~n25924 & n26241 ) ;
  assign n26243 = ( x102 & ~n25916 ) | ( x102 & n26242 ) | ( ~n25916 & n26242 ) ;
  assign n26244 = ( x103 & ~n25908 ) | ( x103 & n26243 ) | ( ~n25908 & n26243 ) ;
  assign n26245 = ( x104 & ~n25900 ) | ( x104 & n26244 ) | ( ~n25900 & n26244 ) ;
  assign n26246 = n7898 | n26245 ;
  assign n26247 = n25900 &  n26246 ;
  assign n26251 = ( n7898 & n25900 ) | ( n7898 & n26244 ) | ( n25900 & n26244 ) ;
  assign n26252 = ( x104 & ~n26251 ) | ( x104 & n25900 ) | ( ~n26251 & n25900 ) ;
  assign n26253 = ~x104 & n26252 ;
  assign n26254 = n26247 | n26253 ;
  assign n26255 = ~x105 & n26254 ;
  assign n26256 = n25908 &  n26246 ;
  assign n26248 = x103 | n25908 ;
  assign n26249 = x103 &  n25908 ;
  assign n26250 = ( n26248 & ~n26249 ) | ( n26248 & 1'b0 ) | ( ~n26249 & 1'b0 ) ;
  assign n26260 = ( n7898 & n26243 ) | ( n7898 & n26250 ) | ( n26243 & n26250 ) ;
  assign n26261 = ( n26243 & ~n26245 ) | ( n26243 & n26250 ) | ( ~n26245 & n26250 ) ;
  assign n26262 = ~n26260 & n26261 ;
  assign n26263 = n26256 | n26262 ;
  assign n26264 = n25916 &  n26246 ;
  assign n26257 = x102 | n25916 ;
  assign n26258 = x102 &  n25916 ;
  assign n26259 = ( n26257 & ~n26258 ) | ( n26257 & 1'b0 ) | ( ~n26258 & 1'b0 ) ;
  assign n26268 = ( n7898 & n26242 ) | ( n7898 & n26259 ) | ( n26242 & n26259 ) ;
  assign n26269 = ( n26242 & ~n26245 ) | ( n26242 & n26259 ) | ( ~n26245 & n26259 ) ;
  assign n26270 = ~n26268 & n26269 ;
  assign n26271 = n26264 | n26270 ;
  assign n26272 = n25924 &  n26246 ;
  assign n26265 = x101 | n25924 ;
  assign n26266 = x101 &  n25924 ;
  assign n26267 = ( n26265 & ~n26266 ) | ( n26265 & 1'b0 ) | ( ~n26266 & 1'b0 ) ;
  assign n26276 = ( n7898 & n26241 ) | ( n7898 & n26267 ) | ( n26241 & n26267 ) ;
  assign n26277 = ( n26241 & ~n26245 ) | ( n26241 & n26267 ) | ( ~n26245 & n26267 ) ;
  assign n26278 = ~n26276 & n26277 ;
  assign n26279 = n26272 | n26278 ;
  assign n26280 = n25932 &  n26246 ;
  assign n26273 = x100 | n25932 ;
  assign n26274 = x100 &  n25932 ;
  assign n26275 = ( n26273 & ~n26274 ) | ( n26273 & 1'b0 ) | ( ~n26274 & 1'b0 ) ;
  assign n26284 = ( n7898 & n26240 ) | ( n7898 & n26275 ) | ( n26240 & n26275 ) ;
  assign n26285 = ( n26240 & ~n26245 ) | ( n26240 & n26275 ) | ( ~n26245 & n26275 ) ;
  assign n26286 = ~n26284 & n26285 ;
  assign n26287 = n26280 | n26286 ;
  assign n26288 = n25940 &  n26246 ;
  assign n26281 = x99 | n25940 ;
  assign n26282 = x99 &  n25940 ;
  assign n26283 = ( n26281 & ~n26282 ) | ( n26281 & 1'b0 ) | ( ~n26282 & 1'b0 ) ;
  assign n26292 = ( n7898 & n26239 ) | ( n7898 & n26283 ) | ( n26239 & n26283 ) ;
  assign n26293 = ( n26239 & ~n26245 ) | ( n26239 & n26283 ) | ( ~n26245 & n26283 ) ;
  assign n26294 = ~n26292 & n26293 ;
  assign n26295 = n26288 | n26294 ;
  assign n26296 = n25948 &  n26246 ;
  assign n26289 = x98 | n25948 ;
  assign n26290 = x98 &  n25948 ;
  assign n26291 = ( n26289 & ~n26290 ) | ( n26289 & 1'b0 ) | ( ~n26290 & 1'b0 ) ;
  assign n26300 = ( n7898 & n26238 ) | ( n7898 & n26291 ) | ( n26238 & n26291 ) ;
  assign n26301 = ( n26238 & ~n26245 ) | ( n26238 & n26291 ) | ( ~n26245 & n26291 ) ;
  assign n26302 = ~n26300 & n26301 ;
  assign n26303 = n26296 | n26302 ;
  assign n26304 = n25956 &  n26246 ;
  assign n26297 = x97 | n25956 ;
  assign n26298 = x97 &  n25956 ;
  assign n26299 = ( n26297 & ~n26298 ) | ( n26297 & 1'b0 ) | ( ~n26298 & 1'b0 ) ;
  assign n26308 = ( n7898 & n26237 ) | ( n7898 & n26299 ) | ( n26237 & n26299 ) ;
  assign n26309 = ( n26237 & ~n26245 ) | ( n26237 & n26299 ) | ( ~n26245 & n26299 ) ;
  assign n26310 = ~n26308 & n26309 ;
  assign n26311 = n26304 | n26310 ;
  assign n26312 = n25964 &  n26246 ;
  assign n26305 = x96 | n25964 ;
  assign n26306 = x96 &  n25964 ;
  assign n26307 = ( n26305 & ~n26306 ) | ( n26305 & 1'b0 ) | ( ~n26306 & 1'b0 ) ;
  assign n26316 = ( n7898 & n26236 ) | ( n7898 & n26307 ) | ( n26236 & n26307 ) ;
  assign n26317 = ( n26236 & ~n26245 ) | ( n26236 & n26307 ) | ( ~n26245 & n26307 ) ;
  assign n26318 = ~n26316 & n26317 ;
  assign n26319 = n26312 | n26318 ;
  assign n26320 = n25972 &  n26246 ;
  assign n26313 = x95 | n25972 ;
  assign n26314 = x95 &  n25972 ;
  assign n26315 = ( n26313 & ~n26314 ) | ( n26313 & 1'b0 ) | ( ~n26314 & 1'b0 ) ;
  assign n26324 = ( n7898 & n26235 ) | ( n7898 & n26315 ) | ( n26235 & n26315 ) ;
  assign n26325 = ( n26235 & ~n26245 ) | ( n26235 & n26315 ) | ( ~n26245 & n26315 ) ;
  assign n26326 = ~n26324 & n26325 ;
  assign n26327 = n26320 | n26326 ;
  assign n26328 = n25980 &  n26246 ;
  assign n26321 = x94 | n25980 ;
  assign n26322 = x94 &  n25980 ;
  assign n26323 = ( n26321 & ~n26322 ) | ( n26321 & 1'b0 ) | ( ~n26322 & 1'b0 ) ;
  assign n26332 = ( n7898 & n26234 ) | ( n7898 & n26323 ) | ( n26234 & n26323 ) ;
  assign n26333 = ( n26234 & ~n26245 ) | ( n26234 & n26323 ) | ( ~n26245 & n26323 ) ;
  assign n26334 = ~n26332 & n26333 ;
  assign n26335 = n26328 | n26334 ;
  assign n26336 = n25988 &  n26246 ;
  assign n26329 = x93 | n25988 ;
  assign n26330 = x93 &  n25988 ;
  assign n26331 = ( n26329 & ~n26330 ) | ( n26329 & 1'b0 ) | ( ~n26330 & 1'b0 ) ;
  assign n26340 = ( n7898 & n26233 ) | ( n7898 & n26331 ) | ( n26233 & n26331 ) ;
  assign n26341 = ( n26233 & ~n26245 ) | ( n26233 & n26331 ) | ( ~n26245 & n26331 ) ;
  assign n26342 = ~n26340 & n26341 ;
  assign n26343 = n26336 | n26342 ;
  assign n26344 = n25996 &  n26246 ;
  assign n26337 = x92 | n25996 ;
  assign n26338 = x92 &  n25996 ;
  assign n26339 = ( n26337 & ~n26338 ) | ( n26337 & 1'b0 ) | ( ~n26338 & 1'b0 ) ;
  assign n26348 = ( n7898 & n26232 ) | ( n7898 & n26339 ) | ( n26232 & n26339 ) ;
  assign n26349 = ( n26232 & ~n26245 ) | ( n26232 & n26339 ) | ( ~n26245 & n26339 ) ;
  assign n26350 = ~n26348 & n26349 ;
  assign n26351 = n26344 | n26350 ;
  assign n26352 = n26004 &  n26246 ;
  assign n26345 = x91 | n26004 ;
  assign n26346 = x91 &  n26004 ;
  assign n26347 = ( n26345 & ~n26346 ) | ( n26345 & 1'b0 ) | ( ~n26346 & 1'b0 ) ;
  assign n26356 = ( n7898 & n26231 ) | ( n7898 & n26347 ) | ( n26231 & n26347 ) ;
  assign n26357 = ( n26231 & ~n26245 ) | ( n26231 & n26347 ) | ( ~n26245 & n26347 ) ;
  assign n26358 = ~n26356 & n26357 ;
  assign n26359 = n26352 | n26358 ;
  assign n26360 = n26012 &  n26246 ;
  assign n26353 = x90 | n26012 ;
  assign n26354 = x90 &  n26012 ;
  assign n26355 = ( n26353 & ~n26354 ) | ( n26353 & 1'b0 ) | ( ~n26354 & 1'b0 ) ;
  assign n26364 = ( n7898 & n26230 ) | ( n7898 & n26355 ) | ( n26230 & n26355 ) ;
  assign n26365 = ( n26230 & ~n26245 ) | ( n26230 & n26355 ) | ( ~n26245 & n26355 ) ;
  assign n26366 = ~n26364 & n26365 ;
  assign n26367 = n26360 | n26366 ;
  assign n26368 = n26020 &  n26246 ;
  assign n26361 = x89 | n26020 ;
  assign n26362 = x89 &  n26020 ;
  assign n26363 = ( n26361 & ~n26362 ) | ( n26361 & 1'b0 ) | ( ~n26362 & 1'b0 ) ;
  assign n26372 = ( n7898 & n26229 ) | ( n7898 & n26363 ) | ( n26229 & n26363 ) ;
  assign n26373 = ( n26229 & ~n26245 ) | ( n26229 & n26363 ) | ( ~n26245 & n26363 ) ;
  assign n26374 = ~n26372 & n26373 ;
  assign n26375 = n26368 | n26374 ;
  assign n26376 = n26028 &  n26246 ;
  assign n26369 = x88 | n26028 ;
  assign n26370 = x88 &  n26028 ;
  assign n26371 = ( n26369 & ~n26370 ) | ( n26369 & 1'b0 ) | ( ~n26370 & 1'b0 ) ;
  assign n26380 = ( n7898 & n26228 ) | ( n7898 & n26371 ) | ( n26228 & n26371 ) ;
  assign n26381 = ( n26228 & ~n26245 ) | ( n26228 & n26371 ) | ( ~n26245 & n26371 ) ;
  assign n26382 = ~n26380 & n26381 ;
  assign n26383 = n26376 | n26382 ;
  assign n26384 = n26036 &  n26246 ;
  assign n26377 = x87 | n26036 ;
  assign n26378 = x87 &  n26036 ;
  assign n26379 = ( n26377 & ~n26378 ) | ( n26377 & 1'b0 ) | ( ~n26378 & 1'b0 ) ;
  assign n26388 = ( n7898 & n26227 ) | ( n7898 & n26379 ) | ( n26227 & n26379 ) ;
  assign n26389 = ( n26227 & ~n26245 ) | ( n26227 & n26379 ) | ( ~n26245 & n26379 ) ;
  assign n26390 = ~n26388 & n26389 ;
  assign n26391 = n26384 | n26390 ;
  assign n26392 = n26044 &  n26246 ;
  assign n26385 = x86 | n26044 ;
  assign n26386 = x86 &  n26044 ;
  assign n26387 = ( n26385 & ~n26386 ) | ( n26385 & 1'b0 ) | ( ~n26386 & 1'b0 ) ;
  assign n26396 = ( n7898 & n26226 ) | ( n7898 & n26387 ) | ( n26226 & n26387 ) ;
  assign n26397 = ( n26226 & ~n26245 ) | ( n26226 & n26387 ) | ( ~n26245 & n26387 ) ;
  assign n26398 = ~n26396 & n26397 ;
  assign n26399 = n26392 | n26398 ;
  assign n26400 = n26052 &  n26246 ;
  assign n26393 = x85 | n26052 ;
  assign n26394 = x85 &  n26052 ;
  assign n26395 = ( n26393 & ~n26394 ) | ( n26393 & 1'b0 ) | ( ~n26394 & 1'b0 ) ;
  assign n26404 = ( n7898 & n26225 ) | ( n7898 & n26395 ) | ( n26225 & n26395 ) ;
  assign n26405 = ( n26225 & ~n26245 ) | ( n26225 & n26395 ) | ( ~n26245 & n26395 ) ;
  assign n26406 = ~n26404 & n26405 ;
  assign n26407 = n26400 | n26406 ;
  assign n26408 = n26060 &  n26246 ;
  assign n26401 = x84 | n26060 ;
  assign n26402 = x84 &  n26060 ;
  assign n26403 = ( n26401 & ~n26402 ) | ( n26401 & 1'b0 ) | ( ~n26402 & 1'b0 ) ;
  assign n26412 = ( n7898 & n26224 ) | ( n7898 & n26403 ) | ( n26224 & n26403 ) ;
  assign n26413 = ( n26224 & ~n26245 ) | ( n26224 & n26403 ) | ( ~n26245 & n26403 ) ;
  assign n26414 = ~n26412 & n26413 ;
  assign n26415 = n26408 | n26414 ;
  assign n26416 = n26068 &  n26246 ;
  assign n26409 = x83 | n26068 ;
  assign n26410 = x83 &  n26068 ;
  assign n26411 = ( n26409 & ~n26410 ) | ( n26409 & 1'b0 ) | ( ~n26410 & 1'b0 ) ;
  assign n26420 = ( n7898 & n26223 ) | ( n7898 & n26411 ) | ( n26223 & n26411 ) ;
  assign n26421 = ( n26223 & ~n26245 ) | ( n26223 & n26411 ) | ( ~n26245 & n26411 ) ;
  assign n26422 = ~n26420 & n26421 ;
  assign n26423 = n26416 | n26422 ;
  assign n26424 = n26076 &  n26246 ;
  assign n26417 = x82 | n26076 ;
  assign n26418 = x82 &  n26076 ;
  assign n26419 = ( n26417 & ~n26418 ) | ( n26417 & 1'b0 ) | ( ~n26418 & 1'b0 ) ;
  assign n26428 = ( n7898 & n26222 ) | ( n7898 & n26419 ) | ( n26222 & n26419 ) ;
  assign n26429 = ( n26222 & ~n26245 ) | ( n26222 & n26419 ) | ( ~n26245 & n26419 ) ;
  assign n26430 = ~n26428 & n26429 ;
  assign n26431 = n26424 | n26430 ;
  assign n26432 = n26084 &  n26246 ;
  assign n26425 = x81 | n26084 ;
  assign n26426 = x81 &  n26084 ;
  assign n26427 = ( n26425 & ~n26426 ) | ( n26425 & 1'b0 ) | ( ~n26426 & 1'b0 ) ;
  assign n26436 = ( n7898 & n26221 ) | ( n7898 & n26427 ) | ( n26221 & n26427 ) ;
  assign n26437 = ( n26221 & ~n26245 ) | ( n26221 & n26427 ) | ( ~n26245 & n26427 ) ;
  assign n26438 = ~n26436 & n26437 ;
  assign n26439 = n26432 | n26438 ;
  assign n26440 = n26092 &  n26246 ;
  assign n26433 = x80 | n26092 ;
  assign n26434 = x80 &  n26092 ;
  assign n26435 = ( n26433 & ~n26434 ) | ( n26433 & 1'b0 ) | ( ~n26434 & 1'b0 ) ;
  assign n26444 = ( n7898 & n26220 ) | ( n7898 & n26435 ) | ( n26220 & n26435 ) ;
  assign n26445 = ( n26220 & ~n26245 ) | ( n26220 & n26435 ) | ( ~n26245 & n26435 ) ;
  assign n26446 = ~n26444 & n26445 ;
  assign n26447 = n26440 | n26446 ;
  assign n26448 = n26100 &  n26246 ;
  assign n26441 = x79 | n26100 ;
  assign n26442 = x79 &  n26100 ;
  assign n26443 = ( n26441 & ~n26442 ) | ( n26441 & 1'b0 ) | ( ~n26442 & 1'b0 ) ;
  assign n26452 = ( n7898 & n26219 ) | ( n7898 & n26443 ) | ( n26219 & n26443 ) ;
  assign n26453 = ( n26219 & ~n26245 ) | ( n26219 & n26443 ) | ( ~n26245 & n26443 ) ;
  assign n26454 = ~n26452 & n26453 ;
  assign n26455 = n26448 | n26454 ;
  assign n26456 = n26108 &  n26246 ;
  assign n26449 = x78 | n26108 ;
  assign n26450 = x78 &  n26108 ;
  assign n26451 = ( n26449 & ~n26450 ) | ( n26449 & 1'b0 ) | ( ~n26450 & 1'b0 ) ;
  assign n26460 = ( n7898 & n26218 ) | ( n7898 & n26451 ) | ( n26218 & n26451 ) ;
  assign n26461 = ( n26218 & ~n26245 ) | ( n26218 & n26451 ) | ( ~n26245 & n26451 ) ;
  assign n26462 = ~n26460 & n26461 ;
  assign n26463 = n26456 | n26462 ;
  assign n26464 = n26116 &  n26246 ;
  assign n26457 = x77 | n26116 ;
  assign n26458 = x77 &  n26116 ;
  assign n26459 = ( n26457 & ~n26458 ) | ( n26457 & 1'b0 ) | ( ~n26458 & 1'b0 ) ;
  assign n26468 = ( n7898 & n26217 ) | ( n7898 & n26459 ) | ( n26217 & n26459 ) ;
  assign n26469 = ( n26217 & ~n26245 ) | ( n26217 & n26459 ) | ( ~n26245 & n26459 ) ;
  assign n26470 = ~n26468 & n26469 ;
  assign n26471 = n26464 | n26470 ;
  assign n26472 = n26124 &  n26246 ;
  assign n26465 = x76 | n26124 ;
  assign n26466 = x76 &  n26124 ;
  assign n26467 = ( n26465 & ~n26466 ) | ( n26465 & 1'b0 ) | ( ~n26466 & 1'b0 ) ;
  assign n26476 = ( n7898 & n26216 ) | ( n7898 & n26467 ) | ( n26216 & n26467 ) ;
  assign n26477 = ( n26216 & ~n26245 ) | ( n26216 & n26467 ) | ( ~n26245 & n26467 ) ;
  assign n26478 = ~n26476 & n26477 ;
  assign n26479 = n26472 | n26478 ;
  assign n26480 = n26132 &  n26246 ;
  assign n26473 = x75 | n26132 ;
  assign n26474 = x75 &  n26132 ;
  assign n26475 = ( n26473 & ~n26474 ) | ( n26473 & 1'b0 ) | ( ~n26474 & 1'b0 ) ;
  assign n26484 = ( n7898 & n26215 ) | ( n7898 & n26475 ) | ( n26215 & n26475 ) ;
  assign n26485 = ( n26215 & ~n26245 ) | ( n26215 & n26475 ) | ( ~n26245 & n26475 ) ;
  assign n26486 = ~n26484 & n26485 ;
  assign n26487 = n26480 | n26486 ;
  assign n26488 = n26140 &  n26246 ;
  assign n26481 = x74 | n26140 ;
  assign n26482 = x74 &  n26140 ;
  assign n26483 = ( n26481 & ~n26482 ) | ( n26481 & 1'b0 ) | ( ~n26482 & 1'b0 ) ;
  assign n26492 = ( n7898 & n26214 ) | ( n7898 & n26483 ) | ( n26214 & n26483 ) ;
  assign n26493 = ( n26214 & ~n26245 ) | ( n26214 & n26483 ) | ( ~n26245 & n26483 ) ;
  assign n26494 = ~n26492 & n26493 ;
  assign n26495 = n26488 | n26494 ;
  assign n26496 = n26148 &  n26246 ;
  assign n26489 = x73 | n26148 ;
  assign n26490 = x73 &  n26148 ;
  assign n26491 = ( n26489 & ~n26490 ) | ( n26489 & 1'b0 ) | ( ~n26490 & 1'b0 ) ;
  assign n26500 = ( n7898 & n26213 ) | ( n7898 & n26491 ) | ( n26213 & n26491 ) ;
  assign n26501 = ( n26213 & ~n26245 ) | ( n26213 & n26491 ) | ( ~n26245 & n26491 ) ;
  assign n26502 = ~n26500 & n26501 ;
  assign n26503 = n26496 | n26502 ;
  assign n26504 = n26156 &  n26246 ;
  assign n26497 = x72 | n26156 ;
  assign n26498 = x72 &  n26156 ;
  assign n26499 = ( n26497 & ~n26498 ) | ( n26497 & 1'b0 ) | ( ~n26498 & 1'b0 ) ;
  assign n26508 = ( n7898 & n26212 ) | ( n7898 & n26499 ) | ( n26212 & n26499 ) ;
  assign n26509 = ( n26212 & ~n26245 ) | ( n26212 & n26499 ) | ( ~n26245 & n26499 ) ;
  assign n26510 = ~n26508 & n26509 ;
  assign n26511 = n26504 | n26510 ;
  assign n26512 = n26164 &  n26246 ;
  assign n26505 = x71 | n26164 ;
  assign n26506 = x71 &  n26164 ;
  assign n26507 = ( n26505 & ~n26506 ) | ( n26505 & 1'b0 ) | ( ~n26506 & 1'b0 ) ;
  assign n26516 = ( n7898 & n26211 ) | ( n7898 & n26507 ) | ( n26211 & n26507 ) ;
  assign n26517 = ( n26211 & ~n26245 ) | ( n26211 & n26507 ) | ( ~n26245 & n26507 ) ;
  assign n26518 = ~n26516 & n26517 ;
  assign n26519 = n26512 | n26518 ;
  assign n26520 = n26172 &  n26246 ;
  assign n26513 = x70 | n26172 ;
  assign n26514 = x70 &  n26172 ;
  assign n26515 = ( n26513 & ~n26514 ) | ( n26513 & 1'b0 ) | ( ~n26514 & 1'b0 ) ;
  assign n26524 = ( n7898 & n26210 ) | ( n7898 & n26515 ) | ( n26210 & n26515 ) ;
  assign n26525 = ( n26210 & ~n26245 ) | ( n26210 & n26515 ) | ( ~n26245 & n26515 ) ;
  assign n26526 = ~n26524 & n26525 ;
  assign n26527 = n26520 | n26526 ;
  assign n26528 = n26180 &  n26246 ;
  assign n26521 = x69 | n26180 ;
  assign n26522 = x69 &  n26180 ;
  assign n26523 = ( n26521 & ~n26522 ) | ( n26521 & 1'b0 ) | ( ~n26522 & 1'b0 ) ;
  assign n26532 = ( n7898 & n26209 ) | ( n7898 & n26523 ) | ( n26209 & n26523 ) ;
  assign n26533 = ( n26209 & ~n26245 ) | ( n26209 & n26523 ) | ( ~n26245 & n26523 ) ;
  assign n26534 = ~n26532 & n26533 ;
  assign n26535 = n26528 | n26534 ;
  assign n26536 = n26188 &  n26246 ;
  assign n26529 = x68 | n26188 ;
  assign n26530 = x68 &  n26188 ;
  assign n26531 = ( n26529 & ~n26530 ) | ( n26529 & 1'b0 ) | ( ~n26530 & 1'b0 ) ;
  assign n26540 = ( n7898 & n26208 ) | ( n7898 & n26531 ) | ( n26208 & n26531 ) ;
  assign n26541 = ( n26208 & ~n26245 ) | ( n26208 & n26531 ) | ( ~n26245 & n26531 ) ;
  assign n26542 = ~n26540 & n26541 ;
  assign n26543 = n26536 | n26542 ;
  assign n26544 = n26193 &  n26246 ;
  assign n26537 = x67 | n26193 ;
  assign n26538 = x67 &  n26193 ;
  assign n26539 = ( n26537 & ~n26538 ) | ( n26537 & 1'b0 ) | ( ~n26538 & 1'b0 ) ;
  assign n26548 = ( n7898 & n26207 ) | ( n7898 & n26539 ) | ( n26207 & n26539 ) ;
  assign n26549 = ( n26207 & ~n26245 ) | ( n26207 & n26539 ) | ( ~n26245 & n26539 ) ;
  assign n26550 = ~n26548 & n26549 ;
  assign n26551 = n26544 | n26550 ;
  assign n26552 = n26201 &  n26246 ;
  assign n26545 = x66 | n26201 ;
  assign n26546 = x66 &  n26201 ;
  assign n26547 = ( n26545 & ~n26546 ) | ( n26545 & 1'b0 ) | ( ~n26546 & 1'b0 ) ;
  assign n26556 = ( n7898 & n26206 ) | ( n7898 & n26547 ) | ( n26206 & n26547 ) ;
  assign n26557 = ( n26206 & ~n26245 ) | ( n26206 & n26547 ) | ( ~n26245 & n26547 ) ;
  assign n26558 = ~n26556 & n26557 ;
  assign n26559 = n26552 | n26558 ;
  assign n26560 = n26205 &  n26246 ;
  assign n26553 = x65 &  n26205 ;
  assign n26554 = x65 | n26204 ;
  assign n26555 = n26203 | n26554 ;
  assign n26561 = ~n26553 & n26555 ;
  assign n26562 = ( n7857 & ~n7898 ) | ( n7857 & n26561 ) | ( ~n7898 & n26561 ) ;
  assign n26563 = ( n7857 & n26245 ) | ( n7857 & n26561 ) | ( n26245 & n26561 ) ;
  assign n26564 = ( n26562 & ~n26563 ) | ( n26562 & 1'b0 ) | ( ~n26563 & 1'b0 ) ;
  assign n26565 = n26560 | n26564 ;
  assign n26566 = ( n8097 & ~n26245 ) | ( n8097 & 1'b0 ) | ( ~n26245 & 1'b0 ) ;
  assign n26567 = ( x23 & ~n26566 ) | ( x23 & 1'b0 ) | ( ~n26566 & 1'b0 ) ;
  assign n26568 = ( n8102 & ~n26245 ) | ( n8102 & 1'b0 ) | ( ~n26245 & 1'b0 ) ;
  assign n26569 = n26567 | n26568 ;
  assign n26570 = ( x65 & ~n26569 ) | ( x65 & n8105 ) | ( ~n26569 & n8105 ) ;
  assign n26571 = ( x66 & ~n26565 ) | ( x66 & n26570 ) | ( ~n26565 & n26570 ) ;
  assign n26572 = ( x67 & ~n26559 ) | ( x67 & n26571 ) | ( ~n26559 & n26571 ) ;
  assign n26573 = ( x68 & ~n26551 ) | ( x68 & n26572 ) | ( ~n26551 & n26572 ) ;
  assign n26574 = ( x69 & ~n26543 ) | ( x69 & n26573 ) | ( ~n26543 & n26573 ) ;
  assign n26575 = ( x70 & ~n26535 ) | ( x70 & n26574 ) | ( ~n26535 & n26574 ) ;
  assign n26576 = ( x71 & ~n26527 ) | ( x71 & n26575 ) | ( ~n26527 & n26575 ) ;
  assign n26577 = ( x72 & ~n26519 ) | ( x72 & n26576 ) | ( ~n26519 & n26576 ) ;
  assign n26578 = ( x73 & ~n26511 ) | ( x73 & n26577 ) | ( ~n26511 & n26577 ) ;
  assign n26579 = ( x74 & ~n26503 ) | ( x74 & n26578 ) | ( ~n26503 & n26578 ) ;
  assign n26580 = ( x75 & ~n26495 ) | ( x75 & n26579 ) | ( ~n26495 & n26579 ) ;
  assign n26581 = ( x76 & ~n26487 ) | ( x76 & n26580 ) | ( ~n26487 & n26580 ) ;
  assign n26582 = ( x77 & ~n26479 ) | ( x77 & n26581 ) | ( ~n26479 & n26581 ) ;
  assign n26583 = ( x78 & ~n26471 ) | ( x78 & n26582 ) | ( ~n26471 & n26582 ) ;
  assign n26584 = ( x79 & ~n26463 ) | ( x79 & n26583 ) | ( ~n26463 & n26583 ) ;
  assign n26585 = ( x80 & ~n26455 ) | ( x80 & n26584 ) | ( ~n26455 & n26584 ) ;
  assign n26586 = ( x81 & ~n26447 ) | ( x81 & n26585 ) | ( ~n26447 & n26585 ) ;
  assign n26587 = ( x82 & ~n26439 ) | ( x82 & n26586 ) | ( ~n26439 & n26586 ) ;
  assign n26588 = ( x83 & ~n26431 ) | ( x83 & n26587 ) | ( ~n26431 & n26587 ) ;
  assign n26589 = ( x84 & ~n26423 ) | ( x84 & n26588 ) | ( ~n26423 & n26588 ) ;
  assign n26590 = ( x85 & ~n26415 ) | ( x85 & n26589 ) | ( ~n26415 & n26589 ) ;
  assign n26591 = ( x86 & ~n26407 ) | ( x86 & n26590 ) | ( ~n26407 & n26590 ) ;
  assign n26592 = ( x87 & ~n26399 ) | ( x87 & n26591 ) | ( ~n26399 & n26591 ) ;
  assign n26593 = ( x88 & ~n26391 ) | ( x88 & n26592 ) | ( ~n26391 & n26592 ) ;
  assign n26594 = ( x89 & ~n26383 ) | ( x89 & n26593 ) | ( ~n26383 & n26593 ) ;
  assign n26595 = ( x90 & ~n26375 ) | ( x90 & n26594 ) | ( ~n26375 & n26594 ) ;
  assign n26596 = ( x91 & ~n26367 ) | ( x91 & n26595 ) | ( ~n26367 & n26595 ) ;
  assign n26597 = ( x92 & ~n26359 ) | ( x92 & n26596 ) | ( ~n26359 & n26596 ) ;
  assign n26598 = ( x93 & ~n26351 ) | ( x93 & n26597 ) | ( ~n26351 & n26597 ) ;
  assign n26599 = ( x94 & ~n26343 ) | ( x94 & n26598 ) | ( ~n26343 & n26598 ) ;
  assign n26600 = ( x95 & ~n26335 ) | ( x95 & n26599 ) | ( ~n26335 & n26599 ) ;
  assign n26601 = ( x96 & ~n26327 ) | ( x96 & n26600 ) | ( ~n26327 & n26600 ) ;
  assign n26602 = ( x97 & ~n26319 ) | ( x97 & n26601 ) | ( ~n26319 & n26601 ) ;
  assign n26603 = ( x98 & ~n26311 ) | ( x98 & n26602 ) | ( ~n26311 & n26602 ) ;
  assign n26604 = ( x99 & ~n26303 ) | ( x99 & n26603 ) | ( ~n26303 & n26603 ) ;
  assign n26605 = ( x100 & ~n26295 ) | ( x100 & n26604 ) | ( ~n26295 & n26604 ) ;
  assign n26606 = ( x101 & ~n26287 ) | ( x101 & n26605 ) | ( ~n26287 & n26605 ) ;
  assign n26607 = ( x102 & ~n26279 ) | ( x102 & n26606 ) | ( ~n26279 & n26606 ) ;
  assign n26608 = ( x103 & ~n26271 ) | ( x103 & n26607 ) | ( ~n26271 & n26607 ) ;
  assign n26609 = ( x104 & ~n26263 ) | ( x104 & n26608 ) | ( ~n26263 & n26608 ) ;
  assign n26610 = ( x105 & ~n26247 ) | ( x105 & 1'b0 ) | ( ~n26247 & 1'b0 ) ;
  assign n26611 = ~n26253 & n26610 ;
  assign n26612 = ( n26609 & ~n26255 ) | ( n26609 & n26611 ) | ( ~n26255 & n26611 ) ;
  assign n26613 = ( n26255 & ~n8276 ) | ( n26255 & n26612 ) | ( ~n8276 & n26612 ) ;
  assign n26614 = n8276 | n26613 ;
  assign n26615 = ~n26254 |  n7898 ;
  assign n26629 = n26263 &  n26615 ;
  assign n26630 = n26614 &  n26629 ;
  assign n26616 = n26614 &  n26615 ;
  assign n26617 = x104 | n26263 ;
  assign n26618 = x104 &  n26263 ;
  assign n26619 = ( n26617 & ~n26618 ) | ( n26617 & 1'b0 ) | ( ~n26618 & 1'b0 ) ;
  assign n26632 = ( n26608 & n26616 ) | ( n26608 & n26619 ) | ( n26616 & n26619 ) ;
  assign n26631 = n26608 | n26619 ;
  assign n26633 = ( n26630 & ~n26632 ) | ( n26630 & n26631 ) | ( ~n26632 & n26631 ) ;
  assign n26621 = n7898 &  n25900 ;
  assign n26622 = n26614 &  n26621 ;
  assign n26620 = n26255 | n26611 ;
  assign n26624 = ( n26609 & n26616 ) | ( n26609 & n26620 ) | ( n26616 & n26620 ) ;
  assign n26623 = n26609 | n26620 ;
  assign n26625 = ( n26622 & ~n26624 ) | ( n26622 & n26623 ) | ( ~n26624 & n26623 ) ;
  assign n26637 = n26271 &  n26615 ;
  assign n26638 = n26614 &  n26637 ;
  assign n26626 = x103 | n26271 ;
  assign n26627 = x103 &  n26271 ;
  assign n26628 = ( n26626 & ~n26627 ) | ( n26626 & 1'b0 ) | ( ~n26627 & 1'b0 ) ;
  assign n26640 = ( n26607 & n26616 ) | ( n26607 & n26628 ) | ( n26616 & n26628 ) ;
  assign n26639 = n26607 | n26628 ;
  assign n26641 = ( n26638 & ~n26640 ) | ( n26638 & n26639 ) | ( ~n26640 & n26639 ) ;
  assign n26645 = n26279 &  n26615 ;
  assign n26646 = n26614 &  n26645 ;
  assign n26634 = x102 | n26279 ;
  assign n26635 = x102 &  n26279 ;
  assign n26636 = ( n26634 & ~n26635 ) | ( n26634 & 1'b0 ) | ( ~n26635 & 1'b0 ) ;
  assign n26648 = ( n26606 & n26616 ) | ( n26606 & n26636 ) | ( n26616 & n26636 ) ;
  assign n26647 = n26606 | n26636 ;
  assign n26649 = ( n26646 & ~n26648 ) | ( n26646 & n26647 ) | ( ~n26648 & n26647 ) ;
  assign n26653 = n26287 &  n26615 ;
  assign n26654 = n26614 &  n26653 ;
  assign n26642 = x101 | n26287 ;
  assign n26643 = x101 &  n26287 ;
  assign n26644 = ( n26642 & ~n26643 ) | ( n26642 & 1'b0 ) | ( ~n26643 & 1'b0 ) ;
  assign n26656 = ( n26605 & n26616 ) | ( n26605 & n26644 ) | ( n26616 & n26644 ) ;
  assign n26655 = n26605 | n26644 ;
  assign n26657 = ( n26654 & ~n26656 ) | ( n26654 & n26655 ) | ( ~n26656 & n26655 ) ;
  assign n26661 = n26295 &  n26615 ;
  assign n26662 = n26614 &  n26661 ;
  assign n26650 = x100 | n26295 ;
  assign n26651 = x100 &  n26295 ;
  assign n26652 = ( n26650 & ~n26651 ) | ( n26650 & 1'b0 ) | ( ~n26651 & 1'b0 ) ;
  assign n26664 = ( n26604 & n26616 ) | ( n26604 & n26652 ) | ( n26616 & n26652 ) ;
  assign n26663 = n26604 | n26652 ;
  assign n26665 = ( n26662 & ~n26664 ) | ( n26662 & n26663 ) | ( ~n26664 & n26663 ) ;
  assign n26669 = n26303 &  n26615 ;
  assign n26670 = n26614 &  n26669 ;
  assign n26658 = x99 | n26303 ;
  assign n26659 = x99 &  n26303 ;
  assign n26660 = ( n26658 & ~n26659 ) | ( n26658 & 1'b0 ) | ( ~n26659 & 1'b0 ) ;
  assign n26672 = ( n26603 & n26616 ) | ( n26603 & n26660 ) | ( n26616 & n26660 ) ;
  assign n26671 = n26603 | n26660 ;
  assign n26673 = ( n26670 & ~n26672 ) | ( n26670 & n26671 ) | ( ~n26672 & n26671 ) ;
  assign n26677 = n26311 &  n26615 ;
  assign n26678 = n26614 &  n26677 ;
  assign n26666 = x98 | n26311 ;
  assign n26667 = x98 &  n26311 ;
  assign n26668 = ( n26666 & ~n26667 ) | ( n26666 & 1'b0 ) | ( ~n26667 & 1'b0 ) ;
  assign n26680 = ( n26602 & n26616 ) | ( n26602 & n26668 ) | ( n26616 & n26668 ) ;
  assign n26679 = n26602 | n26668 ;
  assign n26681 = ( n26678 & ~n26680 ) | ( n26678 & n26679 ) | ( ~n26680 & n26679 ) ;
  assign n26685 = n26319 &  n26615 ;
  assign n26686 = n26614 &  n26685 ;
  assign n26674 = x97 | n26319 ;
  assign n26675 = x97 &  n26319 ;
  assign n26676 = ( n26674 & ~n26675 ) | ( n26674 & 1'b0 ) | ( ~n26675 & 1'b0 ) ;
  assign n26688 = ( n26601 & n26616 ) | ( n26601 & n26676 ) | ( n26616 & n26676 ) ;
  assign n26687 = n26601 | n26676 ;
  assign n26689 = ( n26686 & ~n26688 ) | ( n26686 & n26687 ) | ( ~n26688 & n26687 ) ;
  assign n26693 = n26327 &  n26615 ;
  assign n26694 = n26614 &  n26693 ;
  assign n26682 = x96 | n26327 ;
  assign n26683 = x96 &  n26327 ;
  assign n26684 = ( n26682 & ~n26683 ) | ( n26682 & 1'b0 ) | ( ~n26683 & 1'b0 ) ;
  assign n26696 = ( n26600 & n26616 ) | ( n26600 & n26684 ) | ( n26616 & n26684 ) ;
  assign n26695 = n26600 | n26684 ;
  assign n26697 = ( n26694 & ~n26696 ) | ( n26694 & n26695 ) | ( ~n26696 & n26695 ) ;
  assign n26701 = n26335 &  n26615 ;
  assign n26702 = n26614 &  n26701 ;
  assign n26690 = x95 | n26335 ;
  assign n26691 = x95 &  n26335 ;
  assign n26692 = ( n26690 & ~n26691 ) | ( n26690 & 1'b0 ) | ( ~n26691 & 1'b0 ) ;
  assign n26704 = ( n26599 & n26616 ) | ( n26599 & n26692 ) | ( n26616 & n26692 ) ;
  assign n26703 = n26599 | n26692 ;
  assign n26705 = ( n26702 & ~n26704 ) | ( n26702 & n26703 ) | ( ~n26704 & n26703 ) ;
  assign n26709 = n26343 &  n26615 ;
  assign n26710 = n26614 &  n26709 ;
  assign n26698 = x94 | n26343 ;
  assign n26699 = x94 &  n26343 ;
  assign n26700 = ( n26698 & ~n26699 ) | ( n26698 & 1'b0 ) | ( ~n26699 & 1'b0 ) ;
  assign n26712 = ( n26598 & n26616 ) | ( n26598 & n26700 ) | ( n26616 & n26700 ) ;
  assign n26711 = n26598 | n26700 ;
  assign n26713 = ( n26710 & ~n26712 ) | ( n26710 & n26711 ) | ( ~n26712 & n26711 ) ;
  assign n26717 = n26351 &  n26615 ;
  assign n26718 = n26614 &  n26717 ;
  assign n26706 = x93 | n26351 ;
  assign n26707 = x93 &  n26351 ;
  assign n26708 = ( n26706 & ~n26707 ) | ( n26706 & 1'b0 ) | ( ~n26707 & 1'b0 ) ;
  assign n26720 = ( n26597 & n26616 ) | ( n26597 & n26708 ) | ( n26616 & n26708 ) ;
  assign n26719 = n26597 | n26708 ;
  assign n26721 = ( n26718 & ~n26720 ) | ( n26718 & n26719 ) | ( ~n26720 & n26719 ) ;
  assign n26725 = n26359 &  n26615 ;
  assign n26726 = n26614 &  n26725 ;
  assign n26714 = x92 | n26359 ;
  assign n26715 = x92 &  n26359 ;
  assign n26716 = ( n26714 & ~n26715 ) | ( n26714 & 1'b0 ) | ( ~n26715 & 1'b0 ) ;
  assign n26728 = ( n26596 & n26616 ) | ( n26596 & n26716 ) | ( n26616 & n26716 ) ;
  assign n26727 = n26596 | n26716 ;
  assign n26729 = ( n26726 & ~n26728 ) | ( n26726 & n26727 ) | ( ~n26728 & n26727 ) ;
  assign n26733 = n26367 &  n26615 ;
  assign n26734 = n26614 &  n26733 ;
  assign n26722 = x91 | n26367 ;
  assign n26723 = x91 &  n26367 ;
  assign n26724 = ( n26722 & ~n26723 ) | ( n26722 & 1'b0 ) | ( ~n26723 & 1'b0 ) ;
  assign n26736 = ( n26595 & n26616 ) | ( n26595 & n26724 ) | ( n26616 & n26724 ) ;
  assign n26735 = n26595 | n26724 ;
  assign n26737 = ( n26734 & ~n26736 ) | ( n26734 & n26735 ) | ( ~n26736 & n26735 ) ;
  assign n26741 = n26375 &  n26615 ;
  assign n26742 = n26614 &  n26741 ;
  assign n26730 = x90 | n26375 ;
  assign n26731 = x90 &  n26375 ;
  assign n26732 = ( n26730 & ~n26731 ) | ( n26730 & 1'b0 ) | ( ~n26731 & 1'b0 ) ;
  assign n26744 = ( n26594 & n26616 ) | ( n26594 & n26732 ) | ( n26616 & n26732 ) ;
  assign n26743 = n26594 | n26732 ;
  assign n26745 = ( n26742 & ~n26744 ) | ( n26742 & n26743 ) | ( ~n26744 & n26743 ) ;
  assign n26749 = n26383 &  n26615 ;
  assign n26750 = n26614 &  n26749 ;
  assign n26738 = x89 | n26383 ;
  assign n26739 = x89 &  n26383 ;
  assign n26740 = ( n26738 & ~n26739 ) | ( n26738 & 1'b0 ) | ( ~n26739 & 1'b0 ) ;
  assign n26752 = ( n26593 & n26616 ) | ( n26593 & n26740 ) | ( n26616 & n26740 ) ;
  assign n26751 = n26593 | n26740 ;
  assign n26753 = ( n26750 & ~n26752 ) | ( n26750 & n26751 ) | ( ~n26752 & n26751 ) ;
  assign n26757 = n26391 &  n26615 ;
  assign n26758 = n26614 &  n26757 ;
  assign n26746 = x88 | n26391 ;
  assign n26747 = x88 &  n26391 ;
  assign n26748 = ( n26746 & ~n26747 ) | ( n26746 & 1'b0 ) | ( ~n26747 & 1'b0 ) ;
  assign n26760 = ( n26592 & n26616 ) | ( n26592 & n26748 ) | ( n26616 & n26748 ) ;
  assign n26759 = n26592 | n26748 ;
  assign n26761 = ( n26758 & ~n26760 ) | ( n26758 & n26759 ) | ( ~n26760 & n26759 ) ;
  assign n26765 = n26399 &  n26615 ;
  assign n26766 = n26614 &  n26765 ;
  assign n26754 = x87 | n26399 ;
  assign n26755 = x87 &  n26399 ;
  assign n26756 = ( n26754 & ~n26755 ) | ( n26754 & 1'b0 ) | ( ~n26755 & 1'b0 ) ;
  assign n26768 = ( n26591 & n26616 ) | ( n26591 & n26756 ) | ( n26616 & n26756 ) ;
  assign n26767 = n26591 | n26756 ;
  assign n26769 = ( n26766 & ~n26768 ) | ( n26766 & n26767 ) | ( ~n26768 & n26767 ) ;
  assign n26773 = n26407 &  n26615 ;
  assign n26774 = n26614 &  n26773 ;
  assign n26762 = x86 | n26407 ;
  assign n26763 = x86 &  n26407 ;
  assign n26764 = ( n26762 & ~n26763 ) | ( n26762 & 1'b0 ) | ( ~n26763 & 1'b0 ) ;
  assign n26776 = ( n26590 & n26616 ) | ( n26590 & n26764 ) | ( n26616 & n26764 ) ;
  assign n26775 = n26590 | n26764 ;
  assign n26777 = ( n26774 & ~n26776 ) | ( n26774 & n26775 ) | ( ~n26776 & n26775 ) ;
  assign n26781 = n26415 &  n26615 ;
  assign n26782 = n26614 &  n26781 ;
  assign n26770 = x85 | n26415 ;
  assign n26771 = x85 &  n26415 ;
  assign n26772 = ( n26770 & ~n26771 ) | ( n26770 & 1'b0 ) | ( ~n26771 & 1'b0 ) ;
  assign n26784 = ( n26589 & n26616 ) | ( n26589 & n26772 ) | ( n26616 & n26772 ) ;
  assign n26783 = n26589 | n26772 ;
  assign n26785 = ( n26782 & ~n26784 ) | ( n26782 & n26783 ) | ( ~n26784 & n26783 ) ;
  assign n26789 = n26423 &  n26615 ;
  assign n26790 = n26614 &  n26789 ;
  assign n26778 = x84 | n26423 ;
  assign n26779 = x84 &  n26423 ;
  assign n26780 = ( n26778 & ~n26779 ) | ( n26778 & 1'b0 ) | ( ~n26779 & 1'b0 ) ;
  assign n26792 = ( n26588 & n26616 ) | ( n26588 & n26780 ) | ( n26616 & n26780 ) ;
  assign n26791 = n26588 | n26780 ;
  assign n26793 = ( n26790 & ~n26792 ) | ( n26790 & n26791 ) | ( ~n26792 & n26791 ) ;
  assign n26797 = n26431 &  n26615 ;
  assign n26798 = n26614 &  n26797 ;
  assign n26786 = x83 | n26431 ;
  assign n26787 = x83 &  n26431 ;
  assign n26788 = ( n26786 & ~n26787 ) | ( n26786 & 1'b0 ) | ( ~n26787 & 1'b0 ) ;
  assign n26800 = ( n26587 & n26616 ) | ( n26587 & n26788 ) | ( n26616 & n26788 ) ;
  assign n26799 = n26587 | n26788 ;
  assign n26801 = ( n26798 & ~n26800 ) | ( n26798 & n26799 ) | ( ~n26800 & n26799 ) ;
  assign n26805 = n26439 &  n26615 ;
  assign n26806 = n26614 &  n26805 ;
  assign n26794 = x82 | n26439 ;
  assign n26795 = x82 &  n26439 ;
  assign n26796 = ( n26794 & ~n26795 ) | ( n26794 & 1'b0 ) | ( ~n26795 & 1'b0 ) ;
  assign n26808 = ( n26586 & n26616 ) | ( n26586 & n26796 ) | ( n26616 & n26796 ) ;
  assign n26807 = n26586 | n26796 ;
  assign n26809 = ( n26806 & ~n26808 ) | ( n26806 & n26807 ) | ( ~n26808 & n26807 ) ;
  assign n26813 = n26447 &  n26615 ;
  assign n26814 = n26614 &  n26813 ;
  assign n26802 = x81 | n26447 ;
  assign n26803 = x81 &  n26447 ;
  assign n26804 = ( n26802 & ~n26803 ) | ( n26802 & 1'b0 ) | ( ~n26803 & 1'b0 ) ;
  assign n26816 = ( n26585 & n26616 ) | ( n26585 & n26804 ) | ( n26616 & n26804 ) ;
  assign n26815 = n26585 | n26804 ;
  assign n26817 = ( n26814 & ~n26816 ) | ( n26814 & n26815 ) | ( ~n26816 & n26815 ) ;
  assign n26821 = n26455 &  n26615 ;
  assign n26822 = n26614 &  n26821 ;
  assign n26810 = x80 | n26455 ;
  assign n26811 = x80 &  n26455 ;
  assign n26812 = ( n26810 & ~n26811 ) | ( n26810 & 1'b0 ) | ( ~n26811 & 1'b0 ) ;
  assign n26824 = ( n26584 & n26616 ) | ( n26584 & n26812 ) | ( n26616 & n26812 ) ;
  assign n26823 = n26584 | n26812 ;
  assign n26825 = ( n26822 & ~n26824 ) | ( n26822 & n26823 ) | ( ~n26824 & n26823 ) ;
  assign n26829 = n26463 &  n26615 ;
  assign n26830 = n26614 &  n26829 ;
  assign n26818 = x79 | n26463 ;
  assign n26819 = x79 &  n26463 ;
  assign n26820 = ( n26818 & ~n26819 ) | ( n26818 & 1'b0 ) | ( ~n26819 & 1'b0 ) ;
  assign n26832 = ( n26583 & n26616 ) | ( n26583 & n26820 ) | ( n26616 & n26820 ) ;
  assign n26831 = n26583 | n26820 ;
  assign n26833 = ( n26830 & ~n26832 ) | ( n26830 & n26831 ) | ( ~n26832 & n26831 ) ;
  assign n26837 = n26471 &  n26615 ;
  assign n26838 = n26614 &  n26837 ;
  assign n26826 = x78 | n26471 ;
  assign n26827 = x78 &  n26471 ;
  assign n26828 = ( n26826 & ~n26827 ) | ( n26826 & 1'b0 ) | ( ~n26827 & 1'b0 ) ;
  assign n26840 = ( n26582 & n26616 ) | ( n26582 & n26828 ) | ( n26616 & n26828 ) ;
  assign n26839 = n26582 | n26828 ;
  assign n26841 = ( n26838 & ~n26840 ) | ( n26838 & n26839 ) | ( ~n26840 & n26839 ) ;
  assign n26845 = n26479 &  n26615 ;
  assign n26846 = n26614 &  n26845 ;
  assign n26834 = x77 | n26479 ;
  assign n26835 = x77 &  n26479 ;
  assign n26836 = ( n26834 & ~n26835 ) | ( n26834 & 1'b0 ) | ( ~n26835 & 1'b0 ) ;
  assign n26848 = ( n26581 & n26616 ) | ( n26581 & n26836 ) | ( n26616 & n26836 ) ;
  assign n26847 = n26581 | n26836 ;
  assign n26849 = ( n26846 & ~n26848 ) | ( n26846 & n26847 ) | ( ~n26848 & n26847 ) ;
  assign n26853 = n26487 &  n26615 ;
  assign n26854 = n26614 &  n26853 ;
  assign n26842 = x76 | n26487 ;
  assign n26843 = x76 &  n26487 ;
  assign n26844 = ( n26842 & ~n26843 ) | ( n26842 & 1'b0 ) | ( ~n26843 & 1'b0 ) ;
  assign n26856 = ( n26580 & n26616 ) | ( n26580 & n26844 ) | ( n26616 & n26844 ) ;
  assign n26855 = n26580 | n26844 ;
  assign n26857 = ( n26854 & ~n26856 ) | ( n26854 & n26855 ) | ( ~n26856 & n26855 ) ;
  assign n26861 = n26495 &  n26615 ;
  assign n26862 = n26614 &  n26861 ;
  assign n26850 = x75 | n26495 ;
  assign n26851 = x75 &  n26495 ;
  assign n26852 = ( n26850 & ~n26851 ) | ( n26850 & 1'b0 ) | ( ~n26851 & 1'b0 ) ;
  assign n26864 = ( n26579 & n26616 ) | ( n26579 & n26852 ) | ( n26616 & n26852 ) ;
  assign n26863 = n26579 | n26852 ;
  assign n26865 = ( n26862 & ~n26864 ) | ( n26862 & n26863 ) | ( ~n26864 & n26863 ) ;
  assign n26869 = n26503 &  n26615 ;
  assign n26870 = n26614 &  n26869 ;
  assign n26858 = x74 | n26503 ;
  assign n26859 = x74 &  n26503 ;
  assign n26860 = ( n26858 & ~n26859 ) | ( n26858 & 1'b0 ) | ( ~n26859 & 1'b0 ) ;
  assign n26872 = ( n26578 & n26616 ) | ( n26578 & n26860 ) | ( n26616 & n26860 ) ;
  assign n26871 = n26578 | n26860 ;
  assign n26873 = ( n26870 & ~n26872 ) | ( n26870 & n26871 ) | ( ~n26872 & n26871 ) ;
  assign n26877 = n26511 &  n26615 ;
  assign n26878 = n26614 &  n26877 ;
  assign n26866 = x73 | n26511 ;
  assign n26867 = x73 &  n26511 ;
  assign n26868 = ( n26866 & ~n26867 ) | ( n26866 & 1'b0 ) | ( ~n26867 & 1'b0 ) ;
  assign n26880 = ( n26577 & n26616 ) | ( n26577 & n26868 ) | ( n26616 & n26868 ) ;
  assign n26879 = n26577 | n26868 ;
  assign n26881 = ( n26878 & ~n26880 ) | ( n26878 & n26879 ) | ( ~n26880 & n26879 ) ;
  assign n26885 = n26519 &  n26615 ;
  assign n26886 = n26614 &  n26885 ;
  assign n26874 = x72 | n26519 ;
  assign n26875 = x72 &  n26519 ;
  assign n26876 = ( n26874 & ~n26875 ) | ( n26874 & 1'b0 ) | ( ~n26875 & 1'b0 ) ;
  assign n26888 = ( n26576 & n26616 ) | ( n26576 & n26876 ) | ( n26616 & n26876 ) ;
  assign n26887 = n26576 | n26876 ;
  assign n26889 = ( n26886 & ~n26888 ) | ( n26886 & n26887 ) | ( ~n26888 & n26887 ) ;
  assign n26893 = n26527 &  n26615 ;
  assign n26894 = n26614 &  n26893 ;
  assign n26882 = x71 | n26527 ;
  assign n26883 = x71 &  n26527 ;
  assign n26884 = ( n26882 & ~n26883 ) | ( n26882 & 1'b0 ) | ( ~n26883 & 1'b0 ) ;
  assign n26896 = ( n26575 & n26616 ) | ( n26575 & n26884 ) | ( n26616 & n26884 ) ;
  assign n26895 = n26575 | n26884 ;
  assign n26897 = ( n26894 & ~n26896 ) | ( n26894 & n26895 ) | ( ~n26896 & n26895 ) ;
  assign n26901 = n26535 &  n26615 ;
  assign n26902 = n26614 &  n26901 ;
  assign n26890 = x70 | n26535 ;
  assign n26891 = x70 &  n26535 ;
  assign n26892 = ( n26890 & ~n26891 ) | ( n26890 & 1'b0 ) | ( ~n26891 & 1'b0 ) ;
  assign n26904 = ( n26574 & n26616 ) | ( n26574 & n26892 ) | ( n26616 & n26892 ) ;
  assign n26903 = n26574 | n26892 ;
  assign n26905 = ( n26902 & ~n26904 ) | ( n26902 & n26903 ) | ( ~n26904 & n26903 ) ;
  assign n26909 = n26543 &  n26615 ;
  assign n26910 = n26614 &  n26909 ;
  assign n26898 = x69 | n26543 ;
  assign n26899 = x69 &  n26543 ;
  assign n26900 = ( n26898 & ~n26899 ) | ( n26898 & 1'b0 ) | ( ~n26899 & 1'b0 ) ;
  assign n26912 = ( n26573 & n26616 ) | ( n26573 & n26900 ) | ( n26616 & n26900 ) ;
  assign n26911 = n26573 | n26900 ;
  assign n26913 = ( n26910 & ~n26912 ) | ( n26910 & n26911 ) | ( ~n26912 & n26911 ) ;
  assign n26917 = n26551 &  n26615 ;
  assign n26918 = n26614 &  n26917 ;
  assign n26906 = x68 | n26551 ;
  assign n26907 = x68 &  n26551 ;
  assign n26908 = ( n26906 & ~n26907 ) | ( n26906 & 1'b0 ) | ( ~n26907 & 1'b0 ) ;
  assign n26920 = ( n26572 & n26616 ) | ( n26572 & n26908 ) | ( n26616 & n26908 ) ;
  assign n26919 = n26572 | n26908 ;
  assign n26921 = ( n26918 & ~n26920 ) | ( n26918 & n26919 ) | ( ~n26920 & n26919 ) ;
  assign n26925 = n26559 &  n26615 ;
  assign n26926 = n26614 &  n26925 ;
  assign n26914 = x67 | n26559 ;
  assign n26915 = x67 &  n26559 ;
  assign n26916 = ( n26914 & ~n26915 ) | ( n26914 & 1'b0 ) | ( ~n26915 & 1'b0 ) ;
  assign n26928 = ( n26571 & n26616 ) | ( n26571 & n26916 ) | ( n26616 & n26916 ) ;
  assign n26927 = n26571 | n26916 ;
  assign n26929 = ( n26926 & ~n26928 ) | ( n26926 & n26927 ) | ( ~n26928 & n26927 ) ;
  assign n26930 = n26565 &  n26615 ;
  assign n26931 = n26614 &  n26930 ;
  assign n26922 = x66 | n26565 ;
  assign n26923 = x66 &  n26565 ;
  assign n26924 = ( n26922 & ~n26923 ) | ( n26922 & 1'b0 ) | ( ~n26923 & 1'b0 ) ;
  assign n26933 = ( n26570 & n26616 ) | ( n26570 & n26924 ) | ( n26616 & n26924 ) ;
  assign n26932 = n26570 | n26924 ;
  assign n26934 = ( n26931 & ~n26933 ) | ( n26931 & n26932 ) | ( ~n26933 & n26932 ) ;
  assign n26935 = ( x65 & ~n8105 ) | ( x65 & n26569 ) | ( ~n8105 & n26569 ) ;
  assign n26936 = ( n26570 & ~x65 ) | ( n26570 & n26935 ) | ( ~x65 & n26935 ) ;
  assign n26937 = ~n26616 & n26936 ;
  assign n26938 = n26569 &  n26615 ;
  assign n26939 = n26614 &  n26938 ;
  assign n26940 = n26937 | n26939 ;
  assign n26941 = ( x64 & ~n26616 ) | ( x64 & 1'b0 ) | ( ~n26616 & 1'b0 ) ;
  assign n26942 = ( x22 & ~n26941 ) | ( x22 & 1'b0 ) | ( ~n26941 & 1'b0 ) ;
  assign n26943 = ( n8105 & ~n26616 ) | ( n8105 & 1'b0 ) | ( ~n26616 & 1'b0 ) ;
  assign n26944 = n26942 | n26943 ;
  assign n26945 = ( x65 & ~n26944 ) | ( x65 & n8606 ) | ( ~n26944 & n8606 ) ;
  assign n26946 = ( x66 & ~n26940 ) | ( x66 & n26945 ) | ( ~n26940 & n26945 ) ;
  assign n26947 = ( x67 & ~n26934 ) | ( x67 & n26946 ) | ( ~n26934 & n26946 ) ;
  assign n26948 = ( x68 & ~n26929 ) | ( x68 & n26947 ) | ( ~n26929 & n26947 ) ;
  assign n26949 = ( x69 & ~n26921 ) | ( x69 & n26948 ) | ( ~n26921 & n26948 ) ;
  assign n26950 = ( x70 & ~n26913 ) | ( x70 & n26949 ) | ( ~n26913 & n26949 ) ;
  assign n26951 = ( x71 & ~n26905 ) | ( x71 & n26950 ) | ( ~n26905 & n26950 ) ;
  assign n26952 = ( x72 & ~n26897 ) | ( x72 & n26951 ) | ( ~n26897 & n26951 ) ;
  assign n26953 = ( x73 & ~n26889 ) | ( x73 & n26952 ) | ( ~n26889 & n26952 ) ;
  assign n26954 = ( x74 & ~n26881 ) | ( x74 & n26953 ) | ( ~n26881 & n26953 ) ;
  assign n26955 = ( x75 & ~n26873 ) | ( x75 & n26954 ) | ( ~n26873 & n26954 ) ;
  assign n26956 = ( x76 & ~n26865 ) | ( x76 & n26955 ) | ( ~n26865 & n26955 ) ;
  assign n26957 = ( x77 & ~n26857 ) | ( x77 & n26956 ) | ( ~n26857 & n26956 ) ;
  assign n26958 = ( x78 & ~n26849 ) | ( x78 & n26957 ) | ( ~n26849 & n26957 ) ;
  assign n26959 = ( x79 & ~n26841 ) | ( x79 & n26958 ) | ( ~n26841 & n26958 ) ;
  assign n26960 = ( x80 & ~n26833 ) | ( x80 & n26959 ) | ( ~n26833 & n26959 ) ;
  assign n26961 = ( x81 & ~n26825 ) | ( x81 & n26960 ) | ( ~n26825 & n26960 ) ;
  assign n26962 = ( x82 & ~n26817 ) | ( x82 & n26961 ) | ( ~n26817 & n26961 ) ;
  assign n26963 = ( x83 & ~n26809 ) | ( x83 & n26962 ) | ( ~n26809 & n26962 ) ;
  assign n26964 = ( x84 & ~n26801 ) | ( x84 & n26963 ) | ( ~n26801 & n26963 ) ;
  assign n26965 = ( x85 & ~n26793 ) | ( x85 & n26964 ) | ( ~n26793 & n26964 ) ;
  assign n26966 = ( x86 & ~n26785 ) | ( x86 & n26965 ) | ( ~n26785 & n26965 ) ;
  assign n26967 = ( x87 & ~n26777 ) | ( x87 & n26966 ) | ( ~n26777 & n26966 ) ;
  assign n26968 = ( x88 & ~n26769 ) | ( x88 & n26967 ) | ( ~n26769 & n26967 ) ;
  assign n26969 = ( x89 & ~n26761 ) | ( x89 & n26968 ) | ( ~n26761 & n26968 ) ;
  assign n26970 = ( x90 & ~n26753 ) | ( x90 & n26969 ) | ( ~n26753 & n26969 ) ;
  assign n26971 = ( x91 & ~n26745 ) | ( x91 & n26970 ) | ( ~n26745 & n26970 ) ;
  assign n26972 = ( x92 & ~n26737 ) | ( x92 & n26971 ) | ( ~n26737 & n26971 ) ;
  assign n26973 = ( x93 & ~n26729 ) | ( x93 & n26972 ) | ( ~n26729 & n26972 ) ;
  assign n26974 = ( x94 & ~n26721 ) | ( x94 & n26973 ) | ( ~n26721 & n26973 ) ;
  assign n26975 = ( x95 & ~n26713 ) | ( x95 & n26974 ) | ( ~n26713 & n26974 ) ;
  assign n26976 = ( x96 & ~n26705 ) | ( x96 & n26975 ) | ( ~n26705 & n26975 ) ;
  assign n26977 = ( x97 & ~n26697 ) | ( x97 & n26976 ) | ( ~n26697 & n26976 ) ;
  assign n26978 = ( x98 & ~n26689 ) | ( x98 & n26977 ) | ( ~n26689 & n26977 ) ;
  assign n26979 = ( x99 & ~n26681 ) | ( x99 & n26978 ) | ( ~n26681 & n26978 ) ;
  assign n26980 = ( x100 & ~n26673 ) | ( x100 & n26979 ) | ( ~n26673 & n26979 ) ;
  assign n26981 = ( x101 & ~n26665 ) | ( x101 & n26980 ) | ( ~n26665 & n26980 ) ;
  assign n26982 = ( x102 & ~n26657 ) | ( x102 & n26981 ) | ( ~n26657 & n26981 ) ;
  assign n26983 = ( x103 & ~n26649 ) | ( x103 & n26982 ) | ( ~n26649 & n26982 ) ;
  assign n26984 = ( x104 & ~n26641 ) | ( x104 & n26983 ) | ( ~n26641 & n26983 ) ;
  assign n26985 = ( x105 & ~n26633 ) | ( x105 & n26984 ) | ( ~n26633 & n26984 ) ;
  assign n26986 = ( x106 & ~n26625 ) | ( x106 & n26985 ) | ( ~n26625 & n26985 ) ;
  assign n26987 = n8650 | n26986 ;
  assign n26997 = n26633 &  n26987 ;
  assign n26989 = x105 | n26633 ;
  assign n26990 = x105 &  n26633 ;
  assign n26991 = ( n26989 & ~n26990 ) | ( n26989 & 1'b0 ) | ( ~n26990 & 1'b0 ) ;
  assign n27001 = ( n8650 & n26984 ) | ( n8650 & n26991 ) | ( n26984 & n26991 ) ;
  assign n27002 = ( n26984 & ~n26986 ) | ( n26984 & n26991 ) | ( ~n26986 & n26991 ) ;
  assign n27003 = ~n27001 & n27002 ;
  assign n27004 = n26997 | n27003 ;
  assign n27005 = n26641 &  n26987 ;
  assign n26998 = x104 | n26641 ;
  assign n26999 = x104 &  n26641 ;
  assign n27000 = ( n26998 & ~n26999 ) | ( n26998 & 1'b0 ) | ( ~n26999 & 1'b0 ) ;
  assign n27009 = ( n8650 & n26983 ) | ( n8650 & n27000 ) | ( n26983 & n27000 ) ;
  assign n27010 = ( n26983 & ~n26986 ) | ( n26983 & n27000 ) | ( ~n26986 & n27000 ) ;
  assign n27011 = ~n27009 & n27010 ;
  assign n27012 = n27005 | n27011 ;
  assign n27013 = n26649 &  n26987 ;
  assign n27006 = x103 | n26649 ;
  assign n27007 = x103 &  n26649 ;
  assign n27008 = ( n27006 & ~n27007 ) | ( n27006 & 1'b0 ) | ( ~n27007 & 1'b0 ) ;
  assign n27017 = ( n8650 & n26982 ) | ( n8650 & n27008 ) | ( n26982 & n27008 ) ;
  assign n27018 = ( n26982 & ~n26986 ) | ( n26982 & n27008 ) | ( ~n26986 & n27008 ) ;
  assign n27019 = ~n27017 & n27018 ;
  assign n27020 = n27013 | n27019 ;
  assign n27021 = n26657 &  n26987 ;
  assign n27014 = x102 | n26657 ;
  assign n27015 = x102 &  n26657 ;
  assign n27016 = ( n27014 & ~n27015 ) | ( n27014 & 1'b0 ) | ( ~n27015 & 1'b0 ) ;
  assign n27025 = ( n8650 & n26981 ) | ( n8650 & n27016 ) | ( n26981 & n27016 ) ;
  assign n27026 = ( n26981 & ~n26986 ) | ( n26981 & n27016 ) | ( ~n26986 & n27016 ) ;
  assign n27027 = ~n27025 & n27026 ;
  assign n27028 = n27021 | n27027 ;
  assign n27029 = n26665 &  n26987 ;
  assign n27022 = x101 | n26665 ;
  assign n27023 = x101 &  n26665 ;
  assign n27024 = ( n27022 & ~n27023 ) | ( n27022 & 1'b0 ) | ( ~n27023 & 1'b0 ) ;
  assign n27033 = ( n8650 & n26980 ) | ( n8650 & n27024 ) | ( n26980 & n27024 ) ;
  assign n27034 = ( n26980 & ~n26986 ) | ( n26980 & n27024 ) | ( ~n26986 & n27024 ) ;
  assign n27035 = ~n27033 & n27034 ;
  assign n27036 = n27029 | n27035 ;
  assign n27037 = n26673 &  n26987 ;
  assign n27030 = x100 | n26673 ;
  assign n27031 = x100 &  n26673 ;
  assign n27032 = ( n27030 & ~n27031 ) | ( n27030 & 1'b0 ) | ( ~n27031 & 1'b0 ) ;
  assign n27041 = ( n8650 & n26979 ) | ( n8650 & n27032 ) | ( n26979 & n27032 ) ;
  assign n27042 = ( n26979 & ~n26986 ) | ( n26979 & n27032 ) | ( ~n26986 & n27032 ) ;
  assign n27043 = ~n27041 & n27042 ;
  assign n27044 = n27037 | n27043 ;
  assign n27045 = n26681 &  n26987 ;
  assign n27038 = x99 | n26681 ;
  assign n27039 = x99 &  n26681 ;
  assign n27040 = ( n27038 & ~n27039 ) | ( n27038 & 1'b0 ) | ( ~n27039 & 1'b0 ) ;
  assign n27049 = ( n8650 & n26978 ) | ( n8650 & n27040 ) | ( n26978 & n27040 ) ;
  assign n27050 = ( n26978 & ~n26986 ) | ( n26978 & n27040 ) | ( ~n26986 & n27040 ) ;
  assign n27051 = ~n27049 & n27050 ;
  assign n27052 = n27045 | n27051 ;
  assign n27053 = n26689 &  n26987 ;
  assign n27046 = x98 | n26689 ;
  assign n27047 = x98 &  n26689 ;
  assign n27048 = ( n27046 & ~n27047 ) | ( n27046 & 1'b0 ) | ( ~n27047 & 1'b0 ) ;
  assign n27057 = ( n8650 & n26977 ) | ( n8650 & n27048 ) | ( n26977 & n27048 ) ;
  assign n27058 = ( n26977 & ~n26986 ) | ( n26977 & n27048 ) | ( ~n26986 & n27048 ) ;
  assign n27059 = ~n27057 & n27058 ;
  assign n27060 = n27053 | n27059 ;
  assign n27061 = n26697 &  n26987 ;
  assign n27054 = x97 | n26697 ;
  assign n27055 = x97 &  n26697 ;
  assign n27056 = ( n27054 & ~n27055 ) | ( n27054 & 1'b0 ) | ( ~n27055 & 1'b0 ) ;
  assign n27065 = ( n8650 & n26976 ) | ( n8650 & n27056 ) | ( n26976 & n27056 ) ;
  assign n27066 = ( n26976 & ~n26986 ) | ( n26976 & n27056 ) | ( ~n26986 & n27056 ) ;
  assign n27067 = ~n27065 & n27066 ;
  assign n27068 = n27061 | n27067 ;
  assign n27069 = n26705 &  n26987 ;
  assign n27062 = x96 | n26705 ;
  assign n27063 = x96 &  n26705 ;
  assign n27064 = ( n27062 & ~n27063 ) | ( n27062 & 1'b0 ) | ( ~n27063 & 1'b0 ) ;
  assign n27073 = ( n8650 & n26975 ) | ( n8650 & n27064 ) | ( n26975 & n27064 ) ;
  assign n27074 = ( n26975 & ~n26986 ) | ( n26975 & n27064 ) | ( ~n26986 & n27064 ) ;
  assign n27075 = ~n27073 & n27074 ;
  assign n27076 = n27069 | n27075 ;
  assign n27077 = n26713 &  n26987 ;
  assign n27070 = x95 | n26713 ;
  assign n27071 = x95 &  n26713 ;
  assign n27072 = ( n27070 & ~n27071 ) | ( n27070 & 1'b0 ) | ( ~n27071 & 1'b0 ) ;
  assign n27081 = ( n8650 & n26974 ) | ( n8650 & n27072 ) | ( n26974 & n27072 ) ;
  assign n27082 = ( n26974 & ~n26986 ) | ( n26974 & n27072 ) | ( ~n26986 & n27072 ) ;
  assign n27083 = ~n27081 & n27082 ;
  assign n27084 = n27077 | n27083 ;
  assign n27085 = n26721 &  n26987 ;
  assign n27078 = x94 | n26721 ;
  assign n27079 = x94 &  n26721 ;
  assign n27080 = ( n27078 & ~n27079 ) | ( n27078 & 1'b0 ) | ( ~n27079 & 1'b0 ) ;
  assign n27089 = ( n8650 & n26973 ) | ( n8650 & n27080 ) | ( n26973 & n27080 ) ;
  assign n27090 = ( n26973 & ~n26986 ) | ( n26973 & n27080 ) | ( ~n26986 & n27080 ) ;
  assign n27091 = ~n27089 & n27090 ;
  assign n27092 = n27085 | n27091 ;
  assign n27093 = n26729 &  n26987 ;
  assign n27086 = x93 | n26729 ;
  assign n27087 = x93 &  n26729 ;
  assign n27088 = ( n27086 & ~n27087 ) | ( n27086 & 1'b0 ) | ( ~n27087 & 1'b0 ) ;
  assign n27097 = ( n8650 & n26972 ) | ( n8650 & n27088 ) | ( n26972 & n27088 ) ;
  assign n27098 = ( n26972 & ~n26986 ) | ( n26972 & n27088 ) | ( ~n26986 & n27088 ) ;
  assign n27099 = ~n27097 & n27098 ;
  assign n27100 = n27093 | n27099 ;
  assign n27101 = n26737 &  n26987 ;
  assign n27094 = x92 | n26737 ;
  assign n27095 = x92 &  n26737 ;
  assign n27096 = ( n27094 & ~n27095 ) | ( n27094 & 1'b0 ) | ( ~n27095 & 1'b0 ) ;
  assign n27105 = ( n8650 & n26971 ) | ( n8650 & n27096 ) | ( n26971 & n27096 ) ;
  assign n27106 = ( n26971 & ~n26986 ) | ( n26971 & n27096 ) | ( ~n26986 & n27096 ) ;
  assign n27107 = ~n27105 & n27106 ;
  assign n27108 = n27101 | n27107 ;
  assign n27109 = n26745 &  n26987 ;
  assign n27102 = x91 | n26745 ;
  assign n27103 = x91 &  n26745 ;
  assign n27104 = ( n27102 & ~n27103 ) | ( n27102 & 1'b0 ) | ( ~n27103 & 1'b0 ) ;
  assign n27113 = ( n8650 & n26970 ) | ( n8650 & n27104 ) | ( n26970 & n27104 ) ;
  assign n27114 = ( n26970 & ~n26986 ) | ( n26970 & n27104 ) | ( ~n26986 & n27104 ) ;
  assign n27115 = ~n27113 & n27114 ;
  assign n27116 = n27109 | n27115 ;
  assign n27117 = n26753 &  n26987 ;
  assign n27110 = x90 | n26753 ;
  assign n27111 = x90 &  n26753 ;
  assign n27112 = ( n27110 & ~n27111 ) | ( n27110 & 1'b0 ) | ( ~n27111 & 1'b0 ) ;
  assign n27121 = ( n8650 & n26969 ) | ( n8650 & n27112 ) | ( n26969 & n27112 ) ;
  assign n27122 = ( n26969 & ~n26986 ) | ( n26969 & n27112 ) | ( ~n26986 & n27112 ) ;
  assign n27123 = ~n27121 & n27122 ;
  assign n27124 = n27117 | n27123 ;
  assign n27125 = n26761 &  n26987 ;
  assign n27118 = x89 | n26761 ;
  assign n27119 = x89 &  n26761 ;
  assign n27120 = ( n27118 & ~n27119 ) | ( n27118 & 1'b0 ) | ( ~n27119 & 1'b0 ) ;
  assign n27129 = ( n8650 & n26968 ) | ( n8650 & n27120 ) | ( n26968 & n27120 ) ;
  assign n27130 = ( n26968 & ~n26986 ) | ( n26968 & n27120 ) | ( ~n26986 & n27120 ) ;
  assign n27131 = ~n27129 & n27130 ;
  assign n27132 = n27125 | n27131 ;
  assign n27133 = n26769 &  n26987 ;
  assign n27126 = x88 | n26769 ;
  assign n27127 = x88 &  n26769 ;
  assign n27128 = ( n27126 & ~n27127 ) | ( n27126 & 1'b0 ) | ( ~n27127 & 1'b0 ) ;
  assign n27137 = ( n8650 & n26967 ) | ( n8650 & n27128 ) | ( n26967 & n27128 ) ;
  assign n27138 = ( n26967 & ~n26986 ) | ( n26967 & n27128 ) | ( ~n26986 & n27128 ) ;
  assign n27139 = ~n27137 & n27138 ;
  assign n27140 = n27133 | n27139 ;
  assign n27141 = n26777 &  n26987 ;
  assign n27134 = x87 | n26777 ;
  assign n27135 = x87 &  n26777 ;
  assign n27136 = ( n27134 & ~n27135 ) | ( n27134 & 1'b0 ) | ( ~n27135 & 1'b0 ) ;
  assign n27145 = ( n8650 & n26966 ) | ( n8650 & n27136 ) | ( n26966 & n27136 ) ;
  assign n27146 = ( n26966 & ~n26986 ) | ( n26966 & n27136 ) | ( ~n26986 & n27136 ) ;
  assign n27147 = ~n27145 & n27146 ;
  assign n27148 = n27141 | n27147 ;
  assign n27149 = n26785 &  n26987 ;
  assign n27142 = x86 | n26785 ;
  assign n27143 = x86 &  n26785 ;
  assign n27144 = ( n27142 & ~n27143 ) | ( n27142 & 1'b0 ) | ( ~n27143 & 1'b0 ) ;
  assign n27153 = ( n8650 & n26965 ) | ( n8650 & n27144 ) | ( n26965 & n27144 ) ;
  assign n27154 = ( n26965 & ~n26986 ) | ( n26965 & n27144 ) | ( ~n26986 & n27144 ) ;
  assign n27155 = ~n27153 & n27154 ;
  assign n27156 = n27149 | n27155 ;
  assign n27157 = n26793 &  n26987 ;
  assign n27150 = x85 | n26793 ;
  assign n27151 = x85 &  n26793 ;
  assign n27152 = ( n27150 & ~n27151 ) | ( n27150 & 1'b0 ) | ( ~n27151 & 1'b0 ) ;
  assign n27161 = ( n8650 & n26964 ) | ( n8650 & n27152 ) | ( n26964 & n27152 ) ;
  assign n27162 = ( n26964 & ~n26986 ) | ( n26964 & n27152 ) | ( ~n26986 & n27152 ) ;
  assign n27163 = ~n27161 & n27162 ;
  assign n27164 = n27157 | n27163 ;
  assign n27165 = n26801 &  n26987 ;
  assign n27158 = x84 | n26801 ;
  assign n27159 = x84 &  n26801 ;
  assign n27160 = ( n27158 & ~n27159 ) | ( n27158 & 1'b0 ) | ( ~n27159 & 1'b0 ) ;
  assign n27169 = ( n8650 & n26963 ) | ( n8650 & n27160 ) | ( n26963 & n27160 ) ;
  assign n27170 = ( n26963 & ~n26986 ) | ( n26963 & n27160 ) | ( ~n26986 & n27160 ) ;
  assign n27171 = ~n27169 & n27170 ;
  assign n27172 = n27165 | n27171 ;
  assign n27173 = n26809 &  n26987 ;
  assign n27166 = x83 | n26809 ;
  assign n27167 = x83 &  n26809 ;
  assign n27168 = ( n27166 & ~n27167 ) | ( n27166 & 1'b0 ) | ( ~n27167 & 1'b0 ) ;
  assign n27177 = ( n8650 & n26962 ) | ( n8650 & n27168 ) | ( n26962 & n27168 ) ;
  assign n27178 = ( n26962 & ~n26986 ) | ( n26962 & n27168 ) | ( ~n26986 & n27168 ) ;
  assign n27179 = ~n27177 & n27178 ;
  assign n27180 = n27173 | n27179 ;
  assign n27181 = n26817 &  n26987 ;
  assign n27174 = x82 | n26817 ;
  assign n27175 = x82 &  n26817 ;
  assign n27176 = ( n27174 & ~n27175 ) | ( n27174 & 1'b0 ) | ( ~n27175 & 1'b0 ) ;
  assign n27185 = ( n8650 & n26961 ) | ( n8650 & n27176 ) | ( n26961 & n27176 ) ;
  assign n27186 = ( n26961 & ~n26986 ) | ( n26961 & n27176 ) | ( ~n26986 & n27176 ) ;
  assign n27187 = ~n27185 & n27186 ;
  assign n27188 = n27181 | n27187 ;
  assign n27189 = n26825 &  n26987 ;
  assign n27182 = x81 | n26825 ;
  assign n27183 = x81 &  n26825 ;
  assign n27184 = ( n27182 & ~n27183 ) | ( n27182 & 1'b0 ) | ( ~n27183 & 1'b0 ) ;
  assign n27193 = ( n8650 & n26960 ) | ( n8650 & n27184 ) | ( n26960 & n27184 ) ;
  assign n27194 = ( n26960 & ~n26986 ) | ( n26960 & n27184 ) | ( ~n26986 & n27184 ) ;
  assign n27195 = ~n27193 & n27194 ;
  assign n27196 = n27189 | n27195 ;
  assign n27197 = n26833 &  n26987 ;
  assign n27190 = x80 | n26833 ;
  assign n27191 = x80 &  n26833 ;
  assign n27192 = ( n27190 & ~n27191 ) | ( n27190 & 1'b0 ) | ( ~n27191 & 1'b0 ) ;
  assign n27201 = ( n8650 & n26959 ) | ( n8650 & n27192 ) | ( n26959 & n27192 ) ;
  assign n27202 = ( n26959 & ~n26986 ) | ( n26959 & n27192 ) | ( ~n26986 & n27192 ) ;
  assign n27203 = ~n27201 & n27202 ;
  assign n27204 = n27197 | n27203 ;
  assign n27205 = n26841 &  n26987 ;
  assign n27198 = x79 | n26841 ;
  assign n27199 = x79 &  n26841 ;
  assign n27200 = ( n27198 & ~n27199 ) | ( n27198 & 1'b0 ) | ( ~n27199 & 1'b0 ) ;
  assign n27209 = ( n8650 & n26958 ) | ( n8650 & n27200 ) | ( n26958 & n27200 ) ;
  assign n27210 = ( n26958 & ~n26986 ) | ( n26958 & n27200 ) | ( ~n26986 & n27200 ) ;
  assign n27211 = ~n27209 & n27210 ;
  assign n27212 = n27205 | n27211 ;
  assign n27213 = n26849 &  n26987 ;
  assign n27206 = x78 | n26849 ;
  assign n27207 = x78 &  n26849 ;
  assign n27208 = ( n27206 & ~n27207 ) | ( n27206 & 1'b0 ) | ( ~n27207 & 1'b0 ) ;
  assign n27217 = ( n8650 & n26957 ) | ( n8650 & n27208 ) | ( n26957 & n27208 ) ;
  assign n27218 = ( n26957 & ~n26986 ) | ( n26957 & n27208 ) | ( ~n26986 & n27208 ) ;
  assign n27219 = ~n27217 & n27218 ;
  assign n27220 = n27213 | n27219 ;
  assign n27221 = n26857 &  n26987 ;
  assign n27214 = x77 | n26857 ;
  assign n27215 = x77 &  n26857 ;
  assign n27216 = ( n27214 & ~n27215 ) | ( n27214 & 1'b0 ) | ( ~n27215 & 1'b0 ) ;
  assign n27225 = ( n8650 & n26956 ) | ( n8650 & n27216 ) | ( n26956 & n27216 ) ;
  assign n27226 = ( n26956 & ~n26986 ) | ( n26956 & n27216 ) | ( ~n26986 & n27216 ) ;
  assign n27227 = ~n27225 & n27226 ;
  assign n27228 = n27221 | n27227 ;
  assign n27229 = n26865 &  n26987 ;
  assign n27222 = x76 | n26865 ;
  assign n27223 = x76 &  n26865 ;
  assign n27224 = ( n27222 & ~n27223 ) | ( n27222 & 1'b0 ) | ( ~n27223 & 1'b0 ) ;
  assign n27233 = ( n8650 & n26955 ) | ( n8650 & n27224 ) | ( n26955 & n27224 ) ;
  assign n27234 = ( n26955 & ~n26986 ) | ( n26955 & n27224 ) | ( ~n26986 & n27224 ) ;
  assign n27235 = ~n27233 & n27234 ;
  assign n27236 = n27229 | n27235 ;
  assign n27237 = n26873 &  n26987 ;
  assign n27230 = x75 | n26873 ;
  assign n27231 = x75 &  n26873 ;
  assign n27232 = ( n27230 & ~n27231 ) | ( n27230 & 1'b0 ) | ( ~n27231 & 1'b0 ) ;
  assign n27241 = ( n8650 & n26954 ) | ( n8650 & n27232 ) | ( n26954 & n27232 ) ;
  assign n27242 = ( n26954 & ~n26986 ) | ( n26954 & n27232 ) | ( ~n26986 & n27232 ) ;
  assign n27243 = ~n27241 & n27242 ;
  assign n27244 = n27237 | n27243 ;
  assign n27245 = n26881 &  n26987 ;
  assign n27238 = x74 | n26881 ;
  assign n27239 = x74 &  n26881 ;
  assign n27240 = ( n27238 & ~n27239 ) | ( n27238 & 1'b0 ) | ( ~n27239 & 1'b0 ) ;
  assign n27249 = ( n8650 & n26953 ) | ( n8650 & n27240 ) | ( n26953 & n27240 ) ;
  assign n27250 = ( n26953 & ~n26986 ) | ( n26953 & n27240 ) | ( ~n26986 & n27240 ) ;
  assign n27251 = ~n27249 & n27250 ;
  assign n27252 = n27245 | n27251 ;
  assign n27253 = n26889 &  n26987 ;
  assign n27246 = x73 | n26889 ;
  assign n27247 = x73 &  n26889 ;
  assign n27248 = ( n27246 & ~n27247 ) | ( n27246 & 1'b0 ) | ( ~n27247 & 1'b0 ) ;
  assign n27257 = ( n8650 & n26952 ) | ( n8650 & n27248 ) | ( n26952 & n27248 ) ;
  assign n27258 = ( n26952 & ~n26986 ) | ( n26952 & n27248 ) | ( ~n26986 & n27248 ) ;
  assign n27259 = ~n27257 & n27258 ;
  assign n27260 = n27253 | n27259 ;
  assign n27261 = n26897 &  n26987 ;
  assign n27254 = x72 | n26897 ;
  assign n27255 = x72 &  n26897 ;
  assign n27256 = ( n27254 & ~n27255 ) | ( n27254 & 1'b0 ) | ( ~n27255 & 1'b0 ) ;
  assign n27265 = ( n8650 & n26951 ) | ( n8650 & n27256 ) | ( n26951 & n27256 ) ;
  assign n27266 = ( n26951 & ~n26986 ) | ( n26951 & n27256 ) | ( ~n26986 & n27256 ) ;
  assign n27267 = ~n27265 & n27266 ;
  assign n27268 = n27261 | n27267 ;
  assign n27269 = n26905 &  n26987 ;
  assign n27262 = x71 | n26905 ;
  assign n27263 = x71 &  n26905 ;
  assign n27264 = ( n27262 & ~n27263 ) | ( n27262 & 1'b0 ) | ( ~n27263 & 1'b0 ) ;
  assign n27273 = ( n8650 & n26950 ) | ( n8650 & n27264 ) | ( n26950 & n27264 ) ;
  assign n27274 = ( n26950 & ~n26986 ) | ( n26950 & n27264 ) | ( ~n26986 & n27264 ) ;
  assign n27275 = ~n27273 & n27274 ;
  assign n27276 = n27269 | n27275 ;
  assign n27277 = n26913 &  n26987 ;
  assign n27270 = x70 | n26913 ;
  assign n27271 = x70 &  n26913 ;
  assign n27272 = ( n27270 & ~n27271 ) | ( n27270 & 1'b0 ) | ( ~n27271 & 1'b0 ) ;
  assign n27281 = ( n8650 & n26949 ) | ( n8650 & n27272 ) | ( n26949 & n27272 ) ;
  assign n27282 = ( n26949 & ~n26986 ) | ( n26949 & n27272 ) | ( ~n26986 & n27272 ) ;
  assign n27283 = ~n27281 & n27282 ;
  assign n27284 = n27277 | n27283 ;
  assign n27285 = n26921 &  n26987 ;
  assign n27278 = x69 | n26921 ;
  assign n27279 = x69 &  n26921 ;
  assign n27280 = ( n27278 & ~n27279 ) | ( n27278 & 1'b0 ) | ( ~n27279 & 1'b0 ) ;
  assign n27289 = ( n8650 & n26948 ) | ( n8650 & n27280 ) | ( n26948 & n27280 ) ;
  assign n27290 = ( n26948 & ~n26986 ) | ( n26948 & n27280 ) | ( ~n26986 & n27280 ) ;
  assign n27291 = ~n27289 & n27290 ;
  assign n27292 = n27285 | n27291 ;
  assign n27293 = n26929 &  n26987 ;
  assign n27286 = x68 | n26929 ;
  assign n27287 = x68 &  n26929 ;
  assign n27288 = ( n27286 & ~n27287 ) | ( n27286 & 1'b0 ) | ( ~n27287 & 1'b0 ) ;
  assign n27297 = ( n8650 & n26947 ) | ( n8650 & n27288 ) | ( n26947 & n27288 ) ;
  assign n27298 = ( n26947 & ~n26986 ) | ( n26947 & n27288 ) | ( ~n26986 & n27288 ) ;
  assign n27299 = ~n27297 & n27298 ;
  assign n27300 = n27293 | n27299 ;
  assign n27301 = n26934 &  n26987 ;
  assign n27294 = x67 | n26934 ;
  assign n27295 = x67 &  n26934 ;
  assign n27296 = ( n27294 & ~n27295 ) | ( n27294 & 1'b0 ) | ( ~n27295 & 1'b0 ) ;
  assign n27305 = ( n8650 & n26946 ) | ( n8650 & n27296 ) | ( n26946 & n27296 ) ;
  assign n27306 = ( n26946 & ~n26986 ) | ( n26946 & n27296 ) | ( ~n26986 & n27296 ) ;
  assign n27307 = ~n27305 & n27306 ;
  assign n27308 = n27301 | n27307 ;
  assign n27309 = n26940 &  n26987 ;
  assign n27302 = x66 | n26940 ;
  assign n27303 = x66 &  n26940 ;
  assign n27304 = ( n27302 & ~n27303 ) | ( n27302 & 1'b0 ) | ( ~n27303 & 1'b0 ) ;
  assign n27310 = ( n8650 & n26945 ) | ( n8650 & n27304 ) | ( n26945 & n27304 ) ;
  assign n27311 = ( n26945 & ~n26986 ) | ( n26945 & n27304 ) | ( ~n26986 & n27304 ) ;
  assign n27312 = ~n27310 & n27311 ;
  assign n27313 = n27309 | n27312 ;
  assign n27314 = n26944 &  n26987 ;
  assign n27315 = ( x65 & ~x22 ) | ( x65 & n26941 ) | ( ~x22 & n26941 ) ;
  assign n27316 = ( x22 & ~n26941 ) | ( x22 & x65 ) | ( ~n26941 & x65 ) ;
  assign n27317 = ( n27315 & ~x65 ) | ( n27315 & n27316 ) | ( ~x65 & n27316 ) ;
  assign n27318 = ( n8606 & ~n8650 ) | ( n8606 & n27317 ) | ( ~n8650 & n27317 ) ;
  assign n27319 = ( n8606 & n26986 ) | ( n8606 & n27317 ) | ( n26986 & n27317 ) ;
  assign n27320 = ( n27318 & ~n27319 ) | ( n27318 & 1'b0 ) | ( ~n27319 & 1'b0 ) ;
  assign n27321 = n27314 | n27320 ;
  assign n27322 = ( n8872 & ~n26986 ) | ( n8872 & 1'b0 ) | ( ~n26986 & 1'b0 ) ;
  assign n27323 = ( x21 & ~n27322 ) | ( x21 & 1'b0 ) | ( ~n27322 & 1'b0 ) ;
  assign n27324 = ( n8877 & ~n26986 ) | ( n8877 & 1'b0 ) | ( ~n26986 & 1'b0 ) ;
  assign n27325 = n27323 | n27324 ;
  assign n27326 = ( x65 & ~n27325 ) | ( x65 & n8880 ) | ( ~n27325 & n8880 ) ;
  assign n27327 = ( x66 & ~n27321 ) | ( x66 & n27326 ) | ( ~n27321 & n27326 ) ;
  assign n27328 = ( x67 & ~n27313 ) | ( x67 & n27327 ) | ( ~n27313 & n27327 ) ;
  assign n27329 = ( x68 & ~n27308 ) | ( x68 & n27328 ) | ( ~n27308 & n27328 ) ;
  assign n27330 = ( x69 & ~n27300 ) | ( x69 & n27329 ) | ( ~n27300 & n27329 ) ;
  assign n27331 = ( x70 & ~n27292 ) | ( x70 & n27330 ) | ( ~n27292 & n27330 ) ;
  assign n27332 = ( x71 & ~n27284 ) | ( x71 & n27331 ) | ( ~n27284 & n27331 ) ;
  assign n27333 = ( x72 & ~n27276 ) | ( x72 & n27332 ) | ( ~n27276 & n27332 ) ;
  assign n27334 = ( x73 & ~n27268 ) | ( x73 & n27333 ) | ( ~n27268 & n27333 ) ;
  assign n27335 = ( x74 & ~n27260 ) | ( x74 & n27334 ) | ( ~n27260 & n27334 ) ;
  assign n27336 = ( x75 & ~n27252 ) | ( x75 & n27335 ) | ( ~n27252 & n27335 ) ;
  assign n27337 = ( x76 & ~n27244 ) | ( x76 & n27336 ) | ( ~n27244 & n27336 ) ;
  assign n27338 = ( x77 & ~n27236 ) | ( x77 & n27337 ) | ( ~n27236 & n27337 ) ;
  assign n27339 = ( x78 & ~n27228 ) | ( x78 & n27338 ) | ( ~n27228 & n27338 ) ;
  assign n27340 = ( x79 & ~n27220 ) | ( x79 & n27339 ) | ( ~n27220 & n27339 ) ;
  assign n27341 = ( x80 & ~n27212 ) | ( x80 & n27340 ) | ( ~n27212 & n27340 ) ;
  assign n27342 = ( x81 & ~n27204 ) | ( x81 & n27341 ) | ( ~n27204 & n27341 ) ;
  assign n27343 = ( x82 & ~n27196 ) | ( x82 & n27342 ) | ( ~n27196 & n27342 ) ;
  assign n27344 = ( x83 & ~n27188 ) | ( x83 & n27343 ) | ( ~n27188 & n27343 ) ;
  assign n27345 = ( x84 & ~n27180 ) | ( x84 & n27344 ) | ( ~n27180 & n27344 ) ;
  assign n27346 = ( x85 & ~n27172 ) | ( x85 & n27345 ) | ( ~n27172 & n27345 ) ;
  assign n27347 = ( x86 & ~n27164 ) | ( x86 & n27346 ) | ( ~n27164 & n27346 ) ;
  assign n27348 = ( x87 & ~n27156 ) | ( x87 & n27347 ) | ( ~n27156 & n27347 ) ;
  assign n27349 = ( x88 & ~n27148 ) | ( x88 & n27348 ) | ( ~n27148 & n27348 ) ;
  assign n27350 = ( x89 & ~n27140 ) | ( x89 & n27349 ) | ( ~n27140 & n27349 ) ;
  assign n27351 = ( x90 & ~n27132 ) | ( x90 & n27350 ) | ( ~n27132 & n27350 ) ;
  assign n27352 = ( x91 & ~n27124 ) | ( x91 & n27351 ) | ( ~n27124 & n27351 ) ;
  assign n27353 = ( x92 & ~n27116 ) | ( x92 & n27352 ) | ( ~n27116 & n27352 ) ;
  assign n27354 = ( x93 & ~n27108 ) | ( x93 & n27353 ) | ( ~n27108 & n27353 ) ;
  assign n27355 = ( x94 & ~n27100 ) | ( x94 & n27354 ) | ( ~n27100 & n27354 ) ;
  assign n27356 = ( x95 & ~n27092 ) | ( x95 & n27355 ) | ( ~n27092 & n27355 ) ;
  assign n27357 = ( x96 & ~n27084 ) | ( x96 & n27356 ) | ( ~n27084 & n27356 ) ;
  assign n27358 = ( x97 & ~n27076 ) | ( x97 & n27357 ) | ( ~n27076 & n27357 ) ;
  assign n27359 = ( x98 & ~n27068 ) | ( x98 & n27358 ) | ( ~n27068 & n27358 ) ;
  assign n27360 = ( x99 & ~n27060 ) | ( x99 & n27359 ) | ( ~n27060 & n27359 ) ;
  assign n27361 = ( x100 & ~n27052 ) | ( x100 & n27360 ) | ( ~n27052 & n27360 ) ;
  assign n27362 = ( x101 & ~n27044 ) | ( x101 & n27361 ) | ( ~n27044 & n27361 ) ;
  assign n27363 = ( x102 & ~n27036 ) | ( x102 & n27362 ) | ( ~n27036 & n27362 ) ;
  assign n27364 = ( x103 & ~n27028 ) | ( x103 & n27363 ) | ( ~n27028 & n27363 ) ;
  assign n27365 = ( x104 & ~n27020 ) | ( x104 & n27364 ) | ( ~n27020 & n27364 ) ;
  assign n27366 = ( x105 & ~n27012 ) | ( x105 & n27365 ) | ( ~n27012 & n27365 ) ;
  assign n27367 = ( x106 & ~n27004 ) | ( x106 & n27366 ) | ( ~n27004 & n27366 ) ;
  assign n26988 = n26625 &  n26987 ;
  assign n26992 = ( n8650 & n26625 ) | ( n8650 & n26985 ) | ( n26625 & n26985 ) ;
  assign n26993 = ( x106 & ~n26992 ) | ( x106 & n26625 ) | ( ~n26992 & n26625 ) ;
  assign n26994 = ~x106 & n26993 ;
  assign n26995 = n26988 | n26994 ;
  assign n26996 = ~x107 & n26995 ;
  assign n27368 = ( x107 & ~n26988 ) | ( x107 & 1'b0 ) | ( ~n26988 & 1'b0 ) ;
  assign n27369 = ~n26994 & n27368 ;
  assign n27378 = n26996 | n27369 ;
  assign n27379 = ( n27367 & ~n27378 ) | ( n27367 & 1'b0 ) | ( ~n27378 & 1'b0 ) ;
  assign n27370 = ( n27367 & ~n26996 ) | ( n27367 & n27369 ) | ( ~n26996 & n27369 ) ;
  assign n27371 = ( n26996 & ~n9044 ) | ( n26996 & n27370 ) | ( ~n9044 & n27370 ) ;
  assign n27372 = n9044 | n27371 ;
  assign n27373 = ~n26995 |  n8650 ;
  assign n27374 = n27372 &  n27373 ;
  assign n27380 = ~n27367 & n27378 ;
  assign n27381 = ( n27379 & ~n27374 ) | ( n27379 & n27380 ) | ( ~n27374 & n27380 ) ;
  assign n27382 = n8650 &  n26625 ;
  assign n27383 = n27372 &  n27382 ;
  assign n27384 = n27381 | n27383 ;
  assign n27385 = ~x108 & n27384 ;
  assign n27389 = n27004 &  n27373 ;
  assign n27390 = n27372 &  n27389 ;
  assign n27375 = x106 | n27004 ;
  assign n27376 = x106 &  n27004 ;
  assign n27377 = ( n27375 & ~n27376 ) | ( n27375 & 1'b0 ) | ( ~n27376 & 1'b0 ) ;
  assign n27392 = ( n27366 & n27374 ) | ( n27366 & n27377 ) | ( n27374 & n27377 ) ;
  assign n27391 = n27366 | n27377 ;
  assign n27393 = ( n27390 & ~n27392 ) | ( n27390 & n27391 ) | ( ~n27392 & n27391 ) ;
  assign n27397 = n27012 &  n27373 ;
  assign n27398 = n27372 &  n27397 ;
  assign n27386 = x105 | n27012 ;
  assign n27387 = x105 &  n27012 ;
  assign n27388 = ( n27386 & ~n27387 ) | ( n27386 & 1'b0 ) | ( ~n27387 & 1'b0 ) ;
  assign n27400 = ( n27365 & n27374 ) | ( n27365 & n27388 ) | ( n27374 & n27388 ) ;
  assign n27399 = n27365 | n27388 ;
  assign n27401 = ( n27398 & ~n27400 ) | ( n27398 & n27399 ) | ( ~n27400 & n27399 ) ;
  assign n27405 = n27020 &  n27373 ;
  assign n27406 = n27372 &  n27405 ;
  assign n27394 = x104 | n27020 ;
  assign n27395 = x104 &  n27020 ;
  assign n27396 = ( n27394 & ~n27395 ) | ( n27394 & 1'b0 ) | ( ~n27395 & 1'b0 ) ;
  assign n27408 = ( n27364 & n27374 ) | ( n27364 & n27396 ) | ( n27374 & n27396 ) ;
  assign n27407 = n27364 | n27396 ;
  assign n27409 = ( n27406 & ~n27408 ) | ( n27406 & n27407 ) | ( ~n27408 & n27407 ) ;
  assign n27413 = n27028 &  n27373 ;
  assign n27414 = n27372 &  n27413 ;
  assign n27402 = x103 | n27028 ;
  assign n27403 = x103 &  n27028 ;
  assign n27404 = ( n27402 & ~n27403 ) | ( n27402 & 1'b0 ) | ( ~n27403 & 1'b0 ) ;
  assign n27416 = ( n27363 & n27374 ) | ( n27363 & n27404 ) | ( n27374 & n27404 ) ;
  assign n27415 = n27363 | n27404 ;
  assign n27417 = ( n27414 & ~n27416 ) | ( n27414 & n27415 ) | ( ~n27416 & n27415 ) ;
  assign n27421 = n27036 &  n27373 ;
  assign n27422 = n27372 &  n27421 ;
  assign n27410 = x102 | n27036 ;
  assign n27411 = x102 &  n27036 ;
  assign n27412 = ( n27410 & ~n27411 ) | ( n27410 & 1'b0 ) | ( ~n27411 & 1'b0 ) ;
  assign n27424 = ( n27362 & n27374 ) | ( n27362 & n27412 ) | ( n27374 & n27412 ) ;
  assign n27423 = n27362 | n27412 ;
  assign n27425 = ( n27422 & ~n27424 ) | ( n27422 & n27423 ) | ( ~n27424 & n27423 ) ;
  assign n27429 = n27044 &  n27373 ;
  assign n27430 = n27372 &  n27429 ;
  assign n27418 = x101 | n27044 ;
  assign n27419 = x101 &  n27044 ;
  assign n27420 = ( n27418 & ~n27419 ) | ( n27418 & 1'b0 ) | ( ~n27419 & 1'b0 ) ;
  assign n27432 = ( n27361 & n27374 ) | ( n27361 & n27420 ) | ( n27374 & n27420 ) ;
  assign n27431 = n27361 | n27420 ;
  assign n27433 = ( n27430 & ~n27432 ) | ( n27430 & n27431 ) | ( ~n27432 & n27431 ) ;
  assign n27437 = n27052 &  n27373 ;
  assign n27438 = n27372 &  n27437 ;
  assign n27426 = x100 | n27052 ;
  assign n27427 = x100 &  n27052 ;
  assign n27428 = ( n27426 & ~n27427 ) | ( n27426 & 1'b0 ) | ( ~n27427 & 1'b0 ) ;
  assign n27440 = ( n27360 & n27374 ) | ( n27360 & n27428 ) | ( n27374 & n27428 ) ;
  assign n27439 = n27360 | n27428 ;
  assign n27441 = ( n27438 & ~n27440 ) | ( n27438 & n27439 ) | ( ~n27440 & n27439 ) ;
  assign n27445 = n27060 &  n27373 ;
  assign n27446 = n27372 &  n27445 ;
  assign n27434 = x99 | n27060 ;
  assign n27435 = x99 &  n27060 ;
  assign n27436 = ( n27434 & ~n27435 ) | ( n27434 & 1'b0 ) | ( ~n27435 & 1'b0 ) ;
  assign n27448 = ( n27359 & n27374 ) | ( n27359 & n27436 ) | ( n27374 & n27436 ) ;
  assign n27447 = n27359 | n27436 ;
  assign n27449 = ( n27446 & ~n27448 ) | ( n27446 & n27447 ) | ( ~n27448 & n27447 ) ;
  assign n27453 = n27068 &  n27373 ;
  assign n27454 = n27372 &  n27453 ;
  assign n27442 = x98 | n27068 ;
  assign n27443 = x98 &  n27068 ;
  assign n27444 = ( n27442 & ~n27443 ) | ( n27442 & 1'b0 ) | ( ~n27443 & 1'b0 ) ;
  assign n27456 = ( n27358 & n27374 ) | ( n27358 & n27444 ) | ( n27374 & n27444 ) ;
  assign n27455 = n27358 | n27444 ;
  assign n27457 = ( n27454 & ~n27456 ) | ( n27454 & n27455 ) | ( ~n27456 & n27455 ) ;
  assign n27461 = n27076 &  n27373 ;
  assign n27462 = n27372 &  n27461 ;
  assign n27450 = x97 | n27076 ;
  assign n27451 = x97 &  n27076 ;
  assign n27452 = ( n27450 & ~n27451 ) | ( n27450 & 1'b0 ) | ( ~n27451 & 1'b0 ) ;
  assign n27464 = ( n27357 & n27374 ) | ( n27357 & n27452 ) | ( n27374 & n27452 ) ;
  assign n27463 = n27357 | n27452 ;
  assign n27465 = ( n27462 & ~n27464 ) | ( n27462 & n27463 ) | ( ~n27464 & n27463 ) ;
  assign n27469 = n27084 &  n27373 ;
  assign n27470 = n27372 &  n27469 ;
  assign n27458 = x96 | n27084 ;
  assign n27459 = x96 &  n27084 ;
  assign n27460 = ( n27458 & ~n27459 ) | ( n27458 & 1'b0 ) | ( ~n27459 & 1'b0 ) ;
  assign n27472 = ( n27356 & n27374 ) | ( n27356 & n27460 ) | ( n27374 & n27460 ) ;
  assign n27471 = n27356 | n27460 ;
  assign n27473 = ( n27470 & ~n27472 ) | ( n27470 & n27471 ) | ( ~n27472 & n27471 ) ;
  assign n27477 = n27092 &  n27373 ;
  assign n27478 = n27372 &  n27477 ;
  assign n27466 = x95 | n27092 ;
  assign n27467 = x95 &  n27092 ;
  assign n27468 = ( n27466 & ~n27467 ) | ( n27466 & 1'b0 ) | ( ~n27467 & 1'b0 ) ;
  assign n27480 = ( n27355 & n27374 ) | ( n27355 & n27468 ) | ( n27374 & n27468 ) ;
  assign n27479 = n27355 | n27468 ;
  assign n27481 = ( n27478 & ~n27480 ) | ( n27478 & n27479 ) | ( ~n27480 & n27479 ) ;
  assign n27485 = n27100 &  n27373 ;
  assign n27486 = n27372 &  n27485 ;
  assign n27474 = x94 | n27100 ;
  assign n27475 = x94 &  n27100 ;
  assign n27476 = ( n27474 & ~n27475 ) | ( n27474 & 1'b0 ) | ( ~n27475 & 1'b0 ) ;
  assign n27488 = ( n27354 & n27374 ) | ( n27354 & n27476 ) | ( n27374 & n27476 ) ;
  assign n27487 = n27354 | n27476 ;
  assign n27489 = ( n27486 & ~n27488 ) | ( n27486 & n27487 ) | ( ~n27488 & n27487 ) ;
  assign n27493 = n27108 &  n27373 ;
  assign n27494 = n27372 &  n27493 ;
  assign n27482 = x93 | n27108 ;
  assign n27483 = x93 &  n27108 ;
  assign n27484 = ( n27482 & ~n27483 ) | ( n27482 & 1'b0 ) | ( ~n27483 & 1'b0 ) ;
  assign n27496 = ( n27353 & n27374 ) | ( n27353 & n27484 ) | ( n27374 & n27484 ) ;
  assign n27495 = n27353 | n27484 ;
  assign n27497 = ( n27494 & ~n27496 ) | ( n27494 & n27495 ) | ( ~n27496 & n27495 ) ;
  assign n27501 = n27116 &  n27373 ;
  assign n27502 = n27372 &  n27501 ;
  assign n27490 = x92 | n27116 ;
  assign n27491 = x92 &  n27116 ;
  assign n27492 = ( n27490 & ~n27491 ) | ( n27490 & 1'b0 ) | ( ~n27491 & 1'b0 ) ;
  assign n27504 = ( n27352 & n27374 ) | ( n27352 & n27492 ) | ( n27374 & n27492 ) ;
  assign n27503 = n27352 | n27492 ;
  assign n27505 = ( n27502 & ~n27504 ) | ( n27502 & n27503 ) | ( ~n27504 & n27503 ) ;
  assign n27509 = n27124 &  n27373 ;
  assign n27510 = n27372 &  n27509 ;
  assign n27498 = x91 | n27124 ;
  assign n27499 = x91 &  n27124 ;
  assign n27500 = ( n27498 & ~n27499 ) | ( n27498 & 1'b0 ) | ( ~n27499 & 1'b0 ) ;
  assign n27512 = ( n27351 & n27374 ) | ( n27351 & n27500 ) | ( n27374 & n27500 ) ;
  assign n27511 = n27351 | n27500 ;
  assign n27513 = ( n27510 & ~n27512 ) | ( n27510 & n27511 ) | ( ~n27512 & n27511 ) ;
  assign n27517 = n27132 &  n27373 ;
  assign n27518 = n27372 &  n27517 ;
  assign n27506 = x90 | n27132 ;
  assign n27507 = x90 &  n27132 ;
  assign n27508 = ( n27506 & ~n27507 ) | ( n27506 & 1'b0 ) | ( ~n27507 & 1'b0 ) ;
  assign n27520 = ( n27350 & n27374 ) | ( n27350 & n27508 ) | ( n27374 & n27508 ) ;
  assign n27519 = n27350 | n27508 ;
  assign n27521 = ( n27518 & ~n27520 ) | ( n27518 & n27519 ) | ( ~n27520 & n27519 ) ;
  assign n27525 = n27140 &  n27373 ;
  assign n27526 = n27372 &  n27525 ;
  assign n27514 = x89 | n27140 ;
  assign n27515 = x89 &  n27140 ;
  assign n27516 = ( n27514 & ~n27515 ) | ( n27514 & 1'b0 ) | ( ~n27515 & 1'b0 ) ;
  assign n27528 = ( n27349 & n27374 ) | ( n27349 & n27516 ) | ( n27374 & n27516 ) ;
  assign n27527 = n27349 | n27516 ;
  assign n27529 = ( n27526 & ~n27528 ) | ( n27526 & n27527 ) | ( ~n27528 & n27527 ) ;
  assign n27533 = n27148 &  n27373 ;
  assign n27534 = n27372 &  n27533 ;
  assign n27522 = x88 | n27148 ;
  assign n27523 = x88 &  n27148 ;
  assign n27524 = ( n27522 & ~n27523 ) | ( n27522 & 1'b0 ) | ( ~n27523 & 1'b0 ) ;
  assign n27536 = ( n27348 & n27374 ) | ( n27348 & n27524 ) | ( n27374 & n27524 ) ;
  assign n27535 = n27348 | n27524 ;
  assign n27537 = ( n27534 & ~n27536 ) | ( n27534 & n27535 ) | ( ~n27536 & n27535 ) ;
  assign n27541 = n27156 &  n27373 ;
  assign n27542 = n27372 &  n27541 ;
  assign n27530 = x87 | n27156 ;
  assign n27531 = x87 &  n27156 ;
  assign n27532 = ( n27530 & ~n27531 ) | ( n27530 & 1'b0 ) | ( ~n27531 & 1'b0 ) ;
  assign n27544 = ( n27347 & n27374 ) | ( n27347 & n27532 ) | ( n27374 & n27532 ) ;
  assign n27543 = n27347 | n27532 ;
  assign n27545 = ( n27542 & ~n27544 ) | ( n27542 & n27543 ) | ( ~n27544 & n27543 ) ;
  assign n27549 = n27164 &  n27373 ;
  assign n27550 = n27372 &  n27549 ;
  assign n27538 = x86 | n27164 ;
  assign n27539 = x86 &  n27164 ;
  assign n27540 = ( n27538 & ~n27539 ) | ( n27538 & 1'b0 ) | ( ~n27539 & 1'b0 ) ;
  assign n27552 = ( n27346 & n27374 ) | ( n27346 & n27540 ) | ( n27374 & n27540 ) ;
  assign n27551 = n27346 | n27540 ;
  assign n27553 = ( n27550 & ~n27552 ) | ( n27550 & n27551 ) | ( ~n27552 & n27551 ) ;
  assign n27557 = n27172 &  n27373 ;
  assign n27558 = n27372 &  n27557 ;
  assign n27546 = x85 | n27172 ;
  assign n27547 = x85 &  n27172 ;
  assign n27548 = ( n27546 & ~n27547 ) | ( n27546 & 1'b0 ) | ( ~n27547 & 1'b0 ) ;
  assign n27560 = ( n27345 & n27374 ) | ( n27345 & n27548 ) | ( n27374 & n27548 ) ;
  assign n27559 = n27345 | n27548 ;
  assign n27561 = ( n27558 & ~n27560 ) | ( n27558 & n27559 ) | ( ~n27560 & n27559 ) ;
  assign n27565 = n27180 &  n27373 ;
  assign n27566 = n27372 &  n27565 ;
  assign n27554 = x84 | n27180 ;
  assign n27555 = x84 &  n27180 ;
  assign n27556 = ( n27554 & ~n27555 ) | ( n27554 & 1'b0 ) | ( ~n27555 & 1'b0 ) ;
  assign n27568 = ( n27344 & n27374 ) | ( n27344 & n27556 ) | ( n27374 & n27556 ) ;
  assign n27567 = n27344 | n27556 ;
  assign n27569 = ( n27566 & ~n27568 ) | ( n27566 & n27567 ) | ( ~n27568 & n27567 ) ;
  assign n27573 = n27188 &  n27373 ;
  assign n27574 = n27372 &  n27573 ;
  assign n27562 = x83 | n27188 ;
  assign n27563 = x83 &  n27188 ;
  assign n27564 = ( n27562 & ~n27563 ) | ( n27562 & 1'b0 ) | ( ~n27563 & 1'b0 ) ;
  assign n27576 = ( n27343 & n27374 ) | ( n27343 & n27564 ) | ( n27374 & n27564 ) ;
  assign n27575 = n27343 | n27564 ;
  assign n27577 = ( n27574 & ~n27576 ) | ( n27574 & n27575 ) | ( ~n27576 & n27575 ) ;
  assign n27581 = n27196 &  n27373 ;
  assign n27582 = n27372 &  n27581 ;
  assign n27570 = x82 | n27196 ;
  assign n27571 = x82 &  n27196 ;
  assign n27572 = ( n27570 & ~n27571 ) | ( n27570 & 1'b0 ) | ( ~n27571 & 1'b0 ) ;
  assign n27584 = ( n27342 & n27374 ) | ( n27342 & n27572 ) | ( n27374 & n27572 ) ;
  assign n27583 = n27342 | n27572 ;
  assign n27585 = ( n27582 & ~n27584 ) | ( n27582 & n27583 ) | ( ~n27584 & n27583 ) ;
  assign n27589 = n27204 &  n27373 ;
  assign n27590 = n27372 &  n27589 ;
  assign n27578 = x81 | n27204 ;
  assign n27579 = x81 &  n27204 ;
  assign n27580 = ( n27578 & ~n27579 ) | ( n27578 & 1'b0 ) | ( ~n27579 & 1'b0 ) ;
  assign n27592 = ( n27341 & n27374 ) | ( n27341 & n27580 ) | ( n27374 & n27580 ) ;
  assign n27591 = n27341 | n27580 ;
  assign n27593 = ( n27590 & ~n27592 ) | ( n27590 & n27591 ) | ( ~n27592 & n27591 ) ;
  assign n27597 = n27212 &  n27373 ;
  assign n27598 = n27372 &  n27597 ;
  assign n27586 = x80 | n27212 ;
  assign n27587 = x80 &  n27212 ;
  assign n27588 = ( n27586 & ~n27587 ) | ( n27586 & 1'b0 ) | ( ~n27587 & 1'b0 ) ;
  assign n27600 = ( n27340 & n27374 ) | ( n27340 & n27588 ) | ( n27374 & n27588 ) ;
  assign n27599 = n27340 | n27588 ;
  assign n27601 = ( n27598 & ~n27600 ) | ( n27598 & n27599 ) | ( ~n27600 & n27599 ) ;
  assign n27605 = n27220 &  n27373 ;
  assign n27606 = n27372 &  n27605 ;
  assign n27594 = x79 | n27220 ;
  assign n27595 = x79 &  n27220 ;
  assign n27596 = ( n27594 & ~n27595 ) | ( n27594 & 1'b0 ) | ( ~n27595 & 1'b0 ) ;
  assign n27608 = ( n27339 & n27374 ) | ( n27339 & n27596 ) | ( n27374 & n27596 ) ;
  assign n27607 = n27339 | n27596 ;
  assign n27609 = ( n27606 & ~n27608 ) | ( n27606 & n27607 ) | ( ~n27608 & n27607 ) ;
  assign n27613 = n27228 &  n27373 ;
  assign n27614 = n27372 &  n27613 ;
  assign n27602 = x78 | n27228 ;
  assign n27603 = x78 &  n27228 ;
  assign n27604 = ( n27602 & ~n27603 ) | ( n27602 & 1'b0 ) | ( ~n27603 & 1'b0 ) ;
  assign n27616 = ( n27338 & n27374 ) | ( n27338 & n27604 ) | ( n27374 & n27604 ) ;
  assign n27615 = n27338 | n27604 ;
  assign n27617 = ( n27614 & ~n27616 ) | ( n27614 & n27615 ) | ( ~n27616 & n27615 ) ;
  assign n27621 = n27236 &  n27373 ;
  assign n27622 = n27372 &  n27621 ;
  assign n27610 = x77 | n27236 ;
  assign n27611 = x77 &  n27236 ;
  assign n27612 = ( n27610 & ~n27611 ) | ( n27610 & 1'b0 ) | ( ~n27611 & 1'b0 ) ;
  assign n27624 = ( n27337 & n27374 ) | ( n27337 & n27612 ) | ( n27374 & n27612 ) ;
  assign n27623 = n27337 | n27612 ;
  assign n27625 = ( n27622 & ~n27624 ) | ( n27622 & n27623 ) | ( ~n27624 & n27623 ) ;
  assign n27629 = n27244 &  n27373 ;
  assign n27630 = n27372 &  n27629 ;
  assign n27618 = x76 | n27244 ;
  assign n27619 = x76 &  n27244 ;
  assign n27620 = ( n27618 & ~n27619 ) | ( n27618 & 1'b0 ) | ( ~n27619 & 1'b0 ) ;
  assign n27632 = ( n27336 & n27374 ) | ( n27336 & n27620 ) | ( n27374 & n27620 ) ;
  assign n27631 = n27336 | n27620 ;
  assign n27633 = ( n27630 & ~n27632 ) | ( n27630 & n27631 ) | ( ~n27632 & n27631 ) ;
  assign n27637 = n27252 &  n27373 ;
  assign n27638 = n27372 &  n27637 ;
  assign n27626 = x75 | n27252 ;
  assign n27627 = x75 &  n27252 ;
  assign n27628 = ( n27626 & ~n27627 ) | ( n27626 & 1'b0 ) | ( ~n27627 & 1'b0 ) ;
  assign n27640 = ( n27335 & n27374 ) | ( n27335 & n27628 ) | ( n27374 & n27628 ) ;
  assign n27639 = n27335 | n27628 ;
  assign n27641 = ( n27638 & ~n27640 ) | ( n27638 & n27639 ) | ( ~n27640 & n27639 ) ;
  assign n27645 = n27260 &  n27373 ;
  assign n27646 = n27372 &  n27645 ;
  assign n27634 = x74 | n27260 ;
  assign n27635 = x74 &  n27260 ;
  assign n27636 = ( n27634 & ~n27635 ) | ( n27634 & 1'b0 ) | ( ~n27635 & 1'b0 ) ;
  assign n27648 = ( n27334 & n27374 ) | ( n27334 & n27636 ) | ( n27374 & n27636 ) ;
  assign n27647 = n27334 | n27636 ;
  assign n27649 = ( n27646 & ~n27648 ) | ( n27646 & n27647 ) | ( ~n27648 & n27647 ) ;
  assign n27653 = n27268 &  n27373 ;
  assign n27654 = n27372 &  n27653 ;
  assign n27642 = x73 | n27268 ;
  assign n27643 = x73 &  n27268 ;
  assign n27644 = ( n27642 & ~n27643 ) | ( n27642 & 1'b0 ) | ( ~n27643 & 1'b0 ) ;
  assign n27656 = ( n27333 & n27374 ) | ( n27333 & n27644 ) | ( n27374 & n27644 ) ;
  assign n27655 = n27333 | n27644 ;
  assign n27657 = ( n27654 & ~n27656 ) | ( n27654 & n27655 ) | ( ~n27656 & n27655 ) ;
  assign n27661 = n27276 &  n27373 ;
  assign n27662 = n27372 &  n27661 ;
  assign n27650 = x72 | n27276 ;
  assign n27651 = x72 &  n27276 ;
  assign n27652 = ( n27650 & ~n27651 ) | ( n27650 & 1'b0 ) | ( ~n27651 & 1'b0 ) ;
  assign n27664 = ( n27332 & n27374 ) | ( n27332 & n27652 ) | ( n27374 & n27652 ) ;
  assign n27663 = n27332 | n27652 ;
  assign n27665 = ( n27662 & ~n27664 ) | ( n27662 & n27663 ) | ( ~n27664 & n27663 ) ;
  assign n27669 = n27284 &  n27373 ;
  assign n27670 = n27372 &  n27669 ;
  assign n27658 = x71 | n27284 ;
  assign n27659 = x71 &  n27284 ;
  assign n27660 = ( n27658 & ~n27659 ) | ( n27658 & 1'b0 ) | ( ~n27659 & 1'b0 ) ;
  assign n27672 = ( n27331 & n27374 ) | ( n27331 & n27660 ) | ( n27374 & n27660 ) ;
  assign n27671 = n27331 | n27660 ;
  assign n27673 = ( n27670 & ~n27672 ) | ( n27670 & n27671 ) | ( ~n27672 & n27671 ) ;
  assign n27677 = n27292 &  n27373 ;
  assign n27678 = n27372 &  n27677 ;
  assign n27666 = x70 | n27292 ;
  assign n27667 = x70 &  n27292 ;
  assign n27668 = ( n27666 & ~n27667 ) | ( n27666 & 1'b0 ) | ( ~n27667 & 1'b0 ) ;
  assign n27680 = ( n27330 & n27374 ) | ( n27330 & n27668 ) | ( n27374 & n27668 ) ;
  assign n27679 = n27330 | n27668 ;
  assign n27681 = ( n27678 & ~n27680 ) | ( n27678 & n27679 ) | ( ~n27680 & n27679 ) ;
  assign n27685 = n27300 &  n27373 ;
  assign n27686 = n27372 &  n27685 ;
  assign n27674 = x69 | n27300 ;
  assign n27675 = x69 &  n27300 ;
  assign n27676 = ( n27674 & ~n27675 ) | ( n27674 & 1'b0 ) | ( ~n27675 & 1'b0 ) ;
  assign n27688 = ( n27329 & n27374 ) | ( n27329 & n27676 ) | ( n27374 & n27676 ) ;
  assign n27687 = n27329 | n27676 ;
  assign n27689 = ( n27686 & ~n27688 ) | ( n27686 & n27687 ) | ( ~n27688 & n27687 ) ;
  assign n27693 = n27308 &  n27373 ;
  assign n27694 = n27372 &  n27693 ;
  assign n27682 = x68 | n27308 ;
  assign n27683 = x68 &  n27308 ;
  assign n27684 = ( n27682 & ~n27683 ) | ( n27682 & 1'b0 ) | ( ~n27683 & 1'b0 ) ;
  assign n27696 = ( n27328 & n27374 ) | ( n27328 & n27684 ) | ( n27374 & n27684 ) ;
  assign n27695 = n27328 | n27684 ;
  assign n27697 = ( n27694 & ~n27696 ) | ( n27694 & n27695 ) | ( ~n27696 & n27695 ) ;
  assign n27701 = n27313 &  n27373 ;
  assign n27702 = n27372 &  n27701 ;
  assign n27690 = x67 | n27313 ;
  assign n27691 = x67 &  n27313 ;
  assign n27692 = ( n27690 & ~n27691 ) | ( n27690 & 1'b0 ) | ( ~n27691 & 1'b0 ) ;
  assign n27704 = ( n27327 & n27374 ) | ( n27327 & n27692 ) | ( n27374 & n27692 ) ;
  assign n27703 = n27327 | n27692 ;
  assign n27705 = ( n27702 & ~n27704 ) | ( n27702 & n27703 ) | ( ~n27704 & n27703 ) ;
  assign n27706 = n27321 &  n27373 ;
  assign n27707 = n27372 &  n27706 ;
  assign n27698 = x66 | n27321 ;
  assign n27699 = x66 &  n27321 ;
  assign n27700 = ( n27698 & ~n27699 ) | ( n27698 & 1'b0 ) | ( ~n27699 & 1'b0 ) ;
  assign n27709 = ( n27326 & n27374 ) | ( n27326 & n27700 ) | ( n27374 & n27700 ) ;
  assign n27708 = n27326 | n27700 ;
  assign n27710 = ( n27707 & ~n27709 ) | ( n27707 & n27708 ) | ( ~n27709 & n27708 ) ;
  assign n27711 = ( x65 & ~n8880 ) | ( x65 & n27325 ) | ( ~n8880 & n27325 ) ;
  assign n27712 = ( n27326 & ~x65 ) | ( n27326 & n27711 ) | ( ~x65 & n27711 ) ;
  assign n27713 = ~n27374 & n27712 ;
  assign n27714 = n27325 &  n27373 ;
  assign n27715 = n27372 &  n27714 ;
  assign n27716 = n27713 | n27715 ;
  assign n27717 = ( x64 & ~n27374 ) | ( x64 & 1'b0 ) | ( ~n27374 & 1'b0 ) ;
  assign n27718 = ( x20 & ~n27717 ) | ( x20 & 1'b0 ) | ( ~n27717 & 1'b0 ) ;
  assign n27719 = ( n8880 & ~n27374 ) | ( n8880 & 1'b0 ) | ( ~n27374 & 1'b0 ) ;
  assign n27720 = n27718 | n27719 ;
  assign n27721 = ( x65 & ~n27720 ) | ( x65 & n9279 ) | ( ~n27720 & n9279 ) ;
  assign n27722 = ( x66 & ~n27716 ) | ( x66 & n27721 ) | ( ~n27716 & n27721 ) ;
  assign n27723 = ( x67 & ~n27710 ) | ( x67 & n27722 ) | ( ~n27710 & n27722 ) ;
  assign n27724 = ( x68 & ~n27705 ) | ( x68 & n27723 ) | ( ~n27705 & n27723 ) ;
  assign n27725 = ( x69 & ~n27697 ) | ( x69 & n27724 ) | ( ~n27697 & n27724 ) ;
  assign n27726 = ( x70 & ~n27689 ) | ( x70 & n27725 ) | ( ~n27689 & n27725 ) ;
  assign n27727 = ( x71 & ~n27681 ) | ( x71 & n27726 ) | ( ~n27681 & n27726 ) ;
  assign n27728 = ( x72 & ~n27673 ) | ( x72 & n27727 ) | ( ~n27673 & n27727 ) ;
  assign n27729 = ( x73 & ~n27665 ) | ( x73 & n27728 ) | ( ~n27665 & n27728 ) ;
  assign n27730 = ( x74 & ~n27657 ) | ( x74 & n27729 ) | ( ~n27657 & n27729 ) ;
  assign n27731 = ( x75 & ~n27649 ) | ( x75 & n27730 ) | ( ~n27649 & n27730 ) ;
  assign n27732 = ( x76 & ~n27641 ) | ( x76 & n27731 ) | ( ~n27641 & n27731 ) ;
  assign n27733 = ( x77 & ~n27633 ) | ( x77 & n27732 ) | ( ~n27633 & n27732 ) ;
  assign n27734 = ( x78 & ~n27625 ) | ( x78 & n27733 ) | ( ~n27625 & n27733 ) ;
  assign n27735 = ( x79 & ~n27617 ) | ( x79 & n27734 ) | ( ~n27617 & n27734 ) ;
  assign n27736 = ( x80 & ~n27609 ) | ( x80 & n27735 ) | ( ~n27609 & n27735 ) ;
  assign n27737 = ( x81 & ~n27601 ) | ( x81 & n27736 ) | ( ~n27601 & n27736 ) ;
  assign n27738 = ( x82 & ~n27593 ) | ( x82 & n27737 ) | ( ~n27593 & n27737 ) ;
  assign n27739 = ( x83 & ~n27585 ) | ( x83 & n27738 ) | ( ~n27585 & n27738 ) ;
  assign n27740 = ( x84 & ~n27577 ) | ( x84 & n27739 ) | ( ~n27577 & n27739 ) ;
  assign n27741 = ( x85 & ~n27569 ) | ( x85 & n27740 ) | ( ~n27569 & n27740 ) ;
  assign n27742 = ( x86 & ~n27561 ) | ( x86 & n27741 ) | ( ~n27561 & n27741 ) ;
  assign n27743 = ( x87 & ~n27553 ) | ( x87 & n27742 ) | ( ~n27553 & n27742 ) ;
  assign n27744 = ( x88 & ~n27545 ) | ( x88 & n27743 ) | ( ~n27545 & n27743 ) ;
  assign n27745 = ( x89 & ~n27537 ) | ( x89 & n27744 ) | ( ~n27537 & n27744 ) ;
  assign n27746 = ( x90 & ~n27529 ) | ( x90 & n27745 ) | ( ~n27529 & n27745 ) ;
  assign n27747 = ( x91 & ~n27521 ) | ( x91 & n27746 ) | ( ~n27521 & n27746 ) ;
  assign n27748 = ( x92 & ~n27513 ) | ( x92 & n27747 ) | ( ~n27513 & n27747 ) ;
  assign n27749 = ( x93 & ~n27505 ) | ( x93 & n27748 ) | ( ~n27505 & n27748 ) ;
  assign n27750 = ( x94 & ~n27497 ) | ( x94 & n27749 ) | ( ~n27497 & n27749 ) ;
  assign n27751 = ( x95 & ~n27489 ) | ( x95 & n27750 ) | ( ~n27489 & n27750 ) ;
  assign n27752 = ( x96 & ~n27481 ) | ( x96 & n27751 ) | ( ~n27481 & n27751 ) ;
  assign n27753 = ( x97 & ~n27473 ) | ( x97 & n27752 ) | ( ~n27473 & n27752 ) ;
  assign n27754 = ( x98 & ~n27465 ) | ( x98 & n27753 ) | ( ~n27465 & n27753 ) ;
  assign n27755 = ( x99 & ~n27457 ) | ( x99 & n27754 ) | ( ~n27457 & n27754 ) ;
  assign n27756 = ( x100 & ~n27449 ) | ( x100 & n27755 ) | ( ~n27449 & n27755 ) ;
  assign n27757 = ( x101 & ~n27441 ) | ( x101 & n27756 ) | ( ~n27441 & n27756 ) ;
  assign n27758 = ( x102 & ~n27433 ) | ( x102 & n27757 ) | ( ~n27433 & n27757 ) ;
  assign n27759 = ( x103 & ~n27425 ) | ( x103 & n27758 ) | ( ~n27425 & n27758 ) ;
  assign n27760 = ( x104 & ~n27417 ) | ( x104 & n27759 ) | ( ~n27417 & n27759 ) ;
  assign n27761 = ( x105 & ~n27409 ) | ( x105 & n27760 ) | ( ~n27409 & n27760 ) ;
  assign n27762 = ( x106 & ~n27401 ) | ( x106 & n27761 ) | ( ~n27401 & n27761 ) ;
  assign n27763 = ( x107 & ~n27393 ) | ( x107 & n27762 ) | ( ~n27393 & n27762 ) ;
  assign n27764 = ( x108 & ~n27383 ) | ( x108 & 1'b0 ) | ( ~n27383 & 1'b0 ) ;
  assign n27765 = ~n27381 & n27764 ;
  assign n27766 = ( n27763 & ~n27385 ) | ( n27763 & n27765 ) | ( ~n27385 & n27765 ) ;
  assign n27767 = ( n27385 & ~n9440 ) | ( n27385 & n27766 ) | ( ~n9440 & n27766 ) ;
  assign n27768 = n9440 | n27767 ;
  assign n27769 = ~n27384 |  n9044 ;
  assign n27783 = n27393 &  n27769 ;
  assign n27784 = n27768 &  n27783 ;
  assign n27770 = n27768 &  n27769 ;
  assign n27771 = x107 | n27393 ;
  assign n27772 = x107 &  n27393 ;
  assign n27773 = ( n27771 & ~n27772 ) | ( n27771 & 1'b0 ) | ( ~n27772 & 1'b0 ) ;
  assign n27786 = ( n27762 & n27770 ) | ( n27762 & n27773 ) | ( n27770 & n27773 ) ;
  assign n27785 = n27762 | n27773 ;
  assign n27787 = ( n27784 & ~n27786 ) | ( n27784 & n27785 ) | ( ~n27786 & n27785 ) ;
  assign n27775 = n9044 &  n27384 ;
  assign n27776 = n27768 &  n27775 ;
  assign n27774 = n27385 | n27765 ;
  assign n27778 = ( n27763 & n27770 ) | ( n27763 & n27774 ) | ( n27770 & n27774 ) ;
  assign n27777 = n27763 | n27774 ;
  assign n27779 = ( n27776 & ~n27778 ) | ( n27776 & n27777 ) | ( ~n27778 & n27777 ) ;
  assign n27791 = n27401 &  n27769 ;
  assign n27792 = n27768 &  n27791 ;
  assign n27780 = x106 | n27401 ;
  assign n27781 = x106 &  n27401 ;
  assign n27782 = ( n27780 & ~n27781 ) | ( n27780 & 1'b0 ) | ( ~n27781 & 1'b0 ) ;
  assign n27794 = ( n27761 & n27770 ) | ( n27761 & n27782 ) | ( n27770 & n27782 ) ;
  assign n27793 = n27761 | n27782 ;
  assign n27795 = ( n27792 & ~n27794 ) | ( n27792 & n27793 ) | ( ~n27794 & n27793 ) ;
  assign n27799 = n27409 &  n27769 ;
  assign n27800 = n27768 &  n27799 ;
  assign n27788 = x105 | n27409 ;
  assign n27789 = x105 &  n27409 ;
  assign n27790 = ( n27788 & ~n27789 ) | ( n27788 & 1'b0 ) | ( ~n27789 & 1'b0 ) ;
  assign n27802 = ( n27760 & n27770 ) | ( n27760 & n27790 ) | ( n27770 & n27790 ) ;
  assign n27801 = n27760 | n27790 ;
  assign n27803 = ( n27800 & ~n27802 ) | ( n27800 & n27801 ) | ( ~n27802 & n27801 ) ;
  assign n27807 = n27417 &  n27769 ;
  assign n27808 = n27768 &  n27807 ;
  assign n27796 = x104 | n27417 ;
  assign n27797 = x104 &  n27417 ;
  assign n27798 = ( n27796 & ~n27797 ) | ( n27796 & 1'b0 ) | ( ~n27797 & 1'b0 ) ;
  assign n27810 = ( n27759 & n27770 ) | ( n27759 & n27798 ) | ( n27770 & n27798 ) ;
  assign n27809 = n27759 | n27798 ;
  assign n27811 = ( n27808 & ~n27810 ) | ( n27808 & n27809 ) | ( ~n27810 & n27809 ) ;
  assign n27815 = n27425 &  n27769 ;
  assign n27816 = n27768 &  n27815 ;
  assign n27804 = x103 | n27425 ;
  assign n27805 = x103 &  n27425 ;
  assign n27806 = ( n27804 & ~n27805 ) | ( n27804 & 1'b0 ) | ( ~n27805 & 1'b0 ) ;
  assign n27818 = ( n27758 & n27770 ) | ( n27758 & n27806 ) | ( n27770 & n27806 ) ;
  assign n27817 = n27758 | n27806 ;
  assign n27819 = ( n27816 & ~n27818 ) | ( n27816 & n27817 ) | ( ~n27818 & n27817 ) ;
  assign n27823 = n27433 &  n27769 ;
  assign n27824 = n27768 &  n27823 ;
  assign n27812 = x102 | n27433 ;
  assign n27813 = x102 &  n27433 ;
  assign n27814 = ( n27812 & ~n27813 ) | ( n27812 & 1'b0 ) | ( ~n27813 & 1'b0 ) ;
  assign n27826 = ( n27757 & n27770 ) | ( n27757 & n27814 ) | ( n27770 & n27814 ) ;
  assign n27825 = n27757 | n27814 ;
  assign n27827 = ( n27824 & ~n27826 ) | ( n27824 & n27825 ) | ( ~n27826 & n27825 ) ;
  assign n27831 = n27441 &  n27769 ;
  assign n27832 = n27768 &  n27831 ;
  assign n27820 = x101 | n27441 ;
  assign n27821 = x101 &  n27441 ;
  assign n27822 = ( n27820 & ~n27821 ) | ( n27820 & 1'b0 ) | ( ~n27821 & 1'b0 ) ;
  assign n27834 = ( n27756 & n27770 ) | ( n27756 & n27822 ) | ( n27770 & n27822 ) ;
  assign n27833 = n27756 | n27822 ;
  assign n27835 = ( n27832 & ~n27834 ) | ( n27832 & n27833 ) | ( ~n27834 & n27833 ) ;
  assign n27839 = n27449 &  n27769 ;
  assign n27840 = n27768 &  n27839 ;
  assign n27828 = x100 | n27449 ;
  assign n27829 = x100 &  n27449 ;
  assign n27830 = ( n27828 & ~n27829 ) | ( n27828 & 1'b0 ) | ( ~n27829 & 1'b0 ) ;
  assign n27842 = ( n27755 & n27770 ) | ( n27755 & n27830 ) | ( n27770 & n27830 ) ;
  assign n27841 = n27755 | n27830 ;
  assign n27843 = ( n27840 & ~n27842 ) | ( n27840 & n27841 ) | ( ~n27842 & n27841 ) ;
  assign n27847 = n27457 &  n27769 ;
  assign n27848 = n27768 &  n27847 ;
  assign n27836 = x99 | n27457 ;
  assign n27837 = x99 &  n27457 ;
  assign n27838 = ( n27836 & ~n27837 ) | ( n27836 & 1'b0 ) | ( ~n27837 & 1'b0 ) ;
  assign n27850 = ( n27754 & n27770 ) | ( n27754 & n27838 ) | ( n27770 & n27838 ) ;
  assign n27849 = n27754 | n27838 ;
  assign n27851 = ( n27848 & ~n27850 ) | ( n27848 & n27849 ) | ( ~n27850 & n27849 ) ;
  assign n27855 = n27465 &  n27769 ;
  assign n27856 = n27768 &  n27855 ;
  assign n27844 = x98 | n27465 ;
  assign n27845 = x98 &  n27465 ;
  assign n27846 = ( n27844 & ~n27845 ) | ( n27844 & 1'b0 ) | ( ~n27845 & 1'b0 ) ;
  assign n27858 = ( n27753 & n27770 ) | ( n27753 & n27846 ) | ( n27770 & n27846 ) ;
  assign n27857 = n27753 | n27846 ;
  assign n27859 = ( n27856 & ~n27858 ) | ( n27856 & n27857 ) | ( ~n27858 & n27857 ) ;
  assign n27863 = n27473 &  n27769 ;
  assign n27864 = n27768 &  n27863 ;
  assign n27852 = x97 | n27473 ;
  assign n27853 = x97 &  n27473 ;
  assign n27854 = ( n27852 & ~n27853 ) | ( n27852 & 1'b0 ) | ( ~n27853 & 1'b0 ) ;
  assign n27866 = ( n27752 & n27770 ) | ( n27752 & n27854 ) | ( n27770 & n27854 ) ;
  assign n27865 = n27752 | n27854 ;
  assign n27867 = ( n27864 & ~n27866 ) | ( n27864 & n27865 ) | ( ~n27866 & n27865 ) ;
  assign n27871 = n27481 &  n27769 ;
  assign n27872 = n27768 &  n27871 ;
  assign n27860 = x96 | n27481 ;
  assign n27861 = x96 &  n27481 ;
  assign n27862 = ( n27860 & ~n27861 ) | ( n27860 & 1'b0 ) | ( ~n27861 & 1'b0 ) ;
  assign n27874 = ( n27751 & n27770 ) | ( n27751 & n27862 ) | ( n27770 & n27862 ) ;
  assign n27873 = n27751 | n27862 ;
  assign n27875 = ( n27872 & ~n27874 ) | ( n27872 & n27873 ) | ( ~n27874 & n27873 ) ;
  assign n27879 = n27489 &  n27769 ;
  assign n27880 = n27768 &  n27879 ;
  assign n27868 = x95 | n27489 ;
  assign n27869 = x95 &  n27489 ;
  assign n27870 = ( n27868 & ~n27869 ) | ( n27868 & 1'b0 ) | ( ~n27869 & 1'b0 ) ;
  assign n27882 = ( n27750 & n27770 ) | ( n27750 & n27870 ) | ( n27770 & n27870 ) ;
  assign n27881 = n27750 | n27870 ;
  assign n27883 = ( n27880 & ~n27882 ) | ( n27880 & n27881 ) | ( ~n27882 & n27881 ) ;
  assign n27887 = n27497 &  n27769 ;
  assign n27888 = n27768 &  n27887 ;
  assign n27876 = x94 | n27497 ;
  assign n27877 = x94 &  n27497 ;
  assign n27878 = ( n27876 & ~n27877 ) | ( n27876 & 1'b0 ) | ( ~n27877 & 1'b0 ) ;
  assign n27890 = ( n27749 & n27770 ) | ( n27749 & n27878 ) | ( n27770 & n27878 ) ;
  assign n27889 = n27749 | n27878 ;
  assign n27891 = ( n27888 & ~n27890 ) | ( n27888 & n27889 ) | ( ~n27890 & n27889 ) ;
  assign n27895 = n27505 &  n27769 ;
  assign n27896 = n27768 &  n27895 ;
  assign n27884 = x93 | n27505 ;
  assign n27885 = x93 &  n27505 ;
  assign n27886 = ( n27884 & ~n27885 ) | ( n27884 & 1'b0 ) | ( ~n27885 & 1'b0 ) ;
  assign n27898 = ( n27748 & n27770 ) | ( n27748 & n27886 ) | ( n27770 & n27886 ) ;
  assign n27897 = n27748 | n27886 ;
  assign n27899 = ( n27896 & ~n27898 ) | ( n27896 & n27897 ) | ( ~n27898 & n27897 ) ;
  assign n27903 = n27513 &  n27769 ;
  assign n27904 = n27768 &  n27903 ;
  assign n27892 = x92 | n27513 ;
  assign n27893 = x92 &  n27513 ;
  assign n27894 = ( n27892 & ~n27893 ) | ( n27892 & 1'b0 ) | ( ~n27893 & 1'b0 ) ;
  assign n27906 = ( n27747 & n27770 ) | ( n27747 & n27894 ) | ( n27770 & n27894 ) ;
  assign n27905 = n27747 | n27894 ;
  assign n27907 = ( n27904 & ~n27906 ) | ( n27904 & n27905 ) | ( ~n27906 & n27905 ) ;
  assign n27911 = n27521 &  n27769 ;
  assign n27912 = n27768 &  n27911 ;
  assign n27900 = x91 | n27521 ;
  assign n27901 = x91 &  n27521 ;
  assign n27902 = ( n27900 & ~n27901 ) | ( n27900 & 1'b0 ) | ( ~n27901 & 1'b0 ) ;
  assign n27914 = ( n27746 & n27770 ) | ( n27746 & n27902 ) | ( n27770 & n27902 ) ;
  assign n27913 = n27746 | n27902 ;
  assign n27915 = ( n27912 & ~n27914 ) | ( n27912 & n27913 ) | ( ~n27914 & n27913 ) ;
  assign n27919 = n27529 &  n27769 ;
  assign n27920 = n27768 &  n27919 ;
  assign n27908 = x90 | n27529 ;
  assign n27909 = x90 &  n27529 ;
  assign n27910 = ( n27908 & ~n27909 ) | ( n27908 & 1'b0 ) | ( ~n27909 & 1'b0 ) ;
  assign n27922 = ( n27745 & n27770 ) | ( n27745 & n27910 ) | ( n27770 & n27910 ) ;
  assign n27921 = n27745 | n27910 ;
  assign n27923 = ( n27920 & ~n27922 ) | ( n27920 & n27921 ) | ( ~n27922 & n27921 ) ;
  assign n27927 = n27537 &  n27769 ;
  assign n27928 = n27768 &  n27927 ;
  assign n27916 = x89 | n27537 ;
  assign n27917 = x89 &  n27537 ;
  assign n27918 = ( n27916 & ~n27917 ) | ( n27916 & 1'b0 ) | ( ~n27917 & 1'b0 ) ;
  assign n27930 = ( n27744 & n27770 ) | ( n27744 & n27918 ) | ( n27770 & n27918 ) ;
  assign n27929 = n27744 | n27918 ;
  assign n27931 = ( n27928 & ~n27930 ) | ( n27928 & n27929 ) | ( ~n27930 & n27929 ) ;
  assign n27935 = n27545 &  n27769 ;
  assign n27936 = n27768 &  n27935 ;
  assign n27924 = x88 | n27545 ;
  assign n27925 = x88 &  n27545 ;
  assign n27926 = ( n27924 & ~n27925 ) | ( n27924 & 1'b0 ) | ( ~n27925 & 1'b0 ) ;
  assign n27938 = ( n27743 & n27770 ) | ( n27743 & n27926 ) | ( n27770 & n27926 ) ;
  assign n27937 = n27743 | n27926 ;
  assign n27939 = ( n27936 & ~n27938 ) | ( n27936 & n27937 ) | ( ~n27938 & n27937 ) ;
  assign n27943 = n27553 &  n27769 ;
  assign n27944 = n27768 &  n27943 ;
  assign n27932 = x87 | n27553 ;
  assign n27933 = x87 &  n27553 ;
  assign n27934 = ( n27932 & ~n27933 ) | ( n27932 & 1'b0 ) | ( ~n27933 & 1'b0 ) ;
  assign n27946 = ( n27742 & n27770 ) | ( n27742 & n27934 ) | ( n27770 & n27934 ) ;
  assign n27945 = n27742 | n27934 ;
  assign n27947 = ( n27944 & ~n27946 ) | ( n27944 & n27945 ) | ( ~n27946 & n27945 ) ;
  assign n27951 = n27561 &  n27769 ;
  assign n27952 = n27768 &  n27951 ;
  assign n27940 = x86 | n27561 ;
  assign n27941 = x86 &  n27561 ;
  assign n27942 = ( n27940 & ~n27941 ) | ( n27940 & 1'b0 ) | ( ~n27941 & 1'b0 ) ;
  assign n27954 = ( n27741 & n27770 ) | ( n27741 & n27942 ) | ( n27770 & n27942 ) ;
  assign n27953 = n27741 | n27942 ;
  assign n27955 = ( n27952 & ~n27954 ) | ( n27952 & n27953 ) | ( ~n27954 & n27953 ) ;
  assign n27959 = n27569 &  n27769 ;
  assign n27960 = n27768 &  n27959 ;
  assign n27948 = x85 | n27569 ;
  assign n27949 = x85 &  n27569 ;
  assign n27950 = ( n27948 & ~n27949 ) | ( n27948 & 1'b0 ) | ( ~n27949 & 1'b0 ) ;
  assign n27962 = ( n27740 & n27770 ) | ( n27740 & n27950 ) | ( n27770 & n27950 ) ;
  assign n27961 = n27740 | n27950 ;
  assign n27963 = ( n27960 & ~n27962 ) | ( n27960 & n27961 ) | ( ~n27962 & n27961 ) ;
  assign n27967 = n27577 &  n27769 ;
  assign n27968 = n27768 &  n27967 ;
  assign n27956 = x84 | n27577 ;
  assign n27957 = x84 &  n27577 ;
  assign n27958 = ( n27956 & ~n27957 ) | ( n27956 & 1'b0 ) | ( ~n27957 & 1'b0 ) ;
  assign n27970 = ( n27739 & n27770 ) | ( n27739 & n27958 ) | ( n27770 & n27958 ) ;
  assign n27969 = n27739 | n27958 ;
  assign n27971 = ( n27968 & ~n27970 ) | ( n27968 & n27969 ) | ( ~n27970 & n27969 ) ;
  assign n27975 = n27585 &  n27769 ;
  assign n27976 = n27768 &  n27975 ;
  assign n27964 = x83 | n27585 ;
  assign n27965 = x83 &  n27585 ;
  assign n27966 = ( n27964 & ~n27965 ) | ( n27964 & 1'b0 ) | ( ~n27965 & 1'b0 ) ;
  assign n27978 = ( n27738 & n27770 ) | ( n27738 & n27966 ) | ( n27770 & n27966 ) ;
  assign n27977 = n27738 | n27966 ;
  assign n27979 = ( n27976 & ~n27978 ) | ( n27976 & n27977 ) | ( ~n27978 & n27977 ) ;
  assign n27983 = n27593 &  n27769 ;
  assign n27984 = n27768 &  n27983 ;
  assign n27972 = x82 | n27593 ;
  assign n27973 = x82 &  n27593 ;
  assign n27974 = ( n27972 & ~n27973 ) | ( n27972 & 1'b0 ) | ( ~n27973 & 1'b0 ) ;
  assign n27986 = ( n27737 & n27770 ) | ( n27737 & n27974 ) | ( n27770 & n27974 ) ;
  assign n27985 = n27737 | n27974 ;
  assign n27987 = ( n27984 & ~n27986 ) | ( n27984 & n27985 ) | ( ~n27986 & n27985 ) ;
  assign n27991 = n27601 &  n27769 ;
  assign n27992 = n27768 &  n27991 ;
  assign n27980 = x81 | n27601 ;
  assign n27981 = x81 &  n27601 ;
  assign n27982 = ( n27980 & ~n27981 ) | ( n27980 & 1'b0 ) | ( ~n27981 & 1'b0 ) ;
  assign n27994 = ( n27736 & n27770 ) | ( n27736 & n27982 ) | ( n27770 & n27982 ) ;
  assign n27993 = n27736 | n27982 ;
  assign n27995 = ( n27992 & ~n27994 ) | ( n27992 & n27993 ) | ( ~n27994 & n27993 ) ;
  assign n27999 = n27609 &  n27769 ;
  assign n28000 = n27768 &  n27999 ;
  assign n27988 = x80 | n27609 ;
  assign n27989 = x80 &  n27609 ;
  assign n27990 = ( n27988 & ~n27989 ) | ( n27988 & 1'b0 ) | ( ~n27989 & 1'b0 ) ;
  assign n28002 = ( n27735 & n27770 ) | ( n27735 & n27990 ) | ( n27770 & n27990 ) ;
  assign n28001 = n27735 | n27990 ;
  assign n28003 = ( n28000 & ~n28002 ) | ( n28000 & n28001 ) | ( ~n28002 & n28001 ) ;
  assign n28007 = n27617 &  n27769 ;
  assign n28008 = n27768 &  n28007 ;
  assign n27996 = x79 | n27617 ;
  assign n27997 = x79 &  n27617 ;
  assign n27998 = ( n27996 & ~n27997 ) | ( n27996 & 1'b0 ) | ( ~n27997 & 1'b0 ) ;
  assign n28010 = ( n27734 & n27770 ) | ( n27734 & n27998 ) | ( n27770 & n27998 ) ;
  assign n28009 = n27734 | n27998 ;
  assign n28011 = ( n28008 & ~n28010 ) | ( n28008 & n28009 ) | ( ~n28010 & n28009 ) ;
  assign n28015 = n27625 &  n27769 ;
  assign n28016 = n27768 &  n28015 ;
  assign n28004 = x78 | n27625 ;
  assign n28005 = x78 &  n27625 ;
  assign n28006 = ( n28004 & ~n28005 ) | ( n28004 & 1'b0 ) | ( ~n28005 & 1'b0 ) ;
  assign n28018 = ( n27733 & n27770 ) | ( n27733 & n28006 ) | ( n27770 & n28006 ) ;
  assign n28017 = n27733 | n28006 ;
  assign n28019 = ( n28016 & ~n28018 ) | ( n28016 & n28017 ) | ( ~n28018 & n28017 ) ;
  assign n28023 = n27633 &  n27769 ;
  assign n28024 = n27768 &  n28023 ;
  assign n28012 = x77 | n27633 ;
  assign n28013 = x77 &  n27633 ;
  assign n28014 = ( n28012 & ~n28013 ) | ( n28012 & 1'b0 ) | ( ~n28013 & 1'b0 ) ;
  assign n28026 = ( n27732 & n27770 ) | ( n27732 & n28014 ) | ( n27770 & n28014 ) ;
  assign n28025 = n27732 | n28014 ;
  assign n28027 = ( n28024 & ~n28026 ) | ( n28024 & n28025 ) | ( ~n28026 & n28025 ) ;
  assign n28031 = n27641 &  n27769 ;
  assign n28032 = n27768 &  n28031 ;
  assign n28020 = x76 | n27641 ;
  assign n28021 = x76 &  n27641 ;
  assign n28022 = ( n28020 & ~n28021 ) | ( n28020 & 1'b0 ) | ( ~n28021 & 1'b0 ) ;
  assign n28034 = ( n27731 & n27770 ) | ( n27731 & n28022 ) | ( n27770 & n28022 ) ;
  assign n28033 = n27731 | n28022 ;
  assign n28035 = ( n28032 & ~n28034 ) | ( n28032 & n28033 ) | ( ~n28034 & n28033 ) ;
  assign n28039 = n27649 &  n27769 ;
  assign n28040 = n27768 &  n28039 ;
  assign n28028 = x75 | n27649 ;
  assign n28029 = x75 &  n27649 ;
  assign n28030 = ( n28028 & ~n28029 ) | ( n28028 & 1'b0 ) | ( ~n28029 & 1'b0 ) ;
  assign n28042 = ( n27730 & n27770 ) | ( n27730 & n28030 ) | ( n27770 & n28030 ) ;
  assign n28041 = n27730 | n28030 ;
  assign n28043 = ( n28040 & ~n28042 ) | ( n28040 & n28041 ) | ( ~n28042 & n28041 ) ;
  assign n28047 = n27657 &  n27769 ;
  assign n28048 = n27768 &  n28047 ;
  assign n28036 = x74 | n27657 ;
  assign n28037 = x74 &  n27657 ;
  assign n28038 = ( n28036 & ~n28037 ) | ( n28036 & 1'b0 ) | ( ~n28037 & 1'b0 ) ;
  assign n28050 = ( n27729 & n27770 ) | ( n27729 & n28038 ) | ( n27770 & n28038 ) ;
  assign n28049 = n27729 | n28038 ;
  assign n28051 = ( n28048 & ~n28050 ) | ( n28048 & n28049 ) | ( ~n28050 & n28049 ) ;
  assign n28055 = n27665 &  n27769 ;
  assign n28056 = n27768 &  n28055 ;
  assign n28044 = x73 | n27665 ;
  assign n28045 = x73 &  n27665 ;
  assign n28046 = ( n28044 & ~n28045 ) | ( n28044 & 1'b0 ) | ( ~n28045 & 1'b0 ) ;
  assign n28058 = ( n27728 & n27770 ) | ( n27728 & n28046 ) | ( n27770 & n28046 ) ;
  assign n28057 = n27728 | n28046 ;
  assign n28059 = ( n28056 & ~n28058 ) | ( n28056 & n28057 ) | ( ~n28058 & n28057 ) ;
  assign n28063 = n27673 &  n27769 ;
  assign n28064 = n27768 &  n28063 ;
  assign n28052 = x72 | n27673 ;
  assign n28053 = x72 &  n27673 ;
  assign n28054 = ( n28052 & ~n28053 ) | ( n28052 & 1'b0 ) | ( ~n28053 & 1'b0 ) ;
  assign n28066 = ( n27727 & n27770 ) | ( n27727 & n28054 ) | ( n27770 & n28054 ) ;
  assign n28065 = n27727 | n28054 ;
  assign n28067 = ( n28064 & ~n28066 ) | ( n28064 & n28065 ) | ( ~n28066 & n28065 ) ;
  assign n28071 = n27681 &  n27769 ;
  assign n28072 = n27768 &  n28071 ;
  assign n28060 = x71 | n27681 ;
  assign n28061 = x71 &  n27681 ;
  assign n28062 = ( n28060 & ~n28061 ) | ( n28060 & 1'b0 ) | ( ~n28061 & 1'b0 ) ;
  assign n28074 = ( n27726 & n27770 ) | ( n27726 & n28062 ) | ( n27770 & n28062 ) ;
  assign n28073 = n27726 | n28062 ;
  assign n28075 = ( n28072 & ~n28074 ) | ( n28072 & n28073 ) | ( ~n28074 & n28073 ) ;
  assign n28079 = n27689 &  n27769 ;
  assign n28080 = n27768 &  n28079 ;
  assign n28068 = x70 | n27689 ;
  assign n28069 = x70 &  n27689 ;
  assign n28070 = ( n28068 & ~n28069 ) | ( n28068 & 1'b0 ) | ( ~n28069 & 1'b0 ) ;
  assign n28082 = ( n27725 & n27770 ) | ( n27725 & n28070 ) | ( n27770 & n28070 ) ;
  assign n28081 = n27725 | n28070 ;
  assign n28083 = ( n28080 & ~n28082 ) | ( n28080 & n28081 ) | ( ~n28082 & n28081 ) ;
  assign n28087 = n27697 &  n27769 ;
  assign n28088 = n27768 &  n28087 ;
  assign n28076 = x69 | n27697 ;
  assign n28077 = x69 &  n27697 ;
  assign n28078 = ( n28076 & ~n28077 ) | ( n28076 & 1'b0 ) | ( ~n28077 & 1'b0 ) ;
  assign n28090 = ( n27724 & n27770 ) | ( n27724 & n28078 ) | ( n27770 & n28078 ) ;
  assign n28089 = n27724 | n28078 ;
  assign n28091 = ( n28088 & ~n28090 ) | ( n28088 & n28089 ) | ( ~n28090 & n28089 ) ;
  assign n28095 = n27705 &  n27769 ;
  assign n28096 = n27768 &  n28095 ;
  assign n28084 = x68 | n27705 ;
  assign n28085 = x68 &  n27705 ;
  assign n28086 = ( n28084 & ~n28085 ) | ( n28084 & 1'b0 ) | ( ~n28085 & 1'b0 ) ;
  assign n28098 = ( n27723 & n27770 ) | ( n27723 & n28086 ) | ( n27770 & n28086 ) ;
  assign n28097 = n27723 | n28086 ;
  assign n28099 = ( n28096 & ~n28098 ) | ( n28096 & n28097 ) | ( ~n28098 & n28097 ) ;
  assign n28103 = n27710 &  n27769 ;
  assign n28104 = n27768 &  n28103 ;
  assign n28092 = x67 | n27710 ;
  assign n28093 = x67 &  n27710 ;
  assign n28094 = ( n28092 & ~n28093 ) | ( n28092 & 1'b0 ) | ( ~n28093 & 1'b0 ) ;
  assign n28106 = ( n27722 & n27770 ) | ( n27722 & n28094 ) | ( n27770 & n28094 ) ;
  assign n28105 = n27722 | n28094 ;
  assign n28107 = ( n28104 & ~n28106 ) | ( n28104 & n28105 ) | ( ~n28106 & n28105 ) ;
  assign n28108 = n27716 &  n27769 ;
  assign n28109 = n27768 &  n28108 ;
  assign n28100 = x66 | n27716 ;
  assign n28101 = x66 &  n27716 ;
  assign n28102 = ( n28100 & ~n28101 ) | ( n28100 & 1'b0 ) | ( ~n28101 & 1'b0 ) ;
  assign n28110 = n27721 &  n28102 ;
  assign n28111 = ( n27721 & ~n27770 ) | ( n27721 & n28102 ) | ( ~n27770 & n28102 ) ;
  assign n28112 = ( n28109 & ~n28110 ) | ( n28109 & n28111 ) | ( ~n28110 & n28111 ) ;
  assign n28113 = ( x65 & ~n9279 ) | ( x65 & n27720 ) | ( ~n9279 & n27720 ) ;
  assign n28114 = ( n27721 & ~x65 ) | ( n27721 & n28113 ) | ( ~x65 & n28113 ) ;
  assign n28115 = ~n27770 & n28114 ;
  assign n28116 = n27720 &  n27769 ;
  assign n28117 = n27768 &  n28116 ;
  assign n28118 = n28115 | n28117 ;
  assign n28119 = ( x64 & ~n27770 ) | ( x64 & 1'b0 ) | ( ~n27770 & 1'b0 ) ;
  assign n28120 = ( x19 & ~n28119 ) | ( x19 & 1'b0 ) | ( ~n28119 & 1'b0 ) ;
  assign n28121 = ( n9279 & ~n27770 ) | ( n9279 & 1'b0 ) | ( ~n27770 & 1'b0 ) ;
  assign n28122 = n28120 | n28121 ;
  assign n28123 = ( x65 & ~n28122 ) | ( x65 & n9794 ) | ( ~n28122 & n9794 ) ;
  assign n28124 = ( x66 & ~n28118 ) | ( x66 & n28123 ) | ( ~n28118 & n28123 ) ;
  assign n28125 = ( x67 & ~n28112 ) | ( x67 & n28124 ) | ( ~n28112 & n28124 ) ;
  assign n28126 = ( x68 & ~n28107 ) | ( x68 & n28125 ) | ( ~n28107 & n28125 ) ;
  assign n28127 = ( x69 & ~n28099 ) | ( x69 & n28126 ) | ( ~n28099 & n28126 ) ;
  assign n28128 = ( x70 & ~n28091 ) | ( x70 & n28127 ) | ( ~n28091 & n28127 ) ;
  assign n28129 = ( x71 & ~n28083 ) | ( x71 & n28128 ) | ( ~n28083 & n28128 ) ;
  assign n28130 = ( x72 & ~n28075 ) | ( x72 & n28129 ) | ( ~n28075 & n28129 ) ;
  assign n28131 = ( x73 & ~n28067 ) | ( x73 & n28130 ) | ( ~n28067 & n28130 ) ;
  assign n28132 = ( x74 & ~n28059 ) | ( x74 & n28131 ) | ( ~n28059 & n28131 ) ;
  assign n28133 = ( x75 & ~n28051 ) | ( x75 & n28132 ) | ( ~n28051 & n28132 ) ;
  assign n28134 = ( x76 & ~n28043 ) | ( x76 & n28133 ) | ( ~n28043 & n28133 ) ;
  assign n28135 = ( x77 & ~n28035 ) | ( x77 & n28134 ) | ( ~n28035 & n28134 ) ;
  assign n28136 = ( x78 & ~n28027 ) | ( x78 & n28135 ) | ( ~n28027 & n28135 ) ;
  assign n28137 = ( x79 & ~n28019 ) | ( x79 & n28136 ) | ( ~n28019 & n28136 ) ;
  assign n28138 = ( x80 & ~n28011 ) | ( x80 & n28137 ) | ( ~n28011 & n28137 ) ;
  assign n28139 = ( x81 & ~n28003 ) | ( x81 & n28138 ) | ( ~n28003 & n28138 ) ;
  assign n28140 = ( x82 & ~n27995 ) | ( x82 & n28139 ) | ( ~n27995 & n28139 ) ;
  assign n28141 = ( x83 & ~n27987 ) | ( x83 & n28140 ) | ( ~n27987 & n28140 ) ;
  assign n28142 = ( x84 & ~n27979 ) | ( x84 & n28141 ) | ( ~n27979 & n28141 ) ;
  assign n28143 = ( x85 & ~n27971 ) | ( x85 & n28142 ) | ( ~n27971 & n28142 ) ;
  assign n28144 = ( x86 & ~n27963 ) | ( x86 & n28143 ) | ( ~n27963 & n28143 ) ;
  assign n28145 = ( x87 & ~n27955 ) | ( x87 & n28144 ) | ( ~n27955 & n28144 ) ;
  assign n28146 = ( x88 & ~n27947 ) | ( x88 & n28145 ) | ( ~n27947 & n28145 ) ;
  assign n28147 = ( x89 & ~n27939 ) | ( x89 & n28146 ) | ( ~n27939 & n28146 ) ;
  assign n28148 = ( x90 & ~n27931 ) | ( x90 & n28147 ) | ( ~n27931 & n28147 ) ;
  assign n28149 = ( x91 & ~n27923 ) | ( x91 & n28148 ) | ( ~n27923 & n28148 ) ;
  assign n28150 = ( x92 & ~n27915 ) | ( x92 & n28149 ) | ( ~n27915 & n28149 ) ;
  assign n28151 = ( x93 & ~n27907 ) | ( x93 & n28150 ) | ( ~n27907 & n28150 ) ;
  assign n28152 = ( x94 & ~n27899 ) | ( x94 & n28151 ) | ( ~n27899 & n28151 ) ;
  assign n28153 = ( x95 & ~n27891 ) | ( x95 & n28152 ) | ( ~n27891 & n28152 ) ;
  assign n28154 = ( x96 & ~n27883 ) | ( x96 & n28153 ) | ( ~n27883 & n28153 ) ;
  assign n28155 = ( x97 & ~n27875 ) | ( x97 & n28154 ) | ( ~n27875 & n28154 ) ;
  assign n28156 = ( x98 & ~n27867 ) | ( x98 & n28155 ) | ( ~n27867 & n28155 ) ;
  assign n28157 = ( x99 & ~n27859 ) | ( x99 & n28156 ) | ( ~n27859 & n28156 ) ;
  assign n28158 = ( x100 & ~n27851 ) | ( x100 & n28157 ) | ( ~n27851 & n28157 ) ;
  assign n28159 = ( x101 & ~n27843 ) | ( x101 & n28158 ) | ( ~n27843 & n28158 ) ;
  assign n28160 = ( x102 & ~n27835 ) | ( x102 & n28159 ) | ( ~n27835 & n28159 ) ;
  assign n28161 = ( x103 & ~n27827 ) | ( x103 & n28160 ) | ( ~n27827 & n28160 ) ;
  assign n28162 = ( x104 & ~n27819 ) | ( x104 & n28161 ) | ( ~n27819 & n28161 ) ;
  assign n28163 = ( x105 & ~n27811 ) | ( x105 & n28162 ) | ( ~n27811 & n28162 ) ;
  assign n28164 = ( x106 & ~n27803 ) | ( x106 & n28163 ) | ( ~n27803 & n28163 ) ;
  assign n28165 = ( x107 & ~n27795 ) | ( x107 & n28164 ) | ( ~n27795 & n28164 ) ;
  assign n28166 = ( x108 & ~n27787 ) | ( x108 & n28165 ) | ( ~n27787 & n28165 ) ;
  assign n28167 = ( x109 & ~n27779 ) | ( x109 & n28166 ) | ( ~n27779 & n28166 ) ;
  assign n28168 = n9841 | n28167 ;
  assign n28178 = n27787 &  n28168 ;
  assign n28170 = x108 | n27787 ;
  assign n28171 = x108 &  n27787 ;
  assign n28172 = ( n28170 & ~n28171 ) | ( n28170 & 1'b0 ) | ( ~n28171 & 1'b0 ) ;
  assign n28182 = ( n9841 & n28165 ) | ( n9841 & n28172 ) | ( n28165 & n28172 ) ;
  assign n28183 = ( n28165 & ~n28167 ) | ( n28165 & n28172 ) | ( ~n28167 & n28172 ) ;
  assign n28184 = ~n28182 & n28183 ;
  assign n28185 = n28178 | n28184 ;
  assign n28186 = n27795 &  n28168 ;
  assign n28179 = x107 | n27795 ;
  assign n28180 = x107 &  n27795 ;
  assign n28181 = ( n28179 & ~n28180 ) | ( n28179 & 1'b0 ) | ( ~n28180 & 1'b0 ) ;
  assign n28190 = ( n9841 & n28164 ) | ( n9841 & n28181 ) | ( n28164 & n28181 ) ;
  assign n28191 = ( n28164 & ~n28167 ) | ( n28164 & n28181 ) | ( ~n28167 & n28181 ) ;
  assign n28192 = ~n28190 & n28191 ;
  assign n28193 = n28186 | n28192 ;
  assign n28194 = n27803 &  n28168 ;
  assign n28187 = x106 | n27803 ;
  assign n28188 = x106 &  n27803 ;
  assign n28189 = ( n28187 & ~n28188 ) | ( n28187 & 1'b0 ) | ( ~n28188 & 1'b0 ) ;
  assign n28198 = ( n9841 & n28163 ) | ( n9841 & n28189 ) | ( n28163 & n28189 ) ;
  assign n28199 = ( n28163 & ~n28167 ) | ( n28163 & n28189 ) | ( ~n28167 & n28189 ) ;
  assign n28200 = ~n28198 & n28199 ;
  assign n28201 = n28194 | n28200 ;
  assign n28202 = n27811 &  n28168 ;
  assign n28195 = x105 | n27811 ;
  assign n28196 = x105 &  n27811 ;
  assign n28197 = ( n28195 & ~n28196 ) | ( n28195 & 1'b0 ) | ( ~n28196 & 1'b0 ) ;
  assign n28206 = ( n9841 & n28162 ) | ( n9841 & n28197 ) | ( n28162 & n28197 ) ;
  assign n28207 = ( n28162 & ~n28167 ) | ( n28162 & n28197 ) | ( ~n28167 & n28197 ) ;
  assign n28208 = ~n28206 & n28207 ;
  assign n28209 = n28202 | n28208 ;
  assign n28210 = n27819 &  n28168 ;
  assign n28203 = x104 | n27819 ;
  assign n28204 = x104 &  n27819 ;
  assign n28205 = ( n28203 & ~n28204 ) | ( n28203 & 1'b0 ) | ( ~n28204 & 1'b0 ) ;
  assign n28214 = ( n9841 & n28161 ) | ( n9841 & n28205 ) | ( n28161 & n28205 ) ;
  assign n28215 = ( n28161 & ~n28167 ) | ( n28161 & n28205 ) | ( ~n28167 & n28205 ) ;
  assign n28216 = ~n28214 & n28215 ;
  assign n28217 = n28210 | n28216 ;
  assign n28218 = n27827 &  n28168 ;
  assign n28211 = x103 | n27827 ;
  assign n28212 = x103 &  n27827 ;
  assign n28213 = ( n28211 & ~n28212 ) | ( n28211 & 1'b0 ) | ( ~n28212 & 1'b0 ) ;
  assign n28222 = ( n9841 & n28160 ) | ( n9841 & n28213 ) | ( n28160 & n28213 ) ;
  assign n28223 = ( n28160 & ~n28167 ) | ( n28160 & n28213 ) | ( ~n28167 & n28213 ) ;
  assign n28224 = ~n28222 & n28223 ;
  assign n28225 = n28218 | n28224 ;
  assign n28226 = n27835 &  n28168 ;
  assign n28219 = x102 | n27835 ;
  assign n28220 = x102 &  n27835 ;
  assign n28221 = ( n28219 & ~n28220 ) | ( n28219 & 1'b0 ) | ( ~n28220 & 1'b0 ) ;
  assign n28230 = ( n9841 & n28159 ) | ( n9841 & n28221 ) | ( n28159 & n28221 ) ;
  assign n28231 = ( n28159 & ~n28167 ) | ( n28159 & n28221 ) | ( ~n28167 & n28221 ) ;
  assign n28232 = ~n28230 & n28231 ;
  assign n28233 = n28226 | n28232 ;
  assign n28234 = n27843 &  n28168 ;
  assign n28227 = x101 | n27843 ;
  assign n28228 = x101 &  n27843 ;
  assign n28229 = ( n28227 & ~n28228 ) | ( n28227 & 1'b0 ) | ( ~n28228 & 1'b0 ) ;
  assign n28238 = ( n9841 & n28158 ) | ( n9841 & n28229 ) | ( n28158 & n28229 ) ;
  assign n28239 = ( n28158 & ~n28167 ) | ( n28158 & n28229 ) | ( ~n28167 & n28229 ) ;
  assign n28240 = ~n28238 & n28239 ;
  assign n28241 = n28234 | n28240 ;
  assign n28242 = n27851 &  n28168 ;
  assign n28235 = x100 | n27851 ;
  assign n28236 = x100 &  n27851 ;
  assign n28237 = ( n28235 & ~n28236 ) | ( n28235 & 1'b0 ) | ( ~n28236 & 1'b0 ) ;
  assign n28246 = ( n9841 & n28157 ) | ( n9841 & n28237 ) | ( n28157 & n28237 ) ;
  assign n28247 = ( n28157 & ~n28167 ) | ( n28157 & n28237 ) | ( ~n28167 & n28237 ) ;
  assign n28248 = ~n28246 & n28247 ;
  assign n28249 = n28242 | n28248 ;
  assign n28250 = n27859 &  n28168 ;
  assign n28243 = x99 | n27859 ;
  assign n28244 = x99 &  n27859 ;
  assign n28245 = ( n28243 & ~n28244 ) | ( n28243 & 1'b0 ) | ( ~n28244 & 1'b0 ) ;
  assign n28254 = ( n9841 & n28156 ) | ( n9841 & n28245 ) | ( n28156 & n28245 ) ;
  assign n28255 = ( n28156 & ~n28167 ) | ( n28156 & n28245 ) | ( ~n28167 & n28245 ) ;
  assign n28256 = ~n28254 & n28255 ;
  assign n28257 = n28250 | n28256 ;
  assign n28258 = n27867 &  n28168 ;
  assign n28251 = x98 | n27867 ;
  assign n28252 = x98 &  n27867 ;
  assign n28253 = ( n28251 & ~n28252 ) | ( n28251 & 1'b0 ) | ( ~n28252 & 1'b0 ) ;
  assign n28262 = ( n9841 & n28155 ) | ( n9841 & n28253 ) | ( n28155 & n28253 ) ;
  assign n28263 = ( n28155 & ~n28167 ) | ( n28155 & n28253 ) | ( ~n28167 & n28253 ) ;
  assign n28264 = ~n28262 & n28263 ;
  assign n28265 = n28258 | n28264 ;
  assign n28266 = n27875 &  n28168 ;
  assign n28259 = x97 | n27875 ;
  assign n28260 = x97 &  n27875 ;
  assign n28261 = ( n28259 & ~n28260 ) | ( n28259 & 1'b0 ) | ( ~n28260 & 1'b0 ) ;
  assign n28270 = ( n9841 & n28154 ) | ( n9841 & n28261 ) | ( n28154 & n28261 ) ;
  assign n28271 = ( n28154 & ~n28167 ) | ( n28154 & n28261 ) | ( ~n28167 & n28261 ) ;
  assign n28272 = ~n28270 & n28271 ;
  assign n28273 = n28266 | n28272 ;
  assign n28274 = n27883 &  n28168 ;
  assign n28267 = x96 | n27883 ;
  assign n28268 = x96 &  n27883 ;
  assign n28269 = ( n28267 & ~n28268 ) | ( n28267 & 1'b0 ) | ( ~n28268 & 1'b0 ) ;
  assign n28278 = ( n9841 & n28153 ) | ( n9841 & n28269 ) | ( n28153 & n28269 ) ;
  assign n28279 = ( n28153 & ~n28167 ) | ( n28153 & n28269 ) | ( ~n28167 & n28269 ) ;
  assign n28280 = ~n28278 & n28279 ;
  assign n28281 = n28274 | n28280 ;
  assign n28282 = n27891 &  n28168 ;
  assign n28275 = x95 | n27891 ;
  assign n28276 = x95 &  n27891 ;
  assign n28277 = ( n28275 & ~n28276 ) | ( n28275 & 1'b0 ) | ( ~n28276 & 1'b0 ) ;
  assign n28286 = ( n9841 & n28152 ) | ( n9841 & n28277 ) | ( n28152 & n28277 ) ;
  assign n28287 = ( n28152 & ~n28167 ) | ( n28152 & n28277 ) | ( ~n28167 & n28277 ) ;
  assign n28288 = ~n28286 & n28287 ;
  assign n28289 = n28282 | n28288 ;
  assign n28290 = n27899 &  n28168 ;
  assign n28283 = x94 | n27899 ;
  assign n28284 = x94 &  n27899 ;
  assign n28285 = ( n28283 & ~n28284 ) | ( n28283 & 1'b0 ) | ( ~n28284 & 1'b0 ) ;
  assign n28294 = ( n9841 & n28151 ) | ( n9841 & n28285 ) | ( n28151 & n28285 ) ;
  assign n28295 = ( n28151 & ~n28167 ) | ( n28151 & n28285 ) | ( ~n28167 & n28285 ) ;
  assign n28296 = ~n28294 & n28295 ;
  assign n28297 = n28290 | n28296 ;
  assign n28298 = n27907 &  n28168 ;
  assign n28291 = x93 | n27907 ;
  assign n28292 = x93 &  n27907 ;
  assign n28293 = ( n28291 & ~n28292 ) | ( n28291 & 1'b0 ) | ( ~n28292 & 1'b0 ) ;
  assign n28302 = ( n9841 & n28150 ) | ( n9841 & n28293 ) | ( n28150 & n28293 ) ;
  assign n28303 = ( n28150 & ~n28167 ) | ( n28150 & n28293 ) | ( ~n28167 & n28293 ) ;
  assign n28304 = ~n28302 & n28303 ;
  assign n28305 = n28298 | n28304 ;
  assign n28306 = n27915 &  n28168 ;
  assign n28299 = x92 | n27915 ;
  assign n28300 = x92 &  n27915 ;
  assign n28301 = ( n28299 & ~n28300 ) | ( n28299 & 1'b0 ) | ( ~n28300 & 1'b0 ) ;
  assign n28310 = ( n9841 & n28149 ) | ( n9841 & n28301 ) | ( n28149 & n28301 ) ;
  assign n28311 = ( n28149 & ~n28167 ) | ( n28149 & n28301 ) | ( ~n28167 & n28301 ) ;
  assign n28312 = ~n28310 & n28311 ;
  assign n28313 = n28306 | n28312 ;
  assign n28314 = n27923 &  n28168 ;
  assign n28307 = x91 | n27923 ;
  assign n28308 = x91 &  n27923 ;
  assign n28309 = ( n28307 & ~n28308 ) | ( n28307 & 1'b0 ) | ( ~n28308 & 1'b0 ) ;
  assign n28318 = ( n9841 & n28148 ) | ( n9841 & n28309 ) | ( n28148 & n28309 ) ;
  assign n28319 = ( n28148 & ~n28167 ) | ( n28148 & n28309 ) | ( ~n28167 & n28309 ) ;
  assign n28320 = ~n28318 & n28319 ;
  assign n28321 = n28314 | n28320 ;
  assign n28322 = n27931 &  n28168 ;
  assign n28315 = x90 | n27931 ;
  assign n28316 = x90 &  n27931 ;
  assign n28317 = ( n28315 & ~n28316 ) | ( n28315 & 1'b0 ) | ( ~n28316 & 1'b0 ) ;
  assign n28326 = ( n9841 & n28147 ) | ( n9841 & n28317 ) | ( n28147 & n28317 ) ;
  assign n28327 = ( n28147 & ~n28167 ) | ( n28147 & n28317 ) | ( ~n28167 & n28317 ) ;
  assign n28328 = ~n28326 & n28327 ;
  assign n28329 = n28322 | n28328 ;
  assign n28330 = n27939 &  n28168 ;
  assign n28323 = x89 | n27939 ;
  assign n28324 = x89 &  n27939 ;
  assign n28325 = ( n28323 & ~n28324 ) | ( n28323 & 1'b0 ) | ( ~n28324 & 1'b0 ) ;
  assign n28334 = ( n9841 & n28146 ) | ( n9841 & n28325 ) | ( n28146 & n28325 ) ;
  assign n28335 = ( n28146 & ~n28167 ) | ( n28146 & n28325 ) | ( ~n28167 & n28325 ) ;
  assign n28336 = ~n28334 & n28335 ;
  assign n28337 = n28330 | n28336 ;
  assign n28338 = n27947 &  n28168 ;
  assign n28331 = x88 | n27947 ;
  assign n28332 = x88 &  n27947 ;
  assign n28333 = ( n28331 & ~n28332 ) | ( n28331 & 1'b0 ) | ( ~n28332 & 1'b0 ) ;
  assign n28342 = ( n9841 & n28145 ) | ( n9841 & n28333 ) | ( n28145 & n28333 ) ;
  assign n28343 = ( n28145 & ~n28167 ) | ( n28145 & n28333 ) | ( ~n28167 & n28333 ) ;
  assign n28344 = ~n28342 & n28343 ;
  assign n28345 = n28338 | n28344 ;
  assign n28346 = n27955 &  n28168 ;
  assign n28339 = x87 | n27955 ;
  assign n28340 = x87 &  n27955 ;
  assign n28341 = ( n28339 & ~n28340 ) | ( n28339 & 1'b0 ) | ( ~n28340 & 1'b0 ) ;
  assign n28350 = ( n9841 & n28144 ) | ( n9841 & n28341 ) | ( n28144 & n28341 ) ;
  assign n28351 = ( n28144 & ~n28167 ) | ( n28144 & n28341 ) | ( ~n28167 & n28341 ) ;
  assign n28352 = ~n28350 & n28351 ;
  assign n28353 = n28346 | n28352 ;
  assign n28354 = n27963 &  n28168 ;
  assign n28347 = x86 | n27963 ;
  assign n28348 = x86 &  n27963 ;
  assign n28349 = ( n28347 & ~n28348 ) | ( n28347 & 1'b0 ) | ( ~n28348 & 1'b0 ) ;
  assign n28358 = ( n9841 & n28143 ) | ( n9841 & n28349 ) | ( n28143 & n28349 ) ;
  assign n28359 = ( n28143 & ~n28167 ) | ( n28143 & n28349 ) | ( ~n28167 & n28349 ) ;
  assign n28360 = ~n28358 & n28359 ;
  assign n28361 = n28354 | n28360 ;
  assign n28362 = n27971 &  n28168 ;
  assign n28355 = x85 | n27971 ;
  assign n28356 = x85 &  n27971 ;
  assign n28357 = ( n28355 & ~n28356 ) | ( n28355 & 1'b0 ) | ( ~n28356 & 1'b0 ) ;
  assign n28366 = ( n9841 & n28142 ) | ( n9841 & n28357 ) | ( n28142 & n28357 ) ;
  assign n28367 = ( n28142 & ~n28167 ) | ( n28142 & n28357 ) | ( ~n28167 & n28357 ) ;
  assign n28368 = ~n28366 & n28367 ;
  assign n28369 = n28362 | n28368 ;
  assign n28370 = n27979 &  n28168 ;
  assign n28363 = x84 | n27979 ;
  assign n28364 = x84 &  n27979 ;
  assign n28365 = ( n28363 & ~n28364 ) | ( n28363 & 1'b0 ) | ( ~n28364 & 1'b0 ) ;
  assign n28374 = ( n9841 & n28141 ) | ( n9841 & n28365 ) | ( n28141 & n28365 ) ;
  assign n28375 = ( n28141 & ~n28167 ) | ( n28141 & n28365 ) | ( ~n28167 & n28365 ) ;
  assign n28376 = ~n28374 & n28375 ;
  assign n28377 = n28370 | n28376 ;
  assign n28378 = n27987 &  n28168 ;
  assign n28371 = x83 | n27987 ;
  assign n28372 = x83 &  n27987 ;
  assign n28373 = ( n28371 & ~n28372 ) | ( n28371 & 1'b0 ) | ( ~n28372 & 1'b0 ) ;
  assign n28382 = ( n9841 & n28140 ) | ( n9841 & n28373 ) | ( n28140 & n28373 ) ;
  assign n28383 = ( n28140 & ~n28167 ) | ( n28140 & n28373 ) | ( ~n28167 & n28373 ) ;
  assign n28384 = ~n28382 & n28383 ;
  assign n28385 = n28378 | n28384 ;
  assign n28386 = n27995 &  n28168 ;
  assign n28379 = x82 | n27995 ;
  assign n28380 = x82 &  n27995 ;
  assign n28381 = ( n28379 & ~n28380 ) | ( n28379 & 1'b0 ) | ( ~n28380 & 1'b0 ) ;
  assign n28390 = ( n9841 & n28139 ) | ( n9841 & n28381 ) | ( n28139 & n28381 ) ;
  assign n28391 = ( n28139 & ~n28167 ) | ( n28139 & n28381 ) | ( ~n28167 & n28381 ) ;
  assign n28392 = ~n28390 & n28391 ;
  assign n28393 = n28386 | n28392 ;
  assign n28394 = n28003 &  n28168 ;
  assign n28387 = x81 | n28003 ;
  assign n28388 = x81 &  n28003 ;
  assign n28389 = ( n28387 & ~n28388 ) | ( n28387 & 1'b0 ) | ( ~n28388 & 1'b0 ) ;
  assign n28398 = ( n9841 & n28138 ) | ( n9841 & n28389 ) | ( n28138 & n28389 ) ;
  assign n28399 = ( n28138 & ~n28167 ) | ( n28138 & n28389 ) | ( ~n28167 & n28389 ) ;
  assign n28400 = ~n28398 & n28399 ;
  assign n28401 = n28394 | n28400 ;
  assign n28402 = n28011 &  n28168 ;
  assign n28395 = x80 | n28011 ;
  assign n28396 = x80 &  n28011 ;
  assign n28397 = ( n28395 & ~n28396 ) | ( n28395 & 1'b0 ) | ( ~n28396 & 1'b0 ) ;
  assign n28406 = ( n9841 & n28137 ) | ( n9841 & n28397 ) | ( n28137 & n28397 ) ;
  assign n28407 = ( n28137 & ~n28167 ) | ( n28137 & n28397 ) | ( ~n28167 & n28397 ) ;
  assign n28408 = ~n28406 & n28407 ;
  assign n28409 = n28402 | n28408 ;
  assign n28410 = n28019 &  n28168 ;
  assign n28403 = x79 | n28019 ;
  assign n28404 = x79 &  n28019 ;
  assign n28405 = ( n28403 & ~n28404 ) | ( n28403 & 1'b0 ) | ( ~n28404 & 1'b0 ) ;
  assign n28414 = ( n9841 & n28136 ) | ( n9841 & n28405 ) | ( n28136 & n28405 ) ;
  assign n28415 = ( n28136 & ~n28167 ) | ( n28136 & n28405 ) | ( ~n28167 & n28405 ) ;
  assign n28416 = ~n28414 & n28415 ;
  assign n28417 = n28410 | n28416 ;
  assign n28418 = n28027 &  n28168 ;
  assign n28411 = x78 | n28027 ;
  assign n28412 = x78 &  n28027 ;
  assign n28413 = ( n28411 & ~n28412 ) | ( n28411 & 1'b0 ) | ( ~n28412 & 1'b0 ) ;
  assign n28422 = ( n9841 & n28135 ) | ( n9841 & n28413 ) | ( n28135 & n28413 ) ;
  assign n28423 = ( n28135 & ~n28167 ) | ( n28135 & n28413 ) | ( ~n28167 & n28413 ) ;
  assign n28424 = ~n28422 & n28423 ;
  assign n28425 = n28418 | n28424 ;
  assign n28426 = n28035 &  n28168 ;
  assign n28419 = x77 | n28035 ;
  assign n28420 = x77 &  n28035 ;
  assign n28421 = ( n28419 & ~n28420 ) | ( n28419 & 1'b0 ) | ( ~n28420 & 1'b0 ) ;
  assign n28430 = ( n9841 & n28134 ) | ( n9841 & n28421 ) | ( n28134 & n28421 ) ;
  assign n28431 = ( n28134 & ~n28167 ) | ( n28134 & n28421 ) | ( ~n28167 & n28421 ) ;
  assign n28432 = ~n28430 & n28431 ;
  assign n28433 = n28426 | n28432 ;
  assign n28434 = n28043 &  n28168 ;
  assign n28427 = x76 | n28043 ;
  assign n28428 = x76 &  n28043 ;
  assign n28429 = ( n28427 & ~n28428 ) | ( n28427 & 1'b0 ) | ( ~n28428 & 1'b0 ) ;
  assign n28438 = ( n9841 & n28133 ) | ( n9841 & n28429 ) | ( n28133 & n28429 ) ;
  assign n28439 = ( n28133 & ~n28167 ) | ( n28133 & n28429 ) | ( ~n28167 & n28429 ) ;
  assign n28440 = ~n28438 & n28439 ;
  assign n28441 = n28434 | n28440 ;
  assign n28442 = n28051 &  n28168 ;
  assign n28435 = x75 | n28051 ;
  assign n28436 = x75 &  n28051 ;
  assign n28437 = ( n28435 & ~n28436 ) | ( n28435 & 1'b0 ) | ( ~n28436 & 1'b0 ) ;
  assign n28446 = ( n9841 & n28132 ) | ( n9841 & n28437 ) | ( n28132 & n28437 ) ;
  assign n28447 = ( n28132 & ~n28167 ) | ( n28132 & n28437 ) | ( ~n28167 & n28437 ) ;
  assign n28448 = ~n28446 & n28447 ;
  assign n28449 = n28442 | n28448 ;
  assign n28450 = n28059 &  n28168 ;
  assign n28443 = x74 | n28059 ;
  assign n28444 = x74 &  n28059 ;
  assign n28445 = ( n28443 & ~n28444 ) | ( n28443 & 1'b0 ) | ( ~n28444 & 1'b0 ) ;
  assign n28454 = ( n9841 & n28131 ) | ( n9841 & n28445 ) | ( n28131 & n28445 ) ;
  assign n28455 = ( n28131 & ~n28167 ) | ( n28131 & n28445 ) | ( ~n28167 & n28445 ) ;
  assign n28456 = ~n28454 & n28455 ;
  assign n28457 = n28450 | n28456 ;
  assign n28458 = n28067 &  n28168 ;
  assign n28451 = x73 | n28067 ;
  assign n28452 = x73 &  n28067 ;
  assign n28453 = ( n28451 & ~n28452 ) | ( n28451 & 1'b0 ) | ( ~n28452 & 1'b0 ) ;
  assign n28462 = ( n9841 & n28130 ) | ( n9841 & n28453 ) | ( n28130 & n28453 ) ;
  assign n28463 = ( n28130 & ~n28167 ) | ( n28130 & n28453 ) | ( ~n28167 & n28453 ) ;
  assign n28464 = ~n28462 & n28463 ;
  assign n28465 = n28458 | n28464 ;
  assign n28466 = n28075 &  n28168 ;
  assign n28459 = x72 | n28075 ;
  assign n28460 = x72 &  n28075 ;
  assign n28461 = ( n28459 & ~n28460 ) | ( n28459 & 1'b0 ) | ( ~n28460 & 1'b0 ) ;
  assign n28470 = ( n9841 & n28129 ) | ( n9841 & n28461 ) | ( n28129 & n28461 ) ;
  assign n28471 = ( n28129 & ~n28167 ) | ( n28129 & n28461 ) | ( ~n28167 & n28461 ) ;
  assign n28472 = ~n28470 & n28471 ;
  assign n28473 = n28466 | n28472 ;
  assign n28474 = n28083 &  n28168 ;
  assign n28467 = x71 | n28083 ;
  assign n28468 = x71 &  n28083 ;
  assign n28469 = ( n28467 & ~n28468 ) | ( n28467 & 1'b0 ) | ( ~n28468 & 1'b0 ) ;
  assign n28478 = ( n9841 & n28128 ) | ( n9841 & n28469 ) | ( n28128 & n28469 ) ;
  assign n28479 = ( n28128 & ~n28167 ) | ( n28128 & n28469 ) | ( ~n28167 & n28469 ) ;
  assign n28480 = ~n28478 & n28479 ;
  assign n28481 = n28474 | n28480 ;
  assign n28482 = n28091 &  n28168 ;
  assign n28475 = x70 | n28091 ;
  assign n28476 = x70 &  n28091 ;
  assign n28477 = ( n28475 & ~n28476 ) | ( n28475 & 1'b0 ) | ( ~n28476 & 1'b0 ) ;
  assign n28486 = ( n9841 & n28127 ) | ( n9841 & n28477 ) | ( n28127 & n28477 ) ;
  assign n28487 = ( n28127 & ~n28167 ) | ( n28127 & n28477 ) | ( ~n28167 & n28477 ) ;
  assign n28488 = ~n28486 & n28487 ;
  assign n28489 = n28482 | n28488 ;
  assign n28490 = n28099 &  n28168 ;
  assign n28483 = x69 | n28099 ;
  assign n28484 = x69 &  n28099 ;
  assign n28485 = ( n28483 & ~n28484 ) | ( n28483 & 1'b0 ) | ( ~n28484 & 1'b0 ) ;
  assign n28494 = ( n9841 & n28126 ) | ( n9841 & n28485 ) | ( n28126 & n28485 ) ;
  assign n28495 = ( n28126 & ~n28167 ) | ( n28126 & n28485 ) | ( ~n28167 & n28485 ) ;
  assign n28496 = ~n28494 & n28495 ;
  assign n28497 = n28490 | n28496 ;
  assign n28498 = n28107 &  n28168 ;
  assign n28491 = x68 | n28107 ;
  assign n28492 = x68 &  n28107 ;
  assign n28493 = ( n28491 & ~n28492 ) | ( n28491 & 1'b0 ) | ( ~n28492 & 1'b0 ) ;
  assign n28502 = ( n9841 & n28125 ) | ( n9841 & n28493 ) | ( n28125 & n28493 ) ;
  assign n28503 = ( n28125 & ~n28167 ) | ( n28125 & n28493 ) | ( ~n28167 & n28493 ) ;
  assign n28504 = ~n28502 & n28503 ;
  assign n28505 = n28498 | n28504 ;
  assign n28506 = n28112 &  n28168 ;
  assign n28499 = x67 | n28112 ;
  assign n28500 = x67 &  n28112 ;
  assign n28501 = ( n28499 & ~n28500 ) | ( n28499 & 1'b0 ) | ( ~n28500 & 1'b0 ) ;
  assign n28510 = ( n9841 & n28124 ) | ( n9841 & n28501 ) | ( n28124 & n28501 ) ;
  assign n28511 = ( n28124 & ~n28167 ) | ( n28124 & n28501 ) | ( ~n28167 & n28501 ) ;
  assign n28512 = ~n28510 & n28511 ;
  assign n28513 = n28506 | n28512 ;
  assign n28514 = n28118 &  n28168 ;
  assign n28507 = x66 | n28118 ;
  assign n28508 = x66 &  n28118 ;
  assign n28509 = ( n28507 & ~n28508 ) | ( n28507 & 1'b0 ) | ( ~n28508 & 1'b0 ) ;
  assign n28515 = ( n9841 & n28123 ) | ( n9841 & n28509 ) | ( n28123 & n28509 ) ;
  assign n28516 = ( n28123 & ~n28167 ) | ( n28123 & n28509 ) | ( ~n28167 & n28509 ) ;
  assign n28517 = ~n28515 & n28516 ;
  assign n28518 = n28514 | n28517 ;
  assign n28519 = n28122 &  n28168 ;
  assign n28520 = ( x65 & ~x19 ) | ( x65 & n28119 ) | ( ~x19 & n28119 ) ;
  assign n28521 = ( x19 & ~n28119 ) | ( x19 & x65 ) | ( ~n28119 & x65 ) ;
  assign n28522 = ( n28520 & ~x65 ) | ( n28520 & n28521 ) | ( ~x65 & n28521 ) ;
  assign n28523 = ( n9794 & ~n9841 ) | ( n9794 & n28522 ) | ( ~n9841 & n28522 ) ;
  assign n28524 = ( n9794 & n28167 ) | ( n9794 & n28522 ) | ( n28167 & n28522 ) ;
  assign n28525 = ( n28523 & ~n28524 ) | ( n28523 & 1'b0 ) | ( ~n28524 & 1'b0 ) ;
  assign n28526 = n28519 | n28525 ;
  assign n28527 = ( n10104 & ~n28167 ) | ( n10104 & 1'b0 ) | ( ~n28167 & 1'b0 ) ;
  assign n28528 = ( x18 & ~n28527 ) | ( x18 & 1'b0 ) | ( ~n28527 & 1'b0 ) ;
  assign n28529 = ( n10109 & ~n28167 ) | ( n10109 & 1'b0 ) | ( ~n28167 & 1'b0 ) ;
  assign n28530 = n28528 | n28529 ;
  assign n28531 = ( x65 & ~n28530 ) | ( x65 & n10112 ) | ( ~n28530 & n10112 ) ;
  assign n28532 = ( x66 & ~n28526 ) | ( x66 & n28531 ) | ( ~n28526 & n28531 ) ;
  assign n28533 = ( x67 & ~n28518 ) | ( x67 & n28532 ) | ( ~n28518 & n28532 ) ;
  assign n28534 = ( x68 & ~n28513 ) | ( x68 & n28533 ) | ( ~n28513 & n28533 ) ;
  assign n28535 = ( x69 & ~n28505 ) | ( x69 & n28534 ) | ( ~n28505 & n28534 ) ;
  assign n28536 = ( x70 & ~n28497 ) | ( x70 & n28535 ) | ( ~n28497 & n28535 ) ;
  assign n28537 = ( x71 & ~n28489 ) | ( x71 & n28536 ) | ( ~n28489 & n28536 ) ;
  assign n28538 = ( x72 & ~n28481 ) | ( x72 & n28537 ) | ( ~n28481 & n28537 ) ;
  assign n28539 = ( x73 & ~n28473 ) | ( x73 & n28538 ) | ( ~n28473 & n28538 ) ;
  assign n28540 = ( x74 & ~n28465 ) | ( x74 & n28539 ) | ( ~n28465 & n28539 ) ;
  assign n28541 = ( x75 & ~n28457 ) | ( x75 & n28540 ) | ( ~n28457 & n28540 ) ;
  assign n28542 = ( x76 & ~n28449 ) | ( x76 & n28541 ) | ( ~n28449 & n28541 ) ;
  assign n28543 = ( x77 & ~n28441 ) | ( x77 & n28542 ) | ( ~n28441 & n28542 ) ;
  assign n28544 = ( x78 & ~n28433 ) | ( x78 & n28543 ) | ( ~n28433 & n28543 ) ;
  assign n28545 = ( x79 & ~n28425 ) | ( x79 & n28544 ) | ( ~n28425 & n28544 ) ;
  assign n28546 = ( x80 & ~n28417 ) | ( x80 & n28545 ) | ( ~n28417 & n28545 ) ;
  assign n28547 = ( x81 & ~n28409 ) | ( x81 & n28546 ) | ( ~n28409 & n28546 ) ;
  assign n28548 = ( x82 & ~n28401 ) | ( x82 & n28547 ) | ( ~n28401 & n28547 ) ;
  assign n28549 = ( x83 & ~n28393 ) | ( x83 & n28548 ) | ( ~n28393 & n28548 ) ;
  assign n28550 = ( x84 & ~n28385 ) | ( x84 & n28549 ) | ( ~n28385 & n28549 ) ;
  assign n28551 = ( x85 & ~n28377 ) | ( x85 & n28550 ) | ( ~n28377 & n28550 ) ;
  assign n28552 = ( x86 & ~n28369 ) | ( x86 & n28551 ) | ( ~n28369 & n28551 ) ;
  assign n28553 = ( x87 & ~n28361 ) | ( x87 & n28552 ) | ( ~n28361 & n28552 ) ;
  assign n28554 = ( x88 & ~n28353 ) | ( x88 & n28553 ) | ( ~n28353 & n28553 ) ;
  assign n28555 = ( x89 & ~n28345 ) | ( x89 & n28554 ) | ( ~n28345 & n28554 ) ;
  assign n28556 = ( x90 & ~n28337 ) | ( x90 & n28555 ) | ( ~n28337 & n28555 ) ;
  assign n28557 = ( x91 & ~n28329 ) | ( x91 & n28556 ) | ( ~n28329 & n28556 ) ;
  assign n28558 = ( x92 & ~n28321 ) | ( x92 & n28557 ) | ( ~n28321 & n28557 ) ;
  assign n28559 = ( x93 & ~n28313 ) | ( x93 & n28558 ) | ( ~n28313 & n28558 ) ;
  assign n28560 = ( x94 & ~n28305 ) | ( x94 & n28559 ) | ( ~n28305 & n28559 ) ;
  assign n28561 = ( x95 & ~n28297 ) | ( x95 & n28560 ) | ( ~n28297 & n28560 ) ;
  assign n28562 = ( x96 & ~n28289 ) | ( x96 & n28561 ) | ( ~n28289 & n28561 ) ;
  assign n28563 = ( x97 & ~n28281 ) | ( x97 & n28562 ) | ( ~n28281 & n28562 ) ;
  assign n28564 = ( x98 & ~n28273 ) | ( x98 & n28563 ) | ( ~n28273 & n28563 ) ;
  assign n28565 = ( x99 & ~n28265 ) | ( x99 & n28564 ) | ( ~n28265 & n28564 ) ;
  assign n28566 = ( x100 & ~n28257 ) | ( x100 & n28565 ) | ( ~n28257 & n28565 ) ;
  assign n28567 = ( x101 & ~n28249 ) | ( x101 & n28566 ) | ( ~n28249 & n28566 ) ;
  assign n28568 = ( x102 & ~n28241 ) | ( x102 & n28567 ) | ( ~n28241 & n28567 ) ;
  assign n28569 = ( x103 & ~n28233 ) | ( x103 & n28568 ) | ( ~n28233 & n28568 ) ;
  assign n28570 = ( x104 & ~n28225 ) | ( x104 & n28569 ) | ( ~n28225 & n28569 ) ;
  assign n28571 = ( x105 & ~n28217 ) | ( x105 & n28570 ) | ( ~n28217 & n28570 ) ;
  assign n28572 = ( x106 & ~n28209 ) | ( x106 & n28571 ) | ( ~n28209 & n28571 ) ;
  assign n28573 = ( x107 & ~n28201 ) | ( x107 & n28572 ) | ( ~n28201 & n28572 ) ;
  assign n28574 = ( x108 & ~n28193 ) | ( x108 & n28573 ) | ( ~n28193 & n28573 ) ;
  assign n28575 = ( x109 & ~n28185 ) | ( x109 & n28574 ) | ( ~n28185 & n28574 ) ;
  assign n28169 = n27779 &  n28168 ;
  assign n28173 = ( n9841 & n27779 ) | ( n9841 & n28166 ) | ( n27779 & n28166 ) ;
  assign n28174 = ( x109 & ~n28173 ) | ( x109 & n27779 ) | ( ~n28173 & n27779 ) ;
  assign n28175 = ~x109 & n28174 ;
  assign n28176 = n28169 | n28175 ;
  assign n28177 = ~x110 & n28176 ;
  assign n28576 = ( x110 & ~n28169 ) | ( x110 & 1'b0 ) | ( ~n28169 & 1'b0 ) ;
  assign n28577 = ~n28175 & n28576 ;
  assign n28586 = n28177 | n28577 ;
  assign n28587 = ( n28575 & ~n28586 ) | ( n28575 & 1'b0 ) | ( ~n28586 & 1'b0 ) ;
  assign n28578 = ( n28575 & ~n28177 ) | ( n28575 & n28577 ) | ( ~n28177 & n28577 ) ;
  assign n28579 = ( n28177 & ~n10264 ) | ( n28177 & n28578 ) | ( ~n10264 & n28578 ) ;
  assign n28580 = n10264 | n28579 ;
  assign n28581 = ~n28176 |  n9841 ;
  assign n28582 = n28580 &  n28581 ;
  assign n28588 = ~n28575 & n28586 ;
  assign n28589 = ( n28587 & ~n28582 ) | ( n28587 & n28588 ) | ( ~n28582 & n28588 ) ;
  assign n28590 = n9841 &  n27779 ;
  assign n28591 = n28580 &  n28590 ;
  assign n28592 = n28589 | n28591 ;
  assign n28593 = ~x111 & n28592 ;
  assign n28597 = n28185 &  n28581 ;
  assign n28598 = n28580 &  n28597 ;
  assign n28583 = x109 | n28185 ;
  assign n28584 = x109 &  n28185 ;
  assign n28585 = ( n28583 & ~n28584 ) | ( n28583 & 1'b0 ) | ( ~n28584 & 1'b0 ) ;
  assign n28600 = ( n28574 & n28582 ) | ( n28574 & n28585 ) | ( n28582 & n28585 ) ;
  assign n28599 = n28574 | n28585 ;
  assign n28601 = ( n28598 & ~n28600 ) | ( n28598 & n28599 ) | ( ~n28600 & n28599 ) ;
  assign n28605 = n28193 &  n28581 ;
  assign n28606 = n28580 &  n28605 ;
  assign n28594 = x108 | n28193 ;
  assign n28595 = x108 &  n28193 ;
  assign n28596 = ( n28594 & ~n28595 ) | ( n28594 & 1'b0 ) | ( ~n28595 & 1'b0 ) ;
  assign n28608 = ( n28573 & n28582 ) | ( n28573 & n28596 ) | ( n28582 & n28596 ) ;
  assign n28607 = n28573 | n28596 ;
  assign n28609 = ( n28606 & ~n28608 ) | ( n28606 & n28607 ) | ( ~n28608 & n28607 ) ;
  assign n28613 = n28201 &  n28581 ;
  assign n28614 = n28580 &  n28613 ;
  assign n28602 = x107 | n28201 ;
  assign n28603 = x107 &  n28201 ;
  assign n28604 = ( n28602 & ~n28603 ) | ( n28602 & 1'b0 ) | ( ~n28603 & 1'b0 ) ;
  assign n28616 = ( n28572 & n28582 ) | ( n28572 & n28604 ) | ( n28582 & n28604 ) ;
  assign n28615 = n28572 | n28604 ;
  assign n28617 = ( n28614 & ~n28616 ) | ( n28614 & n28615 ) | ( ~n28616 & n28615 ) ;
  assign n28621 = n28209 &  n28581 ;
  assign n28622 = n28580 &  n28621 ;
  assign n28610 = x106 | n28209 ;
  assign n28611 = x106 &  n28209 ;
  assign n28612 = ( n28610 & ~n28611 ) | ( n28610 & 1'b0 ) | ( ~n28611 & 1'b0 ) ;
  assign n28624 = ( n28571 & n28582 ) | ( n28571 & n28612 ) | ( n28582 & n28612 ) ;
  assign n28623 = n28571 | n28612 ;
  assign n28625 = ( n28622 & ~n28624 ) | ( n28622 & n28623 ) | ( ~n28624 & n28623 ) ;
  assign n28629 = n28217 &  n28581 ;
  assign n28630 = n28580 &  n28629 ;
  assign n28618 = x105 | n28217 ;
  assign n28619 = x105 &  n28217 ;
  assign n28620 = ( n28618 & ~n28619 ) | ( n28618 & 1'b0 ) | ( ~n28619 & 1'b0 ) ;
  assign n28632 = ( n28570 & n28582 ) | ( n28570 & n28620 ) | ( n28582 & n28620 ) ;
  assign n28631 = n28570 | n28620 ;
  assign n28633 = ( n28630 & ~n28632 ) | ( n28630 & n28631 ) | ( ~n28632 & n28631 ) ;
  assign n28637 = n28225 &  n28581 ;
  assign n28638 = n28580 &  n28637 ;
  assign n28626 = x104 | n28225 ;
  assign n28627 = x104 &  n28225 ;
  assign n28628 = ( n28626 & ~n28627 ) | ( n28626 & 1'b0 ) | ( ~n28627 & 1'b0 ) ;
  assign n28640 = ( n28569 & n28582 ) | ( n28569 & n28628 ) | ( n28582 & n28628 ) ;
  assign n28639 = n28569 | n28628 ;
  assign n28641 = ( n28638 & ~n28640 ) | ( n28638 & n28639 ) | ( ~n28640 & n28639 ) ;
  assign n28645 = n28233 &  n28581 ;
  assign n28646 = n28580 &  n28645 ;
  assign n28634 = x103 | n28233 ;
  assign n28635 = x103 &  n28233 ;
  assign n28636 = ( n28634 & ~n28635 ) | ( n28634 & 1'b0 ) | ( ~n28635 & 1'b0 ) ;
  assign n28648 = ( n28568 & n28582 ) | ( n28568 & n28636 ) | ( n28582 & n28636 ) ;
  assign n28647 = n28568 | n28636 ;
  assign n28649 = ( n28646 & ~n28648 ) | ( n28646 & n28647 ) | ( ~n28648 & n28647 ) ;
  assign n28653 = n28241 &  n28581 ;
  assign n28654 = n28580 &  n28653 ;
  assign n28642 = x102 | n28241 ;
  assign n28643 = x102 &  n28241 ;
  assign n28644 = ( n28642 & ~n28643 ) | ( n28642 & 1'b0 ) | ( ~n28643 & 1'b0 ) ;
  assign n28656 = ( n28567 & n28582 ) | ( n28567 & n28644 ) | ( n28582 & n28644 ) ;
  assign n28655 = n28567 | n28644 ;
  assign n28657 = ( n28654 & ~n28656 ) | ( n28654 & n28655 ) | ( ~n28656 & n28655 ) ;
  assign n28661 = n28249 &  n28581 ;
  assign n28662 = n28580 &  n28661 ;
  assign n28650 = x101 | n28249 ;
  assign n28651 = x101 &  n28249 ;
  assign n28652 = ( n28650 & ~n28651 ) | ( n28650 & 1'b0 ) | ( ~n28651 & 1'b0 ) ;
  assign n28664 = ( n28566 & n28582 ) | ( n28566 & n28652 ) | ( n28582 & n28652 ) ;
  assign n28663 = n28566 | n28652 ;
  assign n28665 = ( n28662 & ~n28664 ) | ( n28662 & n28663 ) | ( ~n28664 & n28663 ) ;
  assign n28669 = n28257 &  n28581 ;
  assign n28670 = n28580 &  n28669 ;
  assign n28658 = x100 | n28257 ;
  assign n28659 = x100 &  n28257 ;
  assign n28660 = ( n28658 & ~n28659 ) | ( n28658 & 1'b0 ) | ( ~n28659 & 1'b0 ) ;
  assign n28672 = ( n28565 & n28582 ) | ( n28565 & n28660 ) | ( n28582 & n28660 ) ;
  assign n28671 = n28565 | n28660 ;
  assign n28673 = ( n28670 & ~n28672 ) | ( n28670 & n28671 ) | ( ~n28672 & n28671 ) ;
  assign n28677 = n28265 &  n28581 ;
  assign n28678 = n28580 &  n28677 ;
  assign n28666 = x99 | n28265 ;
  assign n28667 = x99 &  n28265 ;
  assign n28668 = ( n28666 & ~n28667 ) | ( n28666 & 1'b0 ) | ( ~n28667 & 1'b0 ) ;
  assign n28680 = ( n28564 & n28582 ) | ( n28564 & n28668 ) | ( n28582 & n28668 ) ;
  assign n28679 = n28564 | n28668 ;
  assign n28681 = ( n28678 & ~n28680 ) | ( n28678 & n28679 ) | ( ~n28680 & n28679 ) ;
  assign n28685 = n28273 &  n28581 ;
  assign n28686 = n28580 &  n28685 ;
  assign n28674 = x98 | n28273 ;
  assign n28675 = x98 &  n28273 ;
  assign n28676 = ( n28674 & ~n28675 ) | ( n28674 & 1'b0 ) | ( ~n28675 & 1'b0 ) ;
  assign n28688 = ( n28563 & n28582 ) | ( n28563 & n28676 ) | ( n28582 & n28676 ) ;
  assign n28687 = n28563 | n28676 ;
  assign n28689 = ( n28686 & ~n28688 ) | ( n28686 & n28687 ) | ( ~n28688 & n28687 ) ;
  assign n28693 = n28281 &  n28581 ;
  assign n28694 = n28580 &  n28693 ;
  assign n28682 = x97 | n28281 ;
  assign n28683 = x97 &  n28281 ;
  assign n28684 = ( n28682 & ~n28683 ) | ( n28682 & 1'b0 ) | ( ~n28683 & 1'b0 ) ;
  assign n28696 = ( n28562 & n28582 ) | ( n28562 & n28684 ) | ( n28582 & n28684 ) ;
  assign n28695 = n28562 | n28684 ;
  assign n28697 = ( n28694 & ~n28696 ) | ( n28694 & n28695 ) | ( ~n28696 & n28695 ) ;
  assign n28701 = n28289 &  n28581 ;
  assign n28702 = n28580 &  n28701 ;
  assign n28690 = x96 | n28289 ;
  assign n28691 = x96 &  n28289 ;
  assign n28692 = ( n28690 & ~n28691 ) | ( n28690 & 1'b0 ) | ( ~n28691 & 1'b0 ) ;
  assign n28704 = ( n28561 & n28582 ) | ( n28561 & n28692 ) | ( n28582 & n28692 ) ;
  assign n28703 = n28561 | n28692 ;
  assign n28705 = ( n28702 & ~n28704 ) | ( n28702 & n28703 ) | ( ~n28704 & n28703 ) ;
  assign n28709 = n28297 &  n28581 ;
  assign n28710 = n28580 &  n28709 ;
  assign n28698 = x95 | n28297 ;
  assign n28699 = x95 &  n28297 ;
  assign n28700 = ( n28698 & ~n28699 ) | ( n28698 & 1'b0 ) | ( ~n28699 & 1'b0 ) ;
  assign n28712 = ( n28560 & n28582 ) | ( n28560 & n28700 ) | ( n28582 & n28700 ) ;
  assign n28711 = n28560 | n28700 ;
  assign n28713 = ( n28710 & ~n28712 ) | ( n28710 & n28711 ) | ( ~n28712 & n28711 ) ;
  assign n28717 = n28305 &  n28581 ;
  assign n28718 = n28580 &  n28717 ;
  assign n28706 = x94 | n28305 ;
  assign n28707 = x94 &  n28305 ;
  assign n28708 = ( n28706 & ~n28707 ) | ( n28706 & 1'b0 ) | ( ~n28707 & 1'b0 ) ;
  assign n28720 = ( n28559 & n28582 ) | ( n28559 & n28708 ) | ( n28582 & n28708 ) ;
  assign n28719 = n28559 | n28708 ;
  assign n28721 = ( n28718 & ~n28720 ) | ( n28718 & n28719 ) | ( ~n28720 & n28719 ) ;
  assign n28725 = n28313 &  n28581 ;
  assign n28726 = n28580 &  n28725 ;
  assign n28714 = x93 | n28313 ;
  assign n28715 = x93 &  n28313 ;
  assign n28716 = ( n28714 & ~n28715 ) | ( n28714 & 1'b0 ) | ( ~n28715 & 1'b0 ) ;
  assign n28728 = ( n28558 & n28582 ) | ( n28558 & n28716 ) | ( n28582 & n28716 ) ;
  assign n28727 = n28558 | n28716 ;
  assign n28729 = ( n28726 & ~n28728 ) | ( n28726 & n28727 ) | ( ~n28728 & n28727 ) ;
  assign n28733 = n28321 &  n28581 ;
  assign n28734 = n28580 &  n28733 ;
  assign n28722 = x92 | n28321 ;
  assign n28723 = x92 &  n28321 ;
  assign n28724 = ( n28722 & ~n28723 ) | ( n28722 & 1'b0 ) | ( ~n28723 & 1'b0 ) ;
  assign n28736 = ( n28557 & n28582 ) | ( n28557 & n28724 ) | ( n28582 & n28724 ) ;
  assign n28735 = n28557 | n28724 ;
  assign n28737 = ( n28734 & ~n28736 ) | ( n28734 & n28735 ) | ( ~n28736 & n28735 ) ;
  assign n28741 = n28329 &  n28581 ;
  assign n28742 = n28580 &  n28741 ;
  assign n28730 = x91 | n28329 ;
  assign n28731 = x91 &  n28329 ;
  assign n28732 = ( n28730 & ~n28731 ) | ( n28730 & 1'b0 ) | ( ~n28731 & 1'b0 ) ;
  assign n28744 = ( n28556 & n28582 ) | ( n28556 & n28732 ) | ( n28582 & n28732 ) ;
  assign n28743 = n28556 | n28732 ;
  assign n28745 = ( n28742 & ~n28744 ) | ( n28742 & n28743 ) | ( ~n28744 & n28743 ) ;
  assign n28749 = n28337 &  n28581 ;
  assign n28750 = n28580 &  n28749 ;
  assign n28738 = x90 | n28337 ;
  assign n28739 = x90 &  n28337 ;
  assign n28740 = ( n28738 & ~n28739 ) | ( n28738 & 1'b0 ) | ( ~n28739 & 1'b0 ) ;
  assign n28752 = ( n28555 & n28582 ) | ( n28555 & n28740 ) | ( n28582 & n28740 ) ;
  assign n28751 = n28555 | n28740 ;
  assign n28753 = ( n28750 & ~n28752 ) | ( n28750 & n28751 ) | ( ~n28752 & n28751 ) ;
  assign n28757 = n28345 &  n28581 ;
  assign n28758 = n28580 &  n28757 ;
  assign n28746 = x89 | n28345 ;
  assign n28747 = x89 &  n28345 ;
  assign n28748 = ( n28746 & ~n28747 ) | ( n28746 & 1'b0 ) | ( ~n28747 & 1'b0 ) ;
  assign n28760 = ( n28554 & n28582 ) | ( n28554 & n28748 ) | ( n28582 & n28748 ) ;
  assign n28759 = n28554 | n28748 ;
  assign n28761 = ( n28758 & ~n28760 ) | ( n28758 & n28759 ) | ( ~n28760 & n28759 ) ;
  assign n28765 = n28353 &  n28581 ;
  assign n28766 = n28580 &  n28765 ;
  assign n28754 = x88 | n28353 ;
  assign n28755 = x88 &  n28353 ;
  assign n28756 = ( n28754 & ~n28755 ) | ( n28754 & 1'b0 ) | ( ~n28755 & 1'b0 ) ;
  assign n28768 = ( n28553 & n28582 ) | ( n28553 & n28756 ) | ( n28582 & n28756 ) ;
  assign n28767 = n28553 | n28756 ;
  assign n28769 = ( n28766 & ~n28768 ) | ( n28766 & n28767 ) | ( ~n28768 & n28767 ) ;
  assign n28773 = n28361 &  n28581 ;
  assign n28774 = n28580 &  n28773 ;
  assign n28762 = x87 | n28361 ;
  assign n28763 = x87 &  n28361 ;
  assign n28764 = ( n28762 & ~n28763 ) | ( n28762 & 1'b0 ) | ( ~n28763 & 1'b0 ) ;
  assign n28776 = ( n28552 & n28582 ) | ( n28552 & n28764 ) | ( n28582 & n28764 ) ;
  assign n28775 = n28552 | n28764 ;
  assign n28777 = ( n28774 & ~n28776 ) | ( n28774 & n28775 ) | ( ~n28776 & n28775 ) ;
  assign n28781 = n28369 &  n28581 ;
  assign n28782 = n28580 &  n28781 ;
  assign n28770 = x86 | n28369 ;
  assign n28771 = x86 &  n28369 ;
  assign n28772 = ( n28770 & ~n28771 ) | ( n28770 & 1'b0 ) | ( ~n28771 & 1'b0 ) ;
  assign n28784 = ( n28551 & n28582 ) | ( n28551 & n28772 ) | ( n28582 & n28772 ) ;
  assign n28783 = n28551 | n28772 ;
  assign n28785 = ( n28782 & ~n28784 ) | ( n28782 & n28783 ) | ( ~n28784 & n28783 ) ;
  assign n28789 = n28377 &  n28581 ;
  assign n28790 = n28580 &  n28789 ;
  assign n28778 = x85 | n28377 ;
  assign n28779 = x85 &  n28377 ;
  assign n28780 = ( n28778 & ~n28779 ) | ( n28778 & 1'b0 ) | ( ~n28779 & 1'b0 ) ;
  assign n28792 = ( n28550 & n28582 ) | ( n28550 & n28780 ) | ( n28582 & n28780 ) ;
  assign n28791 = n28550 | n28780 ;
  assign n28793 = ( n28790 & ~n28792 ) | ( n28790 & n28791 ) | ( ~n28792 & n28791 ) ;
  assign n28797 = n28385 &  n28581 ;
  assign n28798 = n28580 &  n28797 ;
  assign n28786 = x84 | n28385 ;
  assign n28787 = x84 &  n28385 ;
  assign n28788 = ( n28786 & ~n28787 ) | ( n28786 & 1'b0 ) | ( ~n28787 & 1'b0 ) ;
  assign n28800 = ( n28549 & n28582 ) | ( n28549 & n28788 ) | ( n28582 & n28788 ) ;
  assign n28799 = n28549 | n28788 ;
  assign n28801 = ( n28798 & ~n28800 ) | ( n28798 & n28799 ) | ( ~n28800 & n28799 ) ;
  assign n28805 = n28393 &  n28581 ;
  assign n28806 = n28580 &  n28805 ;
  assign n28794 = x83 | n28393 ;
  assign n28795 = x83 &  n28393 ;
  assign n28796 = ( n28794 & ~n28795 ) | ( n28794 & 1'b0 ) | ( ~n28795 & 1'b0 ) ;
  assign n28808 = ( n28548 & n28582 ) | ( n28548 & n28796 ) | ( n28582 & n28796 ) ;
  assign n28807 = n28548 | n28796 ;
  assign n28809 = ( n28806 & ~n28808 ) | ( n28806 & n28807 ) | ( ~n28808 & n28807 ) ;
  assign n28813 = n28401 &  n28581 ;
  assign n28814 = n28580 &  n28813 ;
  assign n28802 = x82 | n28401 ;
  assign n28803 = x82 &  n28401 ;
  assign n28804 = ( n28802 & ~n28803 ) | ( n28802 & 1'b0 ) | ( ~n28803 & 1'b0 ) ;
  assign n28816 = ( n28547 & n28582 ) | ( n28547 & n28804 ) | ( n28582 & n28804 ) ;
  assign n28815 = n28547 | n28804 ;
  assign n28817 = ( n28814 & ~n28816 ) | ( n28814 & n28815 ) | ( ~n28816 & n28815 ) ;
  assign n28821 = n28409 &  n28581 ;
  assign n28822 = n28580 &  n28821 ;
  assign n28810 = x81 | n28409 ;
  assign n28811 = x81 &  n28409 ;
  assign n28812 = ( n28810 & ~n28811 ) | ( n28810 & 1'b0 ) | ( ~n28811 & 1'b0 ) ;
  assign n28824 = ( n28546 & n28582 ) | ( n28546 & n28812 ) | ( n28582 & n28812 ) ;
  assign n28823 = n28546 | n28812 ;
  assign n28825 = ( n28822 & ~n28824 ) | ( n28822 & n28823 ) | ( ~n28824 & n28823 ) ;
  assign n28829 = n28417 &  n28581 ;
  assign n28830 = n28580 &  n28829 ;
  assign n28818 = x80 | n28417 ;
  assign n28819 = x80 &  n28417 ;
  assign n28820 = ( n28818 & ~n28819 ) | ( n28818 & 1'b0 ) | ( ~n28819 & 1'b0 ) ;
  assign n28832 = ( n28545 & n28582 ) | ( n28545 & n28820 ) | ( n28582 & n28820 ) ;
  assign n28831 = n28545 | n28820 ;
  assign n28833 = ( n28830 & ~n28832 ) | ( n28830 & n28831 ) | ( ~n28832 & n28831 ) ;
  assign n28837 = n28425 &  n28581 ;
  assign n28838 = n28580 &  n28837 ;
  assign n28826 = x79 | n28425 ;
  assign n28827 = x79 &  n28425 ;
  assign n28828 = ( n28826 & ~n28827 ) | ( n28826 & 1'b0 ) | ( ~n28827 & 1'b0 ) ;
  assign n28840 = ( n28544 & n28582 ) | ( n28544 & n28828 ) | ( n28582 & n28828 ) ;
  assign n28839 = n28544 | n28828 ;
  assign n28841 = ( n28838 & ~n28840 ) | ( n28838 & n28839 ) | ( ~n28840 & n28839 ) ;
  assign n28845 = n28433 &  n28581 ;
  assign n28846 = n28580 &  n28845 ;
  assign n28834 = x78 | n28433 ;
  assign n28835 = x78 &  n28433 ;
  assign n28836 = ( n28834 & ~n28835 ) | ( n28834 & 1'b0 ) | ( ~n28835 & 1'b0 ) ;
  assign n28848 = ( n28543 & n28582 ) | ( n28543 & n28836 ) | ( n28582 & n28836 ) ;
  assign n28847 = n28543 | n28836 ;
  assign n28849 = ( n28846 & ~n28848 ) | ( n28846 & n28847 ) | ( ~n28848 & n28847 ) ;
  assign n28853 = n28441 &  n28581 ;
  assign n28854 = n28580 &  n28853 ;
  assign n28842 = x77 | n28441 ;
  assign n28843 = x77 &  n28441 ;
  assign n28844 = ( n28842 & ~n28843 ) | ( n28842 & 1'b0 ) | ( ~n28843 & 1'b0 ) ;
  assign n28856 = ( n28542 & n28582 ) | ( n28542 & n28844 ) | ( n28582 & n28844 ) ;
  assign n28855 = n28542 | n28844 ;
  assign n28857 = ( n28854 & ~n28856 ) | ( n28854 & n28855 ) | ( ~n28856 & n28855 ) ;
  assign n28861 = n28449 &  n28581 ;
  assign n28862 = n28580 &  n28861 ;
  assign n28850 = x76 | n28449 ;
  assign n28851 = x76 &  n28449 ;
  assign n28852 = ( n28850 & ~n28851 ) | ( n28850 & 1'b0 ) | ( ~n28851 & 1'b0 ) ;
  assign n28864 = ( n28541 & n28582 ) | ( n28541 & n28852 ) | ( n28582 & n28852 ) ;
  assign n28863 = n28541 | n28852 ;
  assign n28865 = ( n28862 & ~n28864 ) | ( n28862 & n28863 ) | ( ~n28864 & n28863 ) ;
  assign n28869 = n28457 &  n28581 ;
  assign n28870 = n28580 &  n28869 ;
  assign n28858 = x75 | n28457 ;
  assign n28859 = x75 &  n28457 ;
  assign n28860 = ( n28858 & ~n28859 ) | ( n28858 & 1'b0 ) | ( ~n28859 & 1'b0 ) ;
  assign n28872 = ( n28540 & n28582 ) | ( n28540 & n28860 ) | ( n28582 & n28860 ) ;
  assign n28871 = n28540 | n28860 ;
  assign n28873 = ( n28870 & ~n28872 ) | ( n28870 & n28871 ) | ( ~n28872 & n28871 ) ;
  assign n28877 = n28465 &  n28581 ;
  assign n28878 = n28580 &  n28877 ;
  assign n28866 = x74 | n28465 ;
  assign n28867 = x74 &  n28465 ;
  assign n28868 = ( n28866 & ~n28867 ) | ( n28866 & 1'b0 ) | ( ~n28867 & 1'b0 ) ;
  assign n28880 = ( n28539 & n28582 ) | ( n28539 & n28868 ) | ( n28582 & n28868 ) ;
  assign n28879 = n28539 | n28868 ;
  assign n28881 = ( n28878 & ~n28880 ) | ( n28878 & n28879 ) | ( ~n28880 & n28879 ) ;
  assign n28885 = n28473 &  n28581 ;
  assign n28886 = n28580 &  n28885 ;
  assign n28874 = x73 | n28473 ;
  assign n28875 = x73 &  n28473 ;
  assign n28876 = ( n28874 & ~n28875 ) | ( n28874 & 1'b0 ) | ( ~n28875 & 1'b0 ) ;
  assign n28888 = ( n28538 & n28582 ) | ( n28538 & n28876 ) | ( n28582 & n28876 ) ;
  assign n28887 = n28538 | n28876 ;
  assign n28889 = ( n28886 & ~n28888 ) | ( n28886 & n28887 ) | ( ~n28888 & n28887 ) ;
  assign n28893 = n28481 &  n28581 ;
  assign n28894 = n28580 &  n28893 ;
  assign n28882 = x72 | n28481 ;
  assign n28883 = x72 &  n28481 ;
  assign n28884 = ( n28882 & ~n28883 ) | ( n28882 & 1'b0 ) | ( ~n28883 & 1'b0 ) ;
  assign n28896 = ( n28537 & n28582 ) | ( n28537 & n28884 ) | ( n28582 & n28884 ) ;
  assign n28895 = n28537 | n28884 ;
  assign n28897 = ( n28894 & ~n28896 ) | ( n28894 & n28895 ) | ( ~n28896 & n28895 ) ;
  assign n28901 = n28489 &  n28581 ;
  assign n28902 = n28580 &  n28901 ;
  assign n28890 = x71 | n28489 ;
  assign n28891 = x71 &  n28489 ;
  assign n28892 = ( n28890 & ~n28891 ) | ( n28890 & 1'b0 ) | ( ~n28891 & 1'b0 ) ;
  assign n28904 = ( n28536 & n28582 ) | ( n28536 & n28892 ) | ( n28582 & n28892 ) ;
  assign n28903 = n28536 | n28892 ;
  assign n28905 = ( n28902 & ~n28904 ) | ( n28902 & n28903 ) | ( ~n28904 & n28903 ) ;
  assign n28909 = n28497 &  n28581 ;
  assign n28910 = n28580 &  n28909 ;
  assign n28898 = x70 | n28497 ;
  assign n28899 = x70 &  n28497 ;
  assign n28900 = ( n28898 & ~n28899 ) | ( n28898 & 1'b0 ) | ( ~n28899 & 1'b0 ) ;
  assign n28912 = ( n28535 & n28582 ) | ( n28535 & n28900 ) | ( n28582 & n28900 ) ;
  assign n28911 = n28535 | n28900 ;
  assign n28913 = ( n28910 & ~n28912 ) | ( n28910 & n28911 ) | ( ~n28912 & n28911 ) ;
  assign n28917 = n28505 &  n28581 ;
  assign n28918 = n28580 &  n28917 ;
  assign n28906 = x69 | n28505 ;
  assign n28907 = x69 &  n28505 ;
  assign n28908 = ( n28906 & ~n28907 ) | ( n28906 & 1'b0 ) | ( ~n28907 & 1'b0 ) ;
  assign n28920 = ( n28534 & n28582 ) | ( n28534 & n28908 ) | ( n28582 & n28908 ) ;
  assign n28919 = n28534 | n28908 ;
  assign n28921 = ( n28918 & ~n28920 ) | ( n28918 & n28919 ) | ( ~n28920 & n28919 ) ;
  assign n28925 = n28513 &  n28581 ;
  assign n28926 = n28580 &  n28925 ;
  assign n28914 = x68 | n28513 ;
  assign n28915 = x68 &  n28513 ;
  assign n28916 = ( n28914 & ~n28915 ) | ( n28914 & 1'b0 ) | ( ~n28915 & 1'b0 ) ;
  assign n28928 = ( n28533 & n28582 ) | ( n28533 & n28916 ) | ( n28582 & n28916 ) ;
  assign n28927 = n28533 | n28916 ;
  assign n28929 = ( n28926 & ~n28928 ) | ( n28926 & n28927 ) | ( ~n28928 & n28927 ) ;
  assign n28933 = n28518 &  n28581 ;
  assign n28934 = n28580 &  n28933 ;
  assign n28922 = x67 | n28518 ;
  assign n28923 = x67 &  n28518 ;
  assign n28924 = ( n28922 & ~n28923 ) | ( n28922 & 1'b0 ) | ( ~n28923 & 1'b0 ) ;
  assign n28936 = ( n28532 & n28582 ) | ( n28532 & n28924 ) | ( n28582 & n28924 ) ;
  assign n28935 = n28532 | n28924 ;
  assign n28937 = ( n28934 & ~n28936 ) | ( n28934 & n28935 ) | ( ~n28936 & n28935 ) ;
  assign n28938 = n28526 &  n28581 ;
  assign n28939 = n28580 &  n28938 ;
  assign n28930 = x66 | n28526 ;
  assign n28931 = x66 &  n28526 ;
  assign n28932 = ( n28930 & ~n28931 ) | ( n28930 & 1'b0 ) | ( ~n28931 & 1'b0 ) ;
  assign n28941 = ( n28531 & n28582 ) | ( n28531 & n28932 ) | ( n28582 & n28932 ) ;
  assign n28940 = n28531 | n28932 ;
  assign n28942 = ( n28939 & ~n28941 ) | ( n28939 & n28940 ) | ( ~n28941 & n28940 ) ;
  assign n28943 = ( x65 & ~n10112 ) | ( x65 & n28530 ) | ( ~n10112 & n28530 ) ;
  assign n28944 = ( n28531 & ~x65 ) | ( n28531 & n28943 ) | ( ~x65 & n28943 ) ;
  assign n28945 = ~n28582 & n28944 ;
  assign n28946 = n28530 &  n28581 ;
  assign n28947 = n28580 &  n28946 ;
  assign n28948 = n28945 | n28947 ;
  assign n28949 = ( x64 & ~n28582 ) | ( x64 & 1'b0 ) | ( ~n28582 & 1'b0 ) ;
  assign n28950 = ( x17 & ~n28949 ) | ( x17 & 1'b0 ) | ( ~n28949 & 1'b0 ) ;
  assign n28951 = ( n10112 & ~n28582 ) | ( n10112 & 1'b0 ) | ( ~n28582 & 1'b0 ) ;
  assign n28952 = n28950 | n28951 ;
  assign n28953 = ( x65 & ~n28952 ) | ( x65 & n10539 ) | ( ~n28952 & n10539 ) ;
  assign n28954 = ( x66 & ~n28948 ) | ( x66 & n28953 ) | ( ~n28948 & n28953 ) ;
  assign n28955 = ( x67 & ~n28942 ) | ( x67 & n28954 ) | ( ~n28942 & n28954 ) ;
  assign n28956 = ( x68 & ~n28937 ) | ( x68 & n28955 ) | ( ~n28937 & n28955 ) ;
  assign n28957 = ( x69 & ~n28929 ) | ( x69 & n28956 ) | ( ~n28929 & n28956 ) ;
  assign n28958 = ( x70 & ~n28921 ) | ( x70 & n28957 ) | ( ~n28921 & n28957 ) ;
  assign n28959 = ( x71 & ~n28913 ) | ( x71 & n28958 ) | ( ~n28913 & n28958 ) ;
  assign n28960 = ( x72 & ~n28905 ) | ( x72 & n28959 ) | ( ~n28905 & n28959 ) ;
  assign n28961 = ( x73 & ~n28897 ) | ( x73 & n28960 ) | ( ~n28897 & n28960 ) ;
  assign n28962 = ( x74 & ~n28889 ) | ( x74 & n28961 ) | ( ~n28889 & n28961 ) ;
  assign n28963 = ( x75 & ~n28881 ) | ( x75 & n28962 ) | ( ~n28881 & n28962 ) ;
  assign n28964 = ( x76 & ~n28873 ) | ( x76 & n28963 ) | ( ~n28873 & n28963 ) ;
  assign n28965 = ( x77 & ~n28865 ) | ( x77 & n28964 ) | ( ~n28865 & n28964 ) ;
  assign n28966 = ( x78 & ~n28857 ) | ( x78 & n28965 ) | ( ~n28857 & n28965 ) ;
  assign n28967 = ( x79 & ~n28849 ) | ( x79 & n28966 ) | ( ~n28849 & n28966 ) ;
  assign n28968 = ( x80 & ~n28841 ) | ( x80 & n28967 ) | ( ~n28841 & n28967 ) ;
  assign n28969 = ( x81 & ~n28833 ) | ( x81 & n28968 ) | ( ~n28833 & n28968 ) ;
  assign n28970 = ( x82 & ~n28825 ) | ( x82 & n28969 ) | ( ~n28825 & n28969 ) ;
  assign n28971 = ( x83 & ~n28817 ) | ( x83 & n28970 ) | ( ~n28817 & n28970 ) ;
  assign n28972 = ( x84 & ~n28809 ) | ( x84 & n28971 ) | ( ~n28809 & n28971 ) ;
  assign n28973 = ( x85 & ~n28801 ) | ( x85 & n28972 ) | ( ~n28801 & n28972 ) ;
  assign n28974 = ( x86 & ~n28793 ) | ( x86 & n28973 ) | ( ~n28793 & n28973 ) ;
  assign n28975 = ( x87 & ~n28785 ) | ( x87 & n28974 ) | ( ~n28785 & n28974 ) ;
  assign n28976 = ( x88 & ~n28777 ) | ( x88 & n28975 ) | ( ~n28777 & n28975 ) ;
  assign n28977 = ( x89 & ~n28769 ) | ( x89 & n28976 ) | ( ~n28769 & n28976 ) ;
  assign n28978 = ( x90 & ~n28761 ) | ( x90 & n28977 ) | ( ~n28761 & n28977 ) ;
  assign n28979 = ( x91 & ~n28753 ) | ( x91 & n28978 ) | ( ~n28753 & n28978 ) ;
  assign n28980 = ( x92 & ~n28745 ) | ( x92 & n28979 ) | ( ~n28745 & n28979 ) ;
  assign n28981 = ( x93 & ~n28737 ) | ( x93 & n28980 ) | ( ~n28737 & n28980 ) ;
  assign n28982 = ( x94 & ~n28729 ) | ( x94 & n28981 ) | ( ~n28729 & n28981 ) ;
  assign n28983 = ( x95 & ~n28721 ) | ( x95 & n28982 ) | ( ~n28721 & n28982 ) ;
  assign n28984 = ( x96 & ~n28713 ) | ( x96 & n28983 ) | ( ~n28713 & n28983 ) ;
  assign n28985 = ( x97 & ~n28705 ) | ( x97 & n28984 ) | ( ~n28705 & n28984 ) ;
  assign n28986 = ( x98 & ~n28697 ) | ( x98 & n28985 ) | ( ~n28697 & n28985 ) ;
  assign n28987 = ( x99 & ~n28689 ) | ( x99 & n28986 ) | ( ~n28689 & n28986 ) ;
  assign n28988 = ( x100 & ~n28681 ) | ( x100 & n28987 ) | ( ~n28681 & n28987 ) ;
  assign n28989 = ( x101 & ~n28673 ) | ( x101 & n28988 ) | ( ~n28673 & n28988 ) ;
  assign n28990 = ( x102 & ~n28665 ) | ( x102 & n28989 ) | ( ~n28665 & n28989 ) ;
  assign n28991 = ( x103 & ~n28657 ) | ( x103 & n28990 ) | ( ~n28657 & n28990 ) ;
  assign n28992 = ( x104 & ~n28649 ) | ( x104 & n28991 ) | ( ~n28649 & n28991 ) ;
  assign n28993 = ( x105 & ~n28641 ) | ( x105 & n28992 ) | ( ~n28641 & n28992 ) ;
  assign n28994 = ( x106 & ~n28633 ) | ( x106 & n28993 ) | ( ~n28633 & n28993 ) ;
  assign n28995 = ( x107 & ~n28625 ) | ( x107 & n28994 ) | ( ~n28625 & n28994 ) ;
  assign n28996 = ( x108 & ~n28617 ) | ( x108 & n28995 ) | ( ~n28617 & n28995 ) ;
  assign n28997 = ( x109 & ~n28609 ) | ( x109 & n28996 ) | ( ~n28609 & n28996 ) ;
  assign n28998 = ( x110 & ~n28601 ) | ( x110 & n28997 ) | ( ~n28601 & n28997 ) ;
  assign n28999 = ( x111 & ~n28591 ) | ( x111 & 1'b0 ) | ( ~n28591 & 1'b0 ) ;
  assign n29000 = ~n28589 & n28999 ;
  assign n29001 = ( n28998 & ~n28593 ) | ( n28998 & n29000 ) | ( ~n28593 & n29000 ) ;
  assign n29002 = ( n28593 & ~n270 ) | ( n28593 & n29001 ) | ( ~n270 & n29001 ) ;
  assign n29003 = n270 | n29002 ;
  assign n29004 = ~n28592 |  n10264 ;
  assign n29018 = n28601 &  n29004 ;
  assign n29019 = n29003 &  n29018 ;
  assign n29005 = n29003 &  n29004 ;
  assign n29006 = x110 | n28601 ;
  assign n29007 = x110 &  n28601 ;
  assign n29008 = ( n29006 & ~n29007 ) | ( n29006 & 1'b0 ) | ( ~n29007 & 1'b0 ) ;
  assign n29021 = ( n28997 & n29005 ) | ( n28997 & n29008 ) | ( n29005 & n29008 ) ;
  assign n29020 = n28997 | n29008 ;
  assign n29022 = ( n29019 & ~n29021 ) | ( n29019 & n29020 ) | ( ~n29021 & n29020 ) ;
  assign n29010 = n10264 &  n28592 ;
  assign n29011 = n29003 &  n29010 ;
  assign n29009 = n28593 | n29000 ;
  assign n29013 = ( n28998 & n29005 ) | ( n28998 & n29009 ) | ( n29005 & n29009 ) ;
  assign n29012 = n28998 | n29009 ;
  assign n29014 = ( n29011 & ~n29013 ) | ( n29011 & n29012 ) | ( ~n29013 & n29012 ) ;
  assign n29026 = n28609 &  n29004 ;
  assign n29027 = n29003 &  n29026 ;
  assign n29015 = x109 | n28609 ;
  assign n29016 = x109 &  n28609 ;
  assign n29017 = ( n29015 & ~n29016 ) | ( n29015 & 1'b0 ) | ( ~n29016 & 1'b0 ) ;
  assign n29029 = ( n28996 & n29005 ) | ( n28996 & n29017 ) | ( n29005 & n29017 ) ;
  assign n29028 = n28996 | n29017 ;
  assign n29030 = ( n29027 & ~n29029 ) | ( n29027 & n29028 ) | ( ~n29029 & n29028 ) ;
  assign n29034 = n28617 &  n29004 ;
  assign n29035 = n29003 &  n29034 ;
  assign n29023 = x108 | n28617 ;
  assign n29024 = x108 &  n28617 ;
  assign n29025 = ( n29023 & ~n29024 ) | ( n29023 & 1'b0 ) | ( ~n29024 & 1'b0 ) ;
  assign n29037 = ( n28995 & n29005 ) | ( n28995 & n29025 ) | ( n29005 & n29025 ) ;
  assign n29036 = n28995 | n29025 ;
  assign n29038 = ( n29035 & ~n29037 ) | ( n29035 & n29036 ) | ( ~n29037 & n29036 ) ;
  assign n29042 = n28625 &  n29004 ;
  assign n29043 = n29003 &  n29042 ;
  assign n29031 = x107 | n28625 ;
  assign n29032 = x107 &  n28625 ;
  assign n29033 = ( n29031 & ~n29032 ) | ( n29031 & 1'b0 ) | ( ~n29032 & 1'b0 ) ;
  assign n29045 = ( n28994 & n29005 ) | ( n28994 & n29033 ) | ( n29005 & n29033 ) ;
  assign n29044 = n28994 | n29033 ;
  assign n29046 = ( n29043 & ~n29045 ) | ( n29043 & n29044 ) | ( ~n29045 & n29044 ) ;
  assign n29050 = n28633 &  n29004 ;
  assign n29051 = n29003 &  n29050 ;
  assign n29039 = x106 | n28633 ;
  assign n29040 = x106 &  n28633 ;
  assign n29041 = ( n29039 & ~n29040 ) | ( n29039 & 1'b0 ) | ( ~n29040 & 1'b0 ) ;
  assign n29053 = ( n28993 & n29005 ) | ( n28993 & n29041 ) | ( n29005 & n29041 ) ;
  assign n29052 = n28993 | n29041 ;
  assign n29054 = ( n29051 & ~n29053 ) | ( n29051 & n29052 ) | ( ~n29053 & n29052 ) ;
  assign n29058 = n28641 &  n29004 ;
  assign n29059 = n29003 &  n29058 ;
  assign n29047 = x105 | n28641 ;
  assign n29048 = x105 &  n28641 ;
  assign n29049 = ( n29047 & ~n29048 ) | ( n29047 & 1'b0 ) | ( ~n29048 & 1'b0 ) ;
  assign n29061 = ( n28992 & n29005 ) | ( n28992 & n29049 ) | ( n29005 & n29049 ) ;
  assign n29060 = n28992 | n29049 ;
  assign n29062 = ( n29059 & ~n29061 ) | ( n29059 & n29060 ) | ( ~n29061 & n29060 ) ;
  assign n29066 = n28649 &  n29004 ;
  assign n29067 = n29003 &  n29066 ;
  assign n29055 = x104 | n28649 ;
  assign n29056 = x104 &  n28649 ;
  assign n29057 = ( n29055 & ~n29056 ) | ( n29055 & 1'b0 ) | ( ~n29056 & 1'b0 ) ;
  assign n29069 = ( n28991 & n29005 ) | ( n28991 & n29057 ) | ( n29005 & n29057 ) ;
  assign n29068 = n28991 | n29057 ;
  assign n29070 = ( n29067 & ~n29069 ) | ( n29067 & n29068 ) | ( ~n29069 & n29068 ) ;
  assign n29074 = n28657 &  n29004 ;
  assign n29075 = n29003 &  n29074 ;
  assign n29063 = x103 | n28657 ;
  assign n29064 = x103 &  n28657 ;
  assign n29065 = ( n29063 & ~n29064 ) | ( n29063 & 1'b0 ) | ( ~n29064 & 1'b0 ) ;
  assign n29077 = ( n28990 & n29005 ) | ( n28990 & n29065 ) | ( n29005 & n29065 ) ;
  assign n29076 = n28990 | n29065 ;
  assign n29078 = ( n29075 & ~n29077 ) | ( n29075 & n29076 ) | ( ~n29077 & n29076 ) ;
  assign n29082 = n28665 &  n29004 ;
  assign n29083 = n29003 &  n29082 ;
  assign n29071 = x102 | n28665 ;
  assign n29072 = x102 &  n28665 ;
  assign n29073 = ( n29071 & ~n29072 ) | ( n29071 & 1'b0 ) | ( ~n29072 & 1'b0 ) ;
  assign n29085 = ( n28989 & n29005 ) | ( n28989 & n29073 ) | ( n29005 & n29073 ) ;
  assign n29084 = n28989 | n29073 ;
  assign n29086 = ( n29083 & ~n29085 ) | ( n29083 & n29084 ) | ( ~n29085 & n29084 ) ;
  assign n29090 = n28673 &  n29004 ;
  assign n29091 = n29003 &  n29090 ;
  assign n29079 = x101 | n28673 ;
  assign n29080 = x101 &  n28673 ;
  assign n29081 = ( n29079 & ~n29080 ) | ( n29079 & 1'b0 ) | ( ~n29080 & 1'b0 ) ;
  assign n29093 = ( n28988 & n29005 ) | ( n28988 & n29081 ) | ( n29005 & n29081 ) ;
  assign n29092 = n28988 | n29081 ;
  assign n29094 = ( n29091 & ~n29093 ) | ( n29091 & n29092 ) | ( ~n29093 & n29092 ) ;
  assign n29098 = n28681 &  n29004 ;
  assign n29099 = n29003 &  n29098 ;
  assign n29087 = x100 | n28681 ;
  assign n29088 = x100 &  n28681 ;
  assign n29089 = ( n29087 & ~n29088 ) | ( n29087 & 1'b0 ) | ( ~n29088 & 1'b0 ) ;
  assign n29101 = ( n28987 & n29005 ) | ( n28987 & n29089 ) | ( n29005 & n29089 ) ;
  assign n29100 = n28987 | n29089 ;
  assign n29102 = ( n29099 & ~n29101 ) | ( n29099 & n29100 ) | ( ~n29101 & n29100 ) ;
  assign n29106 = n28689 &  n29004 ;
  assign n29107 = n29003 &  n29106 ;
  assign n29095 = x99 | n28689 ;
  assign n29096 = x99 &  n28689 ;
  assign n29097 = ( n29095 & ~n29096 ) | ( n29095 & 1'b0 ) | ( ~n29096 & 1'b0 ) ;
  assign n29109 = ( n28986 & n29005 ) | ( n28986 & n29097 ) | ( n29005 & n29097 ) ;
  assign n29108 = n28986 | n29097 ;
  assign n29110 = ( n29107 & ~n29109 ) | ( n29107 & n29108 ) | ( ~n29109 & n29108 ) ;
  assign n29114 = n28697 &  n29004 ;
  assign n29115 = n29003 &  n29114 ;
  assign n29103 = x98 | n28697 ;
  assign n29104 = x98 &  n28697 ;
  assign n29105 = ( n29103 & ~n29104 ) | ( n29103 & 1'b0 ) | ( ~n29104 & 1'b0 ) ;
  assign n29117 = ( n28985 & n29005 ) | ( n28985 & n29105 ) | ( n29005 & n29105 ) ;
  assign n29116 = n28985 | n29105 ;
  assign n29118 = ( n29115 & ~n29117 ) | ( n29115 & n29116 ) | ( ~n29117 & n29116 ) ;
  assign n29122 = n28705 &  n29004 ;
  assign n29123 = n29003 &  n29122 ;
  assign n29111 = x97 | n28705 ;
  assign n29112 = x97 &  n28705 ;
  assign n29113 = ( n29111 & ~n29112 ) | ( n29111 & 1'b0 ) | ( ~n29112 & 1'b0 ) ;
  assign n29125 = ( n28984 & n29005 ) | ( n28984 & n29113 ) | ( n29005 & n29113 ) ;
  assign n29124 = n28984 | n29113 ;
  assign n29126 = ( n29123 & ~n29125 ) | ( n29123 & n29124 ) | ( ~n29125 & n29124 ) ;
  assign n29130 = n28713 &  n29004 ;
  assign n29131 = n29003 &  n29130 ;
  assign n29119 = x96 | n28713 ;
  assign n29120 = x96 &  n28713 ;
  assign n29121 = ( n29119 & ~n29120 ) | ( n29119 & 1'b0 ) | ( ~n29120 & 1'b0 ) ;
  assign n29133 = ( n28983 & n29005 ) | ( n28983 & n29121 ) | ( n29005 & n29121 ) ;
  assign n29132 = n28983 | n29121 ;
  assign n29134 = ( n29131 & ~n29133 ) | ( n29131 & n29132 ) | ( ~n29133 & n29132 ) ;
  assign n29138 = n28721 &  n29004 ;
  assign n29139 = n29003 &  n29138 ;
  assign n29127 = x95 | n28721 ;
  assign n29128 = x95 &  n28721 ;
  assign n29129 = ( n29127 & ~n29128 ) | ( n29127 & 1'b0 ) | ( ~n29128 & 1'b0 ) ;
  assign n29141 = ( n28982 & n29005 ) | ( n28982 & n29129 ) | ( n29005 & n29129 ) ;
  assign n29140 = n28982 | n29129 ;
  assign n29142 = ( n29139 & ~n29141 ) | ( n29139 & n29140 ) | ( ~n29141 & n29140 ) ;
  assign n29146 = n28729 &  n29004 ;
  assign n29147 = n29003 &  n29146 ;
  assign n29135 = x94 | n28729 ;
  assign n29136 = x94 &  n28729 ;
  assign n29137 = ( n29135 & ~n29136 ) | ( n29135 & 1'b0 ) | ( ~n29136 & 1'b0 ) ;
  assign n29149 = ( n28981 & n29005 ) | ( n28981 & n29137 ) | ( n29005 & n29137 ) ;
  assign n29148 = n28981 | n29137 ;
  assign n29150 = ( n29147 & ~n29149 ) | ( n29147 & n29148 ) | ( ~n29149 & n29148 ) ;
  assign n29154 = n28737 &  n29004 ;
  assign n29155 = n29003 &  n29154 ;
  assign n29143 = x93 | n28737 ;
  assign n29144 = x93 &  n28737 ;
  assign n29145 = ( n29143 & ~n29144 ) | ( n29143 & 1'b0 ) | ( ~n29144 & 1'b0 ) ;
  assign n29157 = ( n28980 & n29005 ) | ( n28980 & n29145 ) | ( n29005 & n29145 ) ;
  assign n29156 = n28980 | n29145 ;
  assign n29158 = ( n29155 & ~n29157 ) | ( n29155 & n29156 ) | ( ~n29157 & n29156 ) ;
  assign n29162 = n28745 &  n29004 ;
  assign n29163 = n29003 &  n29162 ;
  assign n29151 = x92 | n28745 ;
  assign n29152 = x92 &  n28745 ;
  assign n29153 = ( n29151 & ~n29152 ) | ( n29151 & 1'b0 ) | ( ~n29152 & 1'b0 ) ;
  assign n29165 = ( n28979 & n29005 ) | ( n28979 & n29153 ) | ( n29005 & n29153 ) ;
  assign n29164 = n28979 | n29153 ;
  assign n29166 = ( n29163 & ~n29165 ) | ( n29163 & n29164 ) | ( ~n29165 & n29164 ) ;
  assign n29170 = n28753 &  n29004 ;
  assign n29171 = n29003 &  n29170 ;
  assign n29159 = x91 | n28753 ;
  assign n29160 = x91 &  n28753 ;
  assign n29161 = ( n29159 & ~n29160 ) | ( n29159 & 1'b0 ) | ( ~n29160 & 1'b0 ) ;
  assign n29173 = ( n28978 & n29005 ) | ( n28978 & n29161 ) | ( n29005 & n29161 ) ;
  assign n29172 = n28978 | n29161 ;
  assign n29174 = ( n29171 & ~n29173 ) | ( n29171 & n29172 ) | ( ~n29173 & n29172 ) ;
  assign n29178 = n28761 &  n29004 ;
  assign n29179 = n29003 &  n29178 ;
  assign n29167 = x90 | n28761 ;
  assign n29168 = x90 &  n28761 ;
  assign n29169 = ( n29167 & ~n29168 ) | ( n29167 & 1'b0 ) | ( ~n29168 & 1'b0 ) ;
  assign n29181 = ( n28977 & n29005 ) | ( n28977 & n29169 ) | ( n29005 & n29169 ) ;
  assign n29180 = n28977 | n29169 ;
  assign n29182 = ( n29179 & ~n29181 ) | ( n29179 & n29180 ) | ( ~n29181 & n29180 ) ;
  assign n29186 = n28769 &  n29004 ;
  assign n29187 = n29003 &  n29186 ;
  assign n29175 = x89 | n28769 ;
  assign n29176 = x89 &  n28769 ;
  assign n29177 = ( n29175 & ~n29176 ) | ( n29175 & 1'b0 ) | ( ~n29176 & 1'b0 ) ;
  assign n29189 = ( n28976 & n29005 ) | ( n28976 & n29177 ) | ( n29005 & n29177 ) ;
  assign n29188 = n28976 | n29177 ;
  assign n29190 = ( n29187 & ~n29189 ) | ( n29187 & n29188 ) | ( ~n29189 & n29188 ) ;
  assign n29194 = n28777 &  n29004 ;
  assign n29195 = n29003 &  n29194 ;
  assign n29183 = x88 | n28777 ;
  assign n29184 = x88 &  n28777 ;
  assign n29185 = ( n29183 & ~n29184 ) | ( n29183 & 1'b0 ) | ( ~n29184 & 1'b0 ) ;
  assign n29197 = ( n28975 & n29005 ) | ( n28975 & n29185 ) | ( n29005 & n29185 ) ;
  assign n29196 = n28975 | n29185 ;
  assign n29198 = ( n29195 & ~n29197 ) | ( n29195 & n29196 ) | ( ~n29197 & n29196 ) ;
  assign n29202 = n28785 &  n29004 ;
  assign n29203 = n29003 &  n29202 ;
  assign n29191 = x87 | n28785 ;
  assign n29192 = x87 &  n28785 ;
  assign n29193 = ( n29191 & ~n29192 ) | ( n29191 & 1'b0 ) | ( ~n29192 & 1'b0 ) ;
  assign n29205 = ( n28974 & n29005 ) | ( n28974 & n29193 ) | ( n29005 & n29193 ) ;
  assign n29204 = n28974 | n29193 ;
  assign n29206 = ( n29203 & ~n29205 ) | ( n29203 & n29204 ) | ( ~n29205 & n29204 ) ;
  assign n29210 = n28793 &  n29004 ;
  assign n29211 = n29003 &  n29210 ;
  assign n29199 = x86 | n28793 ;
  assign n29200 = x86 &  n28793 ;
  assign n29201 = ( n29199 & ~n29200 ) | ( n29199 & 1'b0 ) | ( ~n29200 & 1'b0 ) ;
  assign n29213 = ( n28973 & n29005 ) | ( n28973 & n29201 ) | ( n29005 & n29201 ) ;
  assign n29212 = n28973 | n29201 ;
  assign n29214 = ( n29211 & ~n29213 ) | ( n29211 & n29212 ) | ( ~n29213 & n29212 ) ;
  assign n29218 = n28801 &  n29004 ;
  assign n29219 = n29003 &  n29218 ;
  assign n29207 = x85 | n28801 ;
  assign n29208 = x85 &  n28801 ;
  assign n29209 = ( n29207 & ~n29208 ) | ( n29207 & 1'b0 ) | ( ~n29208 & 1'b0 ) ;
  assign n29221 = ( n28972 & n29005 ) | ( n28972 & n29209 ) | ( n29005 & n29209 ) ;
  assign n29220 = n28972 | n29209 ;
  assign n29222 = ( n29219 & ~n29221 ) | ( n29219 & n29220 ) | ( ~n29221 & n29220 ) ;
  assign n29226 = n28809 &  n29004 ;
  assign n29227 = n29003 &  n29226 ;
  assign n29215 = x84 | n28809 ;
  assign n29216 = x84 &  n28809 ;
  assign n29217 = ( n29215 & ~n29216 ) | ( n29215 & 1'b0 ) | ( ~n29216 & 1'b0 ) ;
  assign n29229 = ( n28971 & n29005 ) | ( n28971 & n29217 ) | ( n29005 & n29217 ) ;
  assign n29228 = n28971 | n29217 ;
  assign n29230 = ( n29227 & ~n29229 ) | ( n29227 & n29228 ) | ( ~n29229 & n29228 ) ;
  assign n29234 = n28817 &  n29004 ;
  assign n29235 = n29003 &  n29234 ;
  assign n29223 = x83 | n28817 ;
  assign n29224 = x83 &  n28817 ;
  assign n29225 = ( n29223 & ~n29224 ) | ( n29223 & 1'b0 ) | ( ~n29224 & 1'b0 ) ;
  assign n29237 = ( n28970 & n29005 ) | ( n28970 & n29225 ) | ( n29005 & n29225 ) ;
  assign n29236 = n28970 | n29225 ;
  assign n29238 = ( n29235 & ~n29237 ) | ( n29235 & n29236 ) | ( ~n29237 & n29236 ) ;
  assign n29242 = n28825 &  n29004 ;
  assign n29243 = n29003 &  n29242 ;
  assign n29231 = x82 | n28825 ;
  assign n29232 = x82 &  n28825 ;
  assign n29233 = ( n29231 & ~n29232 ) | ( n29231 & 1'b0 ) | ( ~n29232 & 1'b0 ) ;
  assign n29245 = ( n28969 & n29005 ) | ( n28969 & n29233 ) | ( n29005 & n29233 ) ;
  assign n29244 = n28969 | n29233 ;
  assign n29246 = ( n29243 & ~n29245 ) | ( n29243 & n29244 ) | ( ~n29245 & n29244 ) ;
  assign n29250 = n28833 &  n29004 ;
  assign n29251 = n29003 &  n29250 ;
  assign n29239 = x81 | n28833 ;
  assign n29240 = x81 &  n28833 ;
  assign n29241 = ( n29239 & ~n29240 ) | ( n29239 & 1'b0 ) | ( ~n29240 & 1'b0 ) ;
  assign n29253 = ( n28968 & n29005 ) | ( n28968 & n29241 ) | ( n29005 & n29241 ) ;
  assign n29252 = n28968 | n29241 ;
  assign n29254 = ( n29251 & ~n29253 ) | ( n29251 & n29252 ) | ( ~n29253 & n29252 ) ;
  assign n29258 = n28841 &  n29004 ;
  assign n29259 = n29003 &  n29258 ;
  assign n29247 = x80 | n28841 ;
  assign n29248 = x80 &  n28841 ;
  assign n29249 = ( n29247 & ~n29248 ) | ( n29247 & 1'b0 ) | ( ~n29248 & 1'b0 ) ;
  assign n29261 = ( n28967 & n29005 ) | ( n28967 & n29249 ) | ( n29005 & n29249 ) ;
  assign n29260 = n28967 | n29249 ;
  assign n29262 = ( n29259 & ~n29261 ) | ( n29259 & n29260 ) | ( ~n29261 & n29260 ) ;
  assign n29266 = n28849 &  n29004 ;
  assign n29267 = n29003 &  n29266 ;
  assign n29255 = x79 | n28849 ;
  assign n29256 = x79 &  n28849 ;
  assign n29257 = ( n29255 & ~n29256 ) | ( n29255 & 1'b0 ) | ( ~n29256 & 1'b0 ) ;
  assign n29269 = ( n28966 & n29005 ) | ( n28966 & n29257 ) | ( n29005 & n29257 ) ;
  assign n29268 = n28966 | n29257 ;
  assign n29270 = ( n29267 & ~n29269 ) | ( n29267 & n29268 ) | ( ~n29269 & n29268 ) ;
  assign n29274 = n28857 &  n29004 ;
  assign n29275 = n29003 &  n29274 ;
  assign n29263 = x78 | n28857 ;
  assign n29264 = x78 &  n28857 ;
  assign n29265 = ( n29263 & ~n29264 ) | ( n29263 & 1'b0 ) | ( ~n29264 & 1'b0 ) ;
  assign n29277 = ( n28965 & n29005 ) | ( n28965 & n29265 ) | ( n29005 & n29265 ) ;
  assign n29276 = n28965 | n29265 ;
  assign n29278 = ( n29275 & ~n29277 ) | ( n29275 & n29276 ) | ( ~n29277 & n29276 ) ;
  assign n29282 = n28865 &  n29004 ;
  assign n29283 = n29003 &  n29282 ;
  assign n29271 = x77 | n28865 ;
  assign n29272 = x77 &  n28865 ;
  assign n29273 = ( n29271 & ~n29272 ) | ( n29271 & 1'b0 ) | ( ~n29272 & 1'b0 ) ;
  assign n29285 = ( n28964 & n29005 ) | ( n28964 & n29273 ) | ( n29005 & n29273 ) ;
  assign n29284 = n28964 | n29273 ;
  assign n29286 = ( n29283 & ~n29285 ) | ( n29283 & n29284 ) | ( ~n29285 & n29284 ) ;
  assign n29290 = n28873 &  n29004 ;
  assign n29291 = n29003 &  n29290 ;
  assign n29279 = x76 | n28873 ;
  assign n29280 = x76 &  n28873 ;
  assign n29281 = ( n29279 & ~n29280 ) | ( n29279 & 1'b0 ) | ( ~n29280 & 1'b0 ) ;
  assign n29293 = ( n28963 & n29005 ) | ( n28963 & n29281 ) | ( n29005 & n29281 ) ;
  assign n29292 = n28963 | n29281 ;
  assign n29294 = ( n29291 & ~n29293 ) | ( n29291 & n29292 ) | ( ~n29293 & n29292 ) ;
  assign n29298 = n28881 &  n29004 ;
  assign n29299 = n29003 &  n29298 ;
  assign n29287 = x75 | n28881 ;
  assign n29288 = x75 &  n28881 ;
  assign n29289 = ( n29287 & ~n29288 ) | ( n29287 & 1'b0 ) | ( ~n29288 & 1'b0 ) ;
  assign n29301 = ( n28962 & n29005 ) | ( n28962 & n29289 ) | ( n29005 & n29289 ) ;
  assign n29300 = n28962 | n29289 ;
  assign n29302 = ( n29299 & ~n29301 ) | ( n29299 & n29300 ) | ( ~n29301 & n29300 ) ;
  assign n29306 = n28889 &  n29004 ;
  assign n29307 = n29003 &  n29306 ;
  assign n29295 = x74 | n28889 ;
  assign n29296 = x74 &  n28889 ;
  assign n29297 = ( n29295 & ~n29296 ) | ( n29295 & 1'b0 ) | ( ~n29296 & 1'b0 ) ;
  assign n29309 = ( n28961 & n29005 ) | ( n28961 & n29297 ) | ( n29005 & n29297 ) ;
  assign n29308 = n28961 | n29297 ;
  assign n29310 = ( n29307 & ~n29309 ) | ( n29307 & n29308 ) | ( ~n29309 & n29308 ) ;
  assign n29314 = n28897 &  n29004 ;
  assign n29315 = n29003 &  n29314 ;
  assign n29303 = x73 | n28897 ;
  assign n29304 = x73 &  n28897 ;
  assign n29305 = ( n29303 & ~n29304 ) | ( n29303 & 1'b0 ) | ( ~n29304 & 1'b0 ) ;
  assign n29317 = ( n28960 & n29005 ) | ( n28960 & n29305 ) | ( n29005 & n29305 ) ;
  assign n29316 = n28960 | n29305 ;
  assign n29318 = ( n29315 & ~n29317 ) | ( n29315 & n29316 ) | ( ~n29317 & n29316 ) ;
  assign n29322 = n28905 &  n29004 ;
  assign n29323 = n29003 &  n29322 ;
  assign n29311 = x72 | n28905 ;
  assign n29312 = x72 &  n28905 ;
  assign n29313 = ( n29311 & ~n29312 ) | ( n29311 & 1'b0 ) | ( ~n29312 & 1'b0 ) ;
  assign n29325 = ( n28959 & n29005 ) | ( n28959 & n29313 ) | ( n29005 & n29313 ) ;
  assign n29324 = n28959 | n29313 ;
  assign n29326 = ( n29323 & ~n29325 ) | ( n29323 & n29324 ) | ( ~n29325 & n29324 ) ;
  assign n29330 = n28913 &  n29004 ;
  assign n29331 = n29003 &  n29330 ;
  assign n29319 = x71 | n28913 ;
  assign n29320 = x71 &  n28913 ;
  assign n29321 = ( n29319 & ~n29320 ) | ( n29319 & 1'b0 ) | ( ~n29320 & 1'b0 ) ;
  assign n29333 = ( n28958 & n29005 ) | ( n28958 & n29321 ) | ( n29005 & n29321 ) ;
  assign n29332 = n28958 | n29321 ;
  assign n29334 = ( n29331 & ~n29333 ) | ( n29331 & n29332 ) | ( ~n29333 & n29332 ) ;
  assign n29338 = n28921 &  n29004 ;
  assign n29339 = n29003 &  n29338 ;
  assign n29327 = x70 | n28921 ;
  assign n29328 = x70 &  n28921 ;
  assign n29329 = ( n29327 & ~n29328 ) | ( n29327 & 1'b0 ) | ( ~n29328 & 1'b0 ) ;
  assign n29341 = ( n28957 & n29005 ) | ( n28957 & n29329 ) | ( n29005 & n29329 ) ;
  assign n29340 = n28957 | n29329 ;
  assign n29342 = ( n29339 & ~n29341 ) | ( n29339 & n29340 ) | ( ~n29341 & n29340 ) ;
  assign n29346 = n28929 &  n29004 ;
  assign n29347 = n29003 &  n29346 ;
  assign n29335 = x69 | n28929 ;
  assign n29336 = x69 &  n28929 ;
  assign n29337 = ( n29335 & ~n29336 ) | ( n29335 & 1'b0 ) | ( ~n29336 & 1'b0 ) ;
  assign n29349 = ( n28956 & n29005 ) | ( n28956 & n29337 ) | ( n29005 & n29337 ) ;
  assign n29348 = n28956 | n29337 ;
  assign n29350 = ( n29347 & ~n29349 ) | ( n29347 & n29348 ) | ( ~n29349 & n29348 ) ;
  assign n29354 = n28937 &  n29004 ;
  assign n29355 = n29003 &  n29354 ;
  assign n29343 = x68 | n28937 ;
  assign n29344 = x68 &  n28937 ;
  assign n29345 = ( n29343 & ~n29344 ) | ( n29343 & 1'b0 ) | ( ~n29344 & 1'b0 ) ;
  assign n29357 = ( n28955 & n29005 ) | ( n28955 & n29345 ) | ( n29005 & n29345 ) ;
  assign n29356 = n28955 | n29345 ;
  assign n29358 = ( n29355 & ~n29357 ) | ( n29355 & n29356 ) | ( ~n29357 & n29356 ) ;
  assign n29362 = n28942 &  n29004 ;
  assign n29363 = n29003 &  n29362 ;
  assign n29351 = x67 | n28942 ;
  assign n29352 = x67 &  n28942 ;
  assign n29353 = ( n29351 & ~n29352 ) | ( n29351 & 1'b0 ) | ( ~n29352 & 1'b0 ) ;
  assign n29365 = ( n28954 & n29005 ) | ( n28954 & n29353 ) | ( n29005 & n29353 ) ;
  assign n29364 = n28954 | n29353 ;
  assign n29366 = ( n29363 & ~n29365 ) | ( n29363 & n29364 ) | ( ~n29365 & n29364 ) ;
  assign n29367 = n28948 &  n29004 ;
  assign n29368 = n29003 &  n29367 ;
  assign n29359 = x66 | n28948 ;
  assign n29360 = x66 &  n28948 ;
  assign n29361 = ( n29359 & ~n29360 ) | ( n29359 & 1'b0 ) | ( ~n29360 & 1'b0 ) ;
  assign n29369 = n28953 &  n29361 ;
  assign n29370 = ( n28953 & ~n29005 ) | ( n28953 & n29361 ) | ( ~n29005 & n29361 ) ;
  assign n29371 = ( n29368 & ~n29369 ) | ( n29368 & n29370 ) | ( ~n29369 & n29370 ) ;
  assign n29372 = ( x65 & ~n10539 ) | ( x65 & n28952 ) | ( ~n10539 & n28952 ) ;
  assign n29373 = ( n28953 & ~x65 ) | ( n28953 & n29372 ) | ( ~x65 & n29372 ) ;
  assign n29374 = ~n29005 & n29373 ;
  assign n29375 = n28952 &  n29004 ;
  assign n29376 = n29003 &  n29375 ;
  assign n29377 = n29374 | n29376 ;
  assign n29378 = ( x64 & ~n29005 ) | ( x64 & 1'b0 ) | ( ~n29005 & 1'b0 ) ;
  assign n29379 = ( x16 & ~n29378 ) | ( x16 & 1'b0 ) | ( ~n29378 & 1'b0 ) ;
  assign n29380 = ( n10539 & ~n29005 ) | ( n10539 & 1'b0 ) | ( ~n29005 & 1'b0 ) ;
  assign n29381 = n29379 | n29380 ;
  assign n29382 = ( x65 & ~n29381 ) | ( x65 & n11065 ) | ( ~n29381 & n11065 ) ;
  assign n29383 = ( x66 & ~n29377 ) | ( x66 & n29382 ) | ( ~n29377 & n29382 ) ;
  assign n29384 = ( x67 & ~n29371 ) | ( x67 & n29383 ) | ( ~n29371 & n29383 ) ;
  assign n29385 = ( x68 & ~n29366 ) | ( x68 & n29384 ) | ( ~n29366 & n29384 ) ;
  assign n29386 = ( x69 & ~n29358 ) | ( x69 & n29385 ) | ( ~n29358 & n29385 ) ;
  assign n29387 = ( x70 & ~n29350 ) | ( x70 & n29386 ) | ( ~n29350 & n29386 ) ;
  assign n29388 = ( x71 & ~n29342 ) | ( x71 & n29387 ) | ( ~n29342 & n29387 ) ;
  assign n29389 = ( x72 & ~n29334 ) | ( x72 & n29388 ) | ( ~n29334 & n29388 ) ;
  assign n29390 = ( x73 & ~n29326 ) | ( x73 & n29389 ) | ( ~n29326 & n29389 ) ;
  assign n29391 = ( x74 & ~n29318 ) | ( x74 & n29390 ) | ( ~n29318 & n29390 ) ;
  assign n29392 = ( x75 & ~n29310 ) | ( x75 & n29391 ) | ( ~n29310 & n29391 ) ;
  assign n29393 = ( x76 & ~n29302 ) | ( x76 & n29392 ) | ( ~n29302 & n29392 ) ;
  assign n29394 = ( x77 & ~n29294 ) | ( x77 & n29393 ) | ( ~n29294 & n29393 ) ;
  assign n29395 = ( x78 & ~n29286 ) | ( x78 & n29394 ) | ( ~n29286 & n29394 ) ;
  assign n29396 = ( x79 & ~n29278 ) | ( x79 & n29395 ) | ( ~n29278 & n29395 ) ;
  assign n29397 = ( x80 & ~n29270 ) | ( x80 & n29396 ) | ( ~n29270 & n29396 ) ;
  assign n29398 = ( x81 & ~n29262 ) | ( x81 & n29397 ) | ( ~n29262 & n29397 ) ;
  assign n29399 = ( x82 & ~n29254 ) | ( x82 & n29398 ) | ( ~n29254 & n29398 ) ;
  assign n29400 = ( x83 & ~n29246 ) | ( x83 & n29399 ) | ( ~n29246 & n29399 ) ;
  assign n29401 = ( x84 & ~n29238 ) | ( x84 & n29400 ) | ( ~n29238 & n29400 ) ;
  assign n29402 = ( x85 & ~n29230 ) | ( x85 & n29401 ) | ( ~n29230 & n29401 ) ;
  assign n29403 = ( x86 & ~n29222 ) | ( x86 & n29402 ) | ( ~n29222 & n29402 ) ;
  assign n29404 = ( x87 & ~n29214 ) | ( x87 & n29403 ) | ( ~n29214 & n29403 ) ;
  assign n29405 = ( x88 & ~n29206 ) | ( x88 & n29404 ) | ( ~n29206 & n29404 ) ;
  assign n29406 = ( x89 & ~n29198 ) | ( x89 & n29405 ) | ( ~n29198 & n29405 ) ;
  assign n29407 = ( x90 & ~n29190 ) | ( x90 & n29406 ) | ( ~n29190 & n29406 ) ;
  assign n29408 = ( x91 & ~n29182 ) | ( x91 & n29407 ) | ( ~n29182 & n29407 ) ;
  assign n29409 = ( x92 & ~n29174 ) | ( x92 & n29408 ) | ( ~n29174 & n29408 ) ;
  assign n29410 = ( x93 & ~n29166 ) | ( x93 & n29409 ) | ( ~n29166 & n29409 ) ;
  assign n29411 = ( x94 & ~n29158 ) | ( x94 & n29410 ) | ( ~n29158 & n29410 ) ;
  assign n29412 = ( x95 & ~n29150 ) | ( x95 & n29411 ) | ( ~n29150 & n29411 ) ;
  assign n29413 = ( x96 & ~n29142 ) | ( x96 & n29412 ) | ( ~n29142 & n29412 ) ;
  assign n29414 = ( x97 & ~n29134 ) | ( x97 & n29413 ) | ( ~n29134 & n29413 ) ;
  assign n29415 = ( x98 & ~n29126 ) | ( x98 & n29414 ) | ( ~n29126 & n29414 ) ;
  assign n29416 = ( x99 & ~n29118 ) | ( x99 & n29415 ) | ( ~n29118 & n29415 ) ;
  assign n29417 = ( x100 & ~n29110 ) | ( x100 & n29416 ) | ( ~n29110 & n29416 ) ;
  assign n29418 = ( x101 & ~n29102 ) | ( x101 & n29417 ) | ( ~n29102 & n29417 ) ;
  assign n29419 = ( x102 & ~n29094 ) | ( x102 & n29418 ) | ( ~n29094 & n29418 ) ;
  assign n29420 = ( x103 & ~n29086 ) | ( x103 & n29419 ) | ( ~n29086 & n29419 ) ;
  assign n29421 = ( x104 & ~n29078 ) | ( x104 & n29420 ) | ( ~n29078 & n29420 ) ;
  assign n29422 = ( x105 & ~n29070 ) | ( x105 & n29421 ) | ( ~n29070 & n29421 ) ;
  assign n29423 = ( x106 & ~n29062 ) | ( x106 & n29422 ) | ( ~n29062 & n29422 ) ;
  assign n29424 = ( x107 & ~n29054 ) | ( x107 & n29423 ) | ( ~n29054 & n29423 ) ;
  assign n29425 = ( x108 & ~n29046 ) | ( x108 & n29424 ) | ( ~n29046 & n29424 ) ;
  assign n29426 = ( x109 & ~n29038 ) | ( x109 & n29425 ) | ( ~n29038 & n29425 ) ;
  assign n29427 = ( x110 & ~n29030 ) | ( x110 & n29426 ) | ( ~n29030 & n29426 ) ;
  assign n29428 = ( x111 & ~n29022 ) | ( x111 & n29427 ) | ( ~n29022 & n29427 ) ;
  assign n29429 = ( x112 & ~n29014 ) | ( x112 & n29428 ) | ( ~n29014 & n29428 ) ;
  assign n29430 = n240 | n29429 ;
  assign n29440 = n29022 &  n29430 ;
  assign n29432 = x111 | n29022 ;
  assign n29433 = x111 &  n29022 ;
  assign n29434 = ( n29432 & ~n29433 ) | ( n29432 & 1'b0 ) | ( ~n29433 & 1'b0 ) ;
  assign n29444 = ( n240 & n29427 ) | ( n240 & n29434 ) | ( n29427 & n29434 ) ;
  assign n29445 = ( n29427 & ~n29429 ) | ( n29427 & n29434 ) | ( ~n29429 & n29434 ) ;
  assign n29446 = ~n29444 & n29445 ;
  assign n29447 = n29440 | n29446 ;
  assign n29448 = n29030 &  n29430 ;
  assign n29441 = x110 | n29030 ;
  assign n29442 = x110 &  n29030 ;
  assign n29443 = ( n29441 & ~n29442 ) | ( n29441 & 1'b0 ) | ( ~n29442 & 1'b0 ) ;
  assign n29452 = ( n240 & n29426 ) | ( n240 & n29443 ) | ( n29426 & n29443 ) ;
  assign n29453 = ( n29426 & ~n29429 ) | ( n29426 & n29443 ) | ( ~n29429 & n29443 ) ;
  assign n29454 = ~n29452 & n29453 ;
  assign n29455 = n29448 | n29454 ;
  assign n29456 = n29038 &  n29430 ;
  assign n29449 = x109 | n29038 ;
  assign n29450 = x109 &  n29038 ;
  assign n29451 = ( n29449 & ~n29450 ) | ( n29449 & 1'b0 ) | ( ~n29450 & 1'b0 ) ;
  assign n29460 = ( n240 & n29425 ) | ( n240 & n29451 ) | ( n29425 & n29451 ) ;
  assign n29461 = ( n29425 & ~n29429 ) | ( n29425 & n29451 ) | ( ~n29429 & n29451 ) ;
  assign n29462 = ~n29460 & n29461 ;
  assign n29463 = n29456 | n29462 ;
  assign n29464 = n29046 &  n29430 ;
  assign n29457 = x108 | n29046 ;
  assign n29458 = x108 &  n29046 ;
  assign n29459 = ( n29457 & ~n29458 ) | ( n29457 & 1'b0 ) | ( ~n29458 & 1'b0 ) ;
  assign n29468 = ( n240 & n29424 ) | ( n240 & n29459 ) | ( n29424 & n29459 ) ;
  assign n29469 = ( n29424 & ~n29429 ) | ( n29424 & n29459 ) | ( ~n29429 & n29459 ) ;
  assign n29470 = ~n29468 & n29469 ;
  assign n29471 = n29464 | n29470 ;
  assign n29472 = n29054 &  n29430 ;
  assign n29465 = x107 | n29054 ;
  assign n29466 = x107 &  n29054 ;
  assign n29467 = ( n29465 & ~n29466 ) | ( n29465 & 1'b0 ) | ( ~n29466 & 1'b0 ) ;
  assign n29476 = ( n240 & n29423 ) | ( n240 & n29467 ) | ( n29423 & n29467 ) ;
  assign n29477 = ( n29423 & ~n29429 ) | ( n29423 & n29467 ) | ( ~n29429 & n29467 ) ;
  assign n29478 = ~n29476 & n29477 ;
  assign n29479 = n29472 | n29478 ;
  assign n29480 = n29062 &  n29430 ;
  assign n29473 = x106 | n29062 ;
  assign n29474 = x106 &  n29062 ;
  assign n29475 = ( n29473 & ~n29474 ) | ( n29473 & 1'b0 ) | ( ~n29474 & 1'b0 ) ;
  assign n29484 = ( n240 & n29422 ) | ( n240 & n29475 ) | ( n29422 & n29475 ) ;
  assign n29485 = ( n29422 & ~n29429 ) | ( n29422 & n29475 ) | ( ~n29429 & n29475 ) ;
  assign n29486 = ~n29484 & n29485 ;
  assign n29487 = n29480 | n29486 ;
  assign n29488 = n29070 &  n29430 ;
  assign n29481 = x105 | n29070 ;
  assign n29482 = x105 &  n29070 ;
  assign n29483 = ( n29481 & ~n29482 ) | ( n29481 & 1'b0 ) | ( ~n29482 & 1'b0 ) ;
  assign n29492 = ( n240 & n29421 ) | ( n240 & n29483 ) | ( n29421 & n29483 ) ;
  assign n29493 = ( n29421 & ~n29429 ) | ( n29421 & n29483 ) | ( ~n29429 & n29483 ) ;
  assign n29494 = ~n29492 & n29493 ;
  assign n29495 = n29488 | n29494 ;
  assign n29496 = n29078 &  n29430 ;
  assign n29489 = x104 | n29078 ;
  assign n29490 = x104 &  n29078 ;
  assign n29491 = ( n29489 & ~n29490 ) | ( n29489 & 1'b0 ) | ( ~n29490 & 1'b0 ) ;
  assign n29500 = ( n240 & n29420 ) | ( n240 & n29491 ) | ( n29420 & n29491 ) ;
  assign n29501 = ( n29420 & ~n29429 ) | ( n29420 & n29491 ) | ( ~n29429 & n29491 ) ;
  assign n29502 = ~n29500 & n29501 ;
  assign n29503 = n29496 | n29502 ;
  assign n29504 = n29086 &  n29430 ;
  assign n29497 = x103 | n29086 ;
  assign n29498 = x103 &  n29086 ;
  assign n29499 = ( n29497 & ~n29498 ) | ( n29497 & 1'b0 ) | ( ~n29498 & 1'b0 ) ;
  assign n29508 = ( n240 & n29419 ) | ( n240 & n29499 ) | ( n29419 & n29499 ) ;
  assign n29509 = ( n29419 & ~n29429 ) | ( n29419 & n29499 ) | ( ~n29429 & n29499 ) ;
  assign n29510 = ~n29508 & n29509 ;
  assign n29511 = n29504 | n29510 ;
  assign n29512 = n29094 &  n29430 ;
  assign n29505 = x102 | n29094 ;
  assign n29506 = x102 &  n29094 ;
  assign n29507 = ( n29505 & ~n29506 ) | ( n29505 & 1'b0 ) | ( ~n29506 & 1'b0 ) ;
  assign n29516 = ( n240 & n29418 ) | ( n240 & n29507 ) | ( n29418 & n29507 ) ;
  assign n29517 = ( n29418 & ~n29429 ) | ( n29418 & n29507 ) | ( ~n29429 & n29507 ) ;
  assign n29518 = ~n29516 & n29517 ;
  assign n29519 = n29512 | n29518 ;
  assign n29520 = n29102 &  n29430 ;
  assign n29513 = x101 | n29102 ;
  assign n29514 = x101 &  n29102 ;
  assign n29515 = ( n29513 & ~n29514 ) | ( n29513 & 1'b0 ) | ( ~n29514 & 1'b0 ) ;
  assign n29524 = ( n240 & n29417 ) | ( n240 & n29515 ) | ( n29417 & n29515 ) ;
  assign n29525 = ( n29417 & ~n29429 ) | ( n29417 & n29515 ) | ( ~n29429 & n29515 ) ;
  assign n29526 = ~n29524 & n29525 ;
  assign n29527 = n29520 | n29526 ;
  assign n29528 = n29110 &  n29430 ;
  assign n29521 = x100 | n29110 ;
  assign n29522 = x100 &  n29110 ;
  assign n29523 = ( n29521 & ~n29522 ) | ( n29521 & 1'b0 ) | ( ~n29522 & 1'b0 ) ;
  assign n29532 = ( n240 & n29416 ) | ( n240 & n29523 ) | ( n29416 & n29523 ) ;
  assign n29533 = ( n29416 & ~n29429 ) | ( n29416 & n29523 ) | ( ~n29429 & n29523 ) ;
  assign n29534 = ~n29532 & n29533 ;
  assign n29535 = n29528 | n29534 ;
  assign n29536 = n29118 &  n29430 ;
  assign n29529 = x99 | n29118 ;
  assign n29530 = x99 &  n29118 ;
  assign n29531 = ( n29529 & ~n29530 ) | ( n29529 & 1'b0 ) | ( ~n29530 & 1'b0 ) ;
  assign n29540 = ( n240 & n29415 ) | ( n240 & n29531 ) | ( n29415 & n29531 ) ;
  assign n29541 = ( n29415 & ~n29429 ) | ( n29415 & n29531 ) | ( ~n29429 & n29531 ) ;
  assign n29542 = ~n29540 & n29541 ;
  assign n29543 = n29536 | n29542 ;
  assign n29544 = n29126 &  n29430 ;
  assign n29537 = x98 | n29126 ;
  assign n29538 = x98 &  n29126 ;
  assign n29539 = ( n29537 & ~n29538 ) | ( n29537 & 1'b0 ) | ( ~n29538 & 1'b0 ) ;
  assign n29548 = ( n240 & n29414 ) | ( n240 & n29539 ) | ( n29414 & n29539 ) ;
  assign n29549 = ( n29414 & ~n29429 ) | ( n29414 & n29539 ) | ( ~n29429 & n29539 ) ;
  assign n29550 = ~n29548 & n29549 ;
  assign n29551 = n29544 | n29550 ;
  assign n29552 = n29134 &  n29430 ;
  assign n29545 = x97 | n29134 ;
  assign n29546 = x97 &  n29134 ;
  assign n29547 = ( n29545 & ~n29546 ) | ( n29545 & 1'b0 ) | ( ~n29546 & 1'b0 ) ;
  assign n29556 = ( n240 & n29413 ) | ( n240 & n29547 ) | ( n29413 & n29547 ) ;
  assign n29557 = ( n29413 & ~n29429 ) | ( n29413 & n29547 ) | ( ~n29429 & n29547 ) ;
  assign n29558 = ~n29556 & n29557 ;
  assign n29559 = n29552 | n29558 ;
  assign n29560 = n29142 &  n29430 ;
  assign n29553 = x96 | n29142 ;
  assign n29554 = x96 &  n29142 ;
  assign n29555 = ( n29553 & ~n29554 ) | ( n29553 & 1'b0 ) | ( ~n29554 & 1'b0 ) ;
  assign n29564 = ( n240 & n29412 ) | ( n240 & n29555 ) | ( n29412 & n29555 ) ;
  assign n29565 = ( n29412 & ~n29429 ) | ( n29412 & n29555 ) | ( ~n29429 & n29555 ) ;
  assign n29566 = ~n29564 & n29565 ;
  assign n29567 = n29560 | n29566 ;
  assign n29568 = n29150 &  n29430 ;
  assign n29561 = x95 | n29150 ;
  assign n29562 = x95 &  n29150 ;
  assign n29563 = ( n29561 & ~n29562 ) | ( n29561 & 1'b0 ) | ( ~n29562 & 1'b0 ) ;
  assign n29572 = ( n240 & n29411 ) | ( n240 & n29563 ) | ( n29411 & n29563 ) ;
  assign n29573 = ( n29411 & ~n29429 ) | ( n29411 & n29563 ) | ( ~n29429 & n29563 ) ;
  assign n29574 = ~n29572 & n29573 ;
  assign n29575 = n29568 | n29574 ;
  assign n29576 = n29158 &  n29430 ;
  assign n29569 = x94 | n29158 ;
  assign n29570 = x94 &  n29158 ;
  assign n29571 = ( n29569 & ~n29570 ) | ( n29569 & 1'b0 ) | ( ~n29570 & 1'b0 ) ;
  assign n29580 = ( n240 & n29410 ) | ( n240 & n29571 ) | ( n29410 & n29571 ) ;
  assign n29581 = ( n29410 & ~n29429 ) | ( n29410 & n29571 ) | ( ~n29429 & n29571 ) ;
  assign n29582 = ~n29580 & n29581 ;
  assign n29583 = n29576 | n29582 ;
  assign n29584 = n29166 &  n29430 ;
  assign n29577 = x93 | n29166 ;
  assign n29578 = x93 &  n29166 ;
  assign n29579 = ( n29577 & ~n29578 ) | ( n29577 & 1'b0 ) | ( ~n29578 & 1'b0 ) ;
  assign n29588 = ( n240 & n29409 ) | ( n240 & n29579 ) | ( n29409 & n29579 ) ;
  assign n29589 = ( n29409 & ~n29429 ) | ( n29409 & n29579 ) | ( ~n29429 & n29579 ) ;
  assign n29590 = ~n29588 & n29589 ;
  assign n29591 = n29584 | n29590 ;
  assign n29592 = n29174 &  n29430 ;
  assign n29585 = x92 | n29174 ;
  assign n29586 = x92 &  n29174 ;
  assign n29587 = ( n29585 & ~n29586 ) | ( n29585 & 1'b0 ) | ( ~n29586 & 1'b0 ) ;
  assign n29596 = ( n240 & n29408 ) | ( n240 & n29587 ) | ( n29408 & n29587 ) ;
  assign n29597 = ( n29408 & ~n29429 ) | ( n29408 & n29587 ) | ( ~n29429 & n29587 ) ;
  assign n29598 = ~n29596 & n29597 ;
  assign n29599 = n29592 | n29598 ;
  assign n29600 = n29182 &  n29430 ;
  assign n29593 = x91 | n29182 ;
  assign n29594 = x91 &  n29182 ;
  assign n29595 = ( n29593 & ~n29594 ) | ( n29593 & 1'b0 ) | ( ~n29594 & 1'b0 ) ;
  assign n29604 = ( n240 & n29407 ) | ( n240 & n29595 ) | ( n29407 & n29595 ) ;
  assign n29605 = ( n29407 & ~n29429 ) | ( n29407 & n29595 ) | ( ~n29429 & n29595 ) ;
  assign n29606 = ~n29604 & n29605 ;
  assign n29607 = n29600 | n29606 ;
  assign n29608 = n29190 &  n29430 ;
  assign n29601 = x90 | n29190 ;
  assign n29602 = x90 &  n29190 ;
  assign n29603 = ( n29601 & ~n29602 ) | ( n29601 & 1'b0 ) | ( ~n29602 & 1'b0 ) ;
  assign n29612 = ( n240 & n29406 ) | ( n240 & n29603 ) | ( n29406 & n29603 ) ;
  assign n29613 = ( n29406 & ~n29429 ) | ( n29406 & n29603 ) | ( ~n29429 & n29603 ) ;
  assign n29614 = ~n29612 & n29613 ;
  assign n29615 = n29608 | n29614 ;
  assign n29616 = n29198 &  n29430 ;
  assign n29609 = x89 | n29198 ;
  assign n29610 = x89 &  n29198 ;
  assign n29611 = ( n29609 & ~n29610 ) | ( n29609 & 1'b0 ) | ( ~n29610 & 1'b0 ) ;
  assign n29620 = ( n240 & n29405 ) | ( n240 & n29611 ) | ( n29405 & n29611 ) ;
  assign n29621 = ( n29405 & ~n29429 ) | ( n29405 & n29611 ) | ( ~n29429 & n29611 ) ;
  assign n29622 = ~n29620 & n29621 ;
  assign n29623 = n29616 | n29622 ;
  assign n29624 = n29206 &  n29430 ;
  assign n29617 = x88 | n29206 ;
  assign n29618 = x88 &  n29206 ;
  assign n29619 = ( n29617 & ~n29618 ) | ( n29617 & 1'b0 ) | ( ~n29618 & 1'b0 ) ;
  assign n29628 = ( n240 & n29404 ) | ( n240 & n29619 ) | ( n29404 & n29619 ) ;
  assign n29629 = ( n29404 & ~n29429 ) | ( n29404 & n29619 ) | ( ~n29429 & n29619 ) ;
  assign n29630 = ~n29628 & n29629 ;
  assign n29631 = n29624 | n29630 ;
  assign n29632 = n29214 &  n29430 ;
  assign n29625 = x87 | n29214 ;
  assign n29626 = x87 &  n29214 ;
  assign n29627 = ( n29625 & ~n29626 ) | ( n29625 & 1'b0 ) | ( ~n29626 & 1'b0 ) ;
  assign n29636 = ( n240 & n29403 ) | ( n240 & n29627 ) | ( n29403 & n29627 ) ;
  assign n29637 = ( n29403 & ~n29429 ) | ( n29403 & n29627 ) | ( ~n29429 & n29627 ) ;
  assign n29638 = ~n29636 & n29637 ;
  assign n29639 = n29632 | n29638 ;
  assign n29640 = n29222 &  n29430 ;
  assign n29633 = x86 | n29222 ;
  assign n29634 = x86 &  n29222 ;
  assign n29635 = ( n29633 & ~n29634 ) | ( n29633 & 1'b0 ) | ( ~n29634 & 1'b0 ) ;
  assign n29644 = ( n240 & n29402 ) | ( n240 & n29635 ) | ( n29402 & n29635 ) ;
  assign n29645 = ( n29402 & ~n29429 ) | ( n29402 & n29635 ) | ( ~n29429 & n29635 ) ;
  assign n29646 = ~n29644 & n29645 ;
  assign n29647 = n29640 | n29646 ;
  assign n29648 = n29230 &  n29430 ;
  assign n29641 = x85 | n29230 ;
  assign n29642 = x85 &  n29230 ;
  assign n29643 = ( n29641 & ~n29642 ) | ( n29641 & 1'b0 ) | ( ~n29642 & 1'b0 ) ;
  assign n29652 = ( n240 & n29401 ) | ( n240 & n29643 ) | ( n29401 & n29643 ) ;
  assign n29653 = ( n29401 & ~n29429 ) | ( n29401 & n29643 ) | ( ~n29429 & n29643 ) ;
  assign n29654 = ~n29652 & n29653 ;
  assign n29655 = n29648 | n29654 ;
  assign n29656 = n29238 &  n29430 ;
  assign n29649 = x84 | n29238 ;
  assign n29650 = x84 &  n29238 ;
  assign n29651 = ( n29649 & ~n29650 ) | ( n29649 & 1'b0 ) | ( ~n29650 & 1'b0 ) ;
  assign n29660 = ( n240 & n29400 ) | ( n240 & n29651 ) | ( n29400 & n29651 ) ;
  assign n29661 = ( n29400 & ~n29429 ) | ( n29400 & n29651 ) | ( ~n29429 & n29651 ) ;
  assign n29662 = ~n29660 & n29661 ;
  assign n29663 = n29656 | n29662 ;
  assign n29664 = n29246 &  n29430 ;
  assign n29657 = x83 | n29246 ;
  assign n29658 = x83 &  n29246 ;
  assign n29659 = ( n29657 & ~n29658 ) | ( n29657 & 1'b0 ) | ( ~n29658 & 1'b0 ) ;
  assign n29668 = ( n240 & n29399 ) | ( n240 & n29659 ) | ( n29399 & n29659 ) ;
  assign n29669 = ( n29399 & ~n29429 ) | ( n29399 & n29659 ) | ( ~n29429 & n29659 ) ;
  assign n29670 = ~n29668 & n29669 ;
  assign n29671 = n29664 | n29670 ;
  assign n29672 = n29254 &  n29430 ;
  assign n29665 = x82 | n29254 ;
  assign n29666 = x82 &  n29254 ;
  assign n29667 = ( n29665 & ~n29666 ) | ( n29665 & 1'b0 ) | ( ~n29666 & 1'b0 ) ;
  assign n29676 = ( n240 & n29398 ) | ( n240 & n29667 ) | ( n29398 & n29667 ) ;
  assign n29677 = ( n29398 & ~n29429 ) | ( n29398 & n29667 ) | ( ~n29429 & n29667 ) ;
  assign n29678 = ~n29676 & n29677 ;
  assign n29679 = n29672 | n29678 ;
  assign n29680 = n29262 &  n29430 ;
  assign n29673 = x81 | n29262 ;
  assign n29674 = x81 &  n29262 ;
  assign n29675 = ( n29673 & ~n29674 ) | ( n29673 & 1'b0 ) | ( ~n29674 & 1'b0 ) ;
  assign n29684 = ( n240 & n29397 ) | ( n240 & n29675 ) | ( n29397 & n29675 ) ;
  assign n29685 = ( n29397 & ~n29429 ) | ( n29397 & n29675 ) | ( ~n29429 & n29675 ) ;
  assign n29686 = ~n29684 & n29685 ;
  assign n29687 = n29680 | n29686 ;
  assign n29688 = n29270 &  n29430 ;
  assign n29681 = x80 | n29270 ;
  assign n29682 = x80 &  n29270 ;
  assign n29683 = ( n29681 & ~n29682 ) | ( n29681 & 1'b0 ) | ( ~n29682 & 1'b0 ) ;
  assign n29692 = ( n240 & n29396 ) | ( n240 & n29683 ) | ( n29396 & n29683 ) ;
  assign n29693 = ( n29396 & ~n29429 ) | ( n29396 & n29683 ) | ( ~n29429 & n29683 ) ;
  assign n29694 = ~n29692 & n29693 ;
  assign n29695 = n29688 | n29694 ;
  assign n29696 = n29278 &  n29430 ;
  assign n29689 = x79 | n29278 ;
  assign n29690 = x79 &  n29278 ;
  assign n29691 = ( n29689 & ~n29690 ) | ( n29689 & 1'b0 ) | ( ~n29690 & 1'b0 ) ;
  assign n29700 = ( n240 & n29395 ) | ( n240 & n29691 ) | ( n29395 & n29691 ) ;
  assign n29701 = ( n29395 & ~n29429 ) | ( n29395 & n29691 ) | ( ~n29429 & n29691 ) ;
  assign n29702 = ~n29700 & n29701 ;
  assign n29703 = n29696 | n29702 ;
  assign n29704 = n29286 &  n29430 ;
  assign n29697 = x78 | n29286 ;
  assign n29698 = x78 &  n29286 ;
  assign n29699 = ( n29697 & ~n29698 ) | ( n29697 & 1'b0 ) | ( ~n29698 & 1'b0 ) ;
  assign n29708 = ( n240 & n29394 ) | ( n240 & n29699 ) | ( n29394 & n29699 ) ;
  assign n29709 = ( n29394 & ~n29429 ) | ( n29394 & n29699 ) | ( ~n29429 & n29699 ) ;
  assign n29710 = ~n29708 & n29709 ;
  assign n29711 = n29704 | n29710 ;
  assign n29712 = n29294 &  n29430 ;
  assign n29705 = x77 | n29294 ;
  assign n29706 = x77 &  n29294 ;
  assign n29707 = ( n29705 & ~n29706 ) | ( n29705 & 1'b0 ) | ( ~n29706 & 1'b0 ) ;
  assign n29716 = ( n240 & n29393 ) | ( n240 & n29707 ) | ( n29393 & n29707 ) ;
  assign n29717 = ( n29393 & ~n29429 ) | ( n29393 & n29707 ) | ( ~n29429 & n29707 ) ;
  assign n29718 = ~n29716 & n29717 ;
  assign n29719 = n29712 | n29718 ;
  assign n29720 = n29302 &  n29430 ;
  assign n29713 = x76 | n29302 ;
  assign n29714 = x76 &  n29302 ;
  assign n29715 = ( n29713 & ~n29714 ) | ( n29713 & 1'b0 ) | ( ~n29714 & 1'b0 ) ;
  assign n29724 = ( n240 & n29392 ) | ( n240 & n29715 ) | ( n29392 & n29715 ) ;
  assign n29725 = ( n29392 & ~n29429 ) | ( n29392 & n29715 ) | ( ~n29429 & n29715 ) ;
  assign n29726 = ~n29724 & n29725 ;
  assign n29727 = n29720 | n29726 ;
  assign n29728 = n29310 &  n29430 ;
  assign n29721 = x75 | n29310 ;
  assign n29722 = x75 &  n29310 ;
  assign n29723 = ( n29721 & ~n29722 ) | ( n29721 & 1'b0 ) | ( ~n29722 & 1'b0 ) ;
  assign n29732 = ( n240 & n29391 ) | ( n240 & n29723 ) | ( n29391 & n29723 ) ;
  assign n29733 = ( n29391 & ~n29429 ) | ( n29391 & n29723 ) | ( ~n29429 & n29723 ) ;
  assign n29734 = ~n29732 & n29733 ;
  assign n29735 = n29728 | n29734 ;
  assign n29736 = n29318 &  n29430 ;
  assign n29729 = x74 | n29318 ;
  assign n29730 = x74 &  n29318 ;
  assign n29731 = ( n29729 & ~n29730 ) | ( n29729 & 1'b0 ) | ( ~n29730 & 1'b0 ) ;
  assign n29740 = ( n240 & n29390 ) | ( n240 & n29731 ) | ( n29390 & n29731 ) ;
  assign n29741 = ( n29390 & ~n29429 ) | ( n29390 & n29731 ) | ( ~n29429 & n29731 ) ;
  assign n29742 = ~n29740 & n29741 ;
  assign n29743 = n29736 | n29742 ;
  assign n29744 = n29326 &  n29430 ;
  assign n29737 = x73 | n29326 ;
  assign n29738 = x73 &  n29326 ;
  assign n29739 = ( n29737 & ~n29738 ) | ( n29737 & 1'b0 ) | ( ~n29738 & 1'b0 ) ;
  assign n29748 = ( n240 & n29389 ) | ( n240 & n29739 ) | ( n29389 & n29739 ) ;
  assign n29749 = ( n29389 & ~n29429 ) | ( n29389 & n29739 ) | ( ~n29429 & n29739 ) ;
  assign n29750 = ~n29748 & n29749 ;
  assign n29751 = n29744 | n29750 ;
  assign n29752 = n29334 &  n29430 ;
  assign n29745 = x72 | n29334 ;
  assign n29746 = x72 &  n29334 ;
  assign n29747 = ( n29745 & ~n29746 ) | ( n29745 & 1'b0 ) | ( ~n29746 & 1'b0 ) ;
  assign n29756 = ( n240 & n29388 ) | ( n240 & n29747 ) | ( n29388 & n29747 ) ;
  assign n29757 = ( n29388 & ~n29429 ) | ( n29388 & n29747 ) | ( ~n29429 & n29747 ) ;
  assign n29758 = ~n29756 & n29757 ;
  assign n29759 = n29752 | n29758 ;
  assign n29760 = n29342 &  n29430 ;
  assign n29753 = x71 | n29342 ;
  assign n29754 = x71 &  n29342 ;
  assign n29755 = ( n29753 & ~n29754 ) | ( n29753 & 1'b0 ) | ( ~n29754 & 1'b0 ) ;
  assign n29764 = ( n240 & n29387 ) | ( n240 & n29755 ) | ( n29387 & n29755 ) ;
  assign n29765 = ( n29387 & ~n29429 ) | ( n29387 & n29755 ) | ( ~n29429 & n29755 ) ;
  assign n29766 = ~n29764 & n29765 ;
  assign n29767 = n29760 | n29766 ;
  assign n29768 = n29350 &  n29430 ;
  assign n29761 = x70 | n29350 ;
  assign n29762 = x70 &  n29350 ;
  assign n29763 = ( n29761 & ~n29762 ) | ( n29761 & 1'b0 ) | ( ~n29762 & 1'b0 ) ;
  assign n29772 = ( n240 & n29386 ) | ( n240 & n29763 ) | ( n29386 & n29763 ) ;
  assign n29773 = ( n29386 & ~n29429 ) | ( n29386 & n29763 ) | ( ~n29429 & n29763 ) ;
  assign n29774 = ~n29772 & n29773 ;
  assign n29775 = n29768 | n29774 ;
  assign n29776 = n29358 &  n29430 ;
  assign n29769 = x69 | n29358 ;
  assign n29770 = x69 &  n29358 ;
  assign n29771 = ( n29769 & ~n29770 ) | ( n29769 & 1'b0 ) | ( ~n29770 & 1'b0 ) ;
  assign n29780 = ( n240 & n29385 ) | ( n240 & n29771 ) | ( n29385 & n29771 ) ;
  assign n29781 = ( n29385 & ~n29429 ) | ( n29385 & n29771 ) | ( ~n29429 & n29771 ) ;
  assign n29782 = ~n29780 & n29781 ;
  assign n29783 = n29776 | n29782 ;
  assign n29784 = n29366 &  n29430 ;
  assign n29777 = x68 | n29366 ;
  assign n29778 = x68 &  n29366 ;
  assign n29779 = ( n29777 & ~n29778 ) | ( n29777 & 1'b0 ) | ( ~n29778 & 1'b0 ) ;
  assign n29788 = ( n240 & n29384 ) | ( n240 & n29779 ) | ( n29384 & n29779 ) ;
  assign n29789 = ( n29384 & ~n29429 ) | ( n29384 & n29779 ) | ( ~n29429 & n29779 ) ;
  assign n29790 = ~n29788 & n29789 ;
  assign n29791 = n29784 | n29790 ;
  assign n29792 = n29371 &  n29430 ;
  assign n29785 = x67 | n29371 ;
  assign n29786 = x67 &  n29371 ;
  assign n29787 = ( n29785 & ~n29786 ) | ( n29785 & 1'b0 ) | ( ~n29786 & 1'b0 ) ;
  assign n29796 = ( n240 & n29383 ) | ( n240 & n29787 ) | ( n29383 & n29787 ) ;
  assign n29797 = ( n29383 & ~n29429 ) | ( n29383 & n29787 ) | ( ~n29429 & n29787 ) ;
  assign n29798 = ~n29796 & n29797 ;
  assign n29799 = n29792 | n29798 ;
  assign n29800 = n29377 &  n29430 ;
  assign n29793 = x66 | n29377 ;
  assign n29794 = x66 &  n29377 ;
  assign n29795 = ( n29793 & ~n29794 ) | ( n29793 & 1'b0 ) | ( ~n29794 & 1'b0 ) ;
  assign n29801 = ( n240 & n29382 ) | ( n240 & n29795 ) | ( n29382 & n29795 ) ;
  assign n29802 = ( n29382 & ~n29429 ) | ( n29382 & n29795 ) | ( ~n29429 & n29795 ) ;
  assign n29803 = ~n29801 & n29802 ;
  assign n29804 = n29800 | n29803 ;
  assign n29805 = n29381 &  n29430 ;
  assign n29806 = ( x65 & ~x16 ) | ( x65 & n29378 ) | ( ~x16 & n29378 ) ;
  assign n29807 = ( x16 & ~n29378 ) | ( x16 & x65 ) | ( ~n29378 & x65 ) ;
  assign n29808 = ( n29806 & ~x65 ) | ( n29806 & n29807 ) | ( ~x65 & n29807 ) ;
  assign n29809 = ( n11065 & ~n29429 ) | ( n11065 & n29808 ) | ( ~n29429 & n29808 ) ;
  assign n29810 = ( n240 & n11065 ) | ( n240 & n29808 ) | ( n11065 & n29808 ) ;
  assign n29811 = ( n29809 & ~n29810 ) | ( n29809 & 1'b0 ) | ( ~n29810 & 1'b0 ) ;
  assign n29812 = n29805 | n29811 ;
  assign n29813 = ( n11414 & ~n29429 ) | ( n11414 & 1'b0 ) | ( ~n29429 & 1'b0 ) ;
  assign n29814 = ( x15 & ~n29813 ) | ( x15 & 1'b0 ) | ( ~n29813 & 1'b0 ) ;
  assign n29815 = ( n11418 & ~n29429 ) | ( n11418 & 1'b0 ) | ( ~n29429 & 1'b0 ) ;
  assign n29816 = n29814 | n29815 ;
  assign n29817 = ( x65 & ~n29816 ) | ( x65 & n11421 ) | ( ~n29816 & n11421 ) ;
  assign n29818 = ( x66 & ~n29812 ) | ( x66 & n29817 ) | ( ~n29812 & n29817 ) ;
  assign n29819 = ( x67 & ~n29804 ) | ( x67 & n29818 ) | ( ~n29804 & n29818 ) ;
  assign n29820 = ( x68 & ~n29799 ) | ( x68 & n29819 ) | ( ~n29799 & n29819 ) ;
  assign n29821 = ( x69 & ~n29791 ) | ( x69 & n29820 ) | ( ~n29791 & n29820 ) ;
  assign n29822 = ( x70 & ~n29783 ) | ( x70 & n29821 ) | ( ~n29783 & n29821 ) ;
  assign n29823 = ( x71 & ~n29775 ) | ( x71 & n29822 ) | ( ~n29775 & n29822 ) ;
  assign n29824 = ( x72 & ~n29767 ) | ( x72 & n29823 ) | ( ~n29767 & n29823 ) ;
  assign n29825 = ( x73 & ~n29759 ) | ( x73 & n29824 ) | ( ~n29759 & n29824 ) ;
  assign n29826 = ( x74 & ~n29751 ) | ( x74 & n29825 ) | ( ~n29751 & n29825 ) ;
  assign n29827 = ( x75 & ~n29743 ) | ( x75 & n29826 ) | ( ~n29743 & n29826 ) ;
  assign n29828 = ( x76 & ~n29735 ) | ( x76 & n29827 ) | ( ~n29735 & n29827 ) ;
  assign n29829 = ( x77 & ~n29727 ) | ( x77 & n29828 ) | ( ~n29727 & n29828 ) ;
  assign n29830 = ( x78 & ~n29719 ) | ( x78 & n29829 ) | ( ~n29719 & n29829 ) ;
  assign n29831 = ( x79 & ~n29711 ) | ( x79 & n29830 ) | ( ~n29711 & n29830 ) ;
  assign n29832 = ( x80 & ~n29703 ) | ( x80 & n29831 ) | ( ~n29703 & n29831 ) ;
  assign n29833 = ( x81 & ~n29695 ) | ( x81 & n29832 ) | ( ~n29695 & n29832 ) ;
  assign n29834 = ( x82 & ~n29687 ) | ( x82 & n29833 ) | ( ~n29687 & n29833 ) ;
  assign n29835 = ( x83 & ~n29679 ) | ( x83 & n29834 ) | ( ~n29679 & n29834 ) ;
  assign n29836 = ( x84 & ~n29671 ) | ( x84 & n29835 ) | ( ~n29671 & n29835 ) ;
  assign n29837 = ( x85 & ~n29663 ) | ( x85 & n29836 ) | ( ~n29663 & n29836 ) ;
  assign n29838 = ( x86 & ~n29655 ) | ( x86 & n29837 ) | ( ~n29655 & n29837 ) ;
  assign n29839 = ( x87 & ~n29647 ) | ( x87 & n29838 ) | ( ~n29647 & n29838 ) ;
  assign n29840 = ( x88 & ~n29639 ) | ( x88 & n29839 ) | ( ~n29639 & n29839 ) ;
  assign n29841 = ( x89 & ~n29631 ) | ( x89 & n29840 ) | ( ~n29631 & n29840 ) ;
  assign n29842 = ( x90 & ~n29623 ) | ( x90 & n29841 ) | ( ~n29623 & n29841 ) ;
  assign n29843 = ( x91 & ~n29615 ) | ( x91 & n29842 ) | ( ~n29615 & n29842 ) ;
  assign n29844 = ( x92 & ~n29607 ) | ( x92 & n29843 ) | ( ~n29607 & n29843 ) ;
  assign n29845 = ( x93 & ~n29599 ) | ( x93 & n29844 ) | ( ~n29599 & n29844 ) ;
  assign n29846 = ( x94 & ~n29591 ) | ( x94 & n29845 ) | ( ~n29591 & n29845 ) ;
  assign n29847 = ( x95 & ~n29583 ) | ( x95 & n29846 ) | ( ~n29583 & n29846 ) ;
  assign n29848 = ( x96 & ~n29575 ) | ( x96 & n29847 ) | ( ~n29575 & n29847 ) ;
  assign n29849 = ( x97 & ~n29567 ) | ( x97 & n29848 ) | ( ~n29567 & n29848 ) ;
  assign n29850 = ( x98 & ~n29559 ) | ( x98 & n29849 ) | ( ~n29559 & n29849 ) ;
  assign n29851 = ( x99 & ~n29551 ) | ( x99 & n29850 ) | ( ~n29551 & n29850 ) ;
  assign n29852 = ( x100 & ~n29543 ) | ( x100 & n29851 ) | ( ~n29543 & n29851 ) ;
  assign n29853 = ( x101 & ~n29535 ) | ( x101 & n29852 ) | ( ~n29535 & n29852 ) ;
  assign n29854 = ( x102 & ~n29527 ) | ( x102 & n29853 ) | ( ~n29527 & n29853 ) ;
  assign n29855 = ( x103 & ~n29519 ) | ( x103 & n29854 ) | ( ~n29519 & n29854 ) ;
  assign n29856 = ( x104 & ~n29511 ) | ( x104 & n29855 ) | ( ~n29511 & n29855 ) ;
  assign n29857 = ( x105 & ~n29503 ) | ( x105 & n29856 ) | ( ~n29503 & n29856 ) ;
  assign n29858 = ( x106 & ~n29495 ) | ( x106 & n29857 ) | ( ~n29495 & n29857 ) ;
  assign n29859 = ( x107 & ~n29487 ) | ( x107 & n29858 ) | ( ~n29487 & n29858 ) ;
  assign n29860 = ( x108 & ~n29479 ) | ( x108 & n29859 ) | ( ~n29479 & n29859 ) ;
  assign n29861 = ( x109 & ~n29471 ) | ( x109 & n29860 ) | ( ~n29471 & n29860 ) ;
  assign n29862 = ( x110 & ~n29463 ) | ( x110 & n29861 ) | ( ~n29463 & n29861 ) ;
  assign n29863 = ( x111 & ~n29455 ) | ( x111 & n29862 ) | ( ~n29455 & n29862 ) ;
  assign n29864 = ( x112 & ~n29447 ) | ( x112 & n29863 ) | ( ~n29447 & n29863 ) ;
  assign n29431 = n29014 &  n29430 ;
  assign n29435 = ( n240 & n29014 ) | ( n240 & n29428 ) | ( n29014 & n29428 ) ;
  assign n29436 = ( x112 & ~n29435 ) | ( x112 & n29014 ) | ( ~n29435 & n29014 ) ;
  assign n29437 = ~x112 & n29436 ;
  assign n29438 = n29431 | n29437 ;
  assign n29439 = ~x113 & n29438 ;
  assign n29865 = ( x113 & ~n29431 ) | ( x113 & 1'b0 ) | ( ~n29431 & 1'b0 ) ;
  assign n29866 = ~n29437 & n29865 ;
  assign n29875 = n29439 | n29866 ;
  assign n29876 = ( n29864 & ~n29875 ) | ( n29864 & 1'b0 ) | ( ~n29875 & 1'b0 ) ;
  assign n29867 = ( n29864 & ~n29439 ) | ( n29864 & n29866 ) | ( ~n29439 & n29866 ) ;
  assign n29868 = ( n29439 & ~n11560 ) | ( n29439 & n29867 ) | ( ~n11560 & n29867 ) ;
  assign n29869 = n11560 | n29868 ;
  assign n29870 = ~n29438 |  n240 ;
  assign n29871 = n29869 &  n29870 ;
  assign n29877 = ~n29864 & n29875 ;
  assign n29878 = ( n29876 & ~n29871 ) | ( n29876 & n29877 ) | ( ~n29871 & n29877 ) ;
  assign n29879 = n240 &  n29014 ;
  assign n29880 = n29869 &  n29879 ;
  assign n29881 = n29878 | n29880 ;
  assign n29882 = ~x114 & n29881 ;
  assign n29886 = n29447 &  n29870 ;
  assign n29887 = n29869 &  n29886 ;
  assign n29872 = x112 | n29447 ;
  assign n29873 = x112 &  n29447 ;
  assign n29874 = ( n29872 & ~n29873 ) | ( n29872 & 1'b0 ) | ( ~n29873 & 1'b0 ) ;
  assign n29889 = ( n29863 & n29871 ) | ( n29863 & n29874 ) | ( n29871 & n29874 ) ;
  assign n29888 = n29863 | n29874 ;
  assign n29890 = ( n29887 & ~n29889 ) | ( n29887 & n29888 ) | ( ~n29889 & n29888 ) ;
  assign n29894 = n29455 &  n29870 ;
  assign n29895 = n29869 &  n29894 ;
  assign n29883 = x111 | n29455 ;
  assign n29884 = x111 &  n29455 ;
  assign n29885 = ( n29883 & ~n29884 ) | ( n29883 & 1'b0 ) | ( ~n29884 & 1'b0 ) ;
  assign n29897 = ( n29862 & n29871 ) | ( n29862 & n29885 ) | ( n29871 & n29885 ) ;
  assign n29896 = n29862 | n29885 ;
  assign n29898 = ( n29895 & ~n29897 ) | ( n29895 & n29896 ) | ( ~n29897 & n29896 ) ;
  assign n29902 = n29463 &  n29870 ;
  assign n29903 = n29869 &  n29902 ;
  assign n29891 = x110 | n29463 ;
  assign n29892 = x110 &  n29463 ;
  assign n29893 = ( n29891 & ~n29892 ) | ( n29891 & 1'b0 ) | ( ~n29892 & 1'b0 ) ;
  assign n29905 = ( n29861 & n29871 ) | ( n29861 & n29893 ) | ( n29871 & n29893 ) ;
  assign n29904 = n29861 | n29893 ;
  assign n29906 = ( n29903 & ~n29905 ) | ( n29903 & n29904 ) | ( ~n29905 & n29904 ) ;
  assign n29910 = n29471 &  n29870 ;
  assign n29911 = n29869 &  n29910 ;
  assign n29899 = x109 | n29471 ;
  assign n29900 = x109 &  n29471 ;
  assign n29901 = ( n29899 & ~n29900 ) | ( n29899 & 1'b0 ) | ( ~n29900 & 1'b0 ) ;
  assign n29913 = ( n29860 & n29871 ) | ( n29860 & n29901 ) | ( n29871 & n29901 ) ;
  assign n29912 = n29860 | n29901 ;
  assign n29914 = ( n29911 & ~n29913 ) | ( n29911 & n29912 ) | ( ~n29913 & n29912 ) ;
  assign n29918 = n29479 &  n29870 ;
  assign n29919 = n29869 &  n29918 ;
  assign n29907 = x108 | n29479 ;
  assign n29908 = x108 &  n29479 ;
  assign n29909 = ( n29907 & ~n29908 ) | ( n29907 & 1'b0 ) | ( ~n29908 & 1'b0 ) ;
  assign n29921 = ( n29859 & n29871 ) | ( n29859 & n29909 ) | ( n29871 & n29909 ) ;
  assign n29920 = n29859 | n29909 ;
  assign n29922 = ( n29919 & ~n29921 ) | ( n29919 & n29920 ) | ( ~n29921 & n29920 ) ;
  assign n29926 = n29487 &  n29870 ;
  assign n29927 = n29869 &  n29926 ;
  assign n29915 = x107 | n29487 ;
  assign n29916 = x107 &  n29487 ;
  assign n29917 = ( n29915 & ~n29916 ) | ( n29915 & 1'b0 ) | ( ~n29916 & 1'b0 ) ;
  assign n29929 = ( n29858 & n29871 ) | ( n29858 & n29917 ) | ( n29871 & n29917 ) ;
  assign n29928 = n29858 | n29917 ;
  assign n29930 = ( n29927 & ~n29929 ) | ( n29927 & n29928 ) | ( ~n29929 & n29928 ) ;
  assign n29934 = n29495 &  n29870 ;
  assign n29935 = n29869 &  n29934 ;
  assign n29923 = x106 | n29495 ;
  assign n29924 = x106 &  n29495 ;
  assign n29925 = ( n29923 & ~n29924 ) | ( n29923 & 1'b0 ) | ( ~n29924 & 1'b0 ) ;
  assign n29937 = ( n29857 & n29871 ) | ( n29857 & n29925 ) | ( n29871 & n29925 ) ;
  assign n29936 = n29857 | n29925 ;
  assign n29938 = ( n29935 & ~n29937 ) | ( n29935 & n29936 ) | ( ~n29937 & n29936 ) ;
  assign n29942 = n29503 &  n29870 ;
  assign n29943 = n29869 &  n29942 ;
  assign n29931 = x105 | n29503 ;
  assign n29932 = x105 &  n29503 ;
  assign n29933 = ( n29931 & ~n29932 ) | ( n29931 & 1'b0 ) | ( ~n29932 & 1'b0 ) ;
  assign n29945 = ( n29856 & n29871 ) | ( n29856 & n29933 ) | ( n29871 & n29933 ) ;
  assign n29944 = n29856 | n29933 ;
  assign n29946 = ( n29943 & ~n29945 ) | ( n29943 & n29944 ) | ( ~n29945 & n29944 ) ;
  assign n29950 = n29511 &  n29870 ;
  assign n29951 = n29869 &  n29950 ;
  assign n29939 = x104 | n29511 ;
  assign n29940 = x104 &  n29511 ;
  assign n29941 = ( n29939 & ~n29940 ) | ( n29939 & 1'b0 ) | ( ~n29940 & 1'b0 ) ;
  assign n29953 = ( n29855 & n29871 ) | ( n29855 & n29941 ) | ( n29871 & n29941 ) ;
  assign n29952 = n29855 | n29941 ;
  assign n29954 = ( n29951 & ~n29953 ) | ( n29951 & n29952 ) | ( ~n29953 & n29952 ) ;
  assign n29958 = n29519 &  n29870 ;
  assign n29959 = n29869 &  n29958 ;
  assign n29947 = x103 | n29519 ;
  assign n29948 = x103 &  n29519 ;
  assign n29949 = ( n29947 & ~n29948 ) | ( n29947 & 1'b0 ) | ( ~n29948 & 1'b0 ) ;
  assign n29961 = ( n29854 & n29871 ) | ( n29854 & n29949 ) | ( n29871 & n29949 ) ;
  assign n29960 = n29854 | n29949 ;
  assign n29962 = ( n29959 & ~n29961 ) | ( n29959 & n29960 ) | ( ~n29961 & n29960 ) ;
  assign n29966 = n29527 &  n29870 ;
  assign n29967 = n29869 &  n29966 ;
  assign n29955 = x102 | n29527 ;
  assign n29956 = x102 &  n29527 ;
  assign n29957 = ( n29955 & ~n29956 ) | ( n29955 & 1'b0 ) | ( ~n29956 & 1'b0 ) ;
  assign n29969 = ( n29853 & n29871 ) | ( n29853 & n29957 ) | ( n29871 & n29957 ) ;
  assign n29968 = n29853 | n29957 ;
  assign n29970 = ( n29967 & ~n29969 ) | ( n29967 & n29968 ) | ( ~n29969 & n29968 ) ;
  assign n29974 = n29535 &  n29870 ;
  assign n29975 = n29869 &  n29974 ;
  assign n29963 = x101 | n29535 ;
  assign n29964 = x101 &  n29535 ;
  assign n29965 = ( n29963 & ~n29964 ) | ( n29963 & 1'b0 ) | ( ~n29964 & 1'b0 ) ;
  assign n29977 = ( n29852 & n29871 ) | ( n29852 & n29965 ) | ( n29871 & n29965 ) ;
  assign n29976 = n29852 | n29965 ;
  assign n29978 = ( n29975 & ~n29977 ) | ( n29975 & n29976 ) | ( ~n29977 & n29976 ) ;
  assign n29982 = n29543 &  n29870 ;
  assign n29983 = n29869 &  n29982 ;
  assign n29971 = x100 | n29543 ;
  assign n29972 = x100 &  n29543 ;
  assign n29973 = ( n29971 & ~n29972 ) | ( n29971 & 1'b0 ) | ( ~n29972 & 1'b0 ) ;
  assign n29985 = ( n29851 & n29871 ) | ( n29851 & n29973 ) | ( n29871 & n29973 ) ;
  assign n29984 = n29851 | n29973 ;
  assign n29986 = ( n29983 & ~n29985 ) | ( n29983 & n29984 ) | ( ~n29985 & n29984 ) ;
  assign n29990 = n29551 &  n29870 ;
  assign n29991 = n29869 &  n29990 ;
  assign n29979 = x99 | n29551 ;
  assign n29980 = x99 &  n29551 ;
  assign n29981 = ( n29979 & ~n29980 ) | ( n29979 & 1'b0 ) | ( ~n29980 & 1'b0 ) ;
  assign n29993 = ( n29850 & n29871 ) | ( n29850 & n29981 ) | ( n29871 & n29981 ) ;
  assign n29992 = n29850 | n29981 ;
  assign n29994 = ( n29991 & ~n29993 ) | ( n29991 & n29992 ) | ( ~n29993 & n29992 ) ;
  assign n29998 = n29559 &  n29870 ;
  assign n29999 = n29869 &  n29998 ;
  assign n29987 = x98 | n29559 ;
  assign n29988 = x98 &  n29559 ;
  assign n29989 = ( n29987 & ~n29988 ) | ( n29987 & 1'b0 ) | ( ~n29988 & 1'b0 ) ;
  assign n30001 = ( n29849 & n29871 ) | ( n29849 & n29989 ) | ( n29871 & n29989 ) ;
  assign n30000 = n29849 | n29989 ;
  assign n30002 = ( n29999 & ~n30001 ) | ( n29999 & n30000 ) | ( ~n30001 & n30000 ) ;
  assign n30006 = n29567 &  n29870 ;
  assign n30007 = n29869 &  n30006 ;
  assign n29995 = x97 | n29567 ;
  assign n29996 = x97 &  n29567 ;
  assign n29997 = ( n29995 & ~n29996 ) | ( n29995 & 1'b0 ) | ( ~n29996 & 1'b0 ) ;
  assign n30009 = ( n29848 & n29871 ) | ( n29848 & n29997 ) | ( n29871 & n29997 ) ;
  assign n30008 = n29848 | n29997 ;
  assign n30010 = ( n30007 & ~n30009 ) | ( n30007 & n30008 ) | ( ~n30009 & n30008 ) ;
  assign n30014 = n29575 &  n29870 ;
  assign n30015 = n29869 &  n30014 ;
  assign n30003 = x96 | n29575 ;
  assign n30004 = x96 &  n29575 ;
  assign n30005 = ( n30003 & ~n30004 ) | ( n30003 & 1'b0 ) | ( ~n30004 & 1'b0 ) ;
  assign n30017 = ( n29847 & n29871 ) | ( n29847 & n30005 ) | ( n29871 & n30005 ) ;
  assign n30016 = n29847 | n30005 ;
  assign n30018 = ( n30015 & ~n30017 ) | ( n30015 & n30016 ) | ( ~n30017 & n30016 ) ;
  assign n30022 = n29583 &  n29870 ;
  assign n30023 = n29869 &  n30022 ;
  assign n30011 = x95 | n29583 ;
  assign n30012 = x95 &  n29583 ;
  assign n30013 = ( n30011 & ~n30012 ) | ( n30011 & 1'b0 ) | ( ~n30012 & 1'b0 ) ;
  assign n30025 = ( n29846 & n29871 ) | ( n29846 & n30013 ) | ( n29871 & n30013 ) ;
  assign n30024 = n29846 | n30013 ;
  assign n30026 = ( n30023 & ~n30025 ) | ( n30023 & n30024 ) | ( ~n30025 & n30024 ) ;
  assign n30030 = n29591 &  n29870 ;
  assign n30031 = n29869 &  n30030 ;
  assign n30019 = x94 | n29591 ;
  assign n30020 = x94 &  n29591 ;
  assign n30021 = ( n30019 & ~n30020 ) | ( n30019 & 1'b0 ) | ( ~n30020 & 1'b0 ) ;
  assign n30033 = ( n29845 & n29871 ) | ( n29845 & n30021 ) | ( n29871 & n30021 ) ;
  assign n30032 = n29845 | n30021 ;
  assign n30034 = ( n30031 & ~n30033 ) | ( n30031 & n30032 ) | ( ~n30033 & n30032 ) ;
  assign n30038 = n29599 &  n29870 ;
  assign n30039 = n29869 &  n30038 ;
  assign n30027 = x93 | n29599 ;
  assign n30028 = x93 &  n29599 ;
  assign n30029 = ( n30027 & ~n30028 ) | ( n30027 & 1'b0 ) | ( ~n30028 & 1'b0 ) ;
  assign n30041 = ( n29844 & n29871 ) | ( n29844 & n30029 ) | ( n29871 & n30029 ) ;
  assign n30040 = n29844 | n30029 ;
  assign n30042 = ( n30039 & ~n30041 ) | ( n30039 & n30040 ) | ( ~n30041 & n30040 ) ;
  assign n30046 = n29607 &  n29870 ;
  assign n30047 = n29869 &  n30046 ;
  assign n30035 = x92 | n29607 ;
  assign n30036 = x92 &  n29607 ;
  assign n30037 = ( n30035 & ~n30036 ) | ( n30035 & 1'b0 ) | ( ~n30036 & 1'b0 ) ;
  assign n30049 = ( n29843 & n29871 ) | ( n29843 & n30037 ) | ( n29871 & n30037 ) ;
  assign n30048 = n29843 | n30037 ;
  assign n30050 = ( n30047 & ~n30049 ) | ( n30047 & n30048 ) | ( ~n30049 & n30048 ) ;
  assign n30054 = n29615 &  n29870 ;
  assign n30055 = n29869 &  n30054 ;
  assign n30043 = x91 | n29615 ;
  assign n30044 = x91 &  n29615 ;
  assign n30045 = ( n30043 & ~n30044 ) | ( n30043 & 1'b0 ) | ( ~n30044 & 1'b0 ) ;
  assign n30057 = ( n29842 & n29871 ) | ( n29842 & n30045 ) | ( n29871 & n30045 ) ;
  assign n30056 = n29842 | n30045 ;
  assign n30058 = ( n30055 & ~n30057 ) | ( n30055 & n30056 ) | ( ~n30057 & n30056 ) ;
  assign n30062 = n29623 &  n29870 ;
  assign n30063 = n29869 &  n30062 ;
  assign n30051 = x90 | n29623 ;
  assign n30052 = x90 &  n29623 ;
  assign n30053 = ( n30051 & ~n30052 ) | ( n30051 & 1'b0 ) | ( ~n30052 & 1'b0 ) ;
  assign n30065 = ( n29841 & n29871 ) | ( n29841 & n30053 ) | ( n29871 & n30053 ) ;
  assign n30064 = n29841 | n30053 ;
  assign n30066 = ( n30063 & ~n30065 ) | ( n30063 & n30064 ) | ( ~n30065 & n30064 ) ;
  assign n30070 = n29631 &  n29870 ;
  assign n30071 = n29869 &  n30070 ;
  assign n30059 = x89 | n29631 ;
  assign n30060 = x89 &  n29631 ;
  assign n30061 = ( n30059 & ~n30060 ) | ( n30059 & 1'b0 ) | ( ~n30060 & 1'b0 ) ;
  assign n30073 = ( n29840 & n29871 ) | ( n29840 & n30061 ) | ( n29871 & n30061 ) ;
  assign n30072 = n29840 | n30061 ;
  assign n30074 = ( n30071 & ~n30073 ) | ( n30071 & n30072 ) | ( ~n30073 & n30072 ) ;
  assign n30078 = n29639 &  n29870 ;
  assign n30079 = n29869 &  n30078 ;
  assign n30067 = x88 | n29639 ;
  assign n30068 = x88 &  n29639 ;
  assign n30069 = ( n30067 & ~n30068 ) | ( n30067 & 1'b0 ) | ( ~n30068 & 1'b0 ) ;
  assign n30081 = ( n29839 & n29871 ) | ( n29839 & n30069 ) | ( n29871 & n30069 ) ;
  assign n30080 = n29839 | n30069 ;
  assign n30082 = ( n30079 & ~n30081 ) | ( n30079 & n30080 ) | ( ~n30081 & n30080 ) ;
  assign n30086 = n29647 &  n29870 ;
  assign n30087 = n29869 &  n30086 ;
  assign n30075 = x87 | n29647 ;
  assign n30076 = x87 &  n29647 ;
  assign n30077 = ( n30075 & ~n30076 ) | ( n30075 & 1'b0 ) | ( ~n30076 & 1'b0 ) ;
  assign n30089 = ( n29838 & n29871 ) | ( n29838 & n30077 ) | ( n29871 & n30077 ) ;
  assign n30088 = n29838 | n30077 ;
  assign n30090 = ( n30087 & ~n30089 ) | ( n30087 & n30088 ) | ( ~n30089 & n30088 ) ;
  assign n30094 = n29655 &  n29870 ;
  assign n30095 = n29869 &  n30094 ;
  assign n30083 = x86 | n29655 ;
  assign n30084 = x86 &  n29655 ;
  assign n30085 = ( n30083 & ~n30084 ) | ( n30083 & 1'b0 ) | ( ~n30084 & 1'b0 ) ;
  assign n30097 = ( n29837 & n29871 ) | ( n29837 & n30085 ) | ( n29871 & n30085 ) ;
  assign n30096 = n29837 | n30085 ;
  assign n30098 = ( n30095 & ~n30097 ) | ( n30095 & n30096 ) | ( ~n30097 & n30096 ) ;
  assign n30102 = n29663 &  n29870 ;
  assign n30103 = n29869 &  n30102 ;
  assign n30091 = x85 | n29663 ;
  assign n30092 = x85 &  n29663 ;
  assign n30093 = ( n30091 & ~n30092 ) | ( n30091 & 1'b0 ) | ( ~n30092 & 1'b0 ) ;
  assign n30105 = ( n29836 & n29871 ) | ( n29836 & n30093 ) | ( n29871 & n30093 ) ;
  assign n30104 = n29836 | n30093 ;
  assign n30106 = ( n30103 & ~n30105 ) | ( n30103 & n30104 ) | ( ~n30105 & n30104 ) ;
  assign n30110 = n29671 &  n29870 ;
  assign n30111 = n29869 &  n30110 ;
  assign n30099 = x84 | n29671 ;
  assign n30100 = x84 &  n29671 ;
  assign n30101 = ( n30099 & ~n30100 ) | ( n30099 & 1'b0 ) | ( ~n30100 & 1'b0 ) ;
  assign n30113 = ( n29835 & n29871 ) | ( n29835 & n30101 ) | ( n29871 & n30101 ) ;
  assign n30112 = n29835 | n30101 ;
  assign n30114 = ( n30111 & ~n30113 ) | ( n30111 & n30112 ) | ( ~n30113 & n30112 ) ;
  assign n30118 = n29679 &  n29870 ;
  assign n30119 = n29869 &  n30118 ;
  assign n30107 = x83 | n29679 ;
  assign n30108 = x83 &  n29679 ;
  assign n30109 = ( n30107 & ~n30108 ) | ( n30107 & 1'b0 ) | ( ~n30108 & 1'b0 ) ;
  assign n30121 = ( n29834 & n29871 ) | ( n29834 & n30109 ) | ( n29871 & n30109 ) ;
  assign n30120 = n29834 | n30109 ;
  assign n30122 = ( n30119 & ~n30121 ) | ( n30119 & n30120 ) | ( ~n30121 & n30120 ) ;
  assign n30126 = n29687 &  n29870 ;
  assign n30127 = n29869 &  n30126 ;
  assign n30115 = x82 | n29687 ;
  assign n30116 = x82 &  n29687 ;
  assign n30117 = ( n30115 & ~n30116 ) | ( n30115 & 1'b0 ) | ( ~n30116 & 1'b0 ) ;
  assign n30129 = ( n29833 & n29871 ) | ( n29833 & n30117 ) | ( n29871 & n30117 ) ;
  assign n30128 = n29833 | n30117 ;
  assign n30130 = ( n30127 & ~n30129 ) | ( n30127 & n30128 ) | ( ~n30129 & n30128 ) ;
  assign n30134 = n29695 &  n29870 ;
  assign n30135 = n29869 &  n30134 ;
  assign n30123 = x81 | n29695 ;
  assign n30124 = x81 &  n29695 ;
  assign n30125 = ( n30123 & ~n30124 ) | ( n30123 & 1'b0 ) | ( ~n30124 & 1'b0 ) ;
  assign n30137 = ( n29832 & n29871 ) | ( n29832 & n30125 ) | ( n29871 & n30125 ) ;
  assign n30136 = n29832 | n30125 ;
  assign n30138 = ( n30135 & ~n30137 ) | ( n30135 & n30136 ) | ( ~n30137 & n30136 ) ;
  assign n30142 = n29703 &  n29870 ;
  assign n30143 = n29869 &  n30142 ;
  assign n30131 = x80 | n29703 ;
  assign n30132 = x80 &  n29703 ;
  assign n30133 = ( n30131 & ~n30132 ) | ( n30131 & 1'b0 ) | ( ~n30132 & 1'b0 ) ;
  assign n30145 = ( n29831 & n29871 ) | ( n29831 & n30133 ) | ( n29871 & n30133 ) ;
  assign n30144 = n29831 | n30133 ;
  assign n30146 = ( n30143 & ~n30145 ) | ( n30143 & n30144 ) | ( ~n30145 & n30144 ) ;
  assign n30150 = n29711 &  n29870 ;
  assign n30151 = n29869 &  n30150 ;
  assign n30139 = x79 | n29711 ;
  assign n30140 = x79 &  n29711 ;
  assign n30141 = ( n30139 & ~n30140 ) | ( n30139 & 1'b0 ) | ( ~n30140 & 1'b0 ) ;
  assign n30153 = ( n29830 & n29871 ) | ( n29830 & n30141 ) | ( n29871 & n30141 ) ;
  assign n30152 = n29830 | n30141 ;
  assign n30154 = ( n30151 & ~n30153 ) | ( n30151 & n30152 ) | ( ~n30153 & n30152 ) ;
  assign n30158 = n29719 &  n29870 ;
  assign n30159 = n29869 &  n30158 ;
  assign n30147 = x78 | n29719 ;
  assign n30148 = x78 &  n29719 ;
  assign n30149 = ( n30147 & ~n30148 ) | ( n30147 & 1'b0 ) | ( ~n30148 & 1'b0 ) ;
  assign n30161 = ( n29829 & n29871 ) | ( n29829 & n30149 ) | ( n29871 & n30149 ) ;
  assign n30160 = n29829 | n30149 ;
  assign n30162 = ( n30159 & ~n30161 ) | ( n30159 & n30160 ) | ( ~n30161 & n30160 ) ;
  assign n30166 = n29727 &  n29870 ;
  assign n30167 = n29869 &  n30166 ;
  assign n30155 = x77 | n29727 ;
  assign n30156 = x77 &  n29727 ;
  assign n30157 = ( n30155 & ~n30156 ) | ( n30155 & 1'b0 ) | ( ~n30156 & 1'b0 ) ;
  assign n30169 = ( n29828 & n29871 ) | ( n29828 & n30157 ) | ( n29871 & n30157 ) ;
  assign n30168 = n29828 | n30157 ;
  assign n30170 = ( n30167 & ~n30169 ) | ( n30167 & n30168 ) | ( ~n30169 & n30168 ) ;
  assign n30174 = n29735 &  n29870 ;
  assign n30175 = n29869 &  n30174 ;
  assign n30163 = x76 | n29735 ;
  assign n30164 = x76 &  n29735 ;
  assign n30165 = ( n30163 & ~n30164 ) | ( n30163 & 1'b0 ) | ( ~n30164 & 1'b0 ) ;
  assign n30177 = ( n29827 & n29871 ) | ( n29827 & n30165 ) | ( n29871 & n30165 ) ;
  assign n30176 = n29827 | n30165 ;
  assign n30178 = ( n30175 & ~n30177 ) | ( n30175 & n30176 ) | ( ~n30177 & n30176 ) ;
  assign n30182 = n29743 &  n29870 ;
  assign n30183 = n29869 &  n30182 ;
  assign n30171 = x75 | n29743 ;
  assign n30172 = x75 &  n29743 ;
  assign n30173 = ( n30171 & ~n30172 ) | ( n30171 & 1'b0 ) | ( ~n30172 & 1'b0 ) ;
  assign n30185 = ( n29826 & n29871 ) | ( n29826 & n30173 ) | ( n29871 & n30173 ) ;
  assign n30184 = n29826 | n30173 ;
  assign n30186 = ( n30183 & ~n30185 ) | ( n30183 & n30184 ) | ( ~n30185 & n30184 ) ;
  assign n30190 = n29751 &  n29870 ;
  assign n30191 = n29869 &  n30190 ;
  assign n30179 = x74 | n29751 ;
  assign n30180 = x74 &  n29751 ;
  assign n30181 = ( n30179 & ~n30180 ) | ( n30179 & 1'b0 ) | ( ~n30180 & 1'b0 ) ;
  assign n30193 = ( n29825 & n29871 ) | ( n29825 & n30181 ) | ( n29871 & n30181 ) ;
  assign n30192 = n29825 | n30181 ;
  assign n30194 = ( n30191 & ~n30193 ) | ( n30191 & n30192 ) | ( ~n30193 & n30192 ) ;
  assign n30198 = n29759 &  n29870 ;
  assign n30199 = n29869 &  n30198 ;
  assign n30187 = x73 | n29759 ;
  assign n30188 = x73 &  n29759 ;
  assign n30189 = ( n30187 & ~n30188 ) | ( n30187 & 1'b0 ) | ( ~n30188 & 1'b0 ) ;
  assign n30201 = ( n29824 & n29871 ) | ( n29824 & n30189 ) | ( n29871 & n30189 ) ;
  assign n30200 = n29824 | n30189 ;
  assign n30202 = ( n30199 & ~n30201 ) | ( n30199 & n30200 ) | ( ~n30201 & n30200 ) ;
  assign n30206 = n29767 &  n29870 ;
  assign n30207 = n29869 &  n30206 ;
  assign n30195 = x72 | n29767 ;
  assign n30196 = x72 &  n29767 ;
  assign n30197 = ( n30195 & ~n30196 ) | ( n30195 & 1'b0 ) | ( ~n30196 & 1'b0 ) ;
  assign n30209 = ( n29823 & n29871 ) | ( n29823 & n30197 ) | ( n29871 & n30197 ) ;
  assign n30208 = n29823 | n30197 ;
  assign n30210 = ( n30207 & ~n30209 ) | ( n30207 & n30208 ) | ( ~n30209 & n30208 ) ;
  assign n30214 = n29775 &  n29870 ;
  assign n30215 = n29869 &  n30214 ;
  assign n30203 = x71 | n29775 ;
  assign n30204 = x71 &  n29775 ;
  assign n30205 = ( n30203 & ~n30204 ) | ( n30203 & 1'b0 ) | ( ~n30204 & 1'b0 ) ;
  assign n30217 = ( n29822 & n29871 ) | ( n29822 & n30205 ) | ( n29871 & n30205 ) ;
  assign n30216 = n29822 | n30205 ;
  assign n30218 = ( n30215 & ~n30217 ) | ( n30215 & n30216 ) | ( ~n30217 & n30216 ) ;
  assign n30222 = n29783 &  n29870 ;
  assign n30223 = n29869 &  n30222 ;
  assign n30211 = x70 | n29783 ;
  assign n30212 = x70 &  n29783 ;
  assign n30213 = ( n30211 & ~n30212 ) | ( n30211 & 1'b0 ) | ( ~n30212 & 1'b0 ) ;
  assign n30225 = ( n29821 & n29871 ) | ( n29821 & n30213 ) | ( n29871 & n30213 ) ;
  assign n30224 = n29821 | n30213 ;
  assign n30226 = ( n30223 & ~n30225 ) | ( n30223 & n30224 ) | ( ~n30225 & n30224 ) ;
  assign n30230 = n29791 &  n29870 ;
  assign n30231 = n29869 &  n30230 ;
  assign n30219 = x69 | n29791 ;
  assign n30220 = x69 &  n29791 ;
  assign n30221 = ( n30219 & ~n30220 ) | ( n30219 & 1'b0 ) | ( ~n30220 & 1'b0 ) ;
  assign n30233 = ( n29820 & n29871 ) | ( n29820 & n30221 ) | ( n29871 & n30221 ) ;
  assign n30232 = n29820 | n30221 ;
  assign n30234 = ( n30231 & ~n30233 ) | ( n30231 & n30232 ) | ( ~n30233 & n30232 ) ;
  assign n30238 = n29799 &  n29870 ;
  assign n30239 = n29869 &  n30238 ;
  assign n30227 = x68 | n29799 ;
  assign n30228 = x68 &  n29799 ;
  assign n30229 = ( n30227 & ~n30228 ) | ( n30227 & 1'b0 ) | ( ~n30228 & 1'b0 ) ;
  assign n30241 = ( n29819 & n29871 ) | ( n29819 & n30229 ) | ( n29871 & n30229 ) ;
  assign n30240 = n29819 | n30229 ;
  assign n30242 = ( n30239 & ~n30241 ) | ( n30239 & n30240 ) | ( ~n30241 & n30240 ) ;
  assign n30246 = n29804 &  n29870 ;
  assign n30247 = n29869 &  n30246 ;
  assign n30235 = x67 | n29804 ;
  assign n30236 = x67 &  n29804 ;
  assign n30237 = ( n30235 & ~n30236 ) | ( n30235 & 1'b0 ) | ( ~n30236 & 1'b0 ) ;
  assign n30249 = ( n29818 & n29871 ) | ( n29818 & n30237 ) | ( n29871 & n30237 ) ;
  assign n30248 = n29818 | n30237 ;
  assign n30250 = ( n30247 & ~n30249 ) | ( n30247 & n30248 ) | ( ~n30249 & n30248 ) ;
  assign n30251 = n29812 &  n29870 ;
  assign n30252 = n29869 &  n30251 ;
  assign n30243 = x66 | n29812 ;
  assign n30244 = x66 &  n29812 ;
  assign n30245 = ( n30243 & ~n30244 ) | ( n30243 & 1'b0 ) | ( ~n30244 & 1'b0 ) ;
  assign n30254 = ( n29817 & n29871 ) | ( n29817 & n30245 ) | ( n29871 & n30245 ) ;
  assign n30253 = n29817 | n30245 ;
  assign n30255 = ( n30252 & ~n30254 ) | ( n30252 & n30253 ) | ( ~n30254 & n30253 ) ;
  assign n30256 = ( x65 & ~n11421 ) | ( x65 & n29816 ) | ( ~n11421 & n29816 ) ;
  assign n30257 = ( n29817 & ~x65 ) | ( n29817 & n30256 ) | ( ~x65 & n30256 ) ;
  assign n30258 = ~n29871 & n30257 ;
  assign n30259 = n29816 &  n29870 ;
  assign n30260 = n29869 &  n30259 ;
  assign n30261 = n30258 | n30260 ;
  assign n30262 = ( x64 & ~n29871 ) | ( x64 & 1'b0 ) | ( ~n29871 & 1'b0 ) ;
  assign n30263 = ( x14 & ~n30262 ) | ( x14 & 1'b0 ) | ( ~n30262 & 1'b0 ) ;
  assign n30264 = ( n11421 & ~n29871 ) | ( n11421 & 1'b0 ) | ( ~n29871 & 1'b0 ) ;
  assign n30265 = n30263 | n30264 ;
  assign n30266 = ( x65 & ~n30265 ) | ( x65 & n11875 ) | ( ~n30265 & n11875 ) ;
  assign n30267 = ( x66 & ~n30261 ) | ( x66 & n30266 ) | ( ~n30261 & n30266 ) ;
  assign n30268 = ( x67 & ~n30255 ) | ( x67 & n30267 ) | ( ~n30255 & n30267 ) ;
  assign n30269 = ( x68 & ~n30250 ) | ( x68 & n30268 ) | ( ~n30250 & n30268 ) ;
  assign n30270 = ( x69 & ~n30242 ) | ( x69 & n30269 ) | ( ~n30242 & n30269 ) ;
  assign n30271 = ( x70 & ~n30234 ) | ( x70 & n30270 ) | ( ~n30234 & n30270 ) ;
  assign n30272 = ( x71 & ~n30226 ) | ( x71 & n30271 ) | ( ~n30226 & n30271 ) ;
  assign n30273 = ( x72 & ~n30218 ) | ( x72 & n30272 ) | ( ~n30218 & n30272 ) ;
  assign n30274 = ( x73 & ~n30210 ) | ( x73 & n30273 ) | ( ~n30210 & n30273 ) ;
  assign n30275 = ( x74 & ~n30202 ) | ( x74 & n30274 ) | ( ~n30202 & n30274 ) ;
  assign n30276 = ( x75 & ~n30194 ) | ( x75 & n30275 ) | ( ~n30194 & n30275 ) ;
  assign n30277 = ( x76 & ~n30186 ) | ( x76 & n30276 ) | ( ~n30186 & n30276 ) ;
  assign n30278 = ( x77 & ~n30178 ) | ( x77 & n30277 ) | ( ~n30178 & n30277 ) ;
  assign n30279 = ( x78 & ~n30170 ) | ( x78 & n30278 ) | ( ~n30170 & n30278 ) ;
  assign n30280 = ( x79 & ~n30162 ) | ( x79 & n30279 ) | ( ~n30162 & n30279 ) ;
  assign n30281 = ( x80 & ~n30154 ) | ( x80 & n30280 ) | ( ~n30154 & n30280 ) ;
  assign n30282 = ( x81 & ~n30146 ) | ( x81 & n30281 ) | ( ~n30146 & n30281 ) ;
  assign n30283 = ( x82 & ~n30138 ) | ( x82 & n30282 ) | ( ~n30138 & n30282 ) ;
  assign n30284 = ( x83 & ~n30130 ) | ( x83 & n30283 ) | ( ~n30130 & n30283 ) ;
  assign n30285 = ( x84 & ~n30122 ) | ( x84 & n30284 ) | ( ~n30122 & n30284 ) ;
  assign n30286 = ( x85 & ~n30114 ) | ( x85 & n30285 ) | ( ~n30114 & n30285 ) ;
  assign n30287 = ( x86 & ~n30106 ) | ( x86 & n30286 ) | ( ~n30106 & n30286 ) ;
  assign n30288 = ( x87 & ~n30098 ) | ( x87 & n30287 ) | ( ~n30098 & n30287 ) ;
  assign n30289 = ( x88 & ~n30090 ) | ( x88 & n30288 ) | ( ~n30090 & n30288 ) ;
  assign n30290 = ( x89 & ~n30082 ) | ( x89 & n30289 ) | ( ~n30082 & n30289 ) ;
  assign n30291 = ( x90 & ~n30074 ) | ( x90 & n30290 ) | ( ~n30074 & n30290 ) ;
  assign n30292 = ( x91 & ~n30066 ) | ( x91 & n30291 ) | ( ~n30066 & n30291 ) ;
  assign n30293 = ( x92 & ~n30058 ) | ( x92 & n30292 ) | ( ~n30058 & n30292 ) ;
  assign n30294 = ( x93 & ~n30050 ) | ( x93 & n30293 ) | ( ~n30050 & n30293 ) ;
  assign n30295 = ( x94 & ~n30042 ) | ( x94 & n30294 ) | ( ~n30042 & n30294 ) ;
  assign n30296 = ( x95 & ~n30034 ) | ( x95 & n30295 ) | ( ~n30034 & n30295 ) ;
  assign n30297 = ( x96 & ~n30026 ) | ( x96 & n30296 ) | ( ~n30026 & n30296 ) ;
  assign n30298 = ( x97 & ~n30018 ) | ( x97 & n30297 ) | ( ~n30018 & n30297 ) ;
  assign n30299 = ( x98 & ~n30010 ) | ( x98 & n30298 ) | ( ~n30010 & n30298 ) ;
  assign n30300 = ( x99 & ~n30002 ) | ( x99 & n30299 ) | ( ~n30002 & n30299 ) ;
  assign n30301 = ( x100 & ~n29994 ) | ( x100 & n30300 ) | ( ~n29994 & n30300 ) ;
  assign n30302 = ( x101 & ~n29986 ) | ( x101 & n30301 ) | ( ~n29986 & n30301 ) ;
  assign n30303 = ( x102 & ~n29978 ) | ( x102 & n30302 ) | ( ~n29978 & n30302 ) ;
  assign n30304 = ( x103 & ~n29970 ) | ( x103 & n30303 ) | ( ~n29970 & n30303 ) ;
  assign n30305 = ( x104 & ~n29962 ) | ( x104 & n30304 ) | ( ~n29962 & n30304 ) ;
  assign n30306 = ( x105 & ~n29954 ) | ( x105 & n30305 ) | ( ~n29954 & n30305 ) ;
  assign n30307 = ( x106 & ~n29946 ) | ( x106 & n30306 ) | ( ~n29946 & n30306 ) ;
  assign n30308 = ( x107 & ~n29938 ) | ( x107 & n30307 ) | ( ~n29938 & n30307 ) ;
  assign n30309 = ( x108 & ~n29930 ) | ( x108 & n30308 ) | ( ~n29930 & n30308 ) ;
  assign n30310 = ( x109 & ~n29922 ) | ( x109 & n30309 ) | ( ~n29922 & n30309 ) ;
  assign n30311 = ( x110 & ~n29914 ) | ( x110 & n30310 ) | ( ~n29914 & n30310 ) ;
  assign n30312 = ( x111 & ~n29906 ) | ( x111 & n30311 ) | ( ~n29906 & n30311 ) ;
  assign n30313 = ( x112 & ~n29898 ) | ( x112 & n30312 ) | ( ~n29898 & n30312 ) ;
  assign n30314 = ( x113 & ~n29890 ) | ( x113 & n30313 ) | ( ~n29890 & n30313 ) ;
  assign n30315 = ( x114 & ~n29880 ) | ( x114 & 1'b0 ) | ( ~n29880 & 1'b0 ) ;
  assign n30316 = ~n29878 & n30315 ;
  assign n30317 = ( n30314 & ~n29882 ) | ( n30314 & n30316 ) | ( ~n29882 & n30316 ) ;
  assign n30318 = ( n29882 & ~n12011 ) | ( n29882 & n30317 ) | ( ~n12011 & n30317 ) ;
  assign n30319 = n12011 | n30318 ;
  assign n30320 = ~n29881 |  n11560 ;
  assign n30334 = n29890 &  n30320 ;
  assign n30335 = n30319 &  n30334 ;
  assign n30321 = n30319 &  n30320 ;
  assign n30322 = x113 | n29890 ;
  assign n30323 = x113 &  n29890 ;
  assign n30324 = ( n30322 & ~n30323 ) | ( n30322 & 1'b0 ) | ( ~n30323 & 1'b0 ) ;
  assign n30337 = ( n30313 & n30321 ) | ( n30313 & n30324 ) | ( n30321 & n30324 ) ;
  assign n30336 = n30313 | n30324 ;
  assign n30338 = ( n30335 & ~n30337 ) | ( n30335 & n30336 ) | ( ~n30337 & n30336 ) ;
  assign n30326 = n11560 &  n29881 ;
  assign n30327 = n30319 &  n30326 ;
  assign n30325 = n29882 | n30316 ;
  assign n30329 = ( n30314 & n30321 ) | ( n30314 & n30325 ) | ( n30321 & n30325 ) ;
  assign n30328 = n30314 | n30325 ;
  assign n30330 = ( n30327 & ~n30329 ) | ( n30327 & n30328 ) | ( ~n30329 & n30328 ) ;
  assign n30342 = n29898 &  n30320 ;
  assign n30343 = n30319 &  n30342 ;
  assign n30331 = x112 | n29898 ;
  assign n30332 = x112 &  n29898 ;
  assign n30333 = ( n30331 & ~n30332 ) | ( n30331 & 1'b0 ) | ( ~n30332 & 1'b0 ) ;
  assign n30345 = ( n30312 & n30321 ) | ( n30312 & n30333 ) | ( n30321 & n30333 ) ;
  assign n30344 = n30312 | n30333 ;
  assign n30346 = ( n30343 & ~n30345 ) | ( n30343 & n30344 ) | ( ~n30345 & n30344 ) ;
  assign n30350 = n29906 &  n30320 ;
  assign n30351 = n30319 &  n30350 ;
  assign n30339 = x111 | n29906 ;
  assign n30340 = x111 &  n29906 ;
  assign n30341 = ( n30339 & ~n30340 ) | ( n30339 & 1'b0 ) | ( ~n30340 & 1'b0 ) ;
  assign n30353 = ( n30311 & n30321 ) | ( n30311 & n30341 ) | ( n30321 & n30341 ) ;
  assign n30352 = n30311 | n30341 ;
  assign n30354 = ( n30351 & ~n30353 ) | ( n30351 & n30352 ) | ( ~n30353 & n30352 ) ;
  assign n30358 = n29914 &  n30320 ;
  assign n30359 = n30319 &  n30358 ;
  assign n30347 = x110 | n29914 ;
  assign n30348 = x110 &  n29914 ;
  assign n30349 = ( n30347 & ~n30348 ) | ( n30347 & 1'b0 ) | ( ~n30348 & 1'b0 ) ;
  assign n30361 = ( n30310 & n30321 ) | ( n30310 & n30349 ) | ( n30321 & n30349 ) ;
  assign n30360 = n30310 | n30349 ;
  assign n30362 = ( n30359 & ~n30361 ) | ( n30359 & n30360 ) | ( ~n30361 & n30360 ) ;
  assign n30366 = n29922 &  n30320 ;
  assign n30367 = n30319 &  n30366 ;
  assign n30355 = x109 | n29922 ;
  assign n30356 = x109 &  n29922 ;
  assign n30357 = ( n30355 & ~n30356 ) | ( n30355 & 1'b0 ) | ( ~n30356 & 1'b0 ) ;
  assign n30369 = ( n30309 & n30321 ) | ( n30309 & n30357 ) | ( n30321 & n30357 ) ;
  assign n30368 = n30309 | n30357 ;
  assign n30370 = ( n30367 & ~n30369 ) | ( n30367 & n30368 ) | ( ~n30369 & n30368 ) ;
  assign n30374 = n29930 &  n30320 ;
  assign n30375 = n30319 &  n30374 ;
  assign n30363 = x108 | n29930 ;
  assign n30364 = x108 &  n29930 ;
  assign n30365 = ( n30363 & ~n30364 ) | ( n30363 & 1'b0 ) | ( ~n30364 & 1'b0 ) ;
  assign n30377 = ( n30308 & n30321 ) | ( n30308 & n30365 ) | ( n30321 & n30365 ) ;
  assign n30376 = n30308 | n30365 ;
  assign n30378 = ( n30375 & ~n30377 ) | ( n30375 & n30376 ) | ( ~n30377 & n30376 ) ;
  assign n30382 = n29938 &  n30320 ;
  assign n30383 = n30319 &  n30382 ;
  assign n30371 = x107 | n29938 ;
  assign n30372 = x107 &  n29938 ;
  assign n30373 = ( n30371 & ~n30372 ) | ( n30371 & 1'b0 ) | ( ~n30372 & 1'b0 ) ;
  assign n30385 = ( n30307 & n30321 ) | ( n30307 & n30373 ) | ( n30321 & n30373 ) ;
  assign n30384 = n30307 | n30373 ;
  assign n30386 = ( n30383 & ~n30385 ) | ( n30383 & n30384 ) | ( ~n30385 & n30384 ) ;
  assign n30390 = n29946 &  n30320 ;
  assign n30391 = n30319 &  n30390 ;
  assign n30379 = x106 | n29946 ;
  assign n30380 = x106 &  n29946 ;
  assign n30381 = ( n30379 & ~n30380 ) | ( n30379 & 1'b0 ) | ( ~n30380 & 1'b0 ) ;
  assign n30393 = ( n30306 & n30321 ) | ( n30306 & n30381 ) | ( n30321 & n30381 ) ;
  assign n30392 = n30306 | n30381 ;
  assign n30394 = ( n30391 & ~n30393 ) | ( n30391 & n30392 ) | ( ~n30393 & n30392 ) ;
  assign n30398 = n29954 &  n30320 ;
  assign n30399 = n30319 &  n30398 ;
  assign n30387 = x105 | n29954 ;
  assign n30388 = x105 &  n29954 ;
  assign n30389 = ( n30387 & ~n30388 ) | ( n30387 & 1'b0 ) | ( ~n30388 & 1'b0 ) ;
  assign n30401 = ( n30305 & n30321 ) | ( n30305 & n30389 ) | ( n30321 & n30389 ) ;
  assign n30400 = n30305 | n30389 ;
  assign n30402 = ( n30399 & ~n30401 ) | ( n30399 & n30400 ) | ( ~n30401 & n30400 ) ;
  assign n30406 = n29962 &  n30320 ;
  assign n30407 = n30319 &  n30406 ;
  assign n30395 = x104 | n29962 ;
  assign n30396 = x104 &  n29962 ;
  assign n30397 = ( n30395 & ~n30396 ) | ( n30395 & 1'b0 ) | ( ~n30396 & 1'b0 ) ;
  assign n30409 = ( n30304 & n30321 ) | ( n30304 & n30397 ) | ( n30321 & n30397 ) ;
  assign n30408 = n30304 | n30397 ;
  assign n30410 = ( n30407 & ~n30409 ) | ( n30407 & n30408 ) | ( ~n30409 & n30408 ) ;
  assign n30414 = n29970 &  n30320 ;
  assign n30415 = n30319 &  n30414 ;
  assign n30403 = x103 | n29970 ;
  assign n30404 = x103 &  n29970 ;
  assign n30405 = ( n30403 & ~n30404 ) | ( n30403 & 1'b0 ) | ( ~n30404 & 1'b0 ) ;
  assign n30417 = ( n30303 & n30321 ) | ( n30303 & n30405 ) | ( n30321 & n30405 ) ;
  assign n30416 = n30303 | n30405 ;
  assign n30418 = ( n30415 & ~n30417 ) | ( n30415 & n30416 ) | ( ~n30417 & n30416 ) ;
  assign n30422 = n29978 &  n30320 ;
  assign n30423 = n30319 &  n30422 ;
  assign n30411 = x102 | n29978 ;
  assign n30412 = x102 &  n29978 ;
  assign n30413 = ( n30411 & ~n30412 ) | ( n30411 & 1'b0 ) | ( ~n30412 & 1'b0 ) ;
  assign n30425 = ( n30302 & n30321 ) | ( n30302 & n30413 ) | ( n30321 & n30413 ) ;
  assign n30424 = n30302 | n30413 ;
  assign n30426 = ( n30423 & ~n30425 ) | ( n30423 & n30424 ) | ( ~n30425 & n30424 ) ;
  assign n30430 = n29986 &  n30320 ;
  assign n30431 = n30319 &  n30430 ;
  assign n30419 = x101 | n29986 ;
  assign n30420 = x101 &  n29986 ;
  assign n30421 = ( n30419 & ~n30420 ) | ( n30419 & 1'b0 ) | ( ~n30420 & 1'b0 ) ;
  assign n30433 = ( n30301 & n30321 ) | ( n30301 & n30421 ) | ( n30321 & n30421 ) ;
  assign n30432 = n30301 | n30421 ;
  assign n30434 = ( n30431 & ~n30433 ) | ( n30431 & n30432 ) | ( ~n30433 & n30432 ) ;
  assign n30438 = n29994 &  n30320 ;
  assign n30439 = n30319 &  n30438 ;
  assign n30427 = x100 | n29994 ;
  assign n30428 = x100 &  n29994 ;
  assign n30429 = ( n30427 & ~n30428 ) | ( n30427 & 1'b0 ) | ( ~n30428 & 1'b0 ) ;
  assign n30441 = ( n30300 & n30321 ) | ( n30300 & n30429 ) | ( n30321 & n30429 ) ;
  assign n30440 = n30300 | n30429 ;
  assign n30442 = ( n30439 & ~n30441 ) | ( n30439 & n30440 ) | ( ~n30441 & n30440 ) ;
  assign n30446 = n30002 &  n30320 ;
  assign n30447 = n30319 &  n30446 ;
  assign n30435 = x99 | n30002 ;
  assign n30436 = x99 &  n30002 ;
  assign n30437 = ( n30435 & ~n30436 ) | ( n30435 & 1'b0 ) | ( ~n30436 & 1'b0 ) ;
  assign n30449 = ( n30299 & n30321 ) | ( n30299 & n30437 ) | ( n30321 & n30437 ) ;
  assign n30448 = n30299 | n30437 ;
  assign n30450 = ( n30447 & ~n30449 ) | ( n30447 & n30448 ) | ( ~n30449 & n30448 ) ;
  assign n30454 = n30010 &  n30320 ;
  assign n30455 = n30319 &  n30454 ;
  assign n30443 = x98 | n30010 ;
  assign n30444 = x98 &  n30010 ;
  assign n30445 = ( n30443 & ~n30444 ) | ( n30443 & 1'b0 ) | ( ~n30444 & 1'b0 ) ;
  assign n30457 = ( n30298 & n30321 ) | ( n30298 & n30445 ) | ( n30321 & n30445 ) ;
  assign n30456 = n30298 | n30445 ;
  assign n30458 = ( n30455 & ~n30457 ) | ( n30455 & n30456 ) | ( ~n30457 & n30456 ) ;
  assign n30462 = n30018 &  n30320 ;
  assign n30463 = n30319 &  n30462 ;
  assign n30451 = x97 | n30018 ;
  assign n30452 = x97 &  n30018 ;
  assign n30453 = ( n30451 & ~n30452 ) | ( n30451 & 1'b0 ) | ( ~n30452 & 1'b0 ) ;
  assign n30465 = ( n30297 & n30321 ) | ( n30297 & n30453 ) | ( n30321 & n30453 ) ;
  assign n30464 = n30297 | n30453 ;
  assign n30466 = ( n30463 & ~n30465 ) | ( n30463 & n30464 ) | ( ~n30465 & n30464 ) ;
  assign n30470 = n30026 &  n30320 ;
  assign n30471 = n30319 &  n30470 ;
  assign n30459 = x96 | n30026 ;
  assign n30460 = x96 &  n30026 ;
  assign n30461 = ( n30459 & ~n30460 ) | ( n30459 & 1'b0 ) | ( ~n30460 & 1'b0 ) ;
  assign n30473 = ( n30296 & n30321 ) | ( n30296 & n30461 ) | ( n30321 & n30461 ) ;
  assign n30472 = n30296 | n30461 ;
  assign n30474 = ( n30471 & ~n30473 ) | ( n30471 & n30472 ) | ( ~n30473 & n30472 ) ;
  assign n30478 = n30034 &  n30320 ;
  assign n30479 = n30319 &  n30478 ;
  assign n30467 = x95 | n30034 ;
  assign n30468 = x95 &  n30034 ;
  assign n30469 = ( n30467 & ~n30468 ) | ( n30467 & 1'b0 ) | ( ~n30468 & 1'b0 ) ;
  assign n30481 = ( n30295 & n30321 ) | ( n30295 & n30469 ) | ( n30321 & n30469 ) ;
  assign n30480 = n30295 | n30469 ;
  assign n30482 = ( n30479 & ~n30481 ) | ( n30479 & n30480 ) | ( ~n30481 & n30480 ) ;
  assign n30486 = n30042 &  n30320 ;
  assign n30487 = n30319 &  n30486 ;
  assign n30475 = x94 | n30042 ;
  assign n30476 = x94 &  n30042 ;
  assign n30477 = ( n30475 & ~n30476 ) | ( n30475 & 1'b0 ) | ( ~n30476 & 1'b0 ) ;
  assign n30489 = ( n30294 & n30321 ) | ( n30294 & n30477 ) | ( n30321 & n30477 ) ;
  assign n30488 = n30294 | n30477 ;
  assign n30490 = ( n30487 & ~n30489 ) | ( n30487 & n30488 ) | ( ~n30489 & n30488 ) ;
  assign n30494 = n30050 &  n30320 ;
  assign n30495 = n30319 &  n30494 ;
  assign n30483 = x93 | n30050 ;
  assign n30484 = x93 &  n30050 ;
  assign n30485 = ( n30483 & ~n30484 ) | ( n30483 & 1'b0 ) | ( ~n30484 & 1'b0 ) ;
  assign n30497 = ( n30293 & n30321 ) | ( n30293 & n30485 ) | ( n30321 & n30485 ) ;
  assign n30496 = n30293 | n30485 ;
  assign n30498 = ( n30495 & ~n30497 ) | ( n30495 & n30496 ) | ( ~n30497 & n30496 ) ;
  assign n30502 = n30058 &  n30320 ;
  assign n30503 = n30319 &  n30502 ;
  assign n30491 = x92 | n30058 ;
  assign n30492 = x92 &  n30058 ;
  assign n30493 = ( n30491 & ~n30492 ) | ( n30491 & 1'b0 ) | ( ~n30492 & 1'b0 ) ;
  assign n30505 = ( n30292 & n30321 ) | ( n30292 & n30493 ) | ( n30321 & n30493 ) ;
  assign n30504 = n30292 | n30493 ;
  assign n30506 = ( n30503 & ~n30505 ) | ( n30503 & n30504 ) | ( ~n30505 & n30504 ) ;
  assign n30510 = n30066 &  n30320 ;
  assign n30511 = n30319 &  n30510 ;
  assign n30499 = x91 | n30066 ;
  assign n30500 = x91 &  n30066 ;
  assign n30501 = ( n30499 & ~n30500 ) | ( n30499 & 1'b0 ) | ( ~n30500 & 1'b0 ) ;
  assign n30513 = ( n30291 & n30321 ) | ( n30291 & n30501 ) | ( n30321 & n30501 ) ;
  assign n30512 = n30291 | n30501 ;
  assign n30514 = ( n30511 & ~n30513 ) | ( n30511 & n30512 ) | ( ~n30513 & n30512 ) ;
  assign n30518 = n30074 &  n30320 ;
  assign n30519 = n30319 &  n30518 ;
  assign n30507 = x90 | n30074 ;
  assign n30508 = x90 &  n30074 ;
  assign n30509 = ( n30507 & ~n30508 ) | ( n30507 & 1'b0 ) | ( ~n30508 & 1'b0 ) ;
  assign n30521 = ( n30290 & n30321 ) | ( n30290 & n30509 ) | ( n30321 & n30509 ) ;
  assign n30520 = n30290 | n30509 ;
  assign n30522 = ( n30519 & ~n30521 ) | ( n30519 & n30520 ) | ( ~n30521 & n30520 ) ;
  assign n30526 = n30082 &  n30320 ;
  assign n30527 = n30319 &  n30526 ;
  assign n30515 = x89 | n30082 ;
  assign n30516 = x89 &  n30082 ;
  assign n30517 = ( n30515 & ~n30516 ) | ( n30515 & 1'b0 ) | ( ~n30516 & 1'b0 ) ;
  assign n30529 = ( n30289 & n30321 ) | ( n30289 & n30517 ) | ( n30321 & n30517 ) ;
  assign n30528 = n30289 | n30517 ;
  assign n30530 = ( n30527 & ~n30529 ) | ( n30527 & n30528 ) | ( ~n30529 & n30528 ) ;
  assign n30534 = n30090 &  n30320 ;
  assign n30535 = n30319 &  n30534 ;
  assign n30523 = x88 | n30090 ;
  assign n30524 = x88 &  n30090 ;
  assign n30525 = ( n30523 & ~n30524 ) | ( n30523 & 1'b0 ) | ( ~n30524 & 1'b0 ) ;
  assign n30537 = ( n30288 & n30321 ) | ( n30288 & n30525 ) | ( n30321 & n30525 ) ;
  assign n30536 = n30288 | n30525 ;
  assign n30538 = ( n30535 & ~n30537 ) | ( n30535 & n30536 ) | ( ~n30537 & n30536 ) ;
  assign n30542 = n30098 &  n30320 ;
  assign n30543 = n30319 &  n30542 ;
  assign n30531 = x87 | n30098 ;
  assign n30532 = x87 &  n30098 ;
  assign n30533 = ( n30531 & ~n30532 ) | ( n30531 & 1'b0 ) | ( ~n30532 & 1'b0 ) ;
  assign n30545 = ( n30287 & n30321 ) | ( n30287 & n30533 ) | ( n30321 & n30533 ) ;
  assign n30544 = n30287 | n30533 ;
  assign n30546 = ( n30543 & ~n30545 ) | ( n30543 & n30544 ) | ( ~n30545 & n30544 ) ;
  assign n30550 = n30106 &  n30320 ;
  assign n30551 = n30319 &  n30550 ;
  assign n30539 = x86 | n30106 ;
  assign n30540 = x86 &  n30106 ;
  assign n30541 = ( n30539 & ~n30540 ) | ( n30539 & 1'b0 ) | ( ~n30540 & 1'b0 ) ;
  assign n30553 = ( n30286 & n30321 ) | ( n30286 & n30541 ) | ( n30321 & n30541 ) ;
  assign n30552 = n30286 | n30541 ;
  assign n30554 = ( n30551 & ~n30553 ) | ( n30551 & n30552 ) | ( ~n30553 & n30552 ) ;
  assign n30558 = n30114 &  n30320 ;
  assign n30559 = n30319 &  n30558 ;
  assign n30547 = x85 | n30114 ;
  assign n30548 = x85 &  n30114 ;
  assign n30549 = ( n30547 & ~n30548 ) | ( n30547 & 1'b0 ) | ( ~n30548 & 1'b0 ) ;
  assign n30561 = ( n30285 & n30321 ) | ( n30285 & n30549 ) | ( n30321 & n30549 ) ;
  assign n30560 = n30285 | n30549 ;
  assign n30562 = ( n30559 & ~n30561 ) | ( n30559 & n30560 ) | ( ~n30561 & n30560 ) ;
  assign n30566 = n30122 &  n30320 ;
  assign n30567 = n30319 &  n30566 ;
  assign n30555 = x84 | n30122 ;
  assign n30556 = x84 &  n30122 ;
  assign n30557 = ( n30555 & ~n30556 ) | ( n30555 & 1'b0 ) | ( ~n30556 & 1'b0 ) ;
  assign n30569 = ( n30284 & n30321 ) | ( n30284 & n30557 ) | ( n30321 & n30557 ) ;
  assign n30568 = n30284 | n30557 ;
  assign n30570 = ( n30567 & ~n30569 ) | ( n30567 & n30568 ) | ( ~n30569 & n30568 ) ;
  assign n30574 = n30130 &  n30320 ;
  assign n30575 = n30319 &  n30574 ;
  assign n30563 = x83 | n30130 ;
  assign n30564 = x83 &  n30130 ;
  assign n30565 = ( n30563 & ~n30564 ) | ( n30563 & 1'b0 ) | ( ~n30564 & 1'b0 ) ;
  assign n30577 = ( n30283 & n30321 ) | ( n30283 & n30565 ) | ( n30321 & n30565 ) ;
  assign n30576 = n30283 | n30565 ;
  assign n30578 = ( n30575 & ~n30577 ) | ( n30575 & n30576 ) | ( ~n30577 & n30576 ) ;
  assign n30582 = n30138 &  n30320 ;
  assign n30583 = n30319 &  n30582 ;
  assign n30571 = x82 | n30138 ;
  assign n30572 = x82 &  n30138 ;
  assign n30573 = ( n30571 & ~n30572 ) | ( n30571 & 1'b0 ) | ( ~n30572 & 1'b0 ) ;
  assign n30585 = ( n30282 & n30321 ) | ( n30282 & n30573 ) | ( n30321 & n30573 ) ;
  assign n30584 = n30282 | n30573 ;
  assign n30586 = ( n30583 & ~n30585 ) | ( n30583 & n30584 ) | ( ~n30585 & n30584 ) ;
  assign n30590 = n30146 &  n30320 ;
  assign n30591 = n30319 &  n30590 ;
  assign n30579 = x81 | n30146 ;
  assign n30580 = x81 &  n30146 ;
  assign n30581 = ( n30579 & ~n30580 ) | ( n30579 & 1'b0 ) | ( ~n30580 & 1'b0 ) ;
  assign n30593 = ( n30281 & n30321 ) | ( n30281 & n30581 ) | ( n30321 & n30581 ) ;
  assign n30592 = n30281 | n30581 ;
  assign n30594 = ( n30591 & ~n30593 ) | ( n30591 & n30592 ) | ( ~n30593 & n30592 ) ;
  assign n30598 = n30154 &  n30320 ;
  assign n30599 = n30319 &  n30598 ;
  assign n30587 = x80 | n30154 ;
  assign n30588 = x80 &  n30154 ;
  assign n30589 = ( n30587 & ~n30588 ) | ( n30587 & 1'b0 ) | ( ~n30588 & 1'b0 ) ;
  assign n30601 = ( n30280 & n30321 ) | ( n30280 & n30589 ) | ( n30321 & n30589 ) ;
  assign n30600 = n30280 | n30589 ;
  assign n30602 = ( n30599 & ~n30601 ) | ( n30599 & n30600 ) | ( ~n30601 & n30600 ) ;
  assign n30606 = n30162 &  n30320 ;
  assign n30607 = n30319 &  n30606 ;
  assign n30595 = x79 | n30162 ;
  assign n30596 = x79 &  n30162 ;
  assign n30597 = ( n30595 & ~n30596 ) | ( n30595 & 1'b0 ) | ( ~n30596 & 1'b0 ) ;
  assign n30609 = ( n30279 & n30321 ) | ( n30279 & n30597 ) | ( n30321 & n30597 ) ;
  assign n30608 = n30279 | n30597 ;
  assign n30610 = ( n30607 & ~n30609 ) | ( n30607 & n30608 ) | ( ~n30609 & n30608 ) ;
  assign n30614 = n30170 &  n30320 ;
  assign n30615 = n30319 &  n30614 ;
  assign n30603 = x78 | n30170 ;
  assign n30604 = x78 &  n30170 ;
  assign n30605 = ( n30603 & ~n30604 ) | ( n30603 & 1'b0 ) | ( ~n30604 & 1'b0 ) ;
  assign n30617 = ( n30278 & n30321 ) | ( n30278 & n30605 ) | ( n30321 & n30605 ) ;
  assign n30616 = n30278 | n30605 ;
  assign n30618 = ( n30615 & ~n30617 ) | ( n30615 & n30616 ) | ( ~n30617 & n30616 ) ;
  assign n30622 = n30178 &  n30320 ;
  assign n30623 = n30319 &  n30622 ;
  assign n30611 = x77 | n30178 ;
  assign n30612 = x77 &  n30178 ;
  assign n30613 = ( n30611 & ~n30612 ) | ( n30611 & 1'b0 ) | ( ~n30612 & 1'b0 ) ;
  assign n30625 = ( n30277 & n30321 ) | ( n30277 & n30613 ) | ( n30321 & n30613 ) ;
  assign n30624 = n30277 | n30613 ;
  assign n30626 = ( n30623 & ~n30625 ) | ( n30623 & n30624 ) | ( ~n30625 & n30624 ) ;
  assign n30630 = n30186 &  n30320 ;
  assign n30631 = n30319 &  n30630 ;
  assign n30619 = x76 | n30186 ;
  assign n30620 = x76 &  n30186 ;
  assign n30621 = ( n30619 & ~n30620 ) | ( n30619 & 1'b0 ) | ( ~n30620 & 1'b0 ) ;
  assign n30633 = ( n30276 & n30321 ) | ( n30276 & n30621 ) | ( n30321 & n30621 ) ;
  assign n30632 = n30276 | n30621 ;
  assign n30634 = ( n30631 & ~n30633 ) | ( n30631 & n30632 ) | ( ~n30633 & n30632 ) ;
  assign n30638 = n30194 &  n30320 ;
  assign n30639 = n30319 &  n30638 ;
  assign n30627 = x75 | n30194 ;
  assign n30628 = x75 &  n30194 ;
  assign n30629 = ( n30627 & ~n30628 ) | ( n30627 & 1'b0 ) | ( ~n30628 & 1'b0 ) ;
  assign n30641 = ( n30275 & n30321 ) | ( n30275 & n30629 ) | ( n30321 & n30629 ) ;
  assign n30640 = n30275 | n30629 ;
  assign n30642 = ( n30639 & ~n30641 ) | ( n30639 & n30640 ) | ( ~n30641 & n30640 ) ;
  assign n30646 = n30202 &  n30320 ;
  assign n30647 = n30319 &  n30646 ;
  assign n30635 = x74 | n30202 ;
  assign n30636 = x74 &  n30202 ;
  assign n30637 = ( n30635 & ~n30636 ) | ( n30635 & 1'b0 ) | ( ~n30636 & 1'b0 ) ;
  assign n30649 = ( n30274 & n30321 ) | ( n30274 & n30637 ) | ( n30321 & n30637 ) ;
  assign n30648 = n30274 | n30637 ;
  assign n30650 = ( n30647 & ~n30649 ) | ( n30647 & n30648 ) | ( ~n30649 & n30648 ) ;
  assign n30654 = n30210 &  n30320 ;
  assign n30655 = n30319 &  n30654 ;
  assign n30643 = x73 | n30210 ;
  assign n30644 = x73 &  n30210 ;
  assign n30645 = ( n30643 & ~n30644 ) | ( n30643 & 1'b0 ) | ( ~n30644 & 1'b0 ) ;
  assign n30657 = ( n30273 & n30321 ) | ( n30273 & n30645 ) | ( n30321 & n30645 ) ;
  assign n30656 = n30273 | n30645 ;
  assign n30658 = ( n30655 & ~n30657 ) | ( n30655 & n30656 ) | ( ~n30657 & n30656 ) ;
  assign n30662 = n30218 &  n30320 ;
  assign n30663 = n30319 &  n30662 ;
  assign n30651 = x72 | n30218 ;
  assign n30652 = x72 &  n30218 ;
  assign n30653 = ( n30651 & ~n30652 ) | ( n30651 & 1'b0 ) | ( ~n30652 & 1'b0 ) ;
  assign n30665 = ( n30272 & n30321 ) | ( n30272 & n30653 ) | ( n30321 & n30653 ) ;
  assign n30664 = n30272 | n30653 ;
  assign n30666 = ( n30663 & ~n30665 ) | ( n30663 & n30664 ) | ( ~n30665 & n30664 ) ;
  assign n30670 = n30226 &  n30320 ;
  assign n30671 = n30319 &  n30670 ;
  assign n30659 = x71 | n30226 ;
  assign n30660 = x71 &  n30226 ;
  assign n30661 = ( n30659 & ~n30660 ) | ( n30659 & 1'b0 ) | ( ~n30660 & 1'b0 ) ;
  assign n30673 = ( n30271 & n30321 ) | ( n30271 & n30661 ) | ( n30321 & n30661 ) ;
  assign n30672 = n30271 | n30661 ;
  assign n30674 = ( n30671 & ~n30673 ) | ( n30671 & n30672 ) | ( ~n30673 & n30672 ) ;
  assign n30678 = n30234 &  n30320 ;
  assign n30679 = n30319 &  n30678 ;
  assign n30667 = x70 | n30234 ;
  assign n30668 = x70 &  n30234 ;
  assign n30669 = ( n30667 & ~n30668 ) | ( n30667 & 1'b0 ) | ( ~n30668 & 1'b0 ) ;
  assign n30681 = ( n30270 & n30321 ) | ( n30270 & n30669 ) | ( n30321 & n30669 ) ;
  assign n30680 = n30270 | n30669 ;
  assign n30682 = ( n30679 & ~n30681 ) | ( n30679 & n30680 ) | ( ~n30681 & n30680 ) ;
  assign n30686 = n30242 &  n30320 ;
  assign n30687 = n30319 &  n30686 ;
  assign n30675 = x69 | n30242 ;
  assign n30676 = x69 &  n30242 ;
  assign n30677 = ( n30675 & ~n30676 ) | ( n30675 & 1'b0 ) | ( ~n30676 & 1'b0 ) ;
  assign n30689 = ( n30269 & n30321 ) | ( n30269 & n30677 ) | ( n30321 & n30677 ) ;
  assign n30688 = n30269 | n30677 ;
  assign n30690 = ( n30687 & ~n30689 ) | ( n30687 & n30688 ) | ( ~n30689 & n30688 ) ;
  assign n30694 = n30250 &  n30320 ;
  assign n30695 = n30319 &  n30694 ;
  assign n30683 = x68 | n30250 ;
  assign n30684 = x68 &  n30250 ;
  assign n30685 = ( n30683 & ~n30684 ) | ( n30683 & 1'b0 ) | ( ~n30684 & 1'b0 ) ;
  assign n30697 = ( n30268 & n30321 ) | ( n30268 & n30685 ) | ( n30321 & n30685 ) ;
  assign n30696 = n30268 | n30685 ;
  assign n30698 = ( n30695 & ~n30697 ) | ( n30695 & n30696 ) | ( ~n30697 & n30696 ) ;
  assign n30702 = n30255 &  n30320 ;
  assign n30703 = n30319 &  n30702 ;
  assign n30691 = x67 | n30255 ;
  assign n30692 = x67 &  n30255 ;
  assign n30693 = ( n30691 & ~n30692 ) | ( n30691 & 1'b0 ) | ( ~n30692 & 1'b0 ) ;
  assign n30705 = ( n30267 & n30321 ) | ( n30267 & n30693 ) | ( n30321 & n30693 ) ;
  assign n30704 = n30267 | n30693 ;
  assign n30706 = ( n30703 & ~n30705 ) | ( n30703 & n30704 ) | ( ~n30705 & n30704 ) ;
  assign n30707 = n30261 &  n30320 ;
  assign n30708 = n30319 &  n30707 ;
  assign n30699 = x66 | n30261 ;
  assign n30700 = x66 &  n30261 ;
  assign n30701 = ( n30699 & ~n30700 ) | ( n30699 & 1'b0 ) | ( ~n30700 & 1'b0 ) ;
  assign n30709 = n30266 &  n30701 ;
  assign n30710 = ( n30266 & ~n30321 ) | ( n30266 & n30701 ) | ( ~n30321 & n30701 ) ;
  assign n30711 = ( n30708 & ~n30709 ) | ( n30708 & n30710 ) | ( ~n30709 & n30710 ) ;
  assign n30712 = ( x65 & ~n11875 ) | ( x65 & n30265 ) | ( ~n11875 & n30265 ) ;
  assign n30713 = ( n30266 & ~x65 ) | ( n30266 & n30712 ) | ( ~x65 & n30712 ) ;
  assign n30714 = ~n30321 & n30713 ;
  assign n30715 = n30265 &  n30320 ;
  assign n30716 = n30319 &  n30715 ;
  assign n30717 = n30714 | n30716 ;
  assign n30718 = ( x64 & ~n30321 ) | ( x64 & 1'b0 ) | ( ~n30321 & 1'b0 ) ;
  assign n30719 = ( x13 & ~n30718 ) | ( x13 & 1'b0 ) | ( ~n30718 & 1'b0 ) ;
  assign n30720 = ( n11875 & ~n30321 ) | ( n11875 & 1'b0 ) | ( ~n30321 & 1'b0 ) ;
  assign n30721 = n30719 | n30720 ;
  assign n30722 = ( x65 & ~n30721 ) | ( x65 & n12413 ) | ( ~n30721 & n12413 ) ;
  assign n30723 = ( x66 & ~n30717 ) | ( x66 & n30722 ) | ( ~n30717 & n30722 ) ;
  assign n30724 = ( x67 & ~n30711 ) | ( x67 & n30723 ) | ( ~n30711 & n30723 ) ;
  assign n30725 = ( x68 & ~n30706 ) | ( x68 & n30724 ) | ( ~n30706 & n30724 ) ;
  assign n30726 = ( x69 & ~n30698 ) | ( x69 & n30725 ) | ( ~n30698 & n30725 ) ;
  assign n30727 = ( x70 & ~n30690 ) | ( x70 & n30726 ) | ( ~n30690 & n30726 ) ;
  assign n30728 = ( x71 & ~n30682 ) | ( x71 & n30727 ) | ( ~n30682 & n30727 ) ;
  assign n30729 = ( x72 & ~n30674 ) | ( x72 & n30728 ) | ( ~n30674 & n30728 ) ;
  assign n30730 = ( x73 & ~n30666 ) | ( x73 & n30729 ) | ( ~n30666 & n30729 ) ;
  assign n30731 = ( x74 & ~n30658 ) | ( x74 & n30730 ) | ( ~n30658 & n30730 ) ;
  assign n30732 = ( x75 & ~n30650 ) | ( x75 & n30731 ) | ( ~n30650 & n30731 ) ;
  assign n30733 = ( x76 & ~n30642 ) | ( x76 & n30732 ) | ( ~n30642 & n30732 ) ;
  assign n30734 = ( x77 & ~n30634 ) | ( x77 & n30733 ) | ( ~n30634 & n30733 ) ;
  assign n30735 = ( x78 & ~n30626 ) | ( x78 & n30734 ) | ( ~n30626 & n30734 ) ;
  assign n30736 = ( x79 & ~n30618 ) | ( x79 & n30735 ) | ( ~n30618 & n30735 ) ;
  assign n30737 = ( x80 & ~n30610 ) | ( x80 & n30736 ) | ( ~n30610 & n30736 ) ;
  assign n30738 = ( x81 & ~n30602 ) | ( x81 & n30737 ) | ( ~n30602 & n30737 ) ;
  assign n30739 = ( x82 & ~n30594 ) | ( x82 & n30738 ) | ( ~n30594 & n30738 ) ;
  assign n30740 = ( x83 & ~n30586 ) | ( x83 & n30739 ) | ( ~n30586 & n30739 ) ;
  assign n30741 = ( x84 & ~n30578 ) | ( x84 & n30740 ) | ( ~n30578 & n30740 ) ;
  assign n30742 = ( x85 & ~n30570 ) | ( x85 & n30741 ) | ( ~n30570 & n30741 ) ;
  assign n30743 = ( x86 & ~n30562 ) | ( x86 & n30742 ) | ( ~n30562 & n30742 ) ;
  assign n30744 = ( x87 & ~n30554 ) | ( x87 & n30743 ) | ( ~n30554 & n30743 ) ;
  assign n30745 = ( x88 & ~n30546 ) | ( x88 & n30744 ) | ( ~n30546 & n30744 ) ;
  assign n30746 = ( x89 & ~n30538 ) | ( x89 & n30745 ) | ( ~n30538 & n30745 ) ;
  assign n30747 = ( x90 & ~n30530 ) | ( x90 & n30746 ) | ( ~n30530 & n30746 ) ;
  assign n30748 = ( x91 & ~n30522 ) | ( x91 & n30747 ) | ( ~n30522 & n30747 ) ;
  assign n30749 = ( x92 & ~n30514 ) | ( x92 & n30748 ) | ( ~n30514 & n30748 ) ;
  assign n30750 = ( x93 & ~n30506 ) | ( x93 & n30749 ) | ( ~n30506 & n30749 ) ;
  assign n30751 = ( x94 & ~n30498 ) | ( x94 & n30750 ) | ( ~n30498 & n30750 ) ;
  assign n30752 = ( x95 & ~n30490 ) | ( x95 & n30751 ) | ( ~n30490 & n30751 ) ;
  assign n30753 = ( x96 & ~n30482 ) | ( x96 & n30752 ) | ( ~n30482 & n30752 ) ;
  assign n30754 = ( x97 & ~n30474 ) | ( x97 & n30753 ) | ( ~n30474 & n30753 ) ;
  assign n30755 = ( x98 & ~n30466 ) | ( x98 & n30754 ) | ( ~n30466 & n30754 ) ;
  assign n30756 = ( x99 & ~n30458 ) | ( x99 & n30755 ) | ( ~n30458 & n30755 ) ;
  assign n30757 = ( x100 & ~n30450 ) | ( x100 & n30756 ) | ( ~n30450 & n30756 ) ;
  assign n30758 = ( x101 & ~n30442 ) | ( x101 & n30757 ) | ( ~n30442 & n30757 ) ;
  assign n30759 = ( x102 & ~n30434 ) | ( x102 & n30758 ) | ( ~n30434 & n30758 ) ;
  assign n30760 = ( x103 & ~n30426 ) | ( x103 & n30759 ) | ( ~n30426 & n30759 ) ;
  assign n30761 = ( x104 & ~n30418 ) | ( x104 & n30760 ) | ( ~n30418 & n30760 ) ;
  assign n30762 = ( x105 & ~n30410 ) | ( x105 & n30761 ) | ( ~n30410 & n30761 ) ;
  assign n30763 = ( x106 & ~n30402 ) | ( x106 & n30762 ) | ( ~n30402 & n30762 ) ;
  assign n30764 = ( x107 & ~n30394 ) | ( x107 & n30763 ) | ( ~n30394 & n30763 ) ;
  assign n30765 = ( x108 & ~n30386 ) | ( x108 & n30764 ) | ( ~n30386 & n30764 ) ;
  assign n30766 = ( x109 & ~n30378 ) | ( x109 & n30765 ) | ( ~n30378 & n30765 ) ;
  assign n30767 = ( x110 & ~n30370 ) | ( x110 & n30766 ) | ( ~n30370 & n30766 ) ;
  assign n30768 = ( x111 & ~n30362 ) | ( x111 & n30767 ) | ( ~n30362 & n30767 ) ;
  assign n30769 = ( x112 & ~n30354 ) | ( x112 & n30768 ) | ( ~n30354 & n30768 ) ;
  assign n30770 = ( x113 & ~n30346 ) | ( x113 & n30769 ) | ( ~n30346 & n30769 ) ;
  assign n30771 = ( x114 & ~n30338 ) | ( x114 & n30770 ) | ( ~n30338 & n30770 ) ;
  assign n30772 = ( x115 & ~n30330 ) | ( x115 & n30771 ) | ( ~n30330 & n30771 ) ;
  assign n30773 = n160 | n30772 ;
  assign n30783 = n30338 &  n30773 ;
  assign n30775 = x114 | n30338 ;
  assign n30776 = x114 &  n30338 ;
  assign n30777 = ( n30775 & ~n30776 ) | ( n30775 & 1'b0 ) | ( ~n30776 & 1'b0 ) ;
  assign n30787 = ( n160 & n30770 ) | ( n160 & n30777 ) | ( n30770 & n30777 ) ;
  assign n30788 = ( n30770 & ~n30772 ) | ( n30770 & n30777 ) | ( ~n30772 & n30777 ) ;
  assign n30789 = ~n30787 & n30788 ;
  assign n30790 = n30783 | n30789 ;
  assign n30791 = n30346 &  n30773 ;
  assign n30784 = x113 | n30346 ;
  assign n30785 = x113 &  n30346 ;
  assign n30786 = ( n30784 & ~n30785 ) | ( n30784 & 1'b0 ) | ( ~n30785 & 1'b0 ) ;
  assign n30795 = ( n160 & n30769 ) | ( n160 & n30786 ) | ( n30769 & n30786 ) ;
  assign n30796 = ( n30769 & ~n30772 ) | ( n30769 & n30786 ) | ( ~n30772 & n30786 ) ;
  assign n30797 = ~n30795 & n30796 ;
  assign n30798 = n30791 | n30797 ;
  assign n30799 = n30354 &  n30773 ;
  assign n30792 = x112 | n30354 ;
  assign n30793 = x112 &  n30354 ;
  assign n30794 = ( n30792 & ~n30793 ) | ( n30792 & 1'b0 ) | ( ~n30793 & 1'b0 ) ;
  assign n30803 = ( n160 & n30768 ) | ( n160 & n30794 ) | ( n30768 & n30794 ) ;
  assign n30804 = ( n30768 & ~n30772 ) | ( n30768 & n30794 ) | ( ~n30772 & n30794 ) ;
  assign n30805 = ~n30803 & n30804 ;
  assign n30806 = n30799 | n30805 ;
  assign n30807 = n30362 &  n30773 ;
  assign n30800 = x111 | n30362 ;
  assign n30801 = x111 &  n30362 ;
  assign n30802 = ( n30800 & ~n30801 ) | ( n30800 & 1'b0 ) | ( ~n30801 & 1'b0 ) ;
  assign n30811 = ( n160 & n30767 ) | ( n160 & n30802 ) | ( n30767 & n30802 ) ;
  assign n30812 = ( n30767 & ~n30772 ) | ( n30767 & n30802 ) | ( ~n30772 & n30802 ) ;
  assign n30813 = ~n30811 & n30812 ;
  assign n30814 = n30807 | n30813 ;
  assign n30815 = n30370 &  n30773 ;
  assign n30808 = x110 | n30370 ;
  assign n30809 = x110 &  n30370 ;
  assign n30810 = ( n30808 & ~n30809 ) | ( n30808 & 1'b0 ) | ( ~n30809 & 1'b0 ) ;
  assign n30819 = ( n160 & n30766 ) | ( n160 & n30810 ) | ( n30766 & n30810 ) ;
  assign n30820 = ( n30766 & ~n30772 ) | ( n30766 & n30810 ) | ( ~n30772 & n30810 ) ;
  assign n30821 = ~n30819 & n30820 ;
  assign n30822 = n30815 | n30821 ;
  assign n30823 = n30378 &  n30773 ;
  assign n30816 = x109 | n30378 ;
  assign n30817 = x109 &  n30378 ;
  assign n30818 = ( n30816 & ~n30817 ) | ( n30816 & 1'b0 ) | ( ~n30817 & 1'b0 ) ;
  assign n30827 = ( n160 & n30765 ) | ( n160 & n30818 ) | ( n30765 & n30818 ) ;
  assign n30828 = ( n30765 & ~n30772 ) | ( n30765 & n30818 ) | ( ~n30772 & n30818 ) ;
  assign n30829 = ~n30827 & n30828 ;
  assign n30830 = n30823 | n30829 ;
  assign n30831 = n30386 &  n30773 ;
  assign n30824 = x108 | n30386 ;
  assign n30825 = x108 &  n30386 ;
  assign n30826 = ( n30824 & ~n30825 ) | ( n30824 & 1'b0 ) | ( ~n30825 & 1'b0 ) ;
  assign n30835 = ( n160 & n30764 ) | ( n160 & n30826 ) | ( n30764 & n30826 ) ;
  assign n30836 = ( n30764 & ~n30772 ) | ( n30764 & n30826 ) | ( ~n30772 & n30826 ) ;
  assign n30837 = ~n30835 & n30836 ;
  assign n30838 = n30831 | n30837 ;
  assign n30839 = n30394 &  n30773 ;
  assign n30832 = x107 | n30394 ;
  assign n30833 = x107 &  n30394 ;
  assign n30834 = ( n30832 & ~n30833 ) | ( n30832 & 1'b0 ) | ( ~n30833 & 1'b0 ) ;
  assign n30843 = ( n160 & n30763 ) | ( n160 & n30834 ) | ( n30763 & n30834 ) ;
  assign n30844 = ( n30763 & ~n30772 ) | ( n30763 & n30834 ) | ( ~n30772 & n30834 ) ;
  assign n30845 = ~n30843 & n30844 ;
  assign n30846 = n30839 | n30845 ;
  assign n30847 = n30402 &  n30773 ;
  assign n30840 = x106 | n30402 ;
  assign n30841 = x106 &  n30402 ;
  assign n30842 = ( n30840 & ~n30841 ) | ( n30840 & 1'b0 ) | ( ~n30841 & 1'b0 ) ;
  assign n30851 = ( n160 & n30762 ) | ( n160 & n30842 ) | ( n30762 & n30842 ) ;
  assign n30852 = ( n30762 & ~n30772 ) | ( n30762 & n30842 ) | ( ~n30772 & n30842 ) ;
  assign n30853 = ~n30851 & n30852 ;
  assign n30854 = n30847 | n30853 ;
  assign n30855 = n30410 &  n30773 ;
  assign n30848 = x105 | n30410 ;
  assign n30849 = x105 &  n30410 ;
  assign n30850 = ( n30848 & ~n30849 ) | ( n30848 & 1'b0 ) | ( ~n30849 & 1'b0 ) ;
  assign n30859 = ( n160 & n30761 ) | ( n160 & n30850 ) | ( n30761 & n30850 ) ;
  assign n30860 = ( n30761 & ~n30772 ) | ( n30761 & n30850 ) | ( ~n30772 & n30850 ) ;
  assign n30861 = ~n30859 & n30860 ;
  assign n30862 = n30855 | n30861 ;
  assign n30863 = n30418 &  n30773 ;
  assign n30856 = x104 | n30418 ;
  assign n30857 = x104 &  n30418 ;
  assign n30858 = ( n30856 & ~n30857 ) | ( n30856 & 1'b0 ) | ( ~n30857 & 1'b0 ) ;
  assign n30867 = ( n160 & n30760 ) | ( n160 & n30858 ) | ( n30760 & n30858 ) ;
  assign n30868 = ( n30760 & ~n30772 ) | ( n30760 & n30858 ) | ( ~n30772 & n30858 ) ;
  assign n30869 = ~n30867 & n30868 ;
  assign n30870 = n30863 | n30869 ;
  assign n30871 = n30426 &  n30773 ;
  assign n30864 = x103 | n30426 ;
  assign n30865 = x103 &  n30426 ;
  assign n30866 = ( n30864 & ~n30865 ) | ( n30864 & 1'b0 ) | ( ~n30865 & 1'b0 ) ;
  assign n30875 = ( n160 & n30759 ) | ( n160 & n30866 ) | ( n30759 & n30866 ) ;
  assign n30876 = ( n30759 & ~n30772 ) | ( n30759 & n30866 ) | ( ~n30772 & n30866 ) ;
  assign n30877 = ~n30875 & n30876 ;
  assign n30878 = n30871 | n30877 ;
  assign n30879 = n30434 &  n30773 ;
  assign n30872 = x102 | n30434 ;
  assign n30873 = x102 &  n30434 ;
  assign n30874 = ( n30872 & ~n30873 ) | ( n30872 & 1'b0 ) | ( ~n30873 & 1'b0 ) ;
  assign n30883 = ( n160 & n30758 ) | ( n160 & n30874 ) | ( n30758 & n30874 ) ;
  assign n30884 = ( n30758 & ~n30772 ) | ( n30758 & n30874 ) | ( ~n30772 & n30874 ) ;
  assign n30885 = ~n30883 & n30884 ;
  assign n30886 = n30879 | n30885 ;
  assign n30887 = n30442 &  n30773 ;
  assign n30880 = x101 | n30442 ;
  assign n30881 = x101 &  n30442 ;
  assign n30882 = ( n30880 & ~n30881 ) | ( n30880 & 1'b0 ) | ( ~n30881 & 1'b0 ) ;
  assign n30891 = ( n160 & n30757 ) | ( n160 & n30882 ) | ( n30757 & n30882 ) ;
  assign n30892 = ( n30757 & ~n30772 ) | ( n30757 & n30882 ) | ( ~n30772 & n30882 ) ;
  assign n30893 = ~n30891 & n30892 ;
  assign n30894 = n30887 | n30893 ;
  assign n30895 = n30450 &  n30773 ;
  assign n30888 = x100 | n30450 ;
  assign n30889 = x100 &  n30450 ;
  assign n30890 = ( n30888 & ~n30889 ) | ( n30888 & 1'b0 ) | ( ~n30889 & 1'b0 ) ;
  assign n30899 = ( n160 & n30756 ) | ( n160 & n30890 ) | ( n30756 & n30890 ) ;
  assign n30900 = ( n30756 & ~n30772 ) | ( n30756 & n30890 ) | ( ~n30772 & n30890 ) ;
  assign n30901 = ~n30899 & n30900 ;
  assign n30902 = n30895 | n30901 ;
  assign n30903 = n30458 &  n30773 ;
  assign n30896 = x99 | n30458 ;
  assign n30897 = x99 &  n30458 ;
  assign n30898 = ( n30896 & ~n30897 ) | ( n30896 & 1'b0 ) | ( ~n30897 & 1'b0 ) ;
  assign n30907 = ( n160 & n30755 ) | ( n160 & n30898 ) | ( n30755 & n30898 ) ;
  assign n30908 = ( n30755 & ~n30772 ) | ( n30755 & n30898 ) | ( ~n30772 & n30898 ) ;
  assign n30909 = ~n30907 & n30908 ;
  assign n30910 = n30903 | n30909 ;
  assign n30911 = n30466 &  n30773 ;
  assign n30904 = x98 | n30466 ;
  assign n30905 = x98 &  n30466 ;
  assign n30906 = ( n30904 & ~n30905 ) | ( n30904 & 1'b0 ) | ( ~n30905 & 1'b0 ) ;
  assign n30915 = ( n160 & n30754 ) | ( n160 & n30906 ) | ( n30754 & n30906 ) ;
  assign n30916 = ( n30754 & ~n30772 ) | ( n30754 & n30906 ) | ( ~n30772 & n30906 ) ;
  assign n30917 = ~n30915 & n30916 ;
  assign n30918 = n30911 | n30917 ;
  assign n30919 = n30474 &  n30773 ;
  assign n30912 = x97 | n30474 ;
  assign n30913 = x97 &  n30474 ;
  assign n30914 = ( n30912 & ~n30913 ) | ( n30912 & 1'b0 ) | ( ~n30913 & 1'b0 ) ;
  assign n30923 = ( n160 & n30753 ) | ( n160 & n30914 ) | ( n30753 & n30914 ) ;
  assign n30924 = ( n30753 & ~n30772 ) | ( n30753 & n30914 ) | ( ~n30772 & n30914 ) ;
  assign n30925 = ~n30923 & n30924 ;
  assign n30926 = n30919 | n30925 ;
  assign n30927 = n30482 &  n30773 ;
  assign n30920 = x96 | n30482 ;
  assign n30921 = x96 &  n30482 ;
  assign n30922 = ( n30920 & ~n30921 ) | ( n30920 & 1'b0 ) | ( ~n30921 & 1'b0 ) ;
  assign n30931 = ( n160 & n30752 ) | ( n160 & n30922 ) | ( n30752 & n30922 ) ;
  assign n30932 = ( n30752 & ~n30772 ) | ( n30752 & n30922 ) | ( ~n30772 & n30922 ) ;
  assign n30933 = ~n30931 & n30932 ;
  assign n30934 = n30927 | n30933 ;
  assign n30935 = n30490 &  n30773 ;
  assign n30928 = x95 | n30490 ;
  assign n30929 = x95 &  n30490 ;
  assign n30930 = ( n30928 & ~n30929 ) | ( n30928 & 1'b0 ) | ( ~n30929 & 1'b0 ) ;
  assign n30939 = ( n160 & n30751 ) | ( n160 & n30930 ) | ( n30751 & n30930 ) ;
  assign n30940 = ( n30751 & ~n30772 ) | ( n30751 & n30930 ) | ( ~n30772 & n30930 ) ;
  assign n30941 = ~n30939 & n30940 ;
  assign n30942 = n30935 | n30941 ;
  assign n30943 = n30498 &  n30773 ;
  assign n30936 = x94 | n30498 ;
  assign n30937 = x94 &  n30498 ;
  assign n30938 = ( n30936 & ~n30937 ) | ( n30936 & 1'b0 ) | ( ~n30937 & 1'b0 ) ;
  assign n30947 = ( n160 & n30750 ) | ( n160 & n30938 ) | ( n30750 & n30938 ) ;
  assign n30948 = ( n30750 & ~n30772 ) | ( n30750 & n30938 ) | ( ~n30772 & n30938 ) ;
  assign n30949 = ~n30947 & n30948 ;
  assign n30950 = n30943 | n30949 ;
  assign n30951 = n30506 &  n30773 ;
  assign n30944 = x93 | n30506 ;
  assign n30945 = x93 &  n30506 ;
  assign n30946 = ( n30944 & ~n30945 ) | ( n30944 & 1'b0 ) | ( ~n30945 & 1'b0 ) ;
  assign n30955 = ( n160 & n30749 ) | ( n160 & n30946 ) | ( n30749 & n30946 ) ;
  assign n30956 = ( n30749 & ~n30772 ) | ( n30749 & n30946 ) | ( ~n30772 & n30946 ) ;
  assign n30957 = ~n30955 & n30956 ;
  assign n30958 = n30951 | n30957 ;
  assign n30959 = n30514 &  n30773 ;
  assign n30952 = x92 | n30514 ;
  assign n30953 = x92 &  n30514 ;
  assign n30954 = ( n30952 & ~n30953 ) | ( n30952 & 1'b0 ) | ( ~n30953 & 1'b0 ) ;
  assign n30963 = ( n160 & n30748 ) | ( n160 & n30954 ) | ( n30748 & n30954 ) ;
  assign n30964 = ( n30748 & ~n30772 ) | ( n30748 & n30954 ) | ( ~n30772 & n30954 ) ;
  assign n30965 = ~n30963 & n30964 ;
  assign n30966 = n30959 | n30965 ;
  assign n30967 = n30522 &  n30773 ;
  assign n30960 = x91 | n30522 ;
  assign n30961 = x91 &  n30522 ;
  assign n30962 = ( n30960 & ~n30961 ) | ( n30960 & 1'b0 ) | ( ~n30961 & 1'b0 ) ;
  assign n30971 = ( n160 & n30747 ) | ( n160 & n30962 ) | ( n30747 & n30962 ) ;
  assign n30972 = ( n30747 & ~n30772 ) | ( n30747 & n30962 ) | ( ~n30772 & n30962 ) ;
  assign n30973 = ~n30971 & n30972 ;
  assign n30974 = n30967 | n30973 ;
  assign n30975 = n30530 &  n30773 ;
  assign n30968 = x90 | n30530 ;
  assign n30969 = x90 &  n30530 ;
  assign n30970 = ( n30968 & ~n30969 ) | ( n30968 & 1'b0 ) | ( ~n30969 & 1'b0 ) ;
  assign n30979 = ( n160 & n30746 ) | ( n160 & n30970 ) | ( n30746 & n30970 ) ;
  assign n30980 = ( n30746 & ~n30772 ) | ( n30746 & n30970 ) | ( ~n30772 & n30970 ) ;
  assign n30981 = ~n30979 & n30980 ;
  assign n30982 = n30975 | n30981 ;
  assign n30983 = n30538 &  n30773 ;
  assign n30976 = x89 | n30538 ;
  assign n30977 = x89 &  n30538 ;
  assign n30978 = ( n30976 & ~n30977 ) | ( n30976 & 1'b0 ) | ( ~n30977 & 1'b0 ) ;
  assign n30987 = ( n160 & n30745 ) | ( n160 & n30978 ) | ( n30745 & n30978 ) ;
  assign n30988 = ( n30745 & ~n30772 ) | ( n30745 & n30978 ) | ( ~n30772 & n30978 ) ;
  assign n30989 = ~n30987 & n30988 ;
  assign n30990 = n30983 | n30989 ;
  assign n30991 = n30546 &  n30773 ;
  assign n30984 = x88 | n30546 ;
  assign n30985 = x88 &  n30546 ;
  assign n30986 = ( n30984 & ~n30985 ) | ( n30984 & 1'b0 ) | ( ~n30985 & 1'b0 ) ;
  assign n30995 = ( n160 & n30744 ) | ( n160 & n30986 ) | ( n30744 & n30986 ) ;
  assign n30996 = ( n30744 & ~n30772 ) | ( n30744 & n30986 ) | ( ~n30772 & n30986 ) ;
  assign n30997 = ~n30995 & n30996 ;
  assign n30998 = n30991 | n30997 ;
  assign n30999 = n30554 &  n30773 ;
  assign n30992 = x87 | n30554 ;
  assign n30993 = x87 &  n30554 ;
  assign n30994 = ( n30992 & ~n30993 ) | ( n30992 & 1'b0 ) | ( ~n30993 & 1'b0 ) ;
  assign n31003 = ( n160 & n30743 ) | ( n160 & n30994 ) | ( n30743 & n30994 ) ;
  assign n31004 = ( n30743 & ~n30772 ) | ( n30743 & n30994 ) | ( ~n30772 & n30994 ) ;
  assign n31005 = ~n31003 & n31004 ;
  assign n31006 = n30999 | n31005 ;
  assign n31007 = n30562 &  n30773 ;
  assign n31000 = x86 | n30562 ;
  assign n31001 = x86 &  n30562 ;
  assign n31002 = ( n31000 & ~n31001 ) | ( n31000 & 1'b0 ) | ( ~n31001 & 1'b0 ) ;
  assign n31011 = ( n160 & n30742 ) | ( n160 & n31002 ) | ( n30742 & n31002 ) ;
  assign n31012 = ( n30742 & ~n30772 ) | ( n30742 & n31002 ) | ( ~n30772 & n31002 ) ;
  assign n31013 = ~n31011 & n31012 ;
  assign n31014 = n31007 | n31013 ;
  assign n31015 = n30570 &  n30773 ;
  assign n31008 = x85 | n30570 ;
  assign n31009 = x85 &  n30570 ;
  assign n31010 = ( n31008 & ~n31009 ) | ( n31008 & 1'b0 ) | ( ~n31009 & 1'b0 ) ;
  assign n31019 = ( n160 & n30741 ) | ( n160 & n31010 ) | ( n30741 & n31010 ) ;
  assign n31020 = ( n30741 & ~n30772 ) | ( n30741 & n31010 ) | ( ~n30772 & n31010 ) ;
  assign n31021 = ~n31019 & n31020 ;
  assign n31022 = n31015 | n31021 ;
  assign n31023 = n30578 &  n30773 ;
  assign n31016 = x84 | n30578 ;
  assign n31017 = x84 &  n30578 ;
  assign n31018 = ( n31016 & ~n31017 ) | ( n31016 & 1'b0 ) | ( ~n31017 & 1'b0 ) ;
  assign n31027 = ( n160 & n30740 ) | ( n160 & n31018 ) | ( n30740 & n31018 ) ;
  assign n31028 = ( n30740 & ~n30772 ) | ( n30740 & n31018 ) | ( ~n30772 & n31018 ) ;
  assign n31029 = ~n31027 & n31028 ;
  assign n31030 = n31023 | n31029 ;
  assign n31031 = n30586 &  n30773 ;
  assign n31024 = x83 | n30586 ;
  assign n31025 = x83 &  n30586 ;
  assign n31026 = ( n31024 & ~n31025 ) | ( n31024 & 1'b0 ) | ( ~n31025 & 1'b0 ) ;
  assign n31035 = ( n160 & n30739 ) | ( n160 & n31026 ) | ( n30739 & n31026 ) ;
  assign n31036 = ( n30739 & ~n30772 ) | ( n30739 & n31026 ) | ( ~n30772 & n31026 ) ;
  assign n31037 = ~n31035 & n31036 ;
  assign n31038 = n31031 | n31037 ;
  assign n31039 = n30594 &  n30773 ;
  assign n31032 = x82 | n30594 ;
  assign n31033 = x82 &  n30594 ;
  assign n31034 = ( n31032 & ~n31033 ) | ( n31032 & 1'b0 ) | ( ~n31033 & 1'b0 ) ;
  assign n31043 = ( n160 & n30738 ) | ( n160 & n31034 ) | ( n30738 & n31034 ) ;
  assign n31044 = ( n30738 & ~n30772 ) | ( n30738 & n31034 ) | ( ~n30772 & n31034 ) ;
  assign n31045 = ~n31043 & n31044 ;
  assign n31046 = n31039 | n31045 ;
  assign n31047 = n30602 &  n30773 ;
  assign n31040 = x81 | n30602 ;
  assign n31041 = x81 &  n30602 ;
  assign n31042 = ( n31040 & ~n31041 ) | ( n31040 & 1'b0 ) | ( ~n31041 & 1'b0 ) ;
  assign n31051 = ( n160 & n30737 ) | ( n160 & n31042 ) | ( n30737 & n31042 ) ;
  assign n31052 = ( n30737 & ~n30772 ) | ( n30737 & n31042 ) | ( ~n30772 & n31042 ) ;
  assign n31053 = ~n31051 & n31052 ;
  assign n31054 = n31047 | n31053 ;
  assign n31055 = n30610 &  n30773 ;
  assign n31048 = x80 | n30610 ;
  assign n31049 = x80 &  n30610 ;
  assign n31050 = ( n31048 & ~n31049 ) | ( n31048 & 1'b0 ) | ( ~n31049 & 1'b0 ) ;
  assign n31059 = ( n160 & n30736 ) | ( n160 & n31050 ) | ( n30736 & n31050 ) ;
  assign n31060 = ( n30736 & ~n30772 ) | ( n30736 & n31050 ) | ( ~n30772 & n31050 ) ;
  assign n31061 = ~n31059 & n31060 ;
  assign n31062 = n31055 | n31061 ;
  assign n31063 = n30618 &  n30773 ;
  assign n31056 = x79 | n30618 ;
  assign n31057 = x79 &  n30618 ;
  assign n31058 = ( n31056 & ~n31057 ) | ( n31056 & 1'b0 ) | ( ~n31057 & 1'b0 ) ;
  assign n31067 = ( n160 & n30735 ) | ( n160 & n31058 ) | ( n30735 & n31058 ) ;
  assign n31068 = ( n30735 & ~n30772 ) | ( n30735 & n31058 ) | ( ~n30772 & n31058 ) ;
  assign n31069 = ~n31067 & n31068 ;
  assign n31070 = n31063 | n31069 ;
  assign n31071 = n30626 &  n30773 ;
  assign n31064 = x78 | n30626 ;
  assign n31065 = x78 &  n30626 ;
  assign n31066 = ( n31064 & ~n31065 ) | ( n31064 & 1'b0 ) | ( ~n31065 & 1'b0 ) ;
  assign n31075 = ( n160 & n30734 ) | ( n160 & n31066 ) | ( n30734 & n31066 ) ;
  assign n31076 = ( n30734 & ~n30772 ) | ( n30734 & n31066 ) | ( ~n30772 & n31066 ) ;
  assign n31077 = ~n31075 & n31076 ;
  assign n31078 = n31071 | n31077 ;
  assign n31079 = n30634 &  n30773 ;
  assign n31072 = x77 | n30634 ;
  assign n31073 = x77 &  n30634 ;
  assign n31074 = ( n31072 & ~n31073 ) | ( n31072 & 1'b0 ) | ( ~n31073 & 1'b0 ) ;
  assign n31083 = ( n160 & n30733 ) | ( n160 & n31074 ) | ( n30733 & n31074 ) ;
  assign n31084 = ( n30733 & ~n30772 ) | ( n30733 & n31074 ) | ( ~n30772 & n31074 ) ;
  assign n31085 = ~n31083 & n31084 ;
  assign n31086 = n31079 | n31085 ;
  assign n31087 = n30642 &  n30773 ;
  assign n31080 = x76 | n30642 ;
  assign n31081 = x76 &  n30642 ;
  assign n31082 = ( n31080 & ~n31081 ) | ( n31080 & 1'b0 ) | ( ~n31081 & 1'b0 ) ;
  assign n31091 = ( n160 & n30732 ) | ( n160 & n31082 ) | ( n30732 & n31082 ) ;
  assign n31092 = ( n30732 & ~n30772 ) | ( n30732 & n31082 ) | ( ~n30772 & n31082 ) ;
  assign n31093 = ~n31091 & n31092 ;
  assign n31094 = n31087 | n31093 ;
  assign n31095 = n30650 &  n30773 ;
  assign n31088 = x75 | n30650 ;
  assign n31089 = x75 &  n30650 ;
  assign n31090 = ( n31088 & ~n31089 ) | ( n31088 & 1'b0 ) | ( ~n31089 & 1'b0 ) ;
  assign n31099 = ( n160 & n30731 ) | ( n160 & n31090 ) | ( n30731 & n31090 ) ;
  assign n31100 = ( n30731 & ~n30772 ) | ( n30731 & n31090 ) | ( ~n30772 & n31090 ) ;
  assign n31101 = ~n31099 & n31100 ;
  assign n31102 = n31095 | n31101 ;
  assign n31103 = n30658 &  n30773 ;
  assign n31096 = x74 | n30658 ;
  assign n31097 = x74 &  n30658 ;
  assign n31098 = ( n31096 & ~n31097 ) | ( n31096 & 1'b0 ) | ( ~n31097 & 1'b0 ) ;
  assign n31107 = ( n160 & n30730 ) | ( n160 & n31098 ) | ( n30730 & n31098 ) ;
  assign n31108 = ( n30730 & ~n30772 ) | ( n30730 & n31098 ) | ( ~n30772 & n31098 ) ;
  assign n31109 = ~n31107 & n31108 ;
  assign n31110 = n31103 | n31109 ;
  assign n31111 = n30666 &  n30773 ;
  assign n31104 = x73 | n30666 ;
  assign n31105 = x73 &  n30666 ;
  assign n31106 = ( n31104 & ~n31105 ) | ( n31104 & 1'b0 ) | ( ~n31105 & 1'b0 ) ;
  assign n31115 = ( n160 & n30729 ) | ( n160 & n31106 ) | ( n30729 & n31106 ) ;
  assign n31116 = ( n30729 & ~n30772 ) | ( n30729 & n31106 ) | ( ~n30772 & n31106 ) ;
  assign n31117 = ~n31115 & n31116 ;
  assign n31118 = n31111 | n31117 ;
  assign n31119 = n30674 &  n30773 ;
  assign n31112 = x72 | n30674 ;
  assign n31113 = x72 &  n30674 ;
  assign n31114 = ( n31112 & ~n31113 ) | ( n31112 & 1'b0 ) | ( ~n31113 & 1'b0 ) ;
  assign n31123 = ( n160 & n30728 ) | ( n160 & n31114 ) | ( n30728 & n31114 ) ;
  assign n31124 = ( n30728 & ~n30772 ) | ( n30728 & n31114 ) | ( ~n30772 & n31114 ) ;
  assign n31125 = ~n31123 & n31124 ;
  assign n31126 = n31119 | n31125 ;
  assign n31127 = n30682 &  n30773 ;
  assign n31120 = x71 | n30682 ;
  assign n31121 = x71 &  n30682 ;
  assign n31122 = ( n31120 & ~n31121 ) | ( n31120 & 1'b0 ) | ( ~n31121 & 1'b0 ) ;
  assign n31131 = ( n160 & n30727 ) | ( n160 & n31122 ) | ( n30727 & n31122 ) ;
  assign n31132 = ( n30727 & ~n30772 ) | ( n30727 & n31122 ) | ( ~n30772 & n31122 ) ;
  assign n31133 = ~n31131 & n31132 ;
  assign n31134 = n31127 | n31133 ;
  assign n31135 = n30690 &  n30773 ;
  assign n31128 = x70 | n30690 ;
  assign n31129 = x70 &  n30690 ;
  assign n31130 = ( n31128 & ~n31129 ) | ( n31128 & 1'b0 ) | ( ~n31129 & 1'b0 ) ;
  assign n31139 = ( n160 & n30726 ) | ( n160 & n31130 ) | ( n30726 & n31130 ) ;
  assign n31140 = ( n30726 & ~n30772 ) | ( n30726 & n31130 ) | ( ~n30772 & n31130 ) ;
  assign n31141 = ~n31139 & n31140 ;
  assign n31142 = n31135 | n31141 ;
  assign n31143 = n30698 &  n30773 ;
  assign n31136 = x69 | n30698 ;
  assign n31137 = x69 &  n30698 ;
  assign n31138 = ( n31136 & ~n31137 ) | ( n31136 & 1'b0 ) | ( ~n31137 & 1'b0 ) ;
  assign n31147 = ( n160 & n30725 ) | ( n160 & n31138 ) | ( n30725 & n31138 ) ;
  assign n31148 = ( n30725 & ~n30772 ) | ( n30725 & n31138 ) | ( ~n30772 & n31138 ) ;
  assign n31149 = ~n31147 & n31148 ;
  assign n31150 = n31143 | n31149 ;
  assign n31151 = n30706 &  n30773 ;
  assign n31144 = x68 | n30706 ;
  assign n31145 = x68 &  n30706 ;
  assign n31146 = ( n31144 & ~n31145 ) | ( n31144 & 1'b0 ) | ( ~n31145 & 1'b0 ) ;
  assign n31155 = ( n160 & n30724 ) | ( n160 & n31146 ) | ( n30724 & n31146 ) ;
  assign n31156 = ( n30724 & ~n30772 ) | ( n30724 & n31146 ) | ( ~n30772 & n31146 ) ;
  assign n31157 = ~n31155 & n31156 ;
  assign n31158 = n31151 | n31157 ;
  assign n31159 = n30711 &  n30773 ;
  assign n31152 = x67 | n30711 ;
  assign n31153 = x67 &  n30711 ;
  assign n31154 = ( n31152 & ~n31153 ) | ( n31152 & 1'b0 ) | ( ~n31153 & 1'b0 ) ;
  assign n31163 = ( n160 & n30723 ) | ( n160 & n31154 ) | ( n30723 & n31154 ) ;
  assign n31164 = ( n30723 & ~n30772 ) | ( n30723 & n31154 ) | ( ~n30772 & n31154 ) ;
  assign n31165 = ~n31163 & n31164 ;
  assign n31166 = n31159 | n31165 ;
  assign n31167 = n30717 &  n30773 ;
  assign n31160 = x66 | n30717 ;
  assign n31161 = x66 &  n30717 ;
  assign n31162 = ( n31160 & ~n31161 ) | ( n31160 & 1'b0 ) | ( ~n31161 & 1'b0 ) ;
  assign n31168 = ( n160 & n30722 ) | ( n160 & n31162 ) | ( n30722 & n31162 ) ;
  assign n31169 = ( n30722 & ~n30772 ) | ( n30722 & n31162 ) | ( ~n30772 & n31162 ) ;
  assign n31170 = ~n31168 & n31169 ;
  assign n31171 = n31167 | n31170 ;
  assign n31172 = n30721 &  n30773 ;
  assign n31173 = ( x65 & ~x13 ) | ( x65 & n30718 ) | ( ~x13 & n30718 ) ;
  assign n31174 = ( x13 & ~n30718 ) | ( x13 & x65 ) | ( ~n30718 & x65 ) ;
  assign n31175 = ( n31173 & ~x65 ) | ( n31173 & n31174 ) | ( ~x65 & n31174 ) ;
  assign n31176 = ( n12413 & ~n30772 ) | ( n12413 & n31175 ) | ( ~n30772 & n31175 ) ;
  assign n31177 = ( n160 & n12413 ) | ( n160 & n31175 ) | ( n12413 & n31175 ) ;
  assign n31178 = ( n31176 & ~n31177 ) | ( n31176 & 1'b0 ) | ( ~n31177 & 1'b0 ) ;
  assign n31179 = n31172 | n31178 ;
  assign n31180 = ( n12804 & ~n30772 ) | ( n12804 & 1'b0 ) | ( ~n30772 & 1'b0 ) ;
  assign n31181 = ( x12 & ~n31180 ) | ( x12 & 1'b0 ) | ( ~n31180 & 1'b0 ) ;
  assign n31182 = ( n12808 & ~n30772 ) | ( n12808 & 1'b0 ) | ( ~n30772 & 1'b0 ) ;
  assign n31183 = n31181 | n31182 ;
  assign n31184 = ( x65 & ~n31183 ) | ( x65 & n12811 ) | ( ~n31183 & n12811 ) ;
  assign n31185 = ( x66 & ~n31179 ) | ( x66 & n31184 ) | ( ~n31179 & n31184 ) ;
  assign n31186 = ( x67 & ~n31171 ) | ( x67 & n31185 ) | ( ~n31171 & n31185 ) ;
  assign n31187 = ( x68 & ~n31166 ) | ( x68 & n31186 ) | ( ~n31166 & n31186 ) ;
  assign n31188 = ( x69 & ~n31158 ) | ( x69 & n31187 ) | ( ~n31158 & n31187 ) ;
  assign n31189 = ( x70 & ~n31150 ) | ( x70 & n31188 ) | ( ~n31150 & n31188 ) ;
  assign n31190 = ( x71 & ~n31142 ) | ( x71 & n31189 ) | ( ~n31142 & n31189 ) ;
  assign n31191 = ( x72 & ~n31134 ) | ( x72 & n31190 ) | ( ~n31134 & n31190 ) ;
  assign n31192 = ( x73 & ~n31126 ) | ( x73 & n31191 ) | ( ~n31126 & n31191 ) ;
  assign n31193 = ( x74 & ~n31118 ) | ( x74 & n31192 ) | ( ~n31118 & n31192 ) ;
  assign n31194 = ( x75 & ~n31110 ) | ( x75 & n31193 ) | ( ~n31110 & n31193 ) ;
  assign n31195 = ( x76 & ~n31102 ) | ( x76 & n31194 ) | ( ~n31102 & n31194 ) ;
  assign n31196 = ( x77 & ~n31094 ) | ( x77 & n31195 ) | ( ~n31094 & n31195 ) ;
  assign n31197 = ( x78 & ~n31086 ) | ( x78 & n31196 ) | ( ~n31086 & n31196 ) ;
  assign n31198 = ( x79 & ~n31078 ) | ( x79 & n31197 ) | ( ~n31078 & n31197 ) ;
  assign n31199 = ( x80 & ~n31070 ) | ( x80 & n31198 ) | ( ~n31070 & n31198 ) ;
  assign n31200 = ( x81 & ~n31062 ) | ( x81 & n31199 ) | ( ~n31062 & n31199 ) ;
  assign n31201 = ( x82 & ~n31054 ) | ( x82 & n31200 ) | ( ~n31054 & n31200 ) ;
  assign n31202 = ( x83 & ~n31046 ) | ( x83 & n31201 ) | ( ~n31046 & n31201 ) ;
  assign n31203 = ( x84 & ~n31038 ) | ( x84 & n31202 ) | ( ~n31038 & n31202 ) ;
  assign n31204 = ( x85 & ~n31030 ) | ( x85 & n31203 ) | ( ~n31030 & n31203 ) ;
  assign n31205 = ( x86 & ~n31022 ) | ( x86 & n31204 ) | ( ~n31022 & n31204 ) ;
  assign n31206 = ( x87 & ~n31014 ) | ( x87 & n31205 ) | ( ~n31014 & n31205 ) ;
  assign n31207 = ( x88 & ~n31006 ) | ( x88 & n31206 ) | ( ~n31006 & n31206 ) ;
  assign n31208 = ( x89 & ~n30998 ) | ( x89 & n31207 ) | ( ~n30998 & n31207 ) ;
  assign n31209 = ( x90 & ~n30990 ) | ( x90 & n31208 ) | ( ~n30990 & n31208 ) ;
  assign n31210 = ( x91 & ~n30982 ) | ( x91 & n31209 ) | ( ~n30982 & n31209 ) ;
  assign n31211 = ( x92 & ~n30974 ) | ( x92 & n31210 ) | ( ~n30974 & n31210 ) ;
  assign n31212 = ( x93 & ~n30966 ) | ( x93 & n31211 ) | ( ~n30966 & n31211 ) ;
  assign n31213 = ( x94 & ~n30958 ) | ( x94 & n31212 ) | ( ~n30958 & n31212 ) ;
  assign n31214 = ( x95 & ~n30950 ) | ( x95 & n31213 ) | ( ~n30950 & n31213 ) ;
  assign n31215 = ( x96 & ~n30942 ) | ( x96 & n31214 ) | ( ~n30942 & n31214 ) ;
  assign n31216 = ( x97 & ~n30934 ) | ( x97 & n31215 ) | ( ~n30934 & n31215 ) ;
  assign n31217 = ( x98 & ~n30926 ) | ( x98 & n31216 ) | ( ~n30926 & n31216 ) ;
  assign n31218 = ( x99 & ~n30918 ) | ( x99 & n31217 ) | ( ~n30918 & n31217 ) ;
  assign n31219 = ( x100 & ~n30910 ) | ( x100 & n31218 ) | ( ~n30910 & n31218 ) ;
  assign n31220 = ( x101 & ~n30902 ) | ( x101 & n31219 ) | ( ~n30902 & n31219 ) ;
  assign n31221 = ( x102 & ~n30894 ) | ( x102 & n31220 ) | ( ~n30894 & n31220 ) ;
  assign n31222 = ( x103 & ~n30886 ) | ( x103 & n31221 ) | ( ~n30886 & n31221 ) ;
  assign n31223 = ( x104 & ~n30878 ) | ( x104 & n31222 ) | ( ~n30878 & n31222 ) ;
  assign n31224 = ( x105 & ~n30870 ) | ( x105 & n31223 ) | ( ~n30870 & n31223 ) ;
  assign n31225 = ( x106 & ~n30862 ) | ( x106 & n31224 ) | ( ~n30862 & n31224 ) ;
  assign n31226 = ( x107 & ~n30854 ) | ( x107 & n31225 ) | ( ~n30854 & n31225 ) ;
  assign n31227 = ( x108 & ~n30846 ) | ( x108 & n31226 ) | ( ~n30846 & n31226 ) ;
  assign n31228 = ( x109 & ~n30838 ) | ( x109 & n31227 ) | ( ~n30838 & n31227 ) ;
  assign n31229 = ( x110 & ~n30830 ) | ( x110 & n31228 ) | ( ~n30830 & n31228 ) ;
  assign n31230 = ( x111 & ~n30822 ) | ( x111 & n31229 ) | ( ~n30822 & n31229 ) ;
  assign n31231 = ( x112 & ~n30814 ) | ( x112 & n31230 ) | ( ~n30814 & n31230 ) ;
  assign n31232 = ( x113 & ~n30806 ) | ( x113 & n31231 ) | ( ~n30806 & n31231 ) ;
  assign n31233 = ( x114 & ~n30798 ) | ( x114 & n31232 ) | ( ~n30798 & n31232 ) ;
  assign n31234 = ( x115 & ~n30790 ) | ( x115 & n31233 ) | ( ~n30790 & n31233 ) ;
  assign n30774 = n30330 &  n30773 ;
  assign n30778 = ( n160 & n30330 ) | ( n160 & n30771 ) | ( n30330 & n30771 ) ;
  assign n30779 = ( x115 & ~n30778 ) | ( x115 & n30330 ) | ( ~n30778 & n30330 ) ;
  assign n30780 = ~x115 & n30779 ;
  assign n30781 = n30774 | n30780 ;
  assign n30782 = ~x116 & n30781 ;
  assign n31235 = ( x116 & ~n30774 ) | ( x116 & 1'b0 ) | ( ~n30774 & 1'b0 ) ;
  assign n31236 = ~n30780 & n31235 ;
  assign n31245 = n30782 | n31236 ;
  assign n31246 = ( n31234 & ~n31245 ) | ( n31234 & 1'b0 ) | ( ~n31245 & 1'b0 ) ;
  assign n31237 = ( n31234 & ~n30782 ) | ( n31234 & n31236 ) | ( ~n30782 & n31236 ) ;
  assign n31238 = ( n30782 & ~n425 ) | ( n30782 & n31237 ) | ( ~n425 & n31237 ) ;
  assign n31239 = n425 | n31238 ;
  assign n31240 = ~n30781 |  n160 ;
  assign n31241 = n31239 &  n31240 ;
  assign n31247 = ~n31234 & n31245 ;
  assign n31248 = ( n31246 & ~n31241 ) | ( n31246 & n31247 ) | ( ~n31241 & n31247 ) ;
  assign n31249 = n160 &  n30330 ;
  assign n31250 = n31239 &  n31249 ;
  assign n31251 = n31248 | n31250 ;
  assign n31252 = ~x117 & n31251 ;
  assign n31256 = n30790 &  n31240 ;
  assign n31257 = n31239 &  n31256 ;
  assign n31242 = x115 | n30790 ;
  assign n31243 = x115 &  n30790 ;
  assign n31244 = ( n31242 & ~n31243 ) | ( n31242 & 1'b0 ) | ( ~n31243 & 1'b0 ) ;
  assign n31259 = ( n31233 & n31241 ) | ( n31233 & n31244 ) | ( n31241 & n31244 ) ;
  assign n31258 = n31233 | n31244 ;
  assign n31260 = ( n31257 & ~n31259 ) | ( n31257 & n31258 ) | ( ~n31259 & n31258 ) ;
  assign n31264 = n30798 &  n31240 ;
  assign n31265 = n31239 &  n31264 ;
  assign n31253 = x114 | n30798 ;
  assign n31254 = x114 &  n30798 ;
  assign n31255 = ( n31253 & ~n31254 ) | ( n31253 & 1'b0 ) | ( ~n31254 & 1'b0 ) ;
  assign n31267 = ( n31232 & n31241 ) | ( n31232 & n31255 ) | ( n31241 & n31255 ) ;
  assign n31266 = n31232 | n31255 ;
  assign n31268 = ( n31265 & ~n31267 ) | ( n31265 & n31266 ) | ( ~n31267 & n31266 ) ;
  assign n31272 = n30806 &  n31240 ;
  assign n31273 = n31239 &  n31272 ;
  assign n31261 = x113 | n30806 ;
  assign n31262 = x113 &  n30806 ;
  assign n31263 = ( n31261 & ~n31262 ) | ( n31261 & 1'b0 ) | ( ~n31262 & 1'b0 ) ;
  assign n31275 = ( n31231 & n31241 ) | ( n31231 & n31263 ) | ( n31241 & n31263 ) ;
  assign n31274 = n31231 | n31263 ;
  assign n31276 = ( n31273 & ~n31275 ) | ( n31273 & n31274 ) | ( ~n31275 & n31274 ) ;
  assign n31280 = n30814 &  n31240 ;
  assign n31281 = n31239 &  n31280 ;
  assign n31269 = x112 | n30814 ;
  assign n31270 = x112 &  n30814 ;
  assign n31271 = ( n31269 & ~n31270 ) | ( n31269 & 1'b0 ) | ( ~n31270 & 1'b0 ) ;
  assign n31283 = ( n31230 & n31241 ) | ( n31230 & n31271 ) | ( n31241 & n31271 ) ;
  assign n31282 = n31230 | n31271 ;
  assign n31284 = ( n31281 & ~n31283 ) | ( n31281 & n31282 ) | ( ~n31283 & n31282 ) ;
  assign n31288 = n30822 &  n31240 ;
  assign n31289 = n31239 &  n31288 ;
  assign n31277 = x111 | n30822 ;
  assign n31278 = x111 &  n30822 ;
  assign n31279 = ( n31277 & ~n31278 ) | ( n31277 & 1'b0 ) | ( ~n31278 & 1'b0 ) ;
  assign n31291 = ( n31229 & n31241 ) | ( n31229 & n31279 ) | ( n31241 & n31279 ) ;
  assign n31290 = n31229 | n31279 ;
  assign n31292 = ( n31289 & ~n31291 ) | ( n31289 & n31290 ) | ( ~n31291 & n31290 ) ;
  assign n31296 = n30830 &  n31240 ;
  assign n31297 = n31239 &  n31296 ;
  assign n31285 = x110 | n30830 ;
  assign n31286 = x110 &  n30830 ;
  assign n31287 = ( n31285 & ~n31286 ) | ( n31285 & 1'b0 ) | ( ~n31286 & 1'b0 ) ;
  assign n31299 = ( n31228 & n31241 ) | ( n31228 & n31287 ) | ( n31241 & n31287 ) ;
  assign n31298 = n31228 | n31287 ;
  assign n31300 = ( n31297 & ~n31299 ) | ( n31297 & n31298 ) | ( ~n31299 & n31298 ) ;
  assign n31304 = n30838 &  n31240 ;
  assign n31305 = n31239 &  n31304 ;
  assign n31293 = x109 | n30838 ;
  assign n31294 = x109 &  n30838 ;
  assign n31295 = ( n31293 & ~n31294 ) | ( n31293 & 1'b0 ) | ( ~n31294 & 1'b0 ) ;
  assign n31307 = ( n31227 & n31241 ) | ( n31227 & n31295 ) | ( n31241 & n31295 ) ;
  assign n31306 = n31227 | n31295 ;
  assign n31308 = ( n31305 & ~n31307 ) | ( n31305 & n31306 ) | ( ~n31307 & n31306 ) ;
  assign n31312 = n30846 &  n31240 ;
  assign n31313 = n31239 &  n31312 ;
  assign n31301 = x108 | n30846 ;
  assign n31302 = x108 &  n30846 ;
  assign n31303 = ( n31301 & ~n31302 ) | ( n31301 & 1'b0 ) | ( ~n31302 & 1'b0 ) ;
  assign n31315 = ( n31226 & n31241 ) | ( n31226 & n31303 ) | ( n31241 & n31303 ) ;
  assign n31314 = n31226 | n31303 ;
  assign n31316 = ( n31313 & ~n31315 ) | ( n31313 & n31314 ) | ( ~n31315 & n31314 ) ;
  assign n31320 = n30854 &  n31240 ;
  assign n31321 = n31239 &  n31320 ;
  assign n31309 = x107 | n30854 ;
  assign n31310 = x107 &  n30854 ;
  assign n31311 = ( n31309 & ~n31310 ) | ( n31309 & 1'b0 ) | ( ~n31310 & 1'b0 ) ;
  assign n31323 = ( n31225 & n31241 ) | ( n31225 & n31311 ) | ( n31241 & n31311 ) ;
  assign n31322 = n31225 | n31311 ;
  assign n31324 = ( n31321 & ~n31323 ) | ( n31321 & n31322 ) | ( ~n31323 & n31322 ) ;
  assign n31328 = n30862 &  n31240 ;
  assign n31329 = n31239 &  n31328 ;
  assign n31317 = x106 | n30862 ;
  assign n31318 = x106 &  n30862 ;
  assign n31319 = ( n31317 & ~n31318 ) | ( n31317 & 1'b0 ) | ( ~n31318 & 1'b0 ) ;
  assign n31331 = ( n31224 & n31241 ) | ( n31224 & n31319 ) | ( n31241 & n31319 ) ;
  assign n31330 = n31224 | n31319 ;
  assign n31332 = ( n31329 & ~n31331 ) | ( n31329 & n31330 ) | ( ~n31331 & n31330 ) ;
  assign n31336 = n30870 &  n31240 ;
  assign n31337 = n31239 &  n31336 ;
  assign n31325 = x105 | n30870 ;
  assign n31326 = x105 &  n30870 ;
  assign n31327 = ( n31325 & ~n31326 ) | ( n31325 & 1'b0 ) | ( ~n31326 & 1'b0 ) ;
  assign n31339 = ( n31223 & n31241 ) | ( n31223 & n31327 ) | ( n31241 & n31327 ) ;
  assign n31338 = n31223 | n31327 ;
  assign n31340 = ( n31337 & ~n31339 ) | ( n31337 & n31338 ) | ( ~n31339 & n31338 ) ;
  assign n31344 = n30878 &  n31240 ;
  assign n31345 = n31239 &  n31344 ;
  assign n31333 = x104 | n30878 ;
  assign n31334 = x104 &  n30878 ;
  assign n31335 = ( n31333 & ~n31334 ) | ( n31333 & 1'b0 ) | ( ~n31334 & 1'b0 ) ;
  assign n31347 = ( n31222 & n31241 ) | ( n31222 & n31335 ) | ( n31241 & n31335 ) ;
  assign n31346 = n31222 | n31335 ;
  assign n31348 = ( n31345 & ~n31347 ) | ( n31345 & n31346 ) | ( ~n31347 & n31346 ) ;
  assign n31352 = n30886 &  n31240 ;
  assign n31353 = n31239 &  n31352 ;
  assign n31341 = x103 | n30886 ;
  assign n31342 = x103 &  n30886 ;
  assign n31343 = ( n31341 & ~n31342 ) | ( n31341 & 1'b0 ) | ( ~n31342 & 1'b0 ) ;
  assign n31355 = ( n31221 & n31241 ) | ( n31221 & n31343 ) | ( n31241 & n31343 ) ;
  assign n31354 = n31221 | n31343 ;
  assign n31356 = ( n31353 & ~n31355 ) | ( n31353 & n31354 ) | ( ~n31355 & n31354 ) ;
  assign n31360 = n30894 &  n31240 ;
  assign n31361 = n31239 &  n31360 ;
  assign n31349 = x102 | n30894 ;
  assign n31350 = x102 &  n30894 ;
  assign n31351 = ( n31349 & ~n31350 ) | ( n31349 & 1'b0 ) | ( ~n31350 & 1'b0 ) ;
  assign n31363 = ( n31220 & n31241 ) | ( n31220 & n31351 ) | ( n31241 & n31351 ) ;
  assign n31362 = n31220 | n31351 ;
  assign n31364 = ( n31361 & ~n31363 ) | ( n31361 & n31362 ) | ( ~n31363 & n31362 ) ;
  assign n31368 = n30902 &  n31240 ;
  assign n31369 = n31239 &  n31368 ;
  assign n31357 = x101 | n30902 ;
  assign n31358 = x101 &  n30902 ;
  assign n31359 = ( n31357 & ~n31358 ) | ( n31357 & 1'b0 ) | ( ~n31358 & 1'b0 ) ;
  assign n31371 = ( n31219 & n31241 ) | ( n31219 & n31359 ) | ( n31241 & n31359 ) ;
  assign n31370 = n31219 | n31359 ;
  assign n31372 = ( n31369 & ~n31371 ) | ( n31369 & n31370 ) | ( ~n31371 & n31370 ) ;
  assign n31376 = n30910 &  n31240 ;
  assign n31377 = n31239 &  n31376 ;
  assign n31365 = x100 | n30910 ;
  assign n31366 = x100 &  n30910 ;
  assign n31367 = ( n31365 & ~n31366 ) | ( n31365 & 1'b0 ) | ( ~n31366 & 1'b0 ) ;
  assign n31379 = ( n31218 & n31241 ) | ( n31218 & n31367 ) | ( n31241 & n31367 ) ;
  assign n31378 = n31218 | n31367 ;
  assign n31380 = ( n31377 & ~n31379 ) | ( n31377 & n31378 ) | ( ~n31379 & n31378 ) ;
  assign n31384 = n30918 &  n31240 ;
  assign n31385 = n31239 &  n31384 ;
  assign n31373 = x99 | n30918 ;
  assign n31374 = x99 &  n30918 ;
  assign n31375 = ( n31373 & ~n31374 ) | ( n31373 & 1'b0 ) | ( ~n31374 & 1'b0 ) ;
  assign n31387 = ( n31217 & n31241 ) | ( n31217 & n31375 ) | ( n31241 & n31375 ) ;
  assign n31386 = n31217 | n31375 ;
  assign n31388 = ( n31385 & ~n31387 ) | ( n31385 & n31386 ) | ( ~n31387 & n31386 ) ;
  assign n31392 = n30926 &  n31240 ;
  assign n31393 = n31239 &  n31392 ;
  assign n31381 = x98 | n30926 ;
  assign n31382 = x98 &  n30926 ;
  assign n31383 = ( n31381 & ~n31382 ) | ( n31381 & 1'b0 ) | ( ~n31382 & 1'b0 ) ;
  assign n31395 = ( n31216 & n31241 ) | ( n31216 & n31383 ) | ( n31241 & n31383 ) ;
  assign n31394 = n31216 | n31383 ;
  assign n31396 = ( n31393 & ~n31395 ) | ( n31393 & n31394 ) | ( ~n31395 & n31394 ) ;
  assign n31400 = n30934 &  n31240 ;
  assign n31401 = n31239 &  n31400 ;
  assign n31389 = x97 | n30934 ;
  assign n31390 = x97 &  n30934 ;
  assign n31391 = ( n31389 & ~n31390 ) | ( n31389 & 1'b0 ) | ( ~n31390 & 1'b0 ) ;
  assign n31403 = ( n31215 & n31241 ) | ( n31215 & n31391 ) | ( n31241 & n31391 ) ;
  assign n31402 = n31215 | n31391 ;
  assign n31404 = ( n31401 & ~n31403 ) | ( n31401 & n31402 ) | ( ~n31403 & n31402 ) ;
  assign n31408 = n30942 &  n31240 ;
  assign n31409 = n31239 &  n31408 ;
  assign n31397 = x96 | n30942 ;
  assign n31398 = x96 &  n30942 ;
  assign n31399 = ( n31397 & ~n31398 ) | ( n31397 & 1'b0 ) | ( ~n31398 & 1'b0 ) ;
  assign n31411 = ( n31214 & n31241 ) | ( n31214 & n31399 ) | ( n31241 & n31399 ) ;
  assign n31410 = n31214 | n31399 ;
  assign n31412 = ( n31409 & ~n31411 ) | ( n31409 & n31410 ) | ( ~n31411 & n31410 ) ;
  assign n31416 = n30950 &  n31240 ;
  assign n31417 = n31239 &  n31416 ;
  assign n31405 = x95 | n30950 ;
  assign n31406 = x95 &  n30950 ;
  assign n31407 = ( n31405 & ~n31406 ) | ( n31405 & 1'b0 ) | ( ~n31406 & 1'b0 ) ;
  assign n31419 = ( n31213 & n31241 ) | ( n31213 & n31407 ) | ( n31241 & n31407 ) ;
  assign n31418 = n31213 | n31407 ;
  assign n31420 = ( n31417 & ~n31419 ) | ( n31417 & n31418 ) | ( ~n31419 & n31418 ) ;
  assign n31424 = n30958 &  n31240 ;
  assign n31425 = n31239 &  n31424 ;
  assign n31413 = x94 | n30958 ;
  assign n31414 = x94 &  n30958 ;
  assign n31415 = ( n31413 & ~n31414 ) | ( n31413 & 1'b0 ) | ( ~n31414 & 1'b0 ) ;
  assign n31427 = ( n31212 & n31241 ) | ( n31212 & n31415 ) | ( n31241 & n31415 ) ;
  assign n31426 = n31212 | n31415 ;
  assign n31428 = ( n31425 & ~n31427 ) | ( n31425 & n31426 ) | ( ~n31427 & n31426 ) ;
  assign n31432 = n30966 &  n31240 ;
  assign n31433 = n31239 &  n31432 ;
  assign n31421 = x93 | n30966 ;
  assign n31422 = x93 &  n30966 ;
  assign n31423 = ( n31421 & ~n31422 ) | ( n31421 & 1'b0 ) | ( ~n31422 & 1'b0 ) ;
  assign n31435 = ( n31211 & n31241 ) | ( n31211 & n31423 ) | ( n31241 & n31423 ) ;
  assign n31434 = n31211 | n31423 ;
  assign n31436 = ( n31433 & ~n31435 ) | ( n31433 & n31434 ) | ( ~n31435 & n31434 ) ;
  assign n31440 = n30974 &  n31240 ;
  assign n31441 = n31239 &  n31440 ;
  assign n31429 = x92 | n30974 ;
  assign n31430 = x92 &  n30974 ;
  assign n31431 = ( n31429 & ~n31430 ) | ( n31429 & 1'b0 ) | ( ~n31430 & 1'b0 ) ;
  assign n31443 = ( n31210 & n31241 ) | ( n31210 & n31431 ) | ( n31241 & n31431 ) ;
  assign n31442 = n31210 | n31431 ;
  assign n31444 = ( n31441 & ~n31443 ) | ( n31441 & n31442 ) | ( ~n31443 & n31442 ) ;
  assign n31448 = n30982 &  n31240 ;
  assign n31449 = n31239 &  n31448 ;
  assign n31437 = x91 | n30982 ;
  assign n31438 = x91 &  n30982 ;
  assign n31439 = ( n31437 & ~n31438 ) | ( n31437 & 1'b0 ) | ( ~n31438 & 1'b0 ) ;
  assign n31451 = ( n31209 & n31241 ) | ( n31209 & n31439 ) | ( n31241 & n31439 ) ;
  assign n31450 = n31209 | n31439 ;
  assign n31452 = ( n31449 & ~n31451 ) | ( n31449 & n31450 ) | ( ~n31451 & n31450 ) ;
  assign n31456 = n30990 &  n31240 ;
  assign n31457 = n31239 &  n31456 ;
  assign n31445 = x90 | n30990 ;
  assign n31446 = x90 &  n30990 ;
  assign n31447 = ( n31445 & ~n31446 ) | ( n31445 & 1'b0 ) | ( ~n31446 & 1'b0 ) ;
  assign n31459 = ( n31208 & n31241 ) | ( n31208 & n31447 ) | ( n31241 & n31447 ) ;
  assign n31458 = n31208 | n31447 ;
  assign n31460 = ( n31457 & ~n31459 ) | ( n31457 & n31458 ) | ( ~n31459 & n31458 ) ;
  assign n31464 = n30998 &  n31240 ;
  assign n31465 = n31239 &  n31464 ;
  assign n31453 = x89 | n30998 ;
  assign n31454 = x89 &  n30998 ;
  assign n31455 = ( n31453 & ~n31454 ) | ( n31453 & 1'b0 ) | ( ~n31454 & 1'b0 ) ;
  assign n31467 = ( n31207 & n31241 ) | ( n31207 & n31455 ) | ( n31241 & n31455 ) ;
  assign n31466 = n31207 | n31455 ;
  assign n31468 = ( n31465 & ~n31467 ) | ( n31465 & n31466 ) | ( ~n31467 & n31466 ) ;
  assign n31472 = n31006 &  n31240 ;
  assign n31473 = n31239 &  n31472 ;
  assign n31461 = x88 | n31006 ;
  assign n31462 = x88 &  n31006 ;
  assign n31463 = ( n31461 & ~n31462 ) | ( n31461 & 1'b0 ) | ( ~n31462 & 1'b0 ) ;
  assign n31475 = ( n31206 & n31241 ) | ( n31206 & n31463 ) | ( n31241 & n31463 ) ;
  assign n31474 = n31206 | n31463 ;
  assign n31476 = ( n31473 & ~n31475 ) | ( n31473 & n31474 ) | ( ~n31475 & n31474 ) ;
  assign n31480 = n31014 &  n31240 ;
  assign n31481 = n31239 &  n31480 ;
  assign n31469 = x87 | n31014 ;
  assign n31470 = x87 &  n31014 ;
  assign n31471 = ( n31469 & ~n31470 ) | ( n31469 & 1'b0 ) | ( ~n31470 & 1'b0 ) ;
  assign n31483 = ( n31205 & n31241 ) | ( n31205 & n31471 ) | ( n31241 & n31471 ) ;
  assign n31482 = n31205 | n31471 ;
  assign n31484 = ( n31481 & ~n31483 ) | ( n31481 & n31482 ) | ( ~n31483 & n31482 ) ;
  assign n31488 = n31022 &  n31240 ;
  assign n31489 = n31239 &  n31488 ;
  assign n31477 = x86 | n31022 ;
  assign n31478 = x86 &  n31022 ;
  assign n31479 = ( n31477 & ~n31478 ) | ( n31477 & 1'b0 ) | ( ~n31478 & 1'b0 ) ;
  assign n31491 = ( n31204 & n31241 ) | ( n31204 & n31479 ) | ( n31241 & n31479 ) ;
  assign n31490 = n31204 | n31479 ;
  assign n31492 = ( n31489 & ~n31491 ) | ( n31489 & n31490 ) | ( ~n31491 & n31490 ) ;
  assign n31496 = n31030 &  n31240 ;
  assign n31497 = n31239 &  n31496 ;
  assign n31485 = x85 | n31030 ;
  assign n31486 = x85 &  n31030 ;
  assign n31487 = ( n31485 & ~n31486 ) | ( n31485 & 1'b0 ) | ( ~n31486 & 1'b0 ) ;
  assign n31499 = ( n31203 & n31241 ) | ( n31203 & n31487 ) | ( n31241 & n31487 ) ;
  assign n31498 = n31203 | n31487 ;
  assign n31500 = ( n31497 & ~n31499 ) | ( n31497 & n31498 ) | ( ~n31499 & n31498 ) ;
  assign n31504 = n31038 &  n31240 ;
  assign n31505 = n31239 &  n31504 ;
  assign n31493 = x84 | n31038 ;
  assign n31494 = x84 &  n31038 ;
  assign n31495 = ( n31493 & ~n31494 ) | ( n31493 & 1'b0 ) | ( ~n31494 & 1'b0 ) ;
  assign n31507 = ( n31202 & n31241 ) | ( n31202 & n31495 ) | ( n31241 & n31495 ) ;
  assign n31506 = n31202 | n31495 ;
  assign n31508 = ( n31505 & ~n31507 ) | ( n31505 & n31506 ) | ( ~n31507 & n31506 ) ;
  assign n31512 = n31046 &  n31240 ;
  assign n31513 = n31239 &  n31512 ;
  assign n31501 = x83 | n31046 ;
  assign n31502 = x83 &  n31046 ;
  assign n31503 = ( n31501 & ~n31502 ) | ( n31501 & 1'b0 ) | ( ~n31502 & 1'b0 ) ;
  assign n31515 = ( n31201 & n31241 ) | ( n31201 & n31503 ) | ( n31241 & n31503 ) ;
  assign n31514 = n31201 | n31503 ;
  assign n31516 = ( n31513 & ~n31515 ) | ( n31513 & n31514 ) | ( ~n31515 & n31514 ) ;
  assign n31520 = n31054 &  n31240 ;
  assign n31521 = n31239 &  n31520 ;
  assign n31509 = x82 | n31054 ;
  assign n31510 = x82 &  n31054 ;
  assign n31511 = ( n31509 & ~n31510 ) | ( n31509 & 1'b0 ) | ( ~n31510 & 1'b0 ) ;
  assign n31523 = ( n31200 & n31241 ) | ( n31200 & n31511 ) | ( n31241 & n31511 ) ;
  assign n31522 = n31200 | n31511 ;
  assign n31524 = ( n31521 & ~n31523 ) | ( n31521 & n31522 ) | ( ~n31523 & n31522 ) ;
  assign n31528 = n31062 &  n31240 ;
  assign n31529 = n31239 &  n31528 ;
  assign n31517 = x81 | n31062 ;
  assign n31518 = x81 &  n31062 ;
  assign n31519 = ( n31517 & ~n31518 ) | ( n31517 & 1'b0 ) | ( ~n31518 & 1'b0 ) ;
  assign n31531 = ( n31199 & n31241 ) | ( n31199 & n31519 ) | ( n31241 & n31519 ) ;
  assign n31530 = n31199 | n31519 ;
  assign n31532 = ( n31529 & ~n31531 ) | ( n31529 & n31530 ) | ( ~n31531 & n31530 ) ;
  assign n31536 = n31070 &  n31240 ;
  assign n31537 = n31239 &  n31536 ;
  assign n31525 = x80 | n31070 ;
  assign n31526 = x80 &  n31070 ;
  assign n31527 = ( n31525 & ~n31526 ) | ( n31525 & 1'b0 ) | ( ~n31526 & 1'b0 ) ;
  assign n31539 = ( n31198 & n31241 ) | ( n31198 & n31527 ) | ( n31241 & n31527 ) ;
  assign n31538 = n31198 | n31527 ;
  assign n31540 = ( n31537 & ~n31539 ) | ( n31537 & n31538 ) | ( ~n31539 & n31538 ) ;
  assign n31544 = n31078 &  n31240 ;
  assign n31545 = n31239 &  n31544 ;
  assign n31533 = x79 | n31078 ;
  assign n31534 = x79 &  n31078 ;
  assign n31535 = ( n31533 & ~n31534 ) | ( n31533 & 1'b0 ) | ( ~n31534 & 1'b0 ) ;
  assign n31547 = ( n31197 & n31241 ) | ( n31197 & n31535 ) | ( n31241 & n31535 ) ;
  assign n31546 = n31197 | n31535 ;
  assign n31548 = ( n31545 & ~n31547 ) | ( n31545 & n31546 ) | ( ~n31547 & n31546 ) ;
  assign n31552 = n31086 &  n31240 ;
  assign n31553 = n31239 &  n31552 ;
  assign n31541 = x78 | n31086 ;
  assign n31542 = x78 &  n31086 ;
  assign n31543 = ( n31541 & ~n31542 ) | ( n31541 & 1'b0 ) | ( ~n31542 & 1'b0 ) ;
  assign n31555 = ( n31196 & n31241 ) | ( n31196 & n31543 ) | ( n31241 & n31543 ) ;
  assign n31554 = n31196 | n31543 ;
  assign n31556 = ( n31553 & ~n31555 ) | ( n31553 & n31554 ) | ( ~n31555 & n31554 ) ;
  assign n31560 = n31094 &  n31240 ;
  assign n31561 = n31239 &  n31560 ;
  assign n31549 = x77 | n31094 ;
  assign n31550 = x77 &  n31094 ;
  assign n31551 = ( n31549 & ~n31550 ) | ( n31549 & 1'b0 ) | ( ~n31550 & 1'b0 ) ;
  assign n31563 = ( n31195 & n31241 ) | ( n31195 & n31551 ) | ( n31241 & n31551 ) ;
  assign n31562 = n31195 | n31551 ;
  assign n31564 = ( n31561 & ~n31563 ) | ( n31561 & n31562 ) | ( ~n31563 & n31562 ) ;
  assign n31568 = n31102 &  n31240 ;
  assign n31569 = n31239 &  n31568 ;
  assign n31557 = x76 | n31102 ;
  assign n31558 = x76 &  n31102 ;
  assign n31559 = ( n31557 & ~n31558 ) | ( n31557 & 1'b0 ) | ( ~n31558 & 1'b0 ) ;
  assign n31571 = ( n31194 & n31241 ) | ( n31194 & n31559 ) | ( n31241 & n31559 ) ;
  assign n31570 = n31194 | n31559 ;
  assign n31572 = ( n31569 & ~n31571 ) | ( n31569 & n31570 ) | ( ~n31571 & n31570 ) ;
  assign n31576 = n31110 &  n31240 ;
  assign n31577 = n31239 &  n31576 ;
  assign n31565 = x75 | n31110 ;
  assign n31566 = x75 &  n31110 ;
  assign n31567 = ( n31565 & ~n31566 ) | ( n31565 & 1'b0 ) | ( ~n31566 & 1'b0 ) ;
  assign n31579 = ( n31193 & n31241 ) | ( n31193 & n31567 ) | ( n31241 & n31567 ) ;
  assign n31578 = n31193 | n31567 ;
  assign n31580 = ( n31577 & ~n31579 ) | ( n31577 & n31578 ) | ( ~n31579 & n31578 ) ;
  assign n31584 = n31118 &  n31240 ;
  assign n31585 = n31239 &  n31584 ;
  assign n31573 = x74 | n31118 ;
  assign n31574 = x74 &  n31118 ;
  assign n31575 = ( n31573 & ~n31574 ) | ( n31573 & 1'b0 ) | ( ~n31574 & 1'b0 ) ;
  assign n31587 = ( n31192 & n31241 ) | ( n31192 & n31575 ) | ( n31241 & n31575 ) ;
  assign n31586 = n31192 | n31575 ;
  assign n31588 = ( n31585 & ~n31587 ) | ( n31585 & n31586 ) | ( ~n31587 & n31586 ) ;
  assign n31592 = n31126 &  n31240 ;
  assign n31593 = n31239 &  n31592 ;
  assign n31581 = x73 | n31126 ;
  assign n31582 = x73 &  n31126 ;
  assign n31583 = ( n31581 & ~n31582 ) | ( n31581 & 1'b0 ) | ( ~n31582 & 1'b0 ) ;
  assign n31595 = ( n31191 & n31241 ) | ( n31191 & n31583 ) | ( n31241 & n31583 ) ;
  assign n31594 = n31191 | n31583 ;
  assign n31596 = ( n31593 & ~n31595 ) | ( n31593 & n31594 ) | ( ~n31595 & n31594 ) ;
  assign n31600 = n31134 &  n31240 ;
  assign n31601 = n31239 &  n31600 ;
  assign n31589 = x72 | n31134 ;
  assign n31590 = x72 &  n31134 ;
  assign n31591 = ( n31589 & ~n31590 ) | ( n31589 & 1'b0 ) | ( ~n31590 & 1'b0 ) ;
  assign n31603 = ( n31190 & n31241 ) | ( n31190 & n31591 ) | ( n31241 & n31591 ) ;
  assign n31602 = n31190 | n31591 ;
  assign n31604 = ( n31601 & ~n31603 ) | ( n31601 & n31602 ) | ( ~n31603 & n31602 ) ;
  assign n31608 = n31142 &  n31240 ;
  assign n31609 = n31239 &  n31608 ;
  assign n31597 = x71 | n31142 ;
  assign n31598 = x71 &  n31142 ;
  assign n31599 = ( n31597 & ~n31598 ) | ( n31597 & 1'b0 ) | ( ~n31598 & 1'b0 ) ;
  assign n31611 = ( n31189 & n31241 ) | ( n31189 & n31599 ) | ( n31241 & n31599 ) ;
  assign n31610 = n31189 | n31599 ;
  assign n31612 = ( n31609 & ~n31611 ) | ( n31609 & n31610 ) | ( ~n31611 & n31610 ) ;
  assign n31616 = n31150 &  n31240 ;
  assign n31617 = n31239 &  n31616 ;
  assign n31605 = x70 | n31150 ;
  assign n31606 = x70 &  n31150 ;
  assign n31607 = ( n31605 & ~n31606 ) | ( n31605 & 1'b0 ) | ( ~n31606 & 1'b0 ) ;
  assign n31619 = ( n31188 & n31241 ) | ( n31188 & n31607 ) | ( n31241 & n31607 ) ;
  assign n31618 = n31188 | n31607 ;
  assign n31620 = ( n31617 & ~n31619 ) | ( n31617 & n31618 ) | ( ~n31619 & n31618 ) ;
  assign n31624 = n31158 &  n31240 ;
  assign n31625 = n31239 &  n31624 ;
  assign n31613 = x69 | n31158 ;
  assign n31614 = x69 &  n31158 ;
  assign n31615 = ( n31613 & ~n31614 ) | ( n31613 & 1'b0 ) | ( ~n31614 & 1'b0 ) ;
  assign n31627 = ( n31187 & n31241 ) | ( n31187 & n31615 ) | ( n31241 & n31615 ) ;
  assign n31626 = n31187 | n31615 ;
  assign n31628 = ( n31625 & ~n31627 ) | ( n31625 & n31626 ) | ( ~n31627 & n31626 ) ;
  assign n31632 = n31166 &  n31240 ;
  assign n31633 = n31239 &  n31632 ;
  assign n31621 = x68 | n31166 ;
  assign n31622 = x68 &  n31166 ;
  assign n31623 = ( n31621 & ~n31622 ) | ( n31621 & 1'b0 ) | ( ~n31622 & 1'b0 ) ;
  assign n31635 = ( n31186 & n31241 ) | ( n31186 & n31623 ) | ( n31241 & n31623 ) ;
  assign n31634 = n31186 | n31623 ;
  assign n31636 = ( n31633 & ~n31635 ) | ( n31633 & n31634 ) | ( ~n31635 & n31634 ) ;
  assign n31640 = n31171 &  n31240 ;
  assign n31641 = n31239 &  n31640 ;
  assign n31629 = x67 | n31171 ;
  assign n31630 = x67 &  n31171 ;
  assign n31631 = ( n31629 & ~n31630 ) | ( n31629 & 1'b0 ) | ( ~n31630 & 1'b0 ) ;
  assign n31643 = ( n31185 & n31241 ) | ( n31185 & n31631 ) | ( n31241 & n31631 ) ;
  assign n31642 = n31185 | n31631 ;
  assign n31644 = ( n31641 & ~n31643 ) | ( n31641 & n31642 ) | ( ~n31643 & n31642 ) ;
  assign n31645 = n31179 &  n31240 ;
  assign n31646 = n31239 &  n31645 ;
  assign n31637 = x66 | n31179 ;
  assign n31638 = x66 &  n31179 ;
  assign n31639 = ( n31637 & ~n31638 ) | ( n31637 & 1'b0 ) | ( ~n31638 & 1'b0 ) ;
  assign n31648 = ( n31184 & n31241 ) | ( n31184 & n31639 ) | ( n31241 & n31639 ) ;
  assign n31647 = n31184 | n31639 ;
  assign n31649 = ( n31646 & ~n31648 ) | ( n31646 & n31647 ) | ( ~n31648 & n31647 ) ;
  assign n31650 = ( x65 & ~n12811 ) | ( x65 & n31183 ) | ( ~n12811 & n31183 ) ;
  assign n31651 = ( n31184 & ~x65 ) | ( n31184 & n31650 ) | ( ~x65 & n31650 ) ;
  assign n31652 = ~n31241 & n31651 ;
  assign n31653 = n31183 &  n31240 ;
  assign n31654 = n31239 &  n31653 ;
  assign n31655 = n31652 | n31654 ;
  assign n31656 = ( x64 & ~n31241 ) | ( x64 & 1'b0 ) | ( ~n31241 & 1'b0 ) ;
  assign n31657 = ( x11 & ~n31656 ) | ( x11 & 1'b0 ) | ( ~n31656 & 1'b0 ) ;
  assign n31658 = ( n12811 & ~n31241 ) | ( n12811 & 1'b0 ) | ( ~n31241 & 1'b0 ) ;
  assign n31659 = n31657 | n31658 ;
  assign n31660 = ( x65 & ~n31659 ) | ( x65 & n13294 ) | ( ~n31659 & n13294 ) ;
  assign n31661 = ( x66 & ~n31655 ) | ( x66 & n31660 ) | ( ~n31655 & n31660 ) ;
  assign n31662 = ( x67 & ~n31649 ) | ( x67 & n31661 ) | ( ~n31649 & n31661 ) ;
  assign n31663 = ( x68 & ~n31644 ) | ( x68 & n31662 ) | ( ~n31644 & n31662 ) ;
  assign n31664 = ( x69 & ~n31636 ) | ( x69 & n31663 ) | ( ~n31636 & n31663 ) ;
  assign n31665 = ( x70 & ~n31628 ) | ( x70 & n31664 ) | ( ~n31628 & n31664 ) ;
  assign n31666 = ( x71 & ~n31620 ) | ( x71 & n31665 ) | ( ~n31620 & n31665 ) ;
  assign n31667 = ( x72 & ~n31612 ) | ( x72 & n31666 ) | ( ~n31612 & n31666 ) ;
  assign n31668 = ( x73 & ~n31604 ) | ( x73 & n31667 ) | ( ~n31604 & n31667 ) ;
  assign n31669 = ( x74 & ~n31596 ) | ( x74 & n31668 ) | ( ~n31596 & n31668 ) ;
  assign n31670 = ( x75 & ~n31588 ) | ( x75 & n31669 ) | ( ~n31588 & n31669 ) ;
  assign n31671 = ( x76 & ~n31580 ) | ( x76 & n31670 ) | ( ~n31580 & n31670 ) ;
  assign n31672 = ( x77 & ~n31572 ) | ( x77 & n31671 ) | ( ~n31572 & n31671 ) ;
  assign n31673 = ( x78 & ~n31564 ) | ( x78 & n31672 ) | ( ~n31564 & n31672 ) ;
  assign n31674 = ( x79 & ~n31556 ) | ( x79 & n31673 ) | ( ~n31556 & n31673 ) ;
  assign n31675 = ( x80 & ~n31548 ) | ( x80 & n31674 ) | ( ~n31548 & n31674 ) ;
  assign n31676 = ( x81 & ~n31540 ) | ( x81 & n31675 ) | ( ~n31540 & n31675 ) ;
  assign n31677 = ( x82 & ~n31532 ) | ( x82 & n31676 ) | ( ~n31532 & n31676 ) ;
  assign n31678 = ( x83 & ~n31524 ) | ( x83 & n31677 ) | ( ~n31524 & n31677 ) ;
  assign n31679 = ( x84 & ~n31516 ) | ( x84 & n31678 ) | ( ~n31516 & n31678 ) ;
  assign n31680 = ( x85 & ~n31508 ) | ( x85 & n31679 ) | ( ~n31508 & n31679 ) ;
  assign n31681 = ( x86 & ~n31500 ) | ( x86 & n31680 ) | ( ~n31500 & n31680 ) ;
  assign n31682 = ( x87 & ~n31492 ) | ( x87 & n31681 ) | ( ~n31492 & n31681 ) ;
  assign n31683 = ( x88 & ~n31484 ) | ( x88 & n31682 ) | ( ~n31484 & n31682 ) ;
  assign n31684 = ( x89 & ~n31476 ) | ( x89 & n31683 ) | ( ~n31476 & n31683 ) ;
  assign n31685 = ( x90 & ~n31468 ) | ( x90 & n31684 ) | ( ~n31468 & n31684 ) ;
  assign n31686 = ( x91 & ~n31460 ) | ( x91 & n31685 ) | ( ~n31460 & n31685 ) ;
  assign n31687 = ( x92 & ~n31452 ) | ( x92 & n31686 ) | ( ~n31452 & n31686 ) ;
  assign n31688 = ( x93 & ~n31444 ) | ( x93 & n31687 ) | ( ~n31444 & n31687 ) ;
  assign n31689 = ( x94 & ~n31436 ) | ( x94 & n31688 ) | ( ~n31436 & n31688 ) ;
  assign n31690 = ( x95 & ~n31428 ) | ( x95 & n31689 ) | ( ~n31428 & n31689 ) ;
  assign n31691 = ( x96 & ~n31420 ) | ( x96 & n31690 ) | ( ~n31420 & n31690 ) ;
  assign n31692 = ( x97 & ~n31412 ) | ( x97 & n31691 ) | ( ~n31412 & n31691 ) ;
  assign n31693 = ( x98 & ~n31404 ) | ( x98 & n31692 ) | ( ~n31404 & n31692 ) ;
  assign n31694 = ( x99 & ~n31396 ) | ( x99 & n31693 ) | ( ~n31396 & n31693 ) ;
  assign n31695 = ( x100 & ~n31388 ) | ( x100 & n31694 ) | ( ~n31388 & n31694 ) ;
  assign n31696 = ( x101 & ~n31380 ) | ( x101 & n31695 ) | ( ~n31380 & n31695 ) ;
  assign n31697 = ( x102 & ~n31372 ) | ( x102 & n31696 ) | ( ~n31372 & n31696 ) ;
  assign n31698 = ( x103 & ~n31364 ) | ( x103 & n31697 ) | ( ~n31364 & n31697 ) ;
  assign n31699 = ( x104 & ~n31356 ) | ( x104 & n31698 ) | ( ~n31356 & n31698 ) ;
  assign n31700 = ( x105 & ~n31348 ) | ( x105 & n31699 ) | ( ~n31348 & n31699 ) ;
  assign n31701 = ( x106 & ~n31340 ) | ( x106 & n31700 ) | ( ~n31340 & n31700 ) ;
  assign n31702 = ( x107 & ~n31332 ) | ( x107 & n31701 ) | ( ~n31332 & n31701 ) ;
  assign n31703 = ( x108 & ~n31324 ) | ( x108 & n31702 ) | ( ~n31324 & n31702 ) ;
  assign n31704 = ( x109 & ~n31316 ) | ( x109 & n31703 ) | ( ~n31316 & n31703 ) ;
  assign n31705 = ( x110 & ~n31308 ) | ( x110 & n31704 ) | ( ~n31308 & n31704 ) ;
  assign n31706 = ( x111 & ~n31300 ) | ( x111 & n31705 ) | ( ~n31300 & n31705 ) ;
  assign n31707 = ( x112 & ~n31292 ) | ( x112 & n31706 ) | ( ~n31292 & n31706 ) ;
  assign n31708 = ( x113 & ~n31284 ) | ( x113 & n31707 ) | ( ~n31284 & n31707 ) ;
  assign n31709 = ( x114 & ~n31276 ) | ( x114 & n31708 ) | ( ~n31276 & n31708 ) ;
  assign n31710 = ( x115 & ~n31268 ) | ( x115 & n31709 ) | ( ~n31268 & n31709 ) ;
  assign n31711 = ( x116 & ~n31260 ) | ( x116 & n31710 ) | ( ~n31260 & n31710 ) ;
  assign n31712 = ( x117 & ~n31250 ) | ( x117 & 1'b0 ) | ( ~n31250 & 1'b0 ) ;
  assign n31713 = ~n31248 & n31712 ;
  assign n31714 = ( n31711 & ~n31252 ) | ( n31711 & n31713 ) | ( ~n31252 & n31713 ) ;
  assign n31715 = ( n31252 & ~n13416 ) | ( n31252 & n31714 ) | ( ~n13416 & n31714 ) ;
  assign n31716 = n13416 | n31715 ;
  assign n31717 = ~n31251 |  n425 ;
  assign n31731 = n31260 &  n31717 ;
  assign n31732 = n31716 &  n31731 ;
  assign n31718 = n31716 &  n31717 ;
  assign n31719 = x116 | n31260 ;
  assign n31720 = x116 &  n31260 ;
  assign n31721 = ( n31719 & ~n31720 ) | ( n31719 & 1'b0 ) | ( ~n31720 & 1'b0 ) ;
  assign n31734 = ( n31710 & n31718 ) | ( n31710 & n31721 ) | ( n31718 & n31721 ) ;
  assign n31733 = n31710 | n31721 ;
  assign n31735 = ( n31732 & ~n31734 ) | ( n31732 & n31733 ) | ( ~n31734 & n31733 ) ;
  assign n31723 = n425 &  n31251 ;
  assign n31724 = n31716 &  n31723 ;
  assign n31722 = n31252 | n31713 ;
  assign n31726 = ( n31711 & n31718 ) | ( n31711 & n31722 ) | ( n31718 & n31722 ) ;
  assign n31725 = n31711 | n31722 ;
  assign n31727 = ( n31724 & ~n31726 ) | ( n31724 & n31725 ) | ( ~n31726 & n31725 ) ;
  assign n31739 = n31268 &  n31717 ;
  assign n31740 = n31716 &  n31739 ;
  assign n31728 = x115 | n31268 ;
  assign n31729 = x115 &  n31268 ;
  assign n31730 = ( n31728 & ~n31729 ) | ( n31728 & 1'b0 ) | ( ~n31729 & 1'b0 ) ;
  assign n31742 = ( n31709 & n31718 ) | ( n31709 & n31730 ) | ( n31718 & n31730 ) ;
  assign n31741 = n31709 | n31730 ;
  assign n31743 = ( n31740 & ~n31742 ) | ( n31740 & n31741 ) | ( ~n31742 & n31741 ) ;
  assign n31747 = n31276 &  n31717 ;
  assign n31748 = n31716 &  n31747 ;
  assign n31736 = x114 | n31276 ;
  assign n31737 = x114 &  n31276 ;
  assign n31738 = ( n31736 & ~n31737 ) | ( n31736 & 1'b0 ) | ( ~n31737 & 1'b0 ) ;
  assign n31750 = ( n31708 & n31718 ) | ( n31708 & n31738 ) | ( n31718 & n31738 ) ;
  assign n31749 = n31708 | n31738 ;
  assign n31751 = ( n31748 & ~n31750 ) | ( n31748 & n31749 ) | ( ~n31750 & n31749 ) ;
  assign n31755 = n31284 &  n31717 ;
  assign n31756 = n31716 &  n31755 ;
  assign n31744 = x113 | n31284 ;
  assign n31745 = x113 &  n31284 ;
  assign n31746 = ( n31744 & ~n31745 ) | ( n31744 & 1'b0 ) | ( ~n31745 & 1'b0 ) ;
  assign n31758 = ( n31707 & n31718 ) | ( n31707 & n31746 ) | ( n31718 & n31746 ) ;
  assign n31757 = n31707 | n31746 ;
  assign n31759 = ( n31756 & ~n31758 ) | ( n31756 & n31757 ) | ( ~n31758 & n31757 ) ;
  assign n31763 = n31292 &  n31717 ;
  assign n31764 = n31716 &  n31763 ;
  assign n31752 = x112 | n31292 ;
  assign n31753 = x112 &  n31292 ;
  assign n31754 = ( n31752 & ~n31753 ) | ( n31752 & 1'b0 ) | ( ~n31753 & 1'b0 ) ;
  assign n31766 = ( n31706 & n31718 ) | ( n31706 & n31754 ) | ( n31718 & n31754 ) ;
  assign n31765 = n31706 | n31754 ;
  assign n31767 = ( n31764 & ~n31766 ) | ( n31764 & n31765 ) | ( ~n31766 & n31765 ) ;
  assign n31771 = n31300 &  n31717 ;
  assign n31772 = n31716 &  n31771 ;
  assign n31760 = x111 | n31300 ;
  assign n31761 = x111 &  n31300 ;
  assign n31762 = ( n31760 & ~n31761 ) | ( n31760 & 1'b0 ) | ( ~n31761 & 1'b0 ) ;
  assign n31774 = ( n31705 & n31718 ) | ( n31705 & n31762 ) | ( n31718 & n31762 ) ;
  assign n31773 = n31705 | n31762 ;
  assign n31775 = ( n31772 & ~n31774 ) | ( n31772 & n31773 ) | ( ~n31774 & n31773 ) ;
  assign n31779 = n31308 &  n31717 ;
  assign n31780 = n31716 &  n31779 ;
  assign n31768 = x110 | n31308 ;
  assign n31769 = x110 &  n31308 ;
  assign n31770 = ( n31768 & ~n31769 ) | ( n31768 & 1'b0 ) | ( ~n31769 & 1'b0 ) ;
  assign n31782 = ( n31704 & n31718 ) | ( n31704 & n31770 ) | ( n31718 & n31770 ) ;
  assign n31781 = n31704 | n31770 ;
  assign n31783 = ( n31780 & ~n31782 ) | ( n31780 & n31781 ) | ( ~n31782 & n31781 ) ;
  assign n31787 = n31316 &  n31717 ;
  assign n31788 = n31716 &  n31787 ;
  assign n31776 = x109 | n31316 ;
  assign n31777 = x109 &  n31316 ;
  assign n31778 = ( n31776 & ~n31777 ) | ( n31776 & 1'b0 ) | ( ~n31777 & 1'b0 ) ;
  assign n31790 = ( n31703 & n31718 ) | ( n31703 & n31778 ) | ( n31718 & n31778 ) ;
  assign n31789 = n31703 | n31778 ;
  assign n31791 = ( n31788 & ~n31790 ) | ( n31788 & n31789 ) | ( ~n31790 & n31789 ) ;
  assign n31795 = n31324 &  n31717 ;
  assign n31796 = n31716 &  n31795 ;
  assign n31784 = x108 | n31324 ;
  assign n31785 = x108 &  n31324 ;
  assign n31786 = ( n31784 & ~n31785 ) | ( n31784 & 1'b0 ) | ( ~n31785 & 1'b0 ) ;
  assign n31798 = ( n31702 & n31718 ) | ( n31702 & n31786 ) | ( n31718 & n31786 ) ;
  assign n31797 = n31702 | n31786 ;
  assign n31799 = ( n31796 & ~n31798 ) | ( n31796 & n31797 ) | ( ~n31798 & n31797 ) ;
  assign n31803 = n31332 &  n31717 ;
  assign n31804 = n31716 &  n31803 ;
  assign n31792 = x107 | n31332 ;
  assign n31793 = x107 &  n31332 ;
  assign n31794 = ( n31792 & ~n31793 ) | ( n31792 & 1'b0 ) | ( ~n31793 & 1'b0 ) ;
  assign n31806 = ( n31701 & n31718 ) | ( n31701 & n31794 ) | ( n31718 & n31794 ) ;
  assign n31805 = n31701 | n31794 ;
  assign n31807 = ( n31804 & ~n31806 ) | ( n31804 & n31805 ) | ( ~n31806 & n31805 ) ;
  assign n31811 = n31340 &  n31717 ;
  assign n31812 = n31716 &  n31811 ;
  assign n31800 = x106 | n31340 ;
  assign n31801 = x106 &  n31340 ;
  assign n31802 = ( n31800 & ~n31801 ) | ( n31800 & 1'b0 ) | ( ~n31801 & 1'b0 ) ;
  assign n31814 = ( n31700 & n31718 ) | ( n31700 & n31802 ) | ( n31718 & n31802 ) ;
  assign n31813 = n31700 | n31802 ;
  assign n31815 = ( n31812 & ~n31814 ) | ( n31812 & n31813 ) | ( ~n31814 & n31813 ) ;
  assign n31819 = n31348 &  n31717 ;
  assign n31820 = n31716 &  n31819 ;
  assign n31808 = x105 | n31348 ;
  assign n31809 = x105 &  n31348 ;
  assign n31810 = ( n31808 & ~n31809 ) | ( n31808 & 1'b0 ) | ( ~n31809 & 1'b0 ) ;
  assign n31822 = ( n31699 & n31718 ) | ( n31699 & n31810 ) | ( n31718 & n31810 ) ;
  assign n31821 = n31699 | n31810 ;
  assign n31823 = ( n31820 & ~n31822 ) | ( n31820 & n31821 ) | ( ~n31822 & n31821 ) ;
  assign n31827 = n31356 &  n31717 ;
  assign n31828 = n31716 &  n31827 ;
  assign n31816 = x104 | n31356 ;
  assign n31817 = x104 &  n31356 ;
  assign n31818 = ( n31816 & ~n31817 ) | ( n31816 & 1'b0 ) | ( ~n31817 & 1'b0 ) ;
  assign n31830 = ( n31698 & n31718 ) | ( n31698 & n31818 ) | ( n31718 & n31818 ) ;
  assign n31829 = n31698 | n31818 ;
  assign n31831 = ( n31828 & ~n31830 ) | ( n31828 & n31829 ) | ( ~n31830 & n31829 ) ;
  assign n31835 = n31364 &  n31717 ;
  assign n31836 = n31716 &  n31835 ;
  assign n31824 = x103 | n31364 ;
  assign n31825 = x103 &  n31364 ;
  assign n31826 = ( n31824 & ~n31825 ) | ( n31824 & 1'b0 ) | ( ~n31825 & 1'b0 ) ;
  assign n31838 = ( n31697 & n31718 ) | ( n31697 & n31826 ) | ( n31718 & n31826 ) ;
  assign n31837 = n31697 | n31826 ;
  assign n31839 = ( n31836 & ~n31838 ) | ( n31836 & n31837 ) | ( ~n31838 & n31837 ) ;
  assign n31843 = n31372 &  n31717 ;
  assign n31844 = n31716 &  n31843 ;
  assign n31832 = x102 | n31372 ;
  assign n31833 = x102 &  n31372 ;
  assign n31834 = ( n31832 & ~n31833 ) | ( n31832 & 1'b0 ) | ( ~n31833 & 1'b0 ) ;
  assign n31846 = ( n31696 & n31718 ) | ( n31696 & n31834 ) | ( n31718 & n31834 ) ;
  assign n31845 = n31696 | n31834 ;
  assign n31847 = ( n31844 & ~n31846 ) | ( n31844 & n31845 ) | ( ~n31846 & n31845 ) ;
  assign n31851 = n31380 &  n31717 ;
  assign n31852 = n31716 &  n31851 ;
  assign n31840 = x101 | n31380 ;
  assign n31841 = x101 &  n31380 ;
  assign n31842 = ( n31840 & ~n31841 ) | ( n31840 & 1'b0 ) | ( ~n31841 & 1'b0 ) ;
  assign n31854 = ( n31695 & n31718 ) | ( n31695 & n31842 ) | ( n31718 & n31842 ) ;
  assign n31853 = n31695 | n31842 ;
  assign n31855 = ( n31852 & ~n31854 ) | ( n31852 & n31853 ) | ( ~n31854 & n31853 ) ;
  assign n31859 = n31388 &  n31717 ;
  assign n31860 = n31716 &  n31859 ;
  assign n31848 = x100 | n31388 ;
  assign n31849 = x100 &  n31388 ;
  assign n31850 = ( n31848 & ~n31849 ) | ( n31848 & 1'b0 ) | ( ~n31849 & 1'b0 ) ;
  assign n31862 = ( n31694 & n31718 ) | ( n31694 & n31850 ) | ( n31718 & n31850 ) ;
  assign n31861 = n31694 | n31850 ;
  assign n31863 = ( n31860 & ~n31862 ) | ( n31860 & n31861 ) | ( ~n31862 & n31861 ) ;
  assign n31867 = n31396 &  n31717 ;
  assign n31868 = n31716 &  n31867 ;
  assign n31856 = x99 | n31396 ;
  assign n31857 = x99 &  n31396 ;
  assign n31858 = ( n31856 & ~n31857 ) | ( n31856 & 1'b0 ) | ( ~n31857 & 1'b0 ) ;
  assign n31870 = ( n31693 & n31718 ) | ( n31693 & n31858 ) | ( n31718 & n31858 ) ;
  assign n31869 = n31693 | n31858 ;
  assign n31871 = ( n31868 & ~n31870 ) | ( n31868 & n31869 ) | ( ~n31870 & n31869 ) ;
  assign n31875 = n31404 &  n31717 ;
  assign n31876 = n31716 &  n31875 ;
  assign n31864 = x98 | n31404 ;
  assign n31865 = x98 &  n31404 ;
  assign n31866 = ( n31864 & ~n31865 ) | ( n31864 & 1'b0 ) | ( ~n31865 & 1'b0 ) ;
  assign n31878 = ( n31692 & n31718 ) | ( n31692 & n31866 ) | ( n31718 & n31866 ) ;
  assign n31877 = n31692 | n31866 ;
  assign n31879 = ( n31876 & ~n31878 ) | ( n31876 & n31877 ) | ( ~n31878 & n31877 ) ;
  assign n31883 = n31412 &  n31717 ;
  assign n31884 = n31716 &  n31883 ;
  assign n31872 = x97 | n31412 ;
  assign n31873 = x97 &  n31412 ;
  assign n31874 = ( n31872 & ~n31873 ) | ( n31872 & 1'b0 ) | ( ~n31873 & 1'b0 ) ;
  assign n31886 = ( n31691 & n31718 ) | ( n31691 & n31874 ) | ( n31718 & n31874 ) ;
  assign n31885 = n31691 | n31874 ;
  assign n31887 = ( n31884 & ~n31886 ) | ( n31884 & n31885 ) | ( ~n31886 & n31885 ) ;
  assign n31891 = n31420 &  n31717 ;
  assign n31892 = n31716 &  n31891 ;
  assign n31880 = x96 | n31420 ;
  assign n31881 = x96 &  n31420 ;
  assign n31882 = ( n31880 & ~n31881 ) | ( n31880 & 1'b0 ) | ( ~n31881 & 1'b0 ) ;
  assign n31894 = ( n31690 & n31718 ) | ( n31690 & n31882 ) | ( n31718 & n31882 ) ;
  assign n31893 = n31690 | n31882 ;
  assign n31895 = ( n31892 & ~n31894 ) | ( n31892 & n31893 ) | ( ~n31894 & n31893 ) ;
  assign n31899 = n31428 &  n31717 ;
  assign n31900 = n31716 &  n31899 ;
  assign n31888 = x95 | n31428 ;
  assign n31889 = x95 &  n31428 ;
  assign n31890 = ( n31888 & ~n31889 ) | ( n31888 & 1'b0 ) | ( ~n31889 & 1'b0 ) ;
  assign n31902 = ( n31689 & n31718 ) | ( n31689 & n31890 ) | ( n31718 & n31890 ) ;
  assign n31901 = n31689 | n31890 ;
  assign n31903 = ( n31900 & ~n31902 ) | ( n31900 & n31901 ) | ( ~n31902 & n31901 ) ;
  assign n31907 = n31436 &  n31717 ;
  assign n31908 = n31716 &  n31907 ;
  assign n31896 = x94 | n31436 ;
  assign n31897 = x94 &  n31436 ;
  assign n31898 = ( n31896 & ~n31897 ) | ( n31896 & 1'b0 ) | ( ~n31897 & 1'b0 ) ;
  assign n31910 = ( n31688 & n31718 ) | ( n31688 & n31898 ) | ( n31718 & n31898 ) ;
  assign n31909 = n31688 | n31898 ;
  assign n31911 = ( n31908 & ~n31910 ) | ( n31908 & n31909 ) | ( ~n31910 & n31909 ) ;
  assign n31915 = n31444 &  n31717 ;
  assign n31916 = n31716 &  n31915 ;
  assign n31904 = x93 | n31444 ;
  assign n31905 = x93 &  n31444 ;
  assign n31906 = ( n31904 & ~n31905 ) | ( n31904 & 1'b0 ) | ( ~n31905 & 1'b0 ) ;
  assign n31918 = ( n31687 & n31718 ) | ( n31687 & n31906 ) | ( n31718 & n31906 ) ;
  assign n31917 = n31687 | n31906 ;
  assign n31919 = ( n31916 & ~n31918 ) | ( n31916 & n31917 ) | ( ~n31918 & n31917 ) ;
  assign n31923 = n31452 &  n31717 ;
  assign n31924 = n31716 &  n31923 ;
  assign n31912 = x92 | n31452 ;
  assign n31913 = x92 &  n31452 ;
  assign n31914 = ( n31912 & ~n31913 ) | ( n31912 & 1'b0 ) | ( ~n31913 & 1'b0 ) ;
  assign n31926 = ( n31686 & n31718 ) | ( n31686 & n31914 ) | ( n31718 & n31914 ) ;
  assign n31925 = n31686 | n31914 ;
  assign n31927 = ( n31924 & ~n31926 ) | ( n31924 & n31925 ) | ( ~n31926 & n31925 ) ;
  assign n31931 = n31460 &  n31717 ;
  assign n31932 = n31716 &  n31931 ;
  assign n31920 = x91 | n31460 ;
  assign n31921 = x91 &  n31460 ;
  assign n31922 = ( n31920 & ~n31921 ) | ( n31920 & 1'b0 ) | ( ~n31921 & 1'b0 ) ;
  assign n31934 = ( n31685 & n31718 ) | ( n31685 & n31922 ) | ( n31718 & n31922 ) ;
  assign n31933 = n31685 | n31922 ;
  assign n31935 = ( n31932 & ~n31934 ) | ( n31932 & n31933 ) | ( ~n31934 & n31933 ) ;
  assign n31939 = n31468 &  n31717 ;
  assign n31940 = n31716 &  n31939 ;
  assign n31928 = x90 | n31468 ;
  assign n31929 = x90 &  n31468 ;
  assign n31930 = ( n31928 & ~n31929 ) | ( n31928 & 1'b0 ) | ( ~n31929 & 1'b0 ) ;
  assign n31942 = ( n31684 & n31718 ) | ( n31684 & n31930 ) | ( n31718 & n31930 ) ;
  assign n31941 = n31684 | n31930 ;
  assign n31943 = ( n31940 & ~n31942 ) | ( n31940 & n31941 ) | ( ~n31942 & n31941 ) ;
  assign n31947 = n31476 &  n31717 ;
  assign n31948 = n31716 &  n31947 ;
  assign n31936 = x89 | n31476 ;
  assign n31937 = x89 &  n31476 ;
  assign n31938 = ( n31936 & ~n31937 ) | ( n31936 & 1'b0 ) | ( ~n31937 & 1'b0 ) ;
  assign n31950 = ( n31683 & n31718 ) | ( n31683 & n31938 ) | ( n31718 & n31938 ) ;
  assign n31949 = n31683 | n31938 ;
  assign n31951 = ( n31948 & ~n31950 ) | ( n31948 & n31949 ) | ( ~n31950 & n31949 ) ;
  assign n31955 = n31484 &  n31717 ;
  assign n31956 = n31716 &  n31955 ;
  assign n31944 = x88 | n31484 ;
  assign n31945 = x88 &  n31484 ;
  assign n31946 = ( n31944 & ~n31945 ) | ( n31944 & 1'b0 ) | ( ~n31945 & 1'b0 ) ;
  assign n31958 = ( n31682 & n31718 ) | ( n31682 & n31946 ) | ( n31718 & n31946 ) ;
  assign n31957 = n31682 | n31946 ;
  assign n31959 = ( n31956 & ~n31958 ) | ( n31956 & n31957 ) | ( ~n31958 & n31957 ) ;
  assign n31963 = n31492 &  n31717 ;
  assign n31964 = n31716 &  n31963 ;
  assign n31952 = x87 | n31492 ;
  assign n31953 = x87 &  n31492 ;
  assign n31954 = ( n31952 & ~n31953 ) | ( n31952 & 1'b0 ) | ( ~n31953 & 1'b0 ) ;
  assign n31966 = ( n31681 & n31718 ) | ( n31681 & n31954 ) | ( n31718 & n31954 ) ;
  assign n31965 = n31681 | n31954 ;
  assign n31967 = ( n31964 & ~n31966 ) | ( n31964 & n31965 ) | ( ~n31966 & n31965 ) ;
  assign n31971 = n31500 &  n31717 ;
  assign n31972 = n31716 &  n31971 ;
  assign n31960 = x86 | n31500 ;
  assign n31961 = x86 &  n31500 ;
  assign n31962 = ( n31960 & ~n31961 ) | ( n31960 & 1'b0 ) | ( ~n31961 & 1'b0 ) ;
  assign n31974 = ( n31680 & n31718 ) | ( n31680 & n31962 ) | ( n31718 & n31962 ) ;
  assign n31973 = n31680 | n31962 ;
  assign n31975 = ( n31972 & ~n31974 ) | ( n31972 & n31973 ) | ( ~n31974 & n31973 ) ;
  assign n31979 = n31508 &  n31717 ;
  assign n31980 = n31716 &  n31979 ;
  assign n31968 = x85 | n31508 ;
  assign n31969 = x85 &  n31508 ;
  assign n31970 = ( n31968 & ~n31969 ) | ( n31968 & 1'b0 ) | ( ~n31969 & 1'b0 ) ;
  assign n31982 = ( n31679 & n31718 ) | ( n31679 & n31970 ) | ( n31718 & n31970 ) ;
  assign n31981 = n31679 | n31970 ;
  assign n31983 = ( n31980 & ~n31982 ) | ( n31980 & n31981 ) | ( ~n31982 & n31981 ) ;
  assign n31987 = n31516 &  n31717 ;
  assign n31988 = n31716 &  n31987 ;
  assign n31976 = x84 | n31516 ;
  assign n31977 = x84 &  n31516 ;
  assign n31978 = ( n31976 & ~n31977 ) | ( n31976 & 1'b0 ) | ( ~n31977 & 1'b0 ) ;
  assign n31990 = ( n31678 & n31718 ) | ( n31678 & n31978 ) | ( n31718 & n31978 ) ;
  assign n31989 = n31678 | n31978 ;
  assign n31991 = ( n31988 & ~n31990 ) | ( n31988 & n31989 ) | ( ~n31990 & n31989 ) ;
  assign n31995 = n31524 &  n31717 ;
  assign n31996 = n31716 &  n31995 ;
  assign n31984 = x83 | n31524 ;
  assign n31985 = x83 &  n31524 ;
  assign n31986 = ( n31984 & ~n31985 ) | ( n31984 & 1'b0 ) | ( ~n31985 & 1'b0 ) ;
  assign n31998 = ( n31677 & n31718 ) | ( n31677 & n31986 ) | ( n31718 & n31986 ) ;
  assign n31997 = n31677 | n31986 ;
  assign n31999 = ( n31996 & ~n31998 ) | ( n31996 & n31997 ) | ( ~n31998 & n31997 ) ;
  assign n32003 = n31532 &  n31717 ;
  assign n32004 = n31716 &  n32003 ;
  assign n31992 = x82 | n31532 ;
  assign n31993 = x82 &  n31532 ;
  assign n31994 = ( n31992 & ~n31993 ) | ( n31992 & 1'b0 ) | ( ~n31993 & 1'b0 ) ;
  assign n32006 = ( n31676 & n31718 ) | ( n31676 & n31994 ) | ( n31718 & n31994 ) ;
  assign n32005 = n31676 | n31994 ;
  assign n32007 = ( n32004 & ~n32006 ) | ( n32004 & n32005 ) | ( ~n32006 & n32005 ) ;
  assign n32011 = n31540 &  n31717 ;
  assign n32012 = n31716 &  n32011 ;
  assign n32000 = x81 | n31540 ;
  assign n32001 = x81 &  n31540 ;
  assign n32002 = ( n32000 & ~n32001 ) | ( n32000 & 1'b0 ) | ( ~n32001 & 1'b0 ) ;
  assign n32014 = ( n31675 & n31718 ) | ( n31675 & n32002 ) | ( n31718 & n32002 ) ;
  assign n32013 = n31675 | n32002 ;
  assign n32015 = ( n32012 & ~n32014 ) | ( n32012 & n32013 ) | ( ~n32014 & n32013 ) ;
  assign n32019 = n31548 &  n31717 ;
  assign n32020 = n31716 &  n32019 ;
  assign n32008 = x80 | n31548 ;
  assign n32009 = x80 &  n31548 ;
  assign n32010 = ( n32008 & ~n32009 ) | ( n32008 & 1'b0 ) | ( ~n32009 & 1'b0 ) ;
  assign n32022 = ( n31674 & n31718 ) | ( n31674 & n32010 ) | ( n31718 & n32010 ) ;
  assign n32021 = n31674 | n32010 ;
  assign n32023 = ( n32020 & ~n32022 ) | ( n32020 & n32021 ) | ( ~n32022 & n32021 ) ;
  assign n32027 = n31556 &  n31717 ;
  assign n32028 = n31716 &  n32027 ;
  assign n32016 = x79 | n31556 ;
  assign n32017 = x79 &  n31556 ;
  assign n32018 = ( n32016 & ~n32017 ) | ( n32016 & 1'b0 ) | ( ~n32017 & 1'b0 ) ;
  assign n32030 = ( n31673 & n31718 ) | ( n31673 & n32018 ) | ( n31718 & n32018 ) ;
  assign n32029 = n31673 | n32018 ;
  assign n32031 = ( n32028 & ~n32030 ) | ( n32028 & n32029 ) | ( ~n32030 & n32029 ) ;
  assign n32035 = n31564 &  n31717 ;
  assign n32036 = n31716 &  n32035 ;
  assign n32024 = x78 | n31564 ;
  assign n32025 = x78 &  n31564 ;
  assign n32026 = ( n32024 & ~n32025 ) | ( n32024 & 1'b0 ) | ( ~n32025 & 1'b0 ) ;
  assign n32038 = ( n31672 & n31718 ) | ( n31672 & n32026 ) | ( n31718 & n32026 ) ;
  assign n32037 = n31672 | n32026 ;
  assign n32039 = ( n32036 & ~n32038 ) | ( n32036 & n32037 ) | ( ~n32038 & n32037 ) ;
  assign n32043 = n31572 &  n31717 ;
  assign n32044 = n31716 &  n32043 ;
  assign n32032 = x77 | n31572 ;
  assign n32033 = x77 &  n31572 ;
  assign n32034 = ( n32032 & ~n32033 ) | ( n32032 & 1'b0 ) | ( ~n32033 & 1'b0 ) ;
  assign n32046 = ( n31671 & n31718 ) | ( n31671 & n32034 ) | ( n31718 & n32034 ) ;
  assign n32045 = n31671 | n32034 ;
  assign n32047 = ( n32044 & ~n32046 ) | ( n32044 & n32045 ) | ( ~n32046 & n32045 ) ;
  assign n32051 = n31580 &  n31717 ;
  assign n32052 = n31716 &  n32051 ;
  assign n32040 = x76 | n31580 ;
  assign n32041 = x76 &  n31580 ;
  assign n32042 = ( n32040 & ~n32041 ) | ( n32040 & 1'b0 ) | ( ~n32041 & 1'b0 ) ;
  assign n32054 = ( n31670 & n31718 ) | ( n31670 & n32042 ) | ( n31718 & n32042 ) ;
  assign n32053 = n31670 | n32042 ;
  assign n32055 = ( n32052 & ~n32054 ) | ( n32052 & n32053 ) | ( ~n32054 & n32053 ) ;
  assign n32059 = n31588 &  n31717 ;
  assign n32060 = n31716 &  n32059 ;
  assign n32048 = x75 | n31588 ;
  assign n32049 = x75 &  n31588 ;
  assign n32050 = ( n32048 & ~n32049 ) | ( n32048 & 1'b0 ) | ( ~n32049 & 1'b0 ) ;
  assign n32062 = ( n31669 & n31718 ) | ( n31669 & n32050 ) | ( n31718 & n32050 ) ;
  assign n32061 = n31669 | n32050 ;
  assign n32063 = ( n32060 & ~n32062 ) | ( n32060 & n32061 ) | ( ~n32062 & n32061 ) ;
  assign n32067 = n31596 &  n31717 ;
  assign n32068 = n31716 &  n32067 ;
  assign n32056 = x74 | n31596 ;
  assign n32057 = x74 &  n31596 ;
  assign n32058 = ( n32056 & ~n32057 ) | ( n32056 & 1'b0 ) | ( ~n32057 & 1'b0 ) ;
  assign n32070 = ( n31668 & n31718 ) | ( n31668 & n32058 ) | ( n31718 & n32058 ) ;
  assign n32069 = n31668 | n32058 ;
  assign n32071 = ( n32068 & ~n32070 ) | ( n32068 & n32069 ) | ( ~n32070 & n32069 ) ;
  assign n32075 = n31604 &  n31717 ;
  assign n32076 = n31716 &  n32075 ;
  assign n32064 = x73 | n31604 ;
  assign n32065 = x73 &  n31604 ;
  assign n32066 = ( n32064 & ~n32065 ) | ( n32064 & 1'b0 ) | ( ~n32065 & 1'b0 ) ;
  assign n32078 = ( n31667 & n31718 ) | ( n31667 & n32066 ) | ( n31718 & n32066 ) ;
  assign n32077 = n31667 | n32066 ;
  assign n32079 = ( n32076 & ~n32078 ) | ( n32076 & n32077 ) | ( ~n32078 & n32077 ) ;
  assign n32083 = n31612 &  n31717 ;
  assign n32084 = n31716 &  n32083 ;
  assign n32072 = x72 | n31612 ;
  assign n32073 = x72 &  n31612 ;
  assign n32074 = ( n32072 & ~n32073 ) | ( n32072 & 1'b0 ) | ( ~n32073 & 1'b0 ) ;
  assign n32086 = ( n31666 & n31718 ) | ( n31666 & n32074 ) | ( n31718 & n32074 ) ;
  assign n32085 = n31666 | n32074 ;
  assign n32087 = ( n32084 & ~n32086 ) | ( n32084 & n32085 ) | ( ~n32086 & n32085 ) ;
  assign n32091 = n31620 &  n31717 ;
  assign n32092 = n31716 &  n32091 ;
  assign n32080 = x71 | n31620 ;
  assign n32081 = x71 &  n31620 ;
  assign n32082 = ( n32080 & ~n32081 ) | ( n32080 & 1'b0 ) | ( ~n32081 & 1'b0 ) ;
  assign n32094 = ( n31665 & n31718 ) | ( n31665 & n32082 ) | ( n31718 & n32082 ) ;
  assign n32093 = n31665 | n32082 ;
  assign n32095 = ( n32092 & ~n32094 ) | ( n32092 & n32093 ) | ( ~n32094 & n32093 ) ;
  assign n32099 = n31628 &  n31717 ;
  assign n32100 = n31716 &  n32099 ;
  assign n32088 = x70 | n31628 ;
  assign n32089 = x70 &  n31628 ;
  assign n32090 = ( n32088 & ~n32089 ) | ( n32088 & 1'b0 ) | ( ~n32089 & 1'b0 ) ;
  assign n32102 = ( n31664 & n31718 ) | ( n31664 & n32090 ) | ( n31718 & n32090 ) ;
  assign n32101 = n31664 | n32090 ;
  assign n32103 = ( n32100 & ~n32102 ) | ( n32100 & n32101 ) | ( ~n32102 & n32101 ) ;
  assign n32107 = n31636 &  n31717 ;
  assign n32108 = n31716 &  n32107 ;
  assign n32096 = x69 | n31636 ;
  assign n32097 = x69 &  n31636 ;
  assign n32098 = ( n32096 & ~n32097 ) | ( n32096 & 1'b0 ) | ( ~n32097 & 1'b0 ) ;
  assign n32110 = ( n31663 & n31718 ) | ( n31663 & n32098 ) | ( n31718 & n32098 ) ;
  assign n32109 = n31663 | n32098 ;
  assign n32111 = ( n32108 & ~n32110 ) | ( n32108 & n32109 ) | ( ~n32110 & n32109 ) ;
  assign n32115 = n31644 &  n31717 ;
  assign n32116 = n31716 &  n32115 ;
  assign n32104 = x68 | n31644 ;
  assign n32105 = x68 &  n31644 ;
  assign n32106 = ( n32104 & ~n32105 ) | ( n32104 & 1'b0 ) | ( ~n32105 & 1'b0 ) ;
  assign n32118 = ( n31662 & n31718 ) | ( n31662 & n32106 ) | ( n31718 & n32106 ) ;
  assign n32117 = n31662 | n32106 ;
  assign n32119 = ( n32116 & ~n32118 ) | ( n32116 & n32117 ) | ( ~n32118 & n32117 ) ;
  assign n32123 = n31649 &  n31717 ;
  assign n32124 = n31716 &  n32123 ;
  assign n32112 = x67 | n31649 ;
  assign n32113 = x67 &  n31649 ;
  assign n32114 = ( n32112 & ~n32113 ) | ( n32112 & 1'b0 ) | ( ~n32113 & 1'b0 ) ;
  assign n32126 = ( n31661 & n31718 ) | ( n31661 & n32114 ) | ( n31718 & n32114 ) ;
  assign n32125 = n31661 | n32114 ;
  assign n32127 = ( n32124 & ~n32126 ) | ( n32124 & n32125 ) | ( ~n32126 & n32125 ) ;
  assign n32128 = n31655 &  n31717 ;
  assign n32129 = n31716 &  n32128 ;
  assign n32120 = x66 | n31655 ;
  assign n32121 = x66 &  n31655 ;
  assign n32122 = ( n32120 & ~n32121 ) | ( n32120 & 1'b0 ) | ( ~n32121 & 1'b0 ) ;
  assign n32130 = n31660 &  n32122 ;
  assign n32131 = ( n31660 & ~n31718 ) | ( n31660 & n32122 ) | ( ~n31718 & n32122 ) ;
  assign n32132 = ( n32129 & ~n32130 ) | ( n32129 & n32131 ) | ( ~n32130 & n32131 ) ;
  assign n32133 = ( x65 & ~n13294 ) | ( x65 & n31659 ) | ( ~n13294 & n31659 ) ;
  assign n32134 = ( n31660 & ~x65 ) | ( n31660 & n32133 ) | ( ~x65 & n32133 ) ;
  assign n32135 = ~n31718 & n32134 ;
  assign n32136 = n31659 &  n31717 ;
  assign n32137 = n31716 &  n32136 ;
  assign n32138 = n32135 | n32137 ;
  assign n32139 = ( x64 & ~n31718 ) | ( x64 & 1'b0 ) | ( ~n31718 & 1'b0 ) ;
  assign n32140 = ( x10 & ~n32139 ) | ( x10 & 1'b0 ) | ( ~n32139 & 1'b0 ) ;
  assign n32141 = ( n13294 & ~n31718 ) | ( n13294 & 1'b0 ) | ( ~n31718 & 1'b0 ) ;
  assign n32142 = n32140 | n32141 ;
  assign n32143 = ( x65 & ~n32142 ) | ( x65 & n13842 ) | ( ~n32142 & n13842 ) ;
  assign n32144 = ( x66 & ~n32138 ) | ( x66 & n32143 ) | ( ~n32138 & n32143 ) ;
  assign n32145 = ( x67 & ~n32132 ) | ( x67 & n32144 ) | ( ~n32132 & n32144 ) ;
  assign n32146 = ( x68 & ~n32127 ) | ( x68 & n32145 ) | ( ~n32127 & n32145 ) ;
  assign n32147 = ( x69 & ~n32119 ) | ( x69 & n32146 ) | ( ~n32119 & n32146 ) ;
  assign n32148 = ( x70 & ~n32111 ) | ( x70 & n32147 ) | ( ~n32111 & n32147 ) ;
  assign n32149 = ( x71 & ~n32103 ) | ( x71 & n32148 ) | ( ~n32103 & n32148 ) ;
  assign n32150 = ( x72 & ~n32095 ) | ( x72 & n32149 ) | ( ~n32095 & n32149 ) ;
  assign n32151 = ( x73 & ~n32087 ) | ( x73 & n32150 ) | ( ~n32087 & n32150 ) ;
  assign n32152 = ( x74 & ~n32079 ) | ( x74 & n32151 ) | ( ~n32079 & n32151 ) ;
  assign n32153 = ( x75 & ~n32071 ) | ( x75 & n32152 ) | ( ~n32071 & n32152 ) ;
  assign n32154 = ( x76 & ~n32063 ) | ( x76 & n32153 ) | ( ~n32063 & n32153 ) ;
  assign n32155 = ( x77 & ~n32055 ) | ( x77 & n32154 ) | ( ~n32055 & n32154 ) ;
  assign n32156 = ( x78 & ~n32047 ) | ( x78 & n32155 ) | ( ~n32047 & n32155 ) ;
  assign n32157 = ( x79 & ~n32039 ) | ( x79 & n32156 ) | ( ~n32039 & n32156 ) ;
  assign n32158 = ( x80 & ~n32031 ) | ( x80 & n32157 ) | ( ~n32031 & n32157 ) ;
  assign n32159 = ( x81 & ~n32023 ) | ( x81 & n32158 ) | ( ~n32023 & n32158 ) ;
  assign n32160 = ( x82 & ~n32015 ) | ( x82 & n32159 ) | ( ~n32015 & n32159 ) ;
  assign n32161 = ( x83 & ~n32007 ) | ( x83 & n32160 ) | ( ~n32007 & n32160 ) ;
  assign n32162 = ( x84 & ~n31999 ) | ( x84 & n32161 ) | ( ~n31999 & n32161 ) ;
  assign n32163 = ( x85 & ~n31991 ) | ( x85 & n32162 ) | ( ~n31991 & n32162 ) ;
  assign n32164 = ( x86 & ~n31983 ) | ( x86 & n32163 ) | ( ~n31983 & n32163 ) ;
  assign n32165 = ( x87 & ~n31975 ) | ( x87 & n32164 ) | ( ~n31975 & n32164 ) ;
  assign n32166 = ( x88 & ~n31967 ) | ( x88 & n32165 ) | ( ~n31967 & n32165 ) ;
  assign n32167 = ( x89 & ~n31959 ) | ( x89 & n32166 ) | ( ~n31959 & n32166 ) ;
  assign n32168 = ( x90 & ~n31951 ) | ( x90 & n32167 ) | ( ~n31951 & n32167 ) ;
  assign n32169 = ( x91 & ~n31943 ) | ( x91 & n32168 ) | ( ~n31943 & n32168 ) ;
  assign n32170 = ( x92 & ~n31935 ) | ( x92 & n32169 ) | ( ~n31935 & n32169 ) ;
  assign n32171 = ( x93 & ~n31927 ) | ( x93 & n32170 ) | ( ~n31927 & n32170 ) ;
  assign n32172 = ( x94 & ~n31919 ) | ( x94 & n32171 ) | ( ~n31919 & n32171 ) ;
  assign n32173 = ( x95 & ~n31911 ) | ( x95 & n32172 ) | ( ~n31911 & n32172 ) ;
  assign n32174 = ( x96 & ~n31903 ) | ( x96 & n32173 ) | ( ~n31903 & n32173 ) ;
  assign n32175 = ( x97 & ~n31895 ) | ( x97 & n32174 ) | ( ~n31895 & n32174 ) ;
  assign n32176 = ( x98 & ~n31887 ) | ( x98 & n32175 ) | ( ~n31887 & n32175 ) ;
  assign n32177 = ( x99 & ~n31879 ) | ( x99 & n32176 ) | ( ~n31879 & n32176 ) ;
  assign n32178 = ( x100 & ~n31871 ) | ( x100 & n32177 ) | ( ~n31871 & n32177 ) ;
  assign n32179 = ( x101 & ~n31863 ) | ( x101 & n32178 ) | ( ~n31863 & n32178 ) ;
  assign n32180 = ( x102 & ~n31855 ) | ( x102 & n32179 ) | ( ~n31855 & n32179 ) ;
  assign n32181 = ( x103 & ~n31847 ) | ( x103 & n32180 ) | ( ~n31847 & n32180 ) ;
  assign n32182 = ( x104 & ~n31839 ) | ( x104 & n32181 ) | ( ~n31839 & n32181 ) ;
  assign n32183 = ( x105 & ~n31831 ) | ( x105 & n32182 ) | ( ~n31831 & n32182 ) ;
  assign n32184 = ( x106 & ~n31823 ) | ( x106 & n32183 ) | ( ~n31823 & n32183 ) ;
  assign n32185 = ( x107 & ~n31815 ) | ( x107 & n32184 ) | ( ~n31815 & n32184 ) ;
  assign n32186 = ( x108 & ~n31807 ) | ( x108 & n32185 ) | ( ~n31807 & n32185 ) ;
  assign n32187 = ( x109 & ~n31799 ) | ( x109 & n32186 ) | ( ~n31799 & n32186 ) ;
  assign n32188 = ( x110 & ~n31791 ) | ( x110 & n32187 ) | ( ~n31791 & n32187 ) ;
  assign n32189 = ( x111 & ~n31783 ) | ( x111 & n32188 ) | ( ~n31783 & n32188 ) ;
  assign n32190 = ( x112 & ~n31775 ) | ( x112 & n32189 ) | ( ~n31775 & n32189 ) ;
  assign n32191 = ( x113 & ~n31767 ) | ( x113 & n32190 ) | ( ~n31767 & n32190 ) ;
  assign n32192 = ( x114 & ~n31759 ) | ( x114 & n32191 ) | ( ~n31759 & n32191 ) ;
  assign n32193 = ( x115 & ~n31751 ) | ( x115 & n32192 ) | ( ~n31751 & n32192 ) ;
  assign n32194 = ( x116 & ~n31743 ) | ( x116 & n32193 ) | ( ~n31743 & n32193 ) ;
  assign n32195 = ( x117 & ~n31735 ) | ( x117 & n32194 ) | ( ~n31735 & n32194 ) ;
  assign n32196 = ( x118 & ~n31727 ) | ( x118 & n32195 ) | ( ~n31727 & n32195 ) ;
  assign n32197 = n13898 | n32196 ;
  assign n32207 = n31735 &  n32197 ;
  assign n32199 = x117 | n31735 ;
  assign n32200 = x117 &  n31735 ;
  assign n32201 = ( n32199 & ~n32200 ) | ( n32199 & 1'b0 ) | ( ~n32200 & 1'b0 ) ;
  assign n32211 = ( n13898 & n32194 ) | ( n13898 & n32201 ) | ( n32194 & n32201 ) ;
  assign n32212 = ( n32194 & ~n32196 ) | ( n32194 & n32201 ) | ( ~n32196 & n32201 ) ;
  assign n32213 = ~n32211 & n32212 ;
  assign n32214 = n32207 | n32213 ;
  assign n32215 = n31743 &  n32197 ;
  assign n32208 = x116 | n31743 ;
  assign n32209 = x116 &  n31743 ;
  assign n32210 = ( n32208 & ~n32209 ) | ( n32208 & 1'b0 ) | ( ~n32209 & 1'b0 ) ;
  assign n32219 = ( n13898 & n32193 ) | ( n13898 & n32210 ) | ( n32193 & n32210 ) ;
  assign n32220 = ( n32193 & ~n32196 ) | ( n32193 & n32210 ) | ( ~n32196 & n32210 ) ;
  assign n32221 = ~n32219 & n32220 ;
  assign n32222 = n32215 | n32221 ;
  assign n32223 = n31751 &  n32197 ;
  assign n32216 = x115 | n31751 ;
  assign n32217 = x115 &  n31751 ;
  assign n32218 = ( n32216 & ~n32217 ) | ( n32216 & 1'b0 ) | ( ~n32217 & 1'b0 ) ;
  assign n32227 = ( n13898 & n32192 ) | ( n13898 & n32218 ) | ( n32192 & n32218 ) ;
  assign n32228 = ( n32192 & ~n32196 ) | ( n32192 & n32218 ) | ( ~n32196 & n32218 ) ;
  assign n32229 = ~n32227 & n32228 ;
  assign n32230 = n32223 | n32229 ;
  assign n32231 = n31759 &  n32197 ;
  assign n32224 = x114 | n31759 ;
  assign n32225 = x114 &  n31759 ;
  assign n32226 = ( n32224 & ~n32225 ) | ( n32224 & 1'b0 ) | ( ~n32225 & 1'b0 ) ;
  assign n32235 = ( n13898 & n32191 ) | ( n13898 & n32226 ) | ( n32191 & n32226 ) ;
  assign n32236 = ( n32191 & ~n32196 ) | ( n32191 & n32226 ) | ( ~n32196 & n32226 ) ;
  assign n32237 = ~n32235 & n32236 ;
  assign n32238 = n32231 | n32237 ;
  assign n32239 = n31767 &  n32197 ;
  assign n32232 = x113 | n31767 ;
  assign n32233 = x113 &  n31767 ;
  assign n32234 = ( n32232 & ~n32233 ) | ( n32232 & 1'b0 ) | ( ~n32233 & 1'b0 ) ;
  assign n32243 = ( n13898 & n32190 ) | ( n13898 & n32234 ) | ( n32190 & n32234 ) ;
  assign n32244 = ( n32190 & ~n32196 ) | ( n32190 & n32234 ) | ( ~n32196 & n32234 ) ;
  assign n32245 = ~n32243 & n32244 ;
  assign n32246 = n32239 | n32245 ;
  assign n32247 = n31775 &  n32197 ;
  assign n32240 = x112 | n31775 ;
  assign n32241 = x112 &  n31775 ;
  assign n32242 = ( n32240 & ~n32241 ) | ( n32240 & 1'b0 ) | ( ~n32241 & 1'b0 ) ;
  assign n32251 = ( n13898 & n32189 ) | ( n13898 & n32242 ) | ( n32189 & n32242 ) ;
  assign n32252 = ( n32189 & ~n32196 ) | ( n32189 & n32242 ) | ( ~n32196 & n32242 ) ;
  assign n32253 = ~n32251 & n32252 ;
  assign n32254 = n32247 | n32253 ;
  assign n32255 = n31783 &  n32197 ;
  assign n32248 = x111 | n31783 ;
  assign n32249 = x111 &  n31783 ;
  assign n32250 = ( n32248 & ~n32249 ) | ( n32248 & 1'b0 ) | ( ~n32249 & 1'b0 ) ;
  assign n32259 = ( n13898 & n32188 ) | ( n13898 & n32250 ) | ( n32188 & n32250 ) ;
  assign n32260 = ( n32188 & ~n32196 ) | ( n32188 & n32250 ) | ( ~n32196 & n32250 ) ;
  assign n32261 = ~n32259 & n32260 ;
  assign n32262 = n32255 | n32261 ;
  assign n32263 = n31791 &  n32197 ;
  assign n32256 = x110 | n31791 ;
  assign n32257 = x110 &  n31791 ;
  assign n32258 = ( n32256 & ~n32257 ) | ( n32256 & 1'b0 ) | ( ~n32257 & 1'b0 ) ;
  assign n32267 = ( n13898 & n32187 ) | ( n13898 & n32258 ) | ( n32187 & n32258 ) ;
  assign n32268 = ( n32187 & ~n32196 ) | ( n32187 & n32258 ) | ( ~n32196 & n32258 ) ;
  assign n32269 = ~n32267 & n32268 ;
  assign n32270 = n32263 | n32269 ;
  assign n32271 = n31799 &  n32197 ;
  assign n32264 = x109 | n31799 ;
  assign n32265 = x109 &  n31799 ;
  assign n32266 = ( n32264 & ~n32265 ) | ( n32264 & 1'b0 ) | ( ~n32265 & 1'b0 ) ;
  assign n32275 = ( n13898 & n32186 ) | ( n13898 & n32266 ) | ( n32186 & n32266 ) ;
  assign n32276 = ( n32186 & ~n32196 ) | ( n32186 & n32266 ) | ( ~n32196 & n32266 ) ;
  assign n32277 = ~n32275 & n32276 ;
  assign n32278 = n32271 | n32277 ;
  assign n32279 = n31807 &  n32197 ;
  assign n32272 = x108 | n31807 ;
  assign n32273 = x108 &  n31807 ;
  assign n32274 = ( n32272 & ~n32273 ) | ( n32272 & 1'b0 ) | ( ~n32273 & 1'b0 ) ;
  assign n32283 = ( n13898 & n32185 ) | ( n13898 & n32274 ) | ( n32185 & n32274 ) ;
  assign n32284 = ( n32185 & ~n32196 ) | ( n32185 & n32274 ) | ( ~n32196 & n32274 ) ;
  assign n32285 = ~n32283 & n32284 ;
  assign n32286 = n32279 | n32285 ;
  assign n32287 = n31815 &  n32197 ;
  assign n32280 = x107 | n31815 ;
  assign n32281 = x107 &  n31815 ;
  assign n32282 = ( n32280 & ~n32281 ) | ( n32280 & 1'b0 ) | ( ~n32281 & 1'b0 ) ;
  assign n32291 = ( n13898 & n32184 ) | ( n13898 & n32282 ) | ( n32184 & n32282 ) ;
  assign n32292 = ( n32184 & ~n32196 ) | ( n32184 & n32282 ) | ( ~n32196 & n32282 ) ;
  assign n32293 = ~n32291 & n32292 ;
  assign n32294 = n32287 | n32293 ;
  assign n32295 = n31823 &  n32197 ;
  assign n32288 = x106 | n31823 ;
  assign n32289 = x106 &  n31823 ;
  assign n32290 = ( n32288 & ~n32289 ) | ( n32288 & 1'b0 ) | ( ~n32289 & 1'b0 ) ;
  assign n32299 = ( n13898 & n32183 ) | ( n13898 & n32290 ) | ( n32183 & n32290 ) ;
  assign n32300 = ( n32183 & ~n32196 ) | ( n32183 & n32290 ) | ( ~n32196 & n32290 ) ;
  assign n32301 = ~n32299 & n32300 ;
  assign n32302 = n32295 | n32301 ;
  assign n32303 = n31831 &  n32197 ;
  assign n32296 = x105 | n31831 ;
  assign n32297 = x105 &  n31831 ;
  assign n32298 = ( n32296 & ~n32297 ) | ( n32296 & 1'b0 ) | ( ~n32297 & 1'b0 ) ;
  assign n32307 = ( n13898 & n32182 ) | ( n13898 & n32298 ) | ( n32182 & n32298 ) ;
  assign n32308 = ( n32182 & ~n32196 ) | ( n32182 & n32298 ) | ( ~n32196 & n32298 ) ;
  assign n32309 = ~n32307 & n32308 ;
  assign n32310 = n32303 | n32309 ;
  assign n32311 = n31839 &  n32197 ;
  assign n32304 = x104 | n31839 ;
  assign n32305 = x104 &  n31839 ;
  assign n32306 = ( n32304 & ~n32305 ) | ( n32304 & 1'b0 ) | ( ~n32305 & 1'b0 ) ;
  assign n32315 = ( n13898 & n32181 ) | ( n13898 & n32306 ) | ( n32181 & n32306 ) ;
  assign n32316 = ( n32181 & ~n32196 ) | ( n32181 & n32306 ) | ( ~n32196 & n32306 ) ;
  assign n32317 = ~n32315 & n32316 ;
  assign n32318 = n32311 | n32317 ;
  assign n32319 = n31847 &  n32197 ;
  assign n32312 = x103 | n31847 ;
  assign n32313 = x103 &  n31847 ;
  assign n32314 = ( n32312 & ~n32313 ) | ( n32312 & 1'b0 ) | ( ~n32313 & 1'b0 ) ;
  assign n32323 = ( n13898 & n32180 ) | ( n13898 & n32314 ) | ( n32180 & n32314 ) ;
  assign n32324 = ( n32180 & ~n32196 ) | ( n32180 & n32314 ) | ( ~n32196 & n32314 ) ;
  assign n32325 = ~n32323 & n32324 ;
  assign n32326 = n32319 | n32325 ;
  assign n32327 = n31855 &  n32197 ;
  assign n32320 = x102 | n31855 ;
  assign n32321 = x102 &  n31855 ;
  assign n32322 = ( n32320 & ~n32321 ) | ( n32320 & 1'b0 ) | ( ~n32321 & 1'b0 ) ;
  assign n32331 = ( n13898 & n32179 ) | ( n13898 & n32322 ) | ( n32179 & n32322 ) ;
  assign n32332 = ( n32179 & ~n32196 ) | ( n32179 & n32322 ) | ( ~n32196 & n32322 ) ;
  assign n32333 = ~n32331 & n32332 ;
  assign n32334 = n32327 | n32333 ;
  assign n32335 = n31863 &  n32197 ;
  assign n32328 = x101 | n31863 ;
  assign n32329 = x101 &  n31863 ;
  assign n32330 = ( n32328 & ~n32329 ) | ( n32328 & 1'b0 ) | ( ~n32329 & 1'b0 ) ;
  assign n32339 = ( n13898 & n32178 ) | ( n13898 & n32330 ) | ( n32178 & n32330 ) ;
  assign n32340 = ( n32178 & ~n32196 ) | ( n32178 & n32330 ) | ( ~n32196 & n32330 ) ;
  assign n32341 = ~n32339 & n32340 ;
  assign n32342 = n32335 | n32341 ;
  assign n32343 = n31871 &  n32197 ;
  assign n32336 = x100 | n31871 ;
  assign n32337 = x100 &  n31871 ;
  assign n32338 = ( n32336 & ~n32337 ) | ( n32336 & 1'b0 ) | ( ~n32337 & 1'b0 ) ;
  assign n32347 = ( n13898 & n32177 ) | ( n13898 & n32338 ) | ( n32177 & n32338 ) ;
  assign n32348 = ( n32177 & ~n32196 ) | ( n32177 & n32338 ) | ( ~n32196 & n32338 ) ;
  assign n32349 = ~n32347 & n32348 ;
  assign n32350 = n32343 | n32349 ;
  assign n32351 = n31879 &  n32197 ;
  assign n32344 = x99 | n31879 ;
  assign n32345 = x99 &  n31879 ;
  assign n32346 = ( n32344 & ~n32345 ) | ( n32344 & 1'b0 ) | ( ~n32345 & 1'b0 ) ;
  assign n32355 = ( n13898 & n32176 ) | ( n13898 & n32346 ) | ( n32176 & n32346 ) ;
  assign n32356 = ( n32176 & ~n32196 ) | ( n32176 & n32346 ) | ( ~n32196 & n32346 ) ;
  assign n32357 = ~n32355 & n32356 ;
  assign n32358 = n32351 | n32357 ;
  assign n32359 = n31887 &  n32197 ;
  assign n32352 = x98 | n31887 ;
  assign n32353 = x98 &  n31887 ;
  assign n32354 = ( n32352 & ~n32353 ) | ( n32352 & 1'b0 ) | ( ~n32353 & 1'b0 ) ;
  assign n32363 = ( n13898 & n32175 ) | ( n13898 & n32354 ) | ( n32175 & n32354 ) ;
  assign n32364 = ( n32175 & ~n32196 ) | ( n32175 & n32354 ) | ( ~n32196 & n32354 ) ;
  assign n32365 = ~n32363 & n32364 ;
  assign n32366 = n32359 | n32365 ;
  assign n32367 = n31895 &  n32197 ;
  assign n32360 = x97 | n31895 ;
  assign n32361 = x97 &  n31895 ;
  assign n32362 = ( n32360 & ~n32361 ) | ( n32360 & 1'b0 ) | ( ~n32361 & 1'b0 ) ;
  assign n32371 = ( n13898 & n32174 ) | ( n13898 & n32362 ) | ( n32174 & n32362 ) ;
  assign n32372 = ( n32174 & ~n32196 ) | ( n32174 & n32362 ) | ( ~n32196 & n32362 ) ;
  assign n32373 = ~n32371 & n32372 ;
  assign n32374 = n32367 | n32373 ;
  assign n32375 = n31903 &  n32197 ;
  assign n32368 = x96 | n31903 ;
  assign n32369 = x96 &  n31903 ;
  assign n32370 = ( n32368 & ~n32369 ) | ( n32368 & 1'b0 ) | ( ~n32369 & 1'b0 ) ;
  assign n32379 = ( n13898 & n32173 ) | ( n13898 & n32370 ) | ( n32173 & n32370 ) ;
  assign n32380 = ( n32173 & ~n32196 ) | ( n32173 & n32370 ) | ( ~n32196 & n32370 ) ;
  assign n32381 = ~n32379 & n32380 ;
  assign n32382 = n32375 | n32381 ;
  assign n32383 = n31911 &  n32197 ;
  assign n32376 = x95 | n31911 ;
  assign n32377 = x95 &  n31911 ;
  assign n32378 = ( n32376 & ~n32377 ) | ( n32376 & 1'b0 ) | ( ~n32377 & 1'b0 ) ;
  assign n32387 = ( n13898 & n32172 ) | ( n13898 & n32378 ) | ( n32172 & n32378 ) ;
  assign n32388 = ( n32172 & ~n32196 ) | ( n32172 & n32378 ) | ( ~n32196 & n32378 ) ;
  assign n32389 = ~n32387 & n32388 ;
  assign n32390 = n32383 | n32389 ;
  assign n32391 = n31919 &  n32197 ;
  assign n32384 = x94 | n31919 ;
  assign n32385 = x94 &  n31919 ;
  assign n32386 = ( n32384 & ~n32385 ) | ( n32384 & 1'b0 ) | ( ~n32385 & 1'b0 ) ;
  assign n32395 = ( n13898 & n32171 ) | ( n13898 & n32386 ) | ( n32171 & n32386 ) ;
  assign n32396 = ( n32171 & ~n32196 ) | ( n32171 & n32386 ) | ( ~n32196 & n32386 ) ;
  assign n32397 = ~n32395 & n32396 ;
  assign n32398 = n32391 | n32397 ;
  assign n32399 = n31927 &  n32197 ;
  assign n32392 = x93 | n31927 ;
  assign n32393 = x93 &  n31927 ;
  assign n32394 = ( n32392 & ~n32393 ) | ( n32392 & 1'b0 ) | ( ~n32393 & 1'b0 ) ;
  assign n32403 = ( n13898 & n32170 ) | ( n13898 & n32394 ) | ( n32170 & n32394 ) ;
  assign n32404 = ( n32170 & ~n32196 ) | ( n32170 & n32394 ) | ( ~n32196 & n32394 ) ;
  assign n32405 = ~n32403 & n32404 ;
  assign n32406 = n32399 | n32405 ;
  assign n32407 = n31935 &  n32197 ;
  assign n32400 = x92 | n31935 ;
  assign n32401 = x92 &  n31935 ;
  assign n32402 = ( n32400 & ~n32401 ) | ( n32400 & 1'b0 ) | ( ~n32401 & 1'b0 ) ;
  assign n32411 = ( n13898 & n32169 ) | ( n13898 & n32402 ) | ( n32169 & n32402 ) ;
  assign n32412 = ( n32169 & ~n32196 ) | ( n32169 & n32402 ) | ( ~n32196 & n32402 ) ;
  assign n32413 = ~n32411 & n32412 ;
  assign n32414 = n32407 | n32413 ;
  assign n32415 = n31943 &  n32197 ;
  assign n32408 = x91 | n31943 ;
  assign n32409 = x91 &  n31943 ;
  assign n32410 = ( n32408 & ~n32409 ) | ( n32408 & 1'b0 ) | ( ~n32409 & 1'b0 ) ;
  assign n32419 = ( n13898 & n32168 ) | ( n13898 & n32410 ) | ( n32168 & n32410 ) ;
  assign n32420 = ( n32168 & ~n32196 ) | ( n32168 & n32410 ) | ( ~n32196 & n32410 ) ;
  assign n32421 = ~n32419 & n32420 ;
  assign n32422 = n32415 | n32421 ;
  assign n32423 = n31951 &  n32197 ;
  assign n32416 = x90 | n31951 ;
  assign n32417 = x90 &  n31951 ;
  assign n32418 = ( n32416 & ~n32417 ) | ( n32416 & 1'b0 ) | ( ~n32417 & 1'b0 ) ;
  assign n32427 = ( n13898 & n32167 ) | ( n13898 & n32418 ) | ( n32167 & n32418 ) ;
  assign n32428 = ( n32167 & ~n32196 ) | ( n32167 & n32418 ) | ( ~n32196 & n32418 ) ;
  assign n32429 = ~n32427 & n32428 ;
  assign n32430 = n32423 | n32429 ;
  assign n32431 = n31959 &  n32197 ;
  assign n32424 = x89 | n31959 ;
  assign n32425 = x89 &  n31959 ;
  assign n32426 = ( n32424 & ~n32425 ) | ( n32424 & 1'b0 ) | ( ~n32425 & 1'b0 ) ;
  assign n32435 = ( n13898 & n32166 ) | ( n13898 & n32426 ) | ( n32166 & n32426 ) ;
  assign n32436 = ( n32166 & ~n32196 ) | ( n32166 & n32426 ) | ( ~n32196 & n32426 ) ;
  assign n32437 = ~n32435 & n32436 ;
  assign n32438 = n32431 | n32437 ;
  assign n32439 = n31967 &  n32197 ;
  assign n32432 = x88 | n31967 ;
  assign n32433 = x88 &  n31967 ;
  assign n32434 = ( n32432 & ~n32433 ) | ( n32432 & 1'b0 ) | ( ~n32433 & 1'b0 ) ;
  assign n32443 = ( n13898 & n32165 ) | ( n13898 & n32434 ) | ( n32165 & n32434 ) ;
  assign n32444 = ( n32165 & ~n32196 ) | ( n32165 & n32434 ) | ( ~n32196 & n32434 ) ;
  assign n32445 = ~n32443 & n32444 ;
  assign n32446 = n32439 | n32445 ;
  assign n32447 = n31975 &  n32197 ;
  assign n32440 = x87 | n31975 ;
  assign n32441 = x87 &  n31975 ;
  assign n32442 = ( n32440 & ~n32441 ) | ( n32440 & 1'b0 ) | ( ~n32441 & 1'b0 ) ;
  assign n32451 = ( n13898 & n32164 ) | ( n13898 & n32442 ) | ( n32164 & n32442 ) ;
  assign n32452 = ( n32164 & ~n32196 ) | ( n32164 & n32442 ) | ( ~n32196 & n32442 ) ;
  assign n32453 = ~n32451 & n32452 ;
  assign n32454 = n32447 | n32453 ;
  assign n32455 = n31983 &  n32197 ;
  assign n32448 = x86 | n31983 ;
  assign n32449 = x86 &  n31983 ;
  assign n32450 = ( n32448 & ~n32449 ) | ( n32448 & 1'b0 ) | ( ~n32449 & 1'b0 ) ;
  assign n32459 = ( n13898 & n32163 ) | ( n13898 & n32450 ) | ( n32163 & n32450 ) ;
  assign n32460 = ( n32163 & ~n32196 ) | ( n32163 & n32450 ) | ( ~n32196 & n32450 ) ;
  assign n32461 = ~n32459 & n32460 ;
  assign n32462 = n32455 | n32461 ;
  assign n32463 = n31991 &  n32197 ;
  assign n32456 = x85 | n31991 ;
  assign n32457 = x85 &  n31991 ;
  assign n32458 = ( n32456 & ~n32457 ) | ( n32456 & 1'b0 ) | ( ~n32457 & 1'b0 ) ;
  assign n32467 = ( n13898 & n32162 ) | ( n13898 & n32458 ) | ( n32162 & n32458 ) ;
  assign n32468 = ( n32162 & ~n32196 ) | ( n32162 & n32458 ) | ( ~n32196 & n32458 ) ;
  assign n32469 = ~n32467 & n32468 ;
  assign n32470 = n32463 | n32469 ;
  assign n32471 = n31999 &  n32197 ;
  assign n32464 = x84 | n31999 ;
  assign n32465 = x84 &  n31999 ;
  assign n32466 = ( n32464 & ~n32465 ) | ( n32464 & 1'b0 ) | ( ~n32465 & 1'b0 ) ;
  assign n32475 = ( n13898 & n32161 ) | ( n13898 & n32466 ) | ( n32161 & n32466 ) ;
  assign n32476 = ( n32161 & ~n32196 ) | ( n32161 & n32466 ) | ( ~n32196 & n32466 ) ;
  assign n32477 = ~n32475 & n32476 ;
  assign n32478 = n32471 | n32477 ;
  assign n32479 = n32007 &  n32197 ;
  assign n32472 = x83 | n32007 ;
  assign n32473 = x83 &  n32007 ;
  assign n32474 = ( n32472 & ~n32473 ) | ( n32472 & 1'b0 ) | ( ~n32473 & 1'b0 ) ;
  assign n32483 = ( n13898 & n32160 ) | ( n13898 & n32474 ) | ( n32160 & n32474 ) ;
  assign n32484 = ( n32160 & ~n32196 ) | ( n32160 & n32474 ) | ( ~n32196 & n32474 ) ;
  assign n32485 = ~n32483 & n32484 ;
  assign n32486 = n32479 | n32485 ;
  assign n32487 = n32015 &  n32197 ;
  assign n32480 = x82 | n32015 ;
  assign n32481 = x82 &  n32015 ;
  assign n32482 = ( n32480 & ~n32481 ) | ( n32480 & 1'b0 ) | ( ~n32481 & 1'b0 ) ;
  assign n32491 = ( n13898 & n32159 ) | ( n13898 & n32482 ) | ( n32159 & n32482 ) ;
  assign n32492 = ( n32159 & ~n32196 ) | ( n32159 & n32482 ) | ( ~n32196 & n32482 ) ;
  assign n32493 = ~n32491 & n32492 ;
  assign n32494 = n32487 | n32493 ;
  assign n32495 = n32023 &  n32197 ;
  assign n32488 = x81 | n32023 ;
  assign n32489 = x81 &  n32023 ;
  assign n32490 = ( n32488 & ~n32489 ) | ( n32488 & 1'b0 ) | ( ~n32489 & 1'b0 ) ;
  assign n32499 = ( n13898 & n32158 ) | ( n13898 & n32490 ) | ( n32158 & n32490 ) ;
  assign n32500 = ( n32158 & ~n32196 ) | ( n32158 & n32490 ) | ( ~n32196 & n32490 ) ;
  assign n32501 = ~n32499 & n32500 ;
  assign n32502 = n32495 | n32501 ;
  assign n32503 = n32031 &  n32197 ;
  assign n32496 = x80 | n32031 ;
  assign n32497 = x80 &  n32031 ;
  assign n32498 = ( n32496 & ~n32497 ) | ( n32496 & 1'b0 ) | ( ~n32497 & 1'b0 ) ;
  assign n32507 = ( n13898 & n32157 ) | ( n13898 & n32498 ) | ( n32157 & n32498 ) ;
  assign n32508 = ( n32157 & ~n32196 ) | ( n32157 & n32498 ) | ( ~n32196 & n32498 ) ;
  assign n32509 = ~n32507 & n32508 ;
  assign n32510 = n32503 | n32509 ;
  assign n32511 = n32039 &  n32197 ;
  assign n32504 = x79 | n32039 ;
  assign n32505 = x79 &  n32039 ;
  assign n32506 = ( n32504 & ~n32505 ) | ( n32504 & 1'b0 ) | ( ~n32505 & 1'b0 ) ;
  assign n32515 = ( n13898 & n32156 ) | ( n13898 & n32506 ) | ( n32156 & n32506 ) ;
  assign n32516 = ( n32156 & ~n32196 ) | ( n32156 & n32506 ) | ( ~n32196 & n32506 ) ;
  assign n32517 = ~n32515 & n32516 ;
  assign n32518 = n32511 | n32517 ;
  assign n32519 = n32047 &  n32197 ;
  assign n32512 = x78 | n32047 ;
  assign n32513 = x78 &  n32047 ;
  assign n32514 = ( n32512 & ~n32513 ) | ( n32512 & 1'b0 ) | ( ~n32513 & 1'b0 ) ;
  assign n32523 = ( n13898 & n32155 ) | ( n13898 & n32514 ) | ( n32155 & n32514 ) ;
  assign n32524 = ( n32155 & ~n32196 ) | ( n32155 & n32514 ) | ( ~n32196 & n32514 ) ;
  assign n32525 = ~n32523 & n32524 ;
  assign n32526 = n32519 | n32525 ;
  assign n32527 = n32055 &  n32197 ;
  assign n32520 = x77 | n32055 ;
  assign n32521 = x77 &  n32055 ;
  assign n32522 = ( n32520 & ~n32521 ) | ( n32520 & 1'b0 ) | ( ~n32521 & 1'b0 ) ;
  assign n32531 = ( n13898 & n32154 ) | ( n13898 & n32522 ) | ( n32154 & n32522 ) ;
  assign n32532 = ( n32154 & ~n32196 ) | ( n32154 & n32522 ) | ( ~n32196 & n32522 ) ;
  assign n32533 = ~n32531 & n32532 ;
  assign n32534 = n32527 | n32533 ;
  assign n32535 = n32063 &  n32197 ;
  assign n32528 = x76 | n32063 ;
  assign n32529 = x76 &  n32063 ;
  assign n32530 = ( n32528 & ~n32529 ) | ( n32528 & 1'b0 ) | ( ~n32529 & 1'b0 ) ;
  assign n32539 = ( n13898 & n32153 ) | ( n13898 & n32530 ) | ( n32153 & n32530 ) ;
  assign n32540 = ( n32153 & ~n32196 ) | ( n32153 & n32530 ) | ( ~n32196 & n32530 ) ;
  assign n32541 = ~n32539 & n32540 ;
  assign n32542 = n32535 | n32541 ;
  assign n32543 = n32071 &  n32197 ;
  assign n32536 = x75 | n32071 ;
  assign n32537 = x75 &  n32071 ;
  assign n32538 = ( n32536 & ~n32537 ) | ( n32536 & 1'b0 ) | ( ~n32537 & 1'b0 ) ;
  assign n32547 = ( n13898 & n32152 ) | ( n13898 & n32538 ) | ( n32152 & n32538 ) ;
  assign n32548 = ( n32152 & ~n32196 ) | ( n32152 & n32538 ) | ( ~n32196 & n32538 ) ;
  assign n32549 = ~n32547 & n32548 ;
  assign n32550 = n32543 | n32549 ;
  assign n32551 = n32079 &  n32197 ;
  assign n32544 = x74 | n32079 ;
  assign n32545 = x74 &  n32079 ;
  assign n32546 = ( n32544 & ~n32545 ) | ( n32544 & 1'b0 ) | ( ~n32545 & 1'b0 ) ;
  assign n32555 = ( n13898 & n32151 ) | ( n13898 & n32546 ) | ( n32151 & n32546 ) ;
  assign n32556 = ( n32151 & ~n32196 ) | ( n32151 & n32546 ) | ( ~n32196 & n32546 ) ;
  assign n32557 = ~n32555 & n32556 ;
  assign n32558 = n32551 | n32557 ;
  assign n32559 = n32087 &  n32197 ;
  assign n32552 = x73 | n32087 ;
  assign n32553 = x73 &  n32087 ;
  assign n32554 = ( n32552 & ~n32553 ) | ( n32552 & 1'b0 ) | ( ~n32553 & 1'b0 ) ;
  assign n32563 = ( n13898 & n32150 ) | ( n13898 & n32554 ) | ( n32150 & n32554 ) ;
  assign n32564 = ( n32150 & ~n32196 ) | ( n32150 & n32554 ) | ( ~n32196 & n32554 ) ;
  assign n32565 = ~n32563 & n32564 ;
  assign n32566 = n32559 | n32565 ;
  assign n32567 = n32095 &  n32197 ;
  assign n32560 = x72 | n32095 ;
  assign n32561 = x72 &  n32095 ;
  assign n32562 = ( n32560 & ~n32561 ) | ( n32560 & 1'b0 ) | ( ~n32561 & 1'b0 ) ;
  assign n32571 = ( n13898 & n32149 ) | ( n13898 & n32562 ) | ( n32149 & n32562 ) ;
  assign n32572 = ( n32149 & ~n32196 ) | ( n32149 & n32562 ) | ( ~n32196 & n32562 ) ;
  assign n32573 = ~n32571 & n32572 ;
  assign n32574 = n32567 | n32573 ;
  assign n32575 = n32103 &  n32197 ;
  assign n32568 = x71 | n32103 ;
  assign n32569 = x71 &  n32103 ;
  assign n32570 = ( n32568 & ~n32569 ) | ( n32568 & 1'b0 ) | ( ~n32569 & 1'b0 ) ;
  assign n32579 = ( n13898 & n32148 ) | ( n13898 & n32570 ) | ( n32148 & n32570 ) ;
  assign n32580 = ( n32148 & ~n32196 ) | ( n32148 & n32570 ) | ( ~n32196 & n32570 ) ;
  assign n32581 = ~n32579 & n32580 ;
  assign n32582 = n32575 | n32581 ;
  assign n32583 = n32111 &  n32197 ;
  assign n32576 = x70 | n32111 ;
  assign n32577 = x70 &  n32111 ;
  assign n32578 = ( n32576 & ~n32577 ) | ( n32576 & 1'b0 ) | ( ~n32577 & 1'b0 ) ;
  assign n32587 = ( n13898 & n32147 ) | ( n13898 & n32578 ) | ( n32147 & n32578 ) ;
  assign n32588 = ( n32147 & ~n32196 ) | ( n32147 & n32578 ) | ( ~n32196 & n32578 ) ;
  assign n32589 = ~n32587 & n32588 ;
  assign n32590 = n32583 | n32589 ;
  assign n32591 = n32119 &  n32197 ;
  assign n32584 = x69 | n32119 ;
  assign n32585 = x69 &  n32119 ;
  assign n32586 = ( n32584 & ~n32585 ) | ( n32584 & 1'b0 ) | ( ~n32585 & 1'b0 ) ;
  assign n32595 = ( n13898 & n32146 ) | ( n13898 & n32586 ) | ( n32146 & n32586 ) ;
  assign n32596 = ( n32146 & ~n32196 ) | ( n32146 & n32586 ) | ( ~n32196 & n32586 ) ;
  assign n32597 = ~n32595 & n32596 ;
  assign n32598 = n32591 | n32597 ;
  assign n32599 = n32127 &  n32197 ;
  assign n32592 = x68 | n32127 ;
  assign n32593 = x68 &  n32127 ;
  assign n32594 = ( n32592 & ~n32593 ) | ( n32592 & 1'b0 ) | ( ~n32593 & 1'b0 ) ;
  assign n32603 = ( n13898 & n32145 ) | ( n13898 & n32594 ) | ( n32145 & n32594 ) ;
  assign n32604 = ( n32145 & ~n32196 ) | ( n32145 & n32594 ) | ( ~n32196 & n32594 ) ;
  assign n32605 = ~n32603 & n32604 ;
  assign n32606 = n32599 | n32605 ;
  assign n32607 = n32132 &  n32197 ;
  assign n32600 = x67 | n32132 ;
  assign n32601 = x67 &  n32132 ;
  assign n32602 = ( n32600 & ~n32601 ) | ( n32600 & 1'b0 ) | ( ~n32601 & 1'b0 ) ;
  assign n32611 = ( n13898 & n32144 ) | ( n13898 & n32602 ) | ( n32144 & n32602 ) ;
  assign n32612 = ( n32144 & ~n32196 ) | ( n32144 & n32602 ) | ( ~n32196 & n32602 ) ;
  assign n32613 = ~n32611 & n32612 ;
  assign n32614 = n32607 | n32613 ;
  assign n32615 = n32138 &  n32197 ;
  assign n32608 = x66 | n32138 ;
  assign n32609 = x66 &  n32138 ;
  assign n32610 = ( n32608 & ~n32609 ) | ( n32608 & 1'b0 ) | ( ~n32609 & 1'b0 ) ;
  assign n32616 = ( n13898 & n32143 ) | ( n13898 & n32610 ) | ( n32143 & n32610 ) ;
  assign n32617 = ( n32143 & ~n32196 ) | ( n32143 & n32610 ) | ( ~n32196 & n32610 ) ;
  assign n32618 = ~n32616 & n32617 ;
  assign n32619 = n32615 | n32618 ;
  assign n32620 = n32142 &  n32197 ;
  assign n32621 = ( x65 & ~x10 ) | ( x65 & n32139 ) | ( ~x10 & n32139 ) ;
  assign n32622 = ( x10 & ~n32139 ) | ( x10 & x65 ) | ( ~n32139 & x65 ) ;
  assign n32623 = ( n32621 & ~x65 ) | ( n32621 & n32622 ) | ( ~x65 & n32622 ) ;
  assign n32624 = ( n13842 & ~n13898 ) | ( n13842 & n32623 ) | ( ~n13898 & n32623 ) ;
  assign n32625 = ( n13842 & n32196 ) | ( n13842 & n32623 ) | ( n32196 & n32623 ) ;
  assign n32626 = ( n32624 & ~n32625 ) | ( n32624 & 1'b0 ) | ( ~n32625 & 1'b0 ) ;
  assign n32627 = n32620 | n32626 ;
  assign n32628 = ( n14280 & ~n32196 ) | ( n14280 & 1'b0 ) | ( ~n32196 & 1'b0 ) ;
  assign n32629 = ( x9 & ~n32628 ) | ( x9 & 1'b0 ) | ( ~n32628 & 1'b0 ) ;
  assign n32630 = ( n14285 & ~n32196 ) | ( n14285 & 1'b0 ) | ( ~n32196 & 1'b0 ) ;
  assign n32631 = n32629 | n32630 ;
  assign n32632 = ( x65 & ~n32631 ) | ( x65 & n14288 ) | ( ~n32631 & n14288 ) ;
  assign n32633 = ( x66 & ~n32627 ) | ( x66 & n32632 ) | ( ~n32627 & n32632 ) ;
  assign n32634 = ( x67 & ~n32619 ) | ( x67 & n32633 ) | ( ~n32619 & n32633 ) ;
  assign n32635 = ( x68 & ~n32614 ) | ( x68 & n32634 ) | ( ~n32614 & n32634 ) ;
  assign n32636 = ( x69 & ~n32606 ) | ( x69 & n32635 ) | ( ~n32606 & n32635 ) ;
  assign n32637 = ( x70 & ~n32598 ) | ( x70 & n32636 ) | ( ~n32598 & n32636 ) ;
  assign n32638 = ( x71 & ~n32590 ) | ( x71 & n32637 ) | ( ~n32590 & n32637 ) ;
  assign n32639 = ( x72 & ~n32582 ) | ( x72 & n32638 ) | ( ~n32582 & n32638 ) ;
  assign n32640 = ( x73 & ~n32574 ) | ( x73 & n32639 ) | ( ~n32574 & n32639 ) ;
  assign n32641 = ( x74 & ~n32566 ) | ( x74 & n32640 ) | ( ~n32566 & n32640 ) ;
  assign n32642 = ( x75 & ~n32558 ) | ( x75 & n32641 ) | ( ~n32558 & n32641 ) ;
  assign n32643 = ( x76 & ~n32550 ) | ( x76 & n32642 ) | ( ~n32550 & n32642 ) ;
  assign n32644 = ( x77 & ~n32542 ) | ( x77 & n32643 ) | ( ~n32542 & n32643 ) ;
  assign n32645 = ( x78 & ~n32534 ) | ( x78 & n32644 ) | ( ~n32534 & n32644 ) ;
  assign n32646 = ( x79 & ~n32526 ) | ( x79 & n32645 ) | ( ~n32526 & n32645 ) ;
  assign n32647 = ( x80 & ~n32518 ) | ( x80 & n32646 ) | ( ~n32518 & n32646 ) ;
  assign n32648 = ( x81 & ~n32510 ) | ( x81 & n32647 ) | ( ~n32510 & n32647 ) ;
  assign n32649 = ( x82 & ~n32502 ) | ( x82 & n32648 ) | ( ~n32502 & n32648 ) ;
  assign n32650 = ( x83 & ~n32494 ) | ( x83 & n32649 ) | ( ~n32494 & n32649 ) ;
  assign n32651 = ( x84 & ~n32486 ) | ( x84 & n32650 ) | ( ~n32486 & n32650 ) ;
  assign n32652 = ( x85 & ~n32478 ) | ( x85 & n32651 ) | ( ~n32478 & n32651 ) ;
  assign n32653 = ( x86 & ~n32470 ) | ( x86 & n32652 ) | ( ~n32470 & n32652 ) ;
  assign n32654 = ( x87 & ~n32462 ) | ( x87 & n32653 ) | ( ~n32462 & n32653 ) ;
  assign n32655 = ( x88 & ~n32454 ) | ( x88 & n32654 ) | ( ~n32454 & n32654 ) ;
  assign n32656 = ( x89 & ~n32446 ) | ( x89 & n32655 ) | ( ~n32446 & n32655 ) ;
  assign n32657 = ( x90 & ~n32438 ) | ( x90 & n32656 ) | ( ~n32438 & n32656 ) ;
  assign n32658 = ( x91 & ~n32430 ) | ( x91 & n32657 ) | ( ~n32430 & n32657 ) ;
  assign n32659 = ( x92 & ~n32422 ) | ( x92 & n32658 ) | ( ~n32422 & n32658 ) ;
  assign n32660 = ( x93 & ~n32414 ) | ( x93 & n32659 ) | ( ~n32414 & n32659 ) ;
  assign n32661 = ( x94 & ~n32406 ) | ( x94 & n32660 ) | ( ~n32406 & n32660 ) ;
  assign n32662 = ( x95 & ~n32398 ) | ( x95 & n32661 ) | ( ~n32398 & n32661 ) ;
  assign n32663 = ( x96 & ~n32390 ) | ( x96 & n32662 ) | ( ~n32390 & n32662 ) ;
  assign n32664 = ( x97 & ~n32382 ) | ( x97 & n32663 ) | ( ~n32382 & n32663 ) ;
  assign n32665 = ( x98 & ~n32374 ) | ( x98 & n32664 ) | ( ~n32374 & n32664 ) ;
  assign n32666 = ( x99 & ~n32366 ) | ( x99 & n32665 ) | ( ~n32366 & n32665 ) ;
  assign n32667 = ( x100 & ~n32358 ) | ( x100 & n32666 ) | ( ~n32358 & n32666 ) ;
  assign n32668 = ( x101 & ~n32350 ) | ( x101 & n32667 ) | ( ~n32350 & n32667 ) ;
  assign n32669 = ( x102 & ~n32342 ) | ( x102 & n32668 ) | ( ~n32342 & n32668 ) ;
  assign n32670 = ( x103 & ~n32334 ) | ( x103 & n32669 ) | ( ~n32334 & n32669 ) ;
  assign n32671 = ( x104 & ~n32326 ) | ( x104 & n32670 ) | ( ~n32326 & n32670 ) ;
  assign n32672 = ( x105 & ~n32318 ) | ( x105 & n32671 ) | ( ~n32318 & n32671 ) ;
  assign n32673 = ( x106 & ~n32310 ) | ( x106 & n32672 ) | ( ~n32310 & n32672 ) ;
  assign n32674 = ( x107 & ~n32302 ) | ( x107 & n32673 ) | ( ~n32302 & n32673 ) ;
  assign n32675 = ( x108 & ~n32294 ) | ( x108 & n32674 ) | ( ~n32294 & n32674 ) ;
  assign n32676 = ( x109 & ~n32286 ) | ( x109 & n32675 ) | ( ~n32286 & n32675 ) ;
  assign n32677 = ( x110 & ~n32278 ) | ( x110 & n32676 ) | ( ~n32278 & n32676 ) ;
  assign n32678 = ( x111 & ~n32270 ) | ( x111 & n32677 ) | ( ~n32270 & n32677 ) ;
  assign n32679 = ( x112 & ~n32262 ) | ( x112 & n32678 ) | ( ~n32262 & n32678 ) ;
  assign n32680 = ( x113 & ~n32254 ) | ( x113 & n32679 ) | ( ~n32254 & n32679 ) ;
  assign n32681 = ( x114 & ~n32246 ) | ( x114 & n32680 ) | ( ~n32246 & n32680 ) ;
  assign n32682 = ( x115 & ~n32238 ) | ( x115 & n32681 ) | ( ~n32238 & n32681 ) ;
  assign n32683 = ( x116 & ~n32230 ) | ( x116 & n32682 ) | ( ~n32230 & n32682 ) ;
  assign n32684 = ( x117 & ~n32222 ) | ( x117 & n32683 ) | ( ~n32222 & n32683 ) ;
  assign n32685 = ( x118 & ~n32214 ) | ( x118 & n32684 ) | ( ~n32214 & n32684 ) ;
  assign n32198 = n31727 &  n32197 ;
  assign n32202 = ( n13898 & n31727 ) | ( n13898 & n32195 ) | ( n31727 & n32195 ) ;
  assign n32203 = ( x118 & ~n32202 ) | ( x118 & n31727 ) | ( ~n32202 & n31727 ) ;
  assign n32204 = ~x118 & n32203 ;
  assign n32205 = n32198 | n32204 ;
  assign n32206 = ~x119 & n32205 ;
  assign n32686 = ( x119 & ~n32198 ) | ( x119 & 1'b0 ) | ( ~n32198 & 1'b0 ) ;
  assign n32687 = ~n32204 & n32686 ;
  assign n32696 = n32206 | n32687 ;
  assign n32697 = ( n32685 & ~n32696 ) | ( n32685 & 1'b0 ) | ( ~n32696 & 1'b0 ) ;
  assign n32688 = ( n32685 & ~n32206 ) | ( n32685 & n32687 ) | ( ~n32206 & n32687 ) ;
  assign n32689 = ( n32206 & ~n269 ) | ( n32206 & n32688 ) | ( ~n269 & n32688 ) ;
  assign n32690 = n269 | n32689 ;
  assign n32691 = ~n32205 |  n13898 ;
  assign n32692 = n32690 &  n32691 ;
  assign n32698 = ~n32685 & n32696 ;
  assign n32699 = ( n32697 & ~n32692 ) | ( n32697 & n32698 ) | ( ~n32692 & n32698 ) ;
  assign n32700 = n13898 &  n31727 ;
  assign n32701 = n32690 &  n32700 ;
  assign n32702 = n32699 | n32701 ;
  assign n32703 = ~x120 & n32702 ;
  assign n32707 = n32214 &  n32691 ;
  assign n32708 = n32690 &  n32707 ;
  assign n32693 = x118 | n32214 ;
  assign n32694 = x118 &  n32214 ;
  assign n32695 = ( n32693 & ~n32694 ) | ( n32693 & 1'b0 ) | ( ~n32694 & 1'b0 ) ;
  assign n32710 = ( n32684 & n32692 ) | ( n32684 & n32695 ) | ( n32692 & n32695 ) ;
  assign n32709 = n32684 | n32695 ;
  assign n32711 = ( n32708 & ~n32710 ) | ( n32708 & n32709 ) | ( ~n32710 & n32709 ) ;
  assign n32715 = n32222 &  n32691 ;
  assign n32716 = n32690 &  n32715 ;
  assign n32704 = x117 | n32222 ;
  assign n32705 = x117 &  n32222 ;
  assign n32706 = ( n32704 & ~n32705 ) | ( n32704 & 1'b0 ) | ( ~n32705 & 1'b0 ) ;
  assign n32718 = ( n32683 & n32692 ) | ( n32683 & n32706 ) | ( n32692 & n32706 ) ;
  assign n32717 = n32683 | n32706 ;
  assign n32719 = ( n32716 & ~n32718 ) | ( n32716 & n32717 ) | ( ~n32718 & n32717 ) ;
  assign n32723 = n32230 &  n32691 ;
  assign n32724 = n32690 &  n32723 ;
  assign n32712 = x116 | n32230 ;
  assign n32713 = x116 &  n32230 ;
  assign n32714 = ( n32712 & ~n32713 ) | ( n32712 & 1'b0 ) | ( ~n32713 & 1'b0 ) ;
  assign n32726 = ( n32682 & n32692 ) | ( n32682 & n32714 ) | ( n32692 & n32714 ) ;
  assign n32725 = n32682 | n32714 ;
  assign n32727 = ( n32724 & ~n32726 ) | ( n32724 & n32725 ) | ( ~n32726 & n32725 ) ;
  assign n32731 = n32238 &  n32691 ;
  assign n32732 = n32690 &  n32731 ;
  assign n32720 = x115 | n32238 ;
  assign n32721 = x115 &  n32238 ;
  assign n32722 = ( n32720 & ~n32721 ) | ( n32720 & 1'b0 ) | ( ~n32721 & 1'b0 ) ;
  assign n32734 = ( n32681 & n32692 ) | ( n32681 & n32722 ) | ( n32692 & n32722 ) ;
  assign n32733 = n32681 | n32722 ;
  assign n32735 = ( n32732 & ~n32734 ) | ( n32732 & n32733 ) | ( ~n32734 & n32733 ) ;
  assign n32739 = n32246 &  n32691 ;
  assign n32740 = n32690 &  n32739 ;
  assign n32728 = x114 | n32246 ;
  assign n32729 = x114 &  n32246 ;
  assign n32730 = ( n32728 & ~n32729 ) | ( n32728 & 1'b0 ) | ( ~n32729 & 1'b0 ) ;
  assign n32742 = ( n32680 & n32692 ) | ( n32680 & n32730 ) | ( n32692 & n32730 ) ;
  assign n32741 = n32680 | n32730 ;
  assign n32743 = ( n32740 & ~n32742 ) | ( n32740 & n32741 ) | ( ~n32742 & n32741 ) ;
  assign n32747 = n32254 &  n32691 ;
  assign n32748 = n32690 &  n32747 ;
  assign n32736 = x113 | n32254 ;
  assign n32737 = x113 &  n32254 ;
  assign n32738 = ( n32736 & ~n32737 ) | ( n32736 & 1'b0 ) | ( ~n32737 & 1'b0 ) ;
  assign n32750 = ( n32679 & n32692 ) | ( n32679 & n32738 ) | ( n32692 & n32738 ) ;
  assign n32749 = n32679 | n32738 ;
  assign n32751 = ( n32748 & ~n32750 ) | ( n32748 & n32749 ) | ( ~n32750 & n32749 ) ;
  assign n32755 = n32262 &  n32691 ;
  assign n32756 = n32690 &  n32755 ;
  assign n32744 = x112 | n32262 ;
  assign n32745 = x112 &  n32262 ;
  assign n32746 = ( n32744 & ~n32745 ) | ( n32744 & 1'b0 ) | ( ~n32745 & 1'b0 ) ;
  assign n32758 = ( n32678 & n32692 ) | ( n32678 & n32746 ) | ( n32692 & n32746 ) ;
  assign n32757 = n32678 | n32746 ;
  assign n32759 = ( n32756 & ~n32758 ) | ( n32756 & n32757 ) | ( ~n32758 & n32757 ) ;
  assign n32763 = n32270 &  n32691 ;
  assign n32764 = n32690 &  n32763 ;
  assign n32752 = x111 | n32270 ;
  assign n32753 = x111 &  n32270 ;
  assign n32754 = ( n32752 & ~n32753 ) | ( n32752 & 1'b0 ) | ( ~n32753 & 1'b0 ) ;
  assign n32766 = ( n32677 & n32692 ) | ( n32677 & n32754 ) | ( n32692 & n32754 ) ;
  assign n32765 = n32677 | n32754 ;
  assign n32767 = ( n32764 & ~n32766 ) | ( n32764 & n32765 ) | ( ~n32766 & n32765 ) ;
  assign n32771 = n32278 &  n32691 ;
  assign n32772 = n32690 &  n32771 ;
  assign n32760 = x110 | n32278 ;
  assign n32761 = x110 &  n32278 ;
  assign n32762 = ( n32760 & ~n32761 ) | ( n32760 & 1'b0 ) | ( ~n32761 & 1'b0 ) ;
  assign n32774 = ( n32676 & n32692 ) | ( n32676 & n32762 ) | ( n32692 & n32762 ) ;
  assign n32773 = n32676 | n32762 ;
  assign n32775 = ( n32772 & ~n32774 ) | ( n32772 & n32773 ) | ( ~n32774 & n32773 ) ;
  assign n32779 = n32286 &  n32691 ;
  assign n32780 = n32690 &  n32779 ;
  assign n32768 = x109 | n32286 ;
  assign n32769 = x109 &  n32286 ;
  assign n32770 = ( n32768 & ~n32769 ) | ( n32768 & 1'b0 ) | ( ~n32769 & 1'b0 ) ;
  assign n32782 = ( n32675 & n32692 ) | ( n32675 & n32770 ) | ( n32692 & n32770 ) ;
  assign n32781 = n32675 | n32770 ;
  assign n32783 = ( n32780 & ~n32782 ) | ( n32780 & n32781 ) | ( ~n32782 & n32781 ) ;
  assign n32787 = n32294 &  n32691 ;
  assign n32788 = n32690 &  n32787 ;
  assign n32776 = x108 | n32294 ;
  assign n32777 = x108 &  n32294 ;
  assign n32778 = ( n32776 & ~n32777 ) | ( n32776 & 1'b0 ) | ( ~n32777 & 1'b0 ) ;
  assign n32790 = ( n32674 & n32692 ) | ( n32674 & n32778 ) | ( n32692 & n32778 ) ;
  assign n32789 = n32674 | n32778 ;
  assign n32791 = ( n32788 & ~n32790 ) | ( n32788 & n32789 ) | ( ~n32790 & n32789 ) ;
  assign n32795 = n32302 &  n32691 ;
  assign n32796 = n32690 &  n32795 ;
  assign n32784 = x107 | n32302 ;
  assign n32785 = x107 &  n32302 ;
  assign n32786 = ( n32784 & ~n32785 ) | ( n32784 & 1'b0 ) | ( ~n32785 & 1'b0 ) ;
  assign n32798 = ( n32673 & n32692 ) | ( n32673 & n32786 ) | ( n32692 & n32786 ) ;
  assign n32797 = n32673 | n32786 ;
  assign n32799 = ( n32796 & ~n32798 ) | ( n32796 & n32797 ) | ( ~n32798 & n32797 ) ;
  assign n32803 = n32310 &  n32691 ;
  assign n32804 = n32690 &  n32803 ;
  assign n32792 = x106 | n32310 ;
  assign n32793 = x106 &  n32310 ;
  assign n32794 = ( n32792 & ~n32793 ) | ( n32792 & 1'b0 ) | ( ~n32793 & 1'b0 ) ;
  assign n32806 = ( n32672 & n32692 ) | ( n32672 & n32794 ) | ( n32692 & n32794 ) ;
  assign n32805 = n32672 | n32794 ;
  assign n32807 = ( n32804 & ~n32806 ) | ( n32804 & n32805 ) | ( ~n32806 & n32805 ) ;
  assign n32811 = n32318 &  n32691 ;
  assign n32812 = n32690 &  n32811 ;
  assign n32800 = x105 | n32318 ;
  assign n32801 = x105 &  n32318 ;
  assign n32802 = ( n32800 & ~n32801 ) | ( n32800 & 1'b0 ) | ( ~n32801 & 1'b0 ) ;
  assign n32814 = ( n32671 & n32692 ) | ( n32671 & n32802 ) | ( n32692 & n32802 ) ;
  assign n32813 = n32671 | n32802 ;
  assign n32815 = ( n32812 & ~n32814 ) | ( n32812 & n32813 ) | ( ~n32814 & n32813 ) ;
  assign n32819 = n32326 &  n32691 ;
  assign n32820 = n32690 &  n32819 ;
  assign n32808 = x104 | n32326 ;
  assign n32809 = x104 &  n32326 ;
  assign n32810 = ( n32808 & ~n32809 ) | ( n32808 & 1'b0 ) | ( ~n32809 & 1'b0 ) ;
  assign n32822 = ( n32670 & n32692 ) | ( n32670 & n32810 ) | ( n32692 & n32810 ) ;
  assign n32821 = n32670 | n32810 ;
  assign n32823 = ( n32820 & ~n32822 ) | ( n32820 & n32821 ) | ( ~n32822 & n32821 ) ;
  assign n32827 = n32334 &  n32691 ;
  assign n32828 = n32690 &  n32827 ;
  assign n32816 = x103 | n32334 ;
  assign n32817 = x103 &  n32334 ;
  assign n32818 = ( n32816 & ~n32817 ) | ( n32816 & 1'b0 ) | ( ~n32817 & 1'b0 ) ;
  assign n32830 = ( n32669 & n32692 ) | ( n32669 & n32818 ) | ( n32692 & n32818 ) ;
  assign n32829 = n32669 | n32818 ;
  assign n32831 = ( n32828 & ~n32830 ) | ( n32828 & n32829 ) | ( ~n32830 & n32829 ) ;
  assign n32835 = n32342 &  n32691 ;
  assign n32836 = n32690 &  n32835 ;
  assign n32824 = x102 | n32342 ;
  assign n32825 = x102 &  n32342 ;
  assign n32826 = ( n32824 & ~n32825 ) | ( n32824 & 1'b0 ) | ( ~n32825 & 1'b0 ) ;
  assign n32838 = ( n32668 & n32692 ) | ( n32668 & n32826 ) | ( n32692 & n32826 ) ;
  assign n32837 = n32668 | n32826 ;
  assign n32839 = ( n32836 & ~n32838 ) | ( n32836 & n32837 ) | ( ~n32838 & n32837 ) ;
  assign n32843 = n32350 &  n32691 ;
  assign n32844 = n32690 &  n32843 ;
  assign n32832 = x101 | n32350 ;
  assign n32833 = x101 &  n32350 ;
  assign n32834 = ( n32832 & ~n32833 ) | ( n32832 & 1'b0 ) | ( ~n32833 & 1'b0 ) ;
  assign n32846 = ( n32667 & n32692 ) | ( n32667 & n32834 ) | ( n32692 & n32834 ) ;
  assign n32845 = n32667 | n32834 ;
  assign n32847 = ( n32844 & ~n32846 ) | ( n32844 & n32845 ) | ( ~n32846 & n32845 ) ;
  assign n32851 = n32358 &  n32691 ;
  assign n32852 = n32690 &  n32851 ;
  assign n32840 = x100 | n32358 ;
  assign n32841 = x100 &  n32358 ;
  assign n32842 = ( n32840 & ~n32841 ) | ( n32840 & 1'b0 ) | ( ~n32841 & 1'b0 ) ;
  assign n32854 = ( n32666 & n32692 ) | ( n32666 & n32842 ) | ( n32692 & n32842 ) ;
  assign n32853 = n32666 | n32842 ;
  assign n32855 = ( n32852 & ~n32854 ) | ( n32852 & n32853 ) | ( ~n32854 & n32853 ) ;
  assign n32859 = n32366 &  n32691 ;
  assign n32860 = n32690 &  n32859 ;
  assign n32848 = x99 | n32366 ;
  assign n32849 = x99 &  n32366 ;
  assign n32850 = ( n32848 & ~n32849 ) | ( n32848 & 1'b0 ) | ( ~n32849 & 1'b0 ) ;
  assign n32862 = ( n32665 & n32692 ) | ( n32665 & n32850 ) | ( n32692 & n32850 ) ;
  assign n32861 = n32665 | n32850 ;
  assign n32863 = ( n32860 & ~n32862 ) | ( n32860 & n32861 ) | ( ~n32862 & n32861 ) ;
  assign n32867 = n32374 &  n32691 ;
  assign n32868 = n32690 &  n32867 ;
  assign n32856 = x98 | n32374 ;
  assign n32857 = x98 &  n32374 ;
  assign n32858 = ( n32856 & ~n32857 ) | ( n32856 & 1'b0 ) | ( ~n32857 & 1'b0 ) ;
  assign n32870 = ( n32664 & n32692 ) | ( n32664 & n32858 ) | ( n32692 & n32858 ) ;
  assign n32869 = n32664 | n32858 ;
  assign n32871 = ( n32868 & ~n32870 ) | ( n32868 & n32869 ) | ( ~n32870 & n32869 ) ;
  assign n32875 = n32382 &  n32691 ;
  assign n32876 = n32690 &  n32875 ;
  assign n32864 = x97 | n32382 ;
  assign n32865 = x97 &  n32382 ;
  assign n32866 = ( n32864 & ~n32865 ) | ( n32864 & 1'b0 ) | ( ~n32865 & 1'b0 ) ;
  assign n32878 = ( n32663 & n32692 ) | ( n32663 & n32866 ) | ( n32692 & n32866 ) ;
  assign n32877 = n32663 | n32866 ;
  assign n32879 = ( n32876 & ~n32878 ) | ( n32876 & n32877 ) | ( ~n32878 & n32877 ) ;
  assign n32883 = n32390 &  n32691 ;
  assign n32884 = n32690 &  n32883 ;
  assign n32872 = x96 | n32390 ;
  assign n32873 = x96 &  n32390 ;
  assign n32874 = ( n32872 & ~n32873 ) | ( n32872 & 1'b0 ) | ( ~n32873 & 1'b0 ) ;
  assign n32886 = ( n32662 & n32692 ) | ( n32662 & n32874 ) | ( n32692 & n32874 ) ;
  assign n32885 = n32662 | n32874 ;
  assign n32887 = ( n32884 & ~n32886 ) | ( n32884 & n32885 ) | ( ~n32886 & n32885 ) ;
  assign n32891 = n32398 &  n32691 ;
  assign n32892 = n32690 &  n32891 ;
  assign n32880 = x95 | n32398 ;
  assign n32881 = x95 &  n32398 ;
  assign n32882 = ( n32880 & ~n32881 ) | ( n32880 & 1'b0 ) | ( ~n32881 & 1'b0 ) ;
  assign n32894 = ( n32661 & n32692 ) | ( n32661 & n32882 ) | ( n32692 & n32882 ) ;
  assign n32893 = n32661 | n32882 ;
  assign n32895 = ( n32892 & ~n32894 ) | ( n32892 & n32893 ) | ( ~n32894 & n32893 ) ;
  assign n32899 = n32406 &  n32691 ;
  assign n32900 = n32690 &  n32899 ;
  assign n32888 = x94 | n32406 ;
  assign n32889 = x94 &  n32406 ;
  assign n32890 = ( n32888 & ~n32889 ) | ( n32888 & 1'b0 ) | ( ~n32889 & 1'b0 ) ;
  assign n32902 = ( n32660 & n32692 ) | ( n32660 & n32890 ) | ( n32692 & n32890 ) ;
  assign n32901 = n32660 | n32890 ;
  assign n32903 = ( n32900 & ~n32902 ) | ( n32900 & n32901 ) | ( ~n32902 & n32901 ) ;
  assign n32907 = n32414 &  n32691 ;
  assign n32908 = n32690 &  n32907 ;
  assign n32896 = x93 | n32414 ;
  assign n32897 = x93 &  n32414 ;
  assign n32898 = ( n32896 & ~n32897 ) | ( n32896 & 1'b0 ) | ( ~n32897 & 1'b0 ) ;
  assign n32910 = ( n32659 & n32692 ) | ( n32659 & n32898 ) | ( n32692 & n32898 ) ;
  assign n32909 = n32659 | n32898 ;
  assign n32911 = ( n32908 & ~n32910 ) | ( n32908 & n32909 ) | ( ~n32910 & n32909 ) ;
  assign n32915 = n32422 &  n32691 ;
  assign n32916 = n32690 &  n32915 ;
  assign n32904 = x92 | n32422 ;
  assign n32905 = x92 &  n32422 ;
  assign n32906 = ( n32904 & ~n32905 ) | ( n32904 & 1'b0 ) | ( ~n32905 & 1'b0 ) ;
  assign n32918 = ( n32658 & n32692 ) | ( n32658 & n32906 ) | ( n32692 & n32906 ) ;
  assign n32917 = n32658 | n32906 ;
  assign n32919 = ( n32916 & ~n32918 ) | ( n32916 & n32917 ) | ( ~n32918 & n32917 ) ;
  assign n32923 = n32430 &  n32691 ;
  assign n32924 = n32690 &  n32923 ;
  assign n32912 = x91 | n32430 ;
  assign n32913 = x91 &  n32430 ;
  assign n32914 = ( n32912 & ~n32913 ) | ( n32912 & 1'b0 ) | ( ~n32913 & 1'b0 ) ;
  assign n32926 = ( n32657 & n32692 ) | ( n32657 & n32914 ) | ( n32692 & n32914 ) ;
  assign n32925 = n32657 | n32914 ;
  assign n32927 = ( n32924 & ~n32926 ) | ( n32924 & n32925 ) | ( ~n32926 & n32925 ) ;
  assign n32931 = n32438 &  n32691 ;
  assign n32932 = n32690 &  n32931 ;
  assign n32920 = x90 | n32438 ;
  assign n32921 = x90 &  n32438 ;
  assign n32922 = ( n32920 & ~n32921 ) | ( n32920 & 1'b0 ) | ( ~n32921 & 1'b0 ) ;
  assign n32934 = ( n32656 & n32692 ) | ( n32656 & n32922 ) | ( n32692 & n32922 ) ;
  assign n32933 = n32656 | n32922 ;
  assign n32935 = ( n32932 & ~n32934 ) | ( n32932 & n32933 ) | ( ~n32934 & n32933 ) ;
  assign n32939 = n32446 &  n32691 ;
  assign n32940 = n32690 &  n32939 ;
  assign n32928 = x89 | n32446 ;
  assign n32929 = x89 &  n32446 ;
  assign n32930 = ( n32928 & ~n32929 ) | ( n32928 & 1'b0 ) | ( ~n32929 & 1'b0 ) ;
  assign n32942 = ( n32655 & n32692 ) | ( n32655 & n32930 ) | ( n32692 & n32930 ) ;
  assign n32941 = n32655 | n32930 ;
  assign n32943 = ( n32940 & ~n32942 ) | ( n32940 & n32941 ) | ( ~n32942 & n32941 ) ;
  assign n32947 = n32454 &  n32691 ;
  assign n32948 = n32690 &  n32947 ;
  assign n32936 = x88 | n32454 ;
  assign n32937 = x88 &  n32454 ;
  assign n32938 = ( n32936 & ~n32937 ) | ( n32936 & 1'b0 ) | ( ~n32937 & 1'b0 ) ;
  assign n32950 = ( n32654 & n32692 ) | ( n32654 & n32938 ) | ( n32692 & n32938 ) ;
  assign n32949 = n32654 | n32938 ;
  assign n32951 = ( n32948 & ~n32950 ) | ( n32948 & n32949 ) | ( ~n32950 & n32949 ) ;
  assign n32955 = n32462 &  n32691 ;
  assign n32956 = n32690 &  n32955 ;
  assign n32944 = x87 | n32462 ;
  assign n32945 = x87 &  n32462 ;
  assign n32946 = ( n32944 & ~n32945 ) | ( n32944 & 1'b0 ) | ( ~n32945 & 1'b0 ) ;
  assign n32958 = ( n32653 & n32692 ) | ( n32653 & n32946 ) | ( n32692 & n32946 ) ;
  assign n32957 = n32653 | n32946 ;
  assign n32959 = ( n32956 & ~n32958 ) | ( n32956 & n32957 ) | ( ~n32958 & n32957 ) ;
  assign n32963 = n32470 &  n32691 ;
  assign n32964 = n32690 &  n32963 ;
  assign n32952 = x86 | n32470 ;
  assign n32953 = x86 &  n32470 ;
  assign n32954 = ( n32952 & ~n32953 ) | ( n32952 & 1'b0 ) | ( ~n32953 & 1'b0 ) ;
  assign n32966 = ( n32652 & n32692 ) | ( n32652 & n32954 ) | ( n32692 & n32954 ) ;
  assign n32965 = n32652 | n32954 ;
  assign n32967 = ( n32964 & ~n32966 ) | ( n32964 & n32965 ) | ( ~n32966 & n32965 ) ;
  assign n32971 = n32478 &  n32691 ;
  assign n32972 = n32690 &  n32971 ;
  assign n32960 = x85 | n32478 ;
  assign n32961 = x85 &  n32478 ;
  assign n32962 = ( n32960 & ~n32961 ) | ( n32960 & 1'b0 ) | ( ~n32961 & 1'b0 ) ;
  assign n32974 = ( n32651 & n32692 ) | ( n32651 & n32962 ) | ( n32692 & n32962 ) ;
  assign n32973 = n32651 | n32962 ;
  assign n32975 = ( n32972 & ~n32974 ) | ( n32972 & n32973 ) | ( ~n32974 & n32973 ) ;
  assign n32979 = n32486 &  n32691 ;
  assign n32980 = n32690 &  n32979 ;
  assign n32968 = x84 | n32486 ;
  assign n32969 = x84 &  n32486 ;
  assign n32970 = ( n32968 & ~n32969 ) | ( n32968 & 1'b0 ) | ( ~n32969 & 1'b0 ) ;
  assign n32982 = ( n32650 & n32692 ) | ( n32650 & n32970 ) | ( n32692 & n32970 ) ;
  assign n32981 = n32650 | n32970 ;
  assign n32983 = ( n32980 & ~n32982 ) | ( n32980 & n32981 ) | ( ~n32982 & n32981 ) ;
  assign n32987 = n32494 &  n32691 ;
  assign n32988 = n32690 &  n32987 ;
  assign n32976 = x83 | n32494 ;
  assign n32977 = x83 &  n32494 ;
  assign n32978 = ( n32976 & ~n32977 ) | ( n32976 & 1'b0 ) | ( ~n32977 & 1'b0 ) ;
  assign n32990 = ( n32649 & n32692 ) | ( n32649 & n32978 ) | ( n32692 & n32978 ) ;
  assign n32989 = n32649 | n32978 ;
  assign n32991 = ( n32988 & ~n32990 ) | ( n32988 & n32989 ) | ( ~n32990 & n32989 ) ;
  assign n32995 = n32502 &  n32691 ;
  assign n32996 = n32690 &  n32995 ;
  assign n32984 = x82 | n32502 ;
  assign n32985 = x82 &  n32502 ;
  assign n32986 = ( n32984 & ~n32985 ) | ( n32984 & 1'b0 ) | ( ~n32985 & 1'b0 ) ;
  assign n32998 = ( n32648 & n32692 ) | ( n32648 & n32986 ) | ( n32692 & n32986 ) ;
  assign n32997 = n32648 | n32986 ;
  assign n32999 = ( n32996 & ~n32998 ) | ( n32996 & n32997 ) | ( ~n32998 & n32997 ) ;
  assign n33003 = n32510 &  n32691 ;
  assign n33004 = n32690 &  n33003 ;
  assign n32992 = x81 | n32510 ;
  assign n32993 = x81 &  n32510 ;
  assign n32994 = ( n32992 & ~n32993 ) | ( n32992 & 1'b0 ) | ( ~n32993 & 1'b0 ) ;
  assign n33006 = ( n32647 & n32692 ) | ( n32647 & n32994 ) | ( n32692 & n32994 ) ;
  assign n33005 = n32647 | n32994 ;
  assign n33007 = ( n33004 & ~n33006 ) | ( n33004 & n33005 ) | ( ~n33006 & n33005 ) ;
  assign n33011 = n32518 &  n32691 ;
  assign n33012 = n32690 &  n33011 ;
  assign n33000 = x80 | n32518 ;
  assign n33001 = x80 &  n32518 ;
  assign n33002 = ( n33000 & ~n33001 ) | ( n33000 & 1'b0 ) | ( ~n33001 & 1'b0 ) ;
  assign n33014 = ( n32646 & n32692 ) | ( n32646 & n33002 ) | ( n32692 & n33002 ) ;
  assign n33013 = n32646 | n33002 ;
  assign n33015 = ( n33012 & ~n33014 ) | ( n33012 & n33013 ) | ( ~n33014 & n33013 ) ;
  assign n33019 = n32526 &  n32691 ;
  assign n33020 = n32690 &  n33019 ;
  assign n33008 = x79 | n32526 ;
  assign n33009 = x79 &  n32526 ;
  assign n33010 = ( n33008 & ~n33009 ) | ( n33008 & 1'b0 ) | ( ~n33009 & 1'b0 ) ;
  assign n33022 = ( n32645 & n32692 ) | ( n32645 & n33010 ) | ( n32692 & n33010 ) ;
  assign n33021 = n32645 | n33010 ;
  assign n33023 = ( n33020 & ~n33022 ) | ( n33020 & n33021 ) | ( ~n33022 & n33021 ) ;
  assign n33027 = n32534 &  n32691 ;
  assign n33028 = n32690 &  n33027 ;
  assign n33016 = x78 | n32534 ;
  assign n33017 = x78 &  n32534 ;
  assign n33018 = ( n33016 & ~n33017 ) | ( n33016 & 1'b0 ) | ( ~n33017 & 1'b0 ) ;
  assign n33030 = ( n32644 & n32692 ) | ( n32644 & n33018 ) | ( n32692 & n33018 ) ;
  assign n33029 = n32644 | n33018 ;
  assign n33031 = ( n33028 & ~n33030 ) | ( n33028 & n33029 ) | ( ~n33030 & n33029 ) ;
  assign n33035 = n32542 &  n32691 ;
  assign n33036 = n32690 &  n33035 ;
  assign n33024 = x77 | n32542 ;
  assign n33025 = x77 &  n32542 ;
  assign n33026 = ( n33024 & ~n33025 ) | ( n33024 & 1'b0 ) | ( ~n33025 & 1'b0 ) ;
  assign n33038 = ( n32643 & n32692 ) | ( n32643 & n33026 ) | ( n32692 & n33026 ) ;
  assign n33037 = n32643 | n33026 ;
  assign n33039 = ( n33036 & ~n33038 ) | ( n33036 & n33037 ) | ( ~n33038 & n33037 ) ;
  assign n33043 = n32550 &  n32691 ;
  assign n33044 = n32690 &  n33043 ;
  assign n33032 = x76 | n32550 ;
  assign n33033 = x76 &  n32550 ;
  assign n33034 = ( n33032 & ~n33033 ) | ( n33032 & 1'b0 ) | ( ~n33033 & 1'b0 ) ;
  assign n33046 = ( n32642 & n32692 ) | ( n32642 & n33034 ) | ( n32692 & n33034 ) ;
  assign n33045 = n32642 | n33034 ;
  assign n33047 = ( n33044 & ~n33046 ) | ( n33044 & n33045 ) | ( ~n33046 & n33045 ) ;
  assign n33051 = n32558 &  n32691 ;
  assign n33052 = n32690 &  n33051 ;
  assign n33040 = x75 | n32558 ;
  assign n33041 = x75 &  n32558 ;
  assign n33042 = ( n33040 & ~n33041 ) | ( n33040 & 1'b0 ) | ( ~n33041 & 1'b0 ) ;
  assign n33054 = ( n32641 & n32692 ) | ( n32641 & n33042 ) | ( n32692 & n33042 ) ;
  assign n33053 = n32641 | n33042 ;
  assign n33055 = ( n33052 & ~n33054 ) | ( n33052 & n33053 ) | ( ~n33054 & n33053 ) ;
  assign n33059 = n32566 &  n32691 ;
  assign n33060 = n32690 &  n33059 ;
  assign n33048 = x74 | n32566 ;
  assign n33049 = x74 &  n32566 ;
  assign n33050 = ( n33048 & ~n33049 ) | ( n33048 & 1'b0 ) | ( ~n33049 & 1'b0 ) ;
  assign n33062 = ( n32640 & n32692 ) | ( n32640 & n33050 ) | ( n32692 & n33050 ) ;
  assign n33061 = n32640 | n33050 ;
  assign n33063 = ( n33060 & ~n33062 ) | ( n33060 & n33061 ) | ( ~n33062 & n33061 ) ;
  assign n33067 = n32574 &  n32691 ;
  assign n33068 = n32690 &  n33067 ;
  assign n33056 = x73 | n32574 ;
  assign n33057 = x73 &  n32574 ;
  assign n33058 = ( n33056 & ~n33057 ) | ( n33056 & 1'b0 ) | ( ~n33057 & 1'b0 ) ;
  assign n33070 = ( n32639 & n32692 ) | ( n32639 & n33058 ) | ( n32692 & n33058 ) ;
  assign n33069 = n32639 | n33058 ;
  assign n33071 = ( n33068 & ~n33070 ) | ( n33068 & n33069 ) | ( ~n33070 & n33069 ) ;
  assign n33075 = n32582 &  n32691 ;
  assign n33076 = n32690 &  n33075 ;
  assign n33064 = x72 | n32582 ;
  assign n33065 = x72 &  n32582 ;
  assign n33066 = ( n33064 & ~n33065 ) | ( n33064 & 1'b0 ) | ( ~n33065 & 1'b0 ) ;
  assign n33078 = ( n32638 & n32692 ) | ( n32638 & n33066 ) | ( n32692 & n33066 ) ;
  assign n33077 = n32638 | n33066 ;
  assign n33079 = ( n33076 & ~n33078 ) | ( n33076 & n33077 ) | ( ~n33078 & n33077 ) ;
  assign n33083 = n32590 &  n32691 ;
  assign n33084 = n32690 &  n33083 ;
  assign n33072 = x71 | n32590 ;
  assign n33073 = x71 &  n32590 ;
  assign n33074 = ( n33072 & ~n33073 ) | ( n33072 & 1'b0 ) | ( ~n33073 & 1'b0 ) ;
  assign n33086 = ( n32637 & n32692 ) | ( n32637 & n33074 ) | ( n32692 & n33074 ) ;
  assign n33085 = n32637 | n33074 ;
  assign n33087 = ( n33084 & ~n33086 ) | ( n33084 & n33085 ) | ( ~n33086 & n33085 ) ;
  assign n33091 = n32598 &  n32691 ;
  assign n33092 = n32690 &  n33091 ;
  assign n33080 = x70 | n32598 ;
  assign n33081 = x70 &  n32598 ;
  assign n33082 = ( n33080 & ~n33081 ) | ( n33080 & 1'b0 ) | ( ~n33081 & 1'b0 ) ;
  assign n33094 = ( n32636 & n32692 ) | ( n32636 & n33082 ) | ( n32692 & n33082 ) ;
  assign n33093 = n32636 | n33082 ;
  assign n33095 = ( n33092 & ~n33094 ) | ( n33092 & n33093 ) | ( ~n33094 & n33093 ) ;
  assign n33099 = n32606 &  n32691 ;
  assign n33100 = n32690 &  n33099 ;
  assign n33088 = x69 | n32606 ;
  assign n33089 = x69 &  n32606 ;
  assign n33090 = ( n33088 & ~n33089 ) | ( n33088 & 1'b0 ) | ( ~n33089 & 1'b0 ) ;
  assign n33102 = ( n32635 & n32692 ) | ( n32635 & n33090 ) | ( n32692 & n33090 ) ;
  assign n33101 = n32635 | n33090 ;
  assign n33103 = ( n33100 & ~n33102 ) | ( n33100 & n33101 ) | ( ~n33102 & n33101 ) ;
  assign n33107 = n32614 &  n32691 ;
  assign n33108 = n32690 &  n33107 ;
  assign n33096 = x68 | n32614 ;
  assign n33097 = x68 &  n32614 ;
  assign n33098 = ( n33096 & ~n33097 ) | ( n33096 & 1'b0 ) | ( ~n33097 & 1'b0 ) ;
  assign n33110 = ( n32634 & n32692 ) | ( n32634 & n33098 ) | ( n32692 & n33098 ) ;
  assign n33109 = n32634 | n33098 ;
  assign n33111 = ( n33108 & ~n33110 ) | ( n33108 & n33109 ) | ( ~n33110 & n33109 ) ;
  assign n33115 = n32619 &  n32691 ;
  assign n33116 = n32690 &  n33115 ;
  assign n33104 = x67 | n32619 ;
  assign n33105 = x67 &  n32619 ;
  assign n33106 = ( n33104 & ~n33105 ) | ( n33104 & 1'b0 ) | ( ~n33105 & 1'b0 ) ;
  assign n33118 = ( n32633 & n32692 ) | ( n32633 & n33106 ) | ( n32692 & n33106 ) ;
  assign n33117 = n32633 | n33106 ;
  assign n33119 = ( n33116 & ~n33118 ) | ( n33116 & n33117 ) | ( ~n33118 & n33117 ) ;
  assign n33120 = n32627 &  n32691 ;
  assign n33121 = n32690 &  n33120 ;
  assign n33112 = x66 | n32627 ;
  assign n33113 = x66 &  n32627 ;
  assign n33114 = ( n33112 & ~n33113 ) | ( n33112 & 1'b0 ) | ( ~n33113 & 1'b0 ) ;
  assign n33123 = ( n32632 & n32692 ) | ( n32632 & n33114 ) | ( n32692 & n33114 ) ;
  assign n33122 = n32632 | n33114 ;
  assign n33124 = ( n33121 & ~n33123 ) | ( n33121 & n33122 ) | ( ~n33123 & n33122 ) ;
  assign n33125 = ( x65 & ~n14288 ) | ( x65 & n32631 ) | ( ~n14288 & n32631 ) ;
  assign n33126 = ( n32632 & ~x65 ) | ( n32632 & n33125 ) | ( ~x65 & n33125 ) ;
  assign n33127 = ~n32692 & n33126 ;
  assign n33128 = n32631 &  n32691 ;
  assign n33129 = n32690 &  n33128 ;
  assign n33130 = n33127 | n33129 ;
  assign n33131 = ( x64 & ~n32692 ) | ( x64 & 1'b0 ) | ( ~n32692 & 1'b0 ) ;
  assign n33132 = ( x8 & ~n33131 ) | ( x8 & 1'b0 ) | ( ~n33131 & 1'b0 ) ;
  assign n33133 = ( n14288 & ~n32692 ) | ( n14288 & 1'b0 ) | ( ~n32692 & 1'b0 ) ;
  assign n33134 = n33132 | n33133 ;
  assign n33135 = ( x65 & ~n33134 ) | ( x65 & n14798 ) | ( ~n33134 & n14798 ) ;
  assign n33136 = ( x66 & ~n33130 ) | ( x66 & n33135 ) | ( ~n33130 & n33135 ) ;
  assign n33137 = ( x67 & ~n33124 ) | ( x67 & n33136 ) | ( ~n33124 & n33136 ) ;
  assign n33138 = ( x68 & ~n33119 ) | ( x68 & n33137 ) | ( ~n33119 & n33137 ) ;
  assign n33139 = ( x69 & ~n33111 ) | ( x69 & n33138 ) | ( ~n33111 & n33138 ) ;
  assign n33140 = ( x70 & ~n33103 ) | ( x70 & n33139 ) | ( ~n33103 & n33139 ) ;
  assign n33141 = ( x71 & ~n33095 ) | ( x71 & n33140 ) | ( ~n33095 & n33140 ) ;
  assign n33142 = ( x72 & ~n33087 ) | ( x72 & n33141 ) | ( ~n33087 & n33141 ) ;
  assign n33143 = ( x73 & ~n33079 ) | ( x73 & n33142 ) | ( ~n33079 & n33142 ) ;
  assign n33144 = ( x74 & ~n33071 ) | ( x74 & n33143 ) | ( ~n33071 & n33143 ) ;
  assign n33145 = ( x75 & ~n33063 ) | ( x75 & n33144 ) | ( ~n33063 & n33144 ) ;
  assign n33146 = ( x76 & ~n33055 ) | ( x76 & n33145 ) | ( ~n33055 & n33145 ) ;
  assign n33147 = ( x77 & ~n33047 ) | ( x77 & n33146 ) | ( ~n33047 & n33146 ) ;
  assign n33148 = ( x78 & ~n33039 ) | ( x78 & n33147 ) | ( ~n33039 & n33147 ) ;
  assign n33149 = ( x79 & ~n33031 ) | ( x79 & n33148 ) | ( ~n33031 & n33148 ) ;
  assign n33150 = ( x80 & ~n33023 ) | ( x80 & n33149 ) | ( ~n33023 & n33149 ) ;
  assign n33151 = ( x81 & ~n33015 ) | ( x81 & n33150 ) | ( ~n33015 & n33150 ) ;
  assign n33152 = ( x82 & ~n33007 ) | ( x82 & n33151 ) | ( ~n33007 & n33151 ) ;
  assign n33153 = ( x83 & ~n32999 ) | ( x83 & n33152 ) | ( ~n32999 & n33152 ) ;
  assign n33154 = ( x84 & ~n32991 ) | ( x84 & n33153 ) | ( ~n32991 & n33153 ) ;
  assign n33155 = ( x85 & ~n32983 ) | ( x85 & n33154 ) | ( ~n32983 & n33154 ) ;
  assign n33156 = ( x86 & ~n32975 ) | ( x86 & n33155 ) | ( ~n32975 & n33155 ) ;
  assign n33157 = ( x87 & ~n32967 ) | ( x87 & n33156 ) | ( ~n32967 & n33156 ) ;
  assign n33158 = ( x88 & ~n32959 ) | ( x88 & n33157 ) | ( ~n32959 & n33157 ) ;
  assign n33159 = ( x89 & ~n32951 ) | ( x89 & n33158 ) | ( ~n32951 & n33158 ) ;
  assign n33160 = ( x90 & ~n32943 ) | ( x90 & n33159 ) | ( ~n32943 & n33159 ) ;
  assign n33161 = ( x91 & ~n32935 ) | ( x91 & n33160 ) | ( ~n32935 & n33160 ) ;
  assign n33162 = ( x92 & ~n32927 ) | ( x92 & n33161 ) | ( ~n32927 & n33161 ) ;
  assign n33163 = ( x93 & ~n32919 ) | ( x93 & n33162 ) | ( ~n32919 & n33162 ) ;
  assign n33164 = ( x94 & ~n32911 ) | ( x94 & n33163 ) | ( ~n32911 & n33163 ) ;
  assign n33165 = ( x95 & ~n32903 ) | ( x95 & n33164 ) | ( ~n32903 & n33164 ) ;
  assign n33166 = ( x96 & ~n32895 ) | ( x96 & n33165 ) | ( ~n32895 & n33165 ) ;
  assign n33167 = ( x97 & ~n32887 ) | ( x97 & n33166 ) | ( ~n32887 & n33166 ) ;
  assign n33168 = ( x98 & ~n32879 ) | ( x98 & n33167 ) | ( ~n32879 & n33167 ) ;
  assign n33169 = ( x99 & ~n32871 ) | ( x99 & n33168 ) | ( ~n32871 & n33168 ) ;
  assign n33170 = ( x100 & ~n32863 ) | ( x100 & n33169 ) | ( ~n32863 & n33169 ) ;
  assign n33171 = ( x101 & ~n32855 ) | ( x101 & n33170 ) | ( ~n32855 & n33170 ) ;
  assign n33172 = ( x102 & ~n32847 ) | ( x102 & n33171 ) | ( ~n32847 & n33171 ) ;
  assign n33173 = ( x103 & ~n32839 ) | ( x103 & n33172 ) | ( ~n32839 & n33172 ) ;
  assign n33174 = ( x104 & ~n32831 ) | ( x104 & n33173 ) | ( ~n32831 & n33173 ) ;
  assign n33175 = ( x105 & ~n32823 ) | ( x105 & n33174 ) | ( ~n32823 & n33174 ) ;
  assign n33176 = ( x106 & ~n32815 ) | ( x106 & n33175 ) | ( ~n32815 & n33175 ) ;
  assign n33177 = ( x107 & ~n32807 ) | ( x107 & n33176 ) | ( ~n32807 & n33176 ) ;
  assign n33178 = ( x108 & ~n32799 ) | ( x108 & n33177 ) | ( ~n32799 & n33177 ) ;
  assign n33179 = ( x109 & ~n32791 ) | ( x109 & n33178 ) | ( ~n32791 & n33178 ) ;
  assign n33180 = ( x110 & ~n32783 ) | ( x110 & n33179 ) | ( ~n32783 & n33179 ) ;
  assign n33181 = ( x111 & ~n32775 ) | ( x111 & n33180 ) | ( ~n32775 & n33180 ) ;
  assign n33182 = ( x112 & ~n32767 ) | ( x112 & n33181 ) | ( ~n32767 & n33181 ) ;
  assign n33183 = ( x113 & ~n32759 ) | ( x113 & n33182 ) | ( ~n32759 & n33182 ) ;
  assign n33184 = ( x114 & ~n32751 ) | ( x114 & n33183 ) | ( ~n32751 & n33183 ) ;
  assign n33185 = ( x115 & ~n32743 ) | ( x115 & n33184 ) | ( ~n32743 & n33184 ) ;
  assign n33186 = ( x116 & ~n32735 ) | ( x116 & n33185 ) | ( ~n32735 & n33185 ) ;
  assign n33187 = ( x117 & ~n32727 ) | ( x117 & n33186 ) | ( ~n32727 & n33186 ) ;
  assign n33188 = ( x118 & ~n32719 ) | ( x118 & n33187 ) | ( ~n32719 & n33187 ) ;
  assign n33189 = ( x119 & ~n32711 ) | ( x119 & n33188 ) | ( ~n32711 & n33188 ) ;
  assign n33190 = ( x120 & ~n32701 ) | ( x120 & 1'b0 ) | ( ~n32701 & 1'b0 ) ;
  assign n33191 = ~n32699 & n33190 ;
  assign n33192 = ( n33189 & ~n32703 ) | ( n33189 & n33191 ) | ( ~n32703 & n33191 ) ;
  assign n33193 = ( n32703 & ~n239 ) | ( n32703 & n33192 ) | ( ~n239 & n33192 ) ;
  assign n33194 = n239 | n33193 ;
  assign n33201 = n269 &  n32702 ;
  assign n33202 = n33194 &  n33201 ;
  assign n33195 = ~n32702 |  n269 ;
  assign n33196 = n33194 &  n33195 ;
  assign n33200 = n32703 | n33191 ;
  assign n33204 = ( n33189 & n33196 ) | ( n33189 & n33200 ) | ( n33196 & n33200 ) ;
  assign n33203 = n33189 | n33200 ;
  assign n33205 = ( n33202 & ~n33204 ) | ( n33202 & n33203 ) | ( ~n33204 & n33203 ) ;
  assign n33209 = n32711 &  n33195 ;
  assign n33210 = n33194 &  n33209 ;
  assign n33197 = x119 | n32711 ;
  assign n33198 = x119 &  n32711 ;
  assign n33199 = ( n33197 & ~n33198 ) | ( n33197 & 1'b0 ) | ( ~n33198 & 1'b0 ) ;
  assign n33212 = ( n33188 & n33196 ) | ( n33188 & n33199 ) | ( n33196 & n33199 ) ;
  assign n33211 = n33188 | n33199 ;
  assign n33213 = ( n33210 & ~n33212 ) | ( n33210 & n33211 ) | ( ~n33212 & n33211 ) ;
  assign n33217 = n32719 &  n33195 ;
  assign n33218 = n33194 &  n33217 ;
  assign n33206 = x118 | n32719 ;
  assign n33207 = x118 &  n32719 ;
  assign n33208 = ( n33206 & ~n33207 ) | ( n33206 & 1'b0 ) | ( ~n33207 & 1'b0 ) ;
  assign n33220 = ( n33187 & n33196 ) | ( n33187 & n33208 ) | ( n33196 & n33208 ) ;
  assign n33219 = n33187 | n33208 ;
  assign n33221 = ( n33218 & ~n33220 ) | ( n33218 & n33219 ) | ( ~n33220 & n33219 ) ;
  assign n33225 = n32727 &  n33195 ;
  assign n33226 = n33194 &  n33225 ;
  assign n33214 = x117 | n32727 ;
  assign n33215 = x117 &  n32727 ;
  assign n33216 = ( n33214 & ~n33215 ) | ( n33214 & 1'b0 ) | ( ~n33215 & 1'b0 ) ;
  assign n33228 = ( n33186 & n33196 ) | ( n33186 & n33216 ) | ( n33196 & n33216 ) ;
  assign n33227 = n33186 | n33216 ;
  assign n33229 = ( n33226 & ~n33228 ) | ( n33226 & n33227 ) | ( ~n33228 & n33227 ) ;
  assign n33233 = n32735 &  n33195 ;
  assign n33234 = n33194 &  n33233 ;
  assign n33222 = x116 | n32735 ;
  assign n33223 = x116 &  n32735 ;
  assign n33224 = ( n33222 & ~n33223 ) | ( n33222 & 1'b0 ) | ( ~n33223 & 1'b0 ) ;
  assign n33236 = ( n33185 & n33196 ) | ( n33185 & n33224 ) | ( n33196 & n33224 ) ;
  assign n33235 = n33185 | n33224 ;
  assign n33237 = ( n33234 & ~n33236 ) | ( n33234 & n33235 ) | ( ~n33236 & n33235 ) ;
  assign n33241 = n32743 &  n33195 ;
  assign n33242 = n33194 &  n33241 ;
  assign n33230 = x115 | n32743 ;
  assign n33231 = x115 &  n32743 ;
  assign n33232 = ( n33230 & ~n33231 ) | ( n33230 & 1'b0 ) | ( ~n33231 & 1'b0 ) ;
  assign n33244 = ( n33184 & n33196 ) | ( n33184 & n33232 ) | ( n33196 & n33232 ) ;
  assign n33243 = n33184 | n33232 ;
  assign n33245 = ( n33242 & ~n33244 ) | ( n33242 & n33243 ) | ( ~n33244 & n33243 ) ;
  assign n33249 = n32751 &  n33195 ;
  assign n33250 = n33194 &  n33249 ;
  assign n33238 = x114 | n32751 ;
  assign n33239 = x114 &  n32751 ;
  assign n33240 = ( n33238 & ~n33239 ) | ( n33238 & 1'b0 ) | ( ~n33239 & 1'b0 ) ;
  assign n33252 = ( n33183 & n33196 ) | ( n33183 & n33240 ) | ( n33196 & n33240 ) ;
  assign n33251 = n33183 | n33240 ;
  assign n33253 = ( n33250 & ~n33252 ) | ( n33250 & n33251 ) | ( ~n33252 & n33251 ) ;
  assign n33257 = n32759 &  n33195 ;
  assign n33258 = n33194 &  n33257 ;
  assign n33246 = x113 | n32759 ;
  assign n33247 = x113 &  n32759 ;
  assign n33248 = ( n33246 & ~n33247 ) | ( n33246 & 1'b0 ) | ( ~n33247 & 1'b0 ) ;
  assign n33260 = ( n33182 & n33196 ) | ( n33182 & n33248 ) | ( n33196 & n33248 ) ;
  assign n33259 = n33182 | n33248 ;
  assign n33261 = ( n33258 & ~n33260 ) | ( n33258 & n33259 ) | ( ~n33260 & n33259 ) ;
  assign n33265 = n32767 &  n33195 ;
  assign n33266 = n33194 &  n33265 ;
  assign n33254 = x112 | n32767 ;
  assign n33255 = x112 &  n32767 ;
  assign n33256 = ( n33254 & ~n33255 ) | ( n33254 & 1'b0 ) | ( ~n33255 & 1'b0 ) ;
  assign n33268 = ( n33181 & n33196 ) | ( n33181 & n33256 ) | ( n33196 & n33256 ) ;
  assign n33267 = n33181 | n33256 ;
  assign n33269 = ( n33266 & ~n33268 ) | ( n33266 & n33267 ) | ( ~n33268 & n33267 ) ;
  assign n33273 = n32775 &  n33195 ;
  assign n33274 = n33194 &  n33273 ;
  assign n33262 = x111 | n32775 ;
  assign n33263 = x111 &  n32775 ;
  assign n33264 = ( n33262 & ~n33263 ) | ( n33262 & 1'b0 ) | ( ~n33263 & 1'b0 ) ;
  assign n33276 = ( n33180 & n33196 ) | ( n33180 & n33264 ) | ( n33196 & n33264 ) ;
  assign n33275 = n33180 | n33264 ;
  assign n33277 = ( n33274 & ~n33276 ) | ( n33274 & n33275 ) | ( ~n33276 & n33275 ) ;
  assign n33281 = n32783 &  n33195 ;
  assign n33282 = n33194 &  n33281 ;
  assign n33270 = x110 | n32783 ;
  assign n33271 = x110 &  n32783 ;
  assign n33272 = ( n33270 & ~n33271 ) | ( n33270 & 1'b0 ) | ( ~n33271 & 1'b0 ) ;
  assign n33284 = ( n33179 & n33196 ) | ( n33179 & n33272 ) | ( n33196 & n33272 ) ;
  assign n33283 = n33179 | n33272 ;
  assign n33285 = ( n33282 & ~n33284 ) | ( n33282 & n33283 ) | ( ~n33284 & n33283 ) ;
  assign n33289 = n32791 &  n33195 ;
  assign n33290 = n33194 &  n33289 ;
  assign n33278 = x109 | n32791 ;
  assign n33279 = x109 &  n32791 ;
  assign n33280 = ( n33278 & ~n33279 ) | ( n33278 & 1'b0 ) | ( ~n33279 & 1'b0 ) ;
  assign n33292 = ( n33178 & n33196 ) | ( n33178 & n33280 ) | ( n33196 & n33280 ) ;
  assign n33291 = n33178 | n33280 ;
  assign n33293 = ( n33290 & ~n33292 ) | ( n33290 & n33291 ) | ( ~n33292 & n33291 ) ;
  assign n33297 = n32799 &  n33195 ;
  assign n33298 = n33194 &  n33297 ;
  assign n33286 = x108 | n32799 ;
  assign n33287 = x108 &  n32799 ;
  assign n33288 = ( n33286 & ~n33287 ) | ( n33286 & 1'b0 ) | ( ~n33287 & 1'b0 ) ;
  assign n33300 = ( n33177 & n33196 ) | ( n33177 & n33288 ) | ( n33196 & n33288 ) ;
  assign n33299 = n33177 | n33288 ;
  assign n33301 = ( n33298 & ~n33300 ) | ( n33298 & n33299 ) | ( ~n33300 & n33299 ) ;
  assign n33305 = n32807 &  n33195 ;
  assign n33306 = n33194 &  n33305 ;
  assign n33294 = x107 | n32807 ;
  assign n33295 = x107 &  n32807 ;
  assign n33296 = ( n33294 & ~n33295 ) | ( n33294 & 1'b0 ) | ( ~n33295 & 1'b0 ) ;
  assign n33308 = ( n33176 & n33196 ) | ( n33176 & n33296 ) | ( n33196 & n33296 ) ;
  assign n33307 = n33176 | n33296 ;
  assign n33309 = ( n33306 & ~n33308 ) | ( n33306 & n33307 ) | ( ~n33308 & n33307 ) ;
  assign n33313 = n32815 &  n33195 ;
  assign n33314 = n33194 &  n33313 ;
  assign n33302 = x106 | n32815 ;
  assign n33303 = x106 &  n32815 ;
  assign n33304 = ( n33302 & ~n33303 ) | ( n33302 & 1'b0 ) | ( ~n33303 & 1'b0 ) ;
  assign n33316 = ( n33175 & n33196 ) | ( n33175 & n33304 ) | ( n33196 & n33304 ) ;
  assign n33315 = n33175 | n33304 ;
  assign n33317 = ( n33314 & ~n33316 ) | ( n33314 & n33315 ) | ( ~n33316 & n33315 ) ;
  assign n33321 = n32823 &  n33195 ;
  assign n33322 = n33194 &  n33321 ;
  assign n33310 = x105 | n32823 ;
  assign n33311 = x105 &  n32823 ;
  assign n33312 = ( n33310 & ~n33311 ) | ( n33310 & 1'b0 ) | ( ~n33311 & 1'b0 ) ;
  assign n33324 = ( n33174 & n33196 ) | ( n33174 & n33312 ) | ( n33196 & n33312 ) ;
  assign n33323 = n33174 | n33312 ;
  assign n33325 = ( n33322 & ~n33324 ) | ( n33322 & n33323 ) | ( ~n33324 & n33323 ) ;
  assign n33329 = n32831 &  n33195 ;
  assign n33330 = n33194 &  n33329 ;
  assign n33318 = x104 | n32831 ;
  assign n33319 = x104 &  n32831 ;
  assign n33320 = ( n33318 & ~n33319 ) | ( n33318 & 1'b0 ) | ( ~n33319 & 1'b0 ) ;
  assign n33332 = ( n33173 & n33196 ) | ( n33173 & n33320 ) | ( n33196 & n33320 ) ;
  assign n33331 = n33173 | n33320 ;
  assign n33333 = ( n33330 & ~n33332 ) | ( n33330 & n33331 ) | ( ~n33332 & n33331 ) ;
  assign n33337 = n32839 &  n33195 ;
  assign n33338 = n33194 &  n33337 ;
  assign n33326 = x103 | n32839 ;
  assign n33327 = x103 &  n32839 ;
  assign n33328 = ( n33326 & ~n33327 ) | ( n33326 & 1'b0 ) | ( ~n33327 & 1'b0 ) ;
  assign n33340 = ( n33172 & n33196 ) | ( n33172 & n33328 ) | ( n33196 & n33328 ) ;
  assign n33339 = n33172 | n33328 ;
  assign n33341 = ( n33338 & ~n33340 ) | ( n33338 & n33339 ) | ( ~n33340 & n33339 ) ;
  assign n33345 = n32847 &  n33195 ;
  assign n33346 = n33194 &  n33345 ;
  assign n33334 = x102 | n32847 ;
  assign n33335 = x102 &  n32847 ;
  assign n33336 = ( n33334 & ~n33335 ) | ( n33334 & 1'b0 ) | ( ~n33335 & 1'b0 ) ;
  assign n33348 = ( n33171 & n33196 ) | ( n33171 & n33336 ) | ( n33196 & n33336 ) ;
  assign n33347 = n33171 | n33336 ;
  assign n33349 = ( n33346 & ~n33348 ) | ( n33346 & n33347 ) | ( ~n33348 & n33347 ) ;
  assign n33353 = n32855 &  n33195 ;
  assign n33354 = n33194 &  n33353 ;
  assign n33342 = x101 | n32855 ;
  assign n33343 = x101 &  n32855 ;
  assign n33344 = ( n33342 & ~n33343 ) | ( n33342 & 1'b0 ) | ( ~n33343 & 1'b0 ) ;
  assign n33356 = ( n33170 & n33196 ) | ( n33170 & n33344 ) | ( n33196 & n33344 ) ;
  assign n33355 = n33170 | n33344 ;
  assign n33357 = ( n33354 & ~n33356 ) | ( n33354 & n33355 ) | ( ~n33356 & n33355 ) ;
  assign n33361 = n32863 &  n33195 ;
  assign n33362 = n33194 &  n33361 ;
  assign n33350 = x100 | n32863 ;
  assign n33351 = x100 &  n32863 ;
  assign n33352 = ( n33350 & ~n33351 ) | ( n33350 & 1'b0 ) | ( ~n33351 & 1'b0 ) ;
  assign n33364 = ( n33169 & n33196 ) | ( n33169 & n33352 ) | ( n33196 & n33352 ) ;
  assign n33363 = n33169 | n33352 ;
  assign n33365 = ( n33362 & ~n33364 ) | ( n33362 & n33363 ) | ( ~n33364 & n33363 ) ;
  assign n33369 = n32871 &  n33195 ;
  assign n33370 = n33194 &  n33369 ;
  assign n33358 = x99 | n32871 ;
  assign n33359 = x99 &  n32871 ;
  assign n33360 = ( n33358 & ~n33359 ) | ( n33358 & 1'b0 ) | ( ~n33359 & 1'b0 ) ;
  assign n33372 = ( n33168 & n33196 ) | ( n33168 & n33360 ) | ( n33196 & n33360 ) ;
  assign n33371 = n33168 | n33360 ;
  assign n33373 = ( n33370 & ~n33372 ) | ( n33370 & n33371 ) | ( ~n33372 & n33371 ) ;
  assign n33377 = n32879 &  n33195 ;
  assign n33378 = n33194 &  n33377 ;
  assign n33366 = x98 | n32879 ;
  assign n33367 = x98 &  n32879 ;
  assign n33368 = ( n33366 & ~n33367 ) | ( n33366 & 1'b0 ) | ( ~n33367 & 1'b0 ) ;
  assign n33380 = ( n33167 & n33196 ) | ( n33167 & n33368 ) | ( n33196 & n33368 ) ;
  assign n33379 = n33167 | n33368 ;
  assign n33381 = ( n33378 & ~n33380 ) | ( n33378 & n33379 ) | ( ~n33380 & n33379 ) ;
  assign n33385 = n32887 &  n33195 ;
  assign n33386 = n33194 &  n33385 ;
  assign n33374 = x97 | n32887 ;
  assign n33375 = x97 &  n32887 ;
  assign n33376 = ( n33374 & ~n33375 ) | ( n33374 & 1'b0 ) | ( ~n33375 & 1'b0 ) ;
  assign n33388 = ( n33166 & n33196 ) | ( n33166 & n33376 ) | ( n33196 & n33376 ) ;
  assign n33387 = n33166 | n33376 ;
  assign n33389 = ( n33386 & ~n33388 ) | ( n33386 & n33387 ) | ( ~n33388 & n33387 ) ;
  assign n33393 = n32895 &  n33195 ;
  assign n33394 = n33194 &  n33393 ;
  assign n33382 = x96 | n32895 ;
  assign n33383 = x96 &  n32895 ;
  assign n33384 = ( n33382 & ~n33383 ) | ( n33382 & 1'b0 ) | ( ~n33383 & 1'b0 ) ;
  assign n33396 = ( n33165 & n33196 ) | ( n33165 & n33384 ) | ( n33196 & n33384 ) ;
  assign n33395 = n33165 | n33384 ;
  assign n33397 = ( n33394 & ~n33396 ) | ( n33394 & n33395 ) | ( ~n33396 & n33395 ) ;
  assign n33401 = n32903 &  n33195 ;
  assign n33402 = n33194 &  n33401 ;
  assign n33390 = x95 | n32903 ;
  assign n33391 = x95 &  n32903 ;
  assign n33392 = ( n33390 & ~n33391 ) | ( n33390 & 1'b0 ) | ( ~n33391 & 1'b0 ) ;
  assign n33404 = ( n33164 & n33196 ) | ( n33164 & n33392 ) | ( n33196 & n33392 ) ;
  assign n33403 = n33164 | n33392 ;
  assign n33405 = ( n33402 & ~n33404 ) | ( n33402 & n33403 ) | ( ~n33404 & n33403 ) ;
  assign n33409 = n32911 &  n33195 ;
  assign n33410 = n33194 &  n33409 ;
  assign n33398 = x94 | n32911 ;
  assign n33399 = x94 &  n32911 ;
  assign n33400 = ( n33398 & ~n33399 ) | ( n33398 & 1'b0 ) | ( ~n33399 & 1'b0 ) ;
  assign n33412 = ( n33163 & n33196 ) | ( n33163 & n33400 ) | ( n33196 & n33400 ) ;
  assign n33411 = n33163 | n33400 ;
  assign n33413 = ( n33410 & ~n33412 ) | ( n33410 & n33411 ) | ( ~n33412 & n33411 ) ;
  assign n33417 = n32919 &  n33195 ;
  assign n33418 = n33194 &  n33417 ;
  assign n33406 = x93 | n32919 ;
  assign n33407 = x93 &  n32919 ;
  assign n33408 = ( n33406 & ~n33407 ) | ( n33406 & 1'b0 ) | ( ~n33407 & 1'b0 ) ;
  assign n33420 = ( n33162 & n33196 ) | ( n33162 & n33408 ) | ( n33196 & n33408 ) ;
  assign n33419 = n33162 | n33408 ;
  assign n33421 = ( n33418 & ~n33420 ) | ( n33418 & n33419 ) | ( ~n33420 & n33419 ) ;
  assign n33425 = n32927 &  n33195 ;
  assign n33426 = n33194 &  n33425 ;
  assign n33414 = x92 | n32927 ;
  assign n33415 = x92 &  n32927 ;
  assign n33416 = ( n33414 & ~n33415 ) | ( n33414 & 1'b0 ) | ( ~n33415 & 1'b0 ) ;
  assign n33428 = ( n33161 & n33196 ) | ( n33161 & n33416 ) | ( n33196 & n33416 ) ;
  assign n33427 = n33161 | n33416 ;
  assign n33429 = ( n33426 & ~n33428 ) | ( n33426 & n33427 ) | ( ~n33428 & n33427 ) ;
  assign n33433 = n32935 &  n33195 ;
  assign n33434 = n33194 &  n33433 ;
  assign n33422 = x91 | n32935 ;
  assign n33423 = x91 &  n32935 ;
  assign n33424 = ( n33422 & ~n33423 ) | ( n33422 & 1'b0 ) | ( ~n33423 & 1'b0 ) ;
  assign n33436 = ( n33160 & n33196 ) | ( n33160 & n33424 ) | ( n33196 & n33424 ) ;
  assign n33435 = n33160 | n33424 ;
  assign n33437 = ( n33434 & ~n33436 ) | ( n33434 & n33435 ) | ( ~n33436 & n33435 ) ;
  assign n33441 = n32943 &  n33195 ;
  assign n33442 = n33194 &  n33441 ;
  assign n33430 = x90 | n32943 ;
  assign n33431 = x90 &  n32943 ;
  assign n33432 = ( n33430 & ~n33431 ) | ( n33430 & 1'b0 ) | ( ~n33431 & 1'b0 ) ;
  assign n33444 = ( n33159 & n33196 ) | ( n33159 & n33432 ) | ( n33196 & n33432 ) ;
  assign n33443 = n33159 | n33432 ;
  assign n33445 = ( n33442 & ~n33444 ) | ( n33442 & n33443 ) | ( ~n33444 & n33443 ) ;
  assign n33449 = n32951 &  n33195 ;
  assign n33450 = n33194 &  n33449 ;
  assign n33438 = x89 | n32951 ;
  assign n33439 = x89 &  n32951 ;
  assign n33440 = ( n33438 & ~n33439 ) | ( n33438 & 1'b0 ) | ( ~n33439 & 1'b0 ) ;
  assign n33452 = ( n33158 & n33196 ) | ( n33158 & n33440 ) | ( n33196 & n33440 ) ;
  assign n33451 = n33158 | n33440 ;
  assign n33453 = ( n33450 & ~n33452 ) | ( n33450 & n33451 ) | ( ~n33452 & n33451 ) ;
  assign n33457 = n32959 &  n33195 ;
  assign n33458 = n33194 &  n33457 ;
  assign n33446 = x88 | n32959 ;
  assign n33447 = x88 &  n32959 ;
  assign n33448 = ( n33446 & ~n33447 ) | ( n33446 & 1'b0 ) | ( ~n33447 & 1'b0 ) ;
  assign n33460 = ( n33157 & n33196 ) | ( n33157 & n33448 ) | ( n33196 & n33448 ) ;
  assign n33459 = n33157 | n33448 ;
  assign n33461 = ( n33458 & ~n33460 ) | ( n33458 & n33459 ) | ( ~n33460 & n33459 ) ;
  assign n33465 = n32967 &  n33195 ;
  assign n33466 = n33194 &  n33465 ;
  assign n33454 = x87 | n32967 ;
  assign n33455 = x87 &  n32967 ;
  assign n33456 = ( n33454 & ~n33455 ) | ( n33454 & 1'b0 ) | ( ~n33455 & 1'b0 ) ;
  assign n33468 = ( n33156 & n33196 ) | ( n33156 & n33456 ) | ( n33196 & n33456 ) ;
  assign n33467 = n33156 | n33456 ;
  assign n33469 = ( n33466 & ~n33468 ) | ( n33466 & n33467 ) | ( ~n33468 & n33467 ) ;
  assign n33473 = n32975 &  n33195 ;
  assign n33474 = n33194 &  n33473 ;
  assign n33462 = x86 | n32975 ;
  assign n33463 = x86 &  n32975 ;
  assign n33464 = ( n33462 & ~n33463 ) | ( n33462 & 1'b0 ) | ( ~n33463 & 1'b0 ) ;
  assign n33476 = ( n33155 & n33196 ) | ( n33155 & n33464 ) | ( n33196 & n33464 ) ;
  assign n33475 = n33155 | n33464 ;
  assign n33477 = ( n33474 & ~n33476 ) | ( n33474 & n33475 ) | ( ~n33476 & n33475 ) ;
  assign n33481 = n32983 &  n33195 ;
  assign n33482 = n33194 &  n33481 ;
  assign n33470 = x85 | n32983 ;
  assign n33471 = x85 &  n32983 ;
  assign n33472 = ( n33470 & ~n33471 ) | ( n33470 & 1'b0 ) | ( ~n33471 & 1'b0 ) ;
  assign n33484 = ( n33154 & n33196 ) | ( n33154 & n33472 ) | ( n33196 & n33472 ) ;
  assign n33483 = n33154 | n33472 ;
  assign n33485 = ( n33482 & ~n33484 ) | ( n33482 & n33483 ) | ( ~n33484 & n33483 ) ;
  assign n33489 = n32991 &  n33195 ;
  assign n33490 = n33194 &  n33489 ;
  assign n33478 = x84 | n32991 ;
  assign n33479 = x84 &  n32991 ;
  assign n33480 = ( n33478 & ~n33479 ) | ( n33478 & 1'b0 ) | ( ~n33479 & 1'b0 ) ;
  assign n33492 = ( n33153 & n33196 ) | ( n33153 & n33480 ) | ( n33196 & n33480 ) ;
  assign n33491 = n33153 | n33480 ;
  assign n33493 = ( n33490 & ~n33492 ) | ( n33490 & n33491 ) | ( ~n33492 & n33491 ) ;
  assign n33497 = n32999 &  n33195 ;
  assign n33498 = n33194 &  n33497 ;
  assign n33486 = x83 | n32999 ;
  assign n33487 = x83 &  n32999 ;
  assign n33488 = ( n33486 & ~n33487 ) | ( n33486 & 1'b0 ) | ( ~n33487 & 1'b0 ) ;
  assign n33500 = ( n33152 & n33196 ) | ( n33152 & n33488 ) | ( n33196 & n33488 ) ;
  assign n33499 = n33152 | n33488 ;
  assign n33501 = ( n33498 & ~n33500 ) | ( n33498 & n33499 ) | ( ~n33500 & n33499 ) ;
  assign n33505 = n33007 &  n33195 ;
  assign n33506 = n33194 &  n33505 ;
  assign n33494 = x82 | n33007 ;
  assign n33495 = x82 &  n33007 ;
  assign n33496 = ( n33494 & ~n33495 ) | ( n33494 & 1'b0 ) | ( ~n33495 & 1'b0 ) ;
  assign n33508 = ( n33151 & n33196 ) | ( n33151 & n33496 ) | ( n33196 & n33496 ) ;
  assign n33507 = n33151 | n33496 ;
  assign n33509 = ( n33506 & ~n33508 ) | ( n33506 & n33507 ) | ( ~n33508 & n33507 ) ;
  assign n33513 = n33015 &  n33195 ;
  assign n33514 = n33194 &  n33513 ;
  assign n33502 = x81 | n33015 ;
  assign n33503 = x81 &  n33015 ;
  assign n33504 = ( n33502 & ~n33503 ) | ( n33502 & 1'b0 ) | ( ~n33503 & 1'b0 ) ;
  assign n33516 = ( n33150 & n33196 ) | ( n33150 & n33504 ) | ( n33196 & n33504 ) ;
  assign n33515 = n33150 | n33504 ;
  assign n33517 = ( n33514 & ~n33516 ) | ( n33514 & n33515 ) | ( ~n33516 & n33515 ) ;
  assign n33521 = n33023 &  n33195 ;
  assign n33522 = n33194 &  n33521 ;
  assign n33510 = x80 | n33023 ;
  assign n33511 = x80 &  n33023 ;
  assign n33512 = ( n33510 & ~n33511 ) | ( n33510 & 1'b0 ) | ( ~n33511 & 1'b0 ) ;
  assign n33524 = ( n33149 & n33196 ) | ( n33149 & n33512 ) | ( n33196 & n33512 ) ;
  assign n33523 = n33149 | n33512 ;
  assign n33525 = ( n33522 & ~n33524 ) | ( n33522 & n33523 ) | ( ~n33524 & n33523 ) ;
  assign n33529 = n33031 &  n33195 ;
  assign n33530 = n33194 &  n33529 ;
  assign n33518 = x79 | n33031 ;
  assign n33519 = x79 &  n33031 ;
  assign n33520 = ( n33518 & ~n33519 ) | ( n33518 & 1'b0 ) | ( ~n33519 & 1'b0 ) ;
  assign n33532 = ( n33148 & n33196 ) | ( n33148 & n33520 ) | ( n33196 & n33520 ) ;
  assign n33531 = n33148 | n33520 ;
  assign n33533 = ( n33530 & ~n33532 ) | ( n33530 & n33531 ) | ( ~n33532 & n33531 ) ;
  assign n33537 = n33039 &  n33195 ;
  assign n33538 = n33194 &  n33537 ;
  assign n33526 = x78 | n33039 ;
  assign n33527 = x78 &  n33039 ;
  assign n33528 = ( n33526 & ~n33527 ) | ( n33526 & 1'b0 ) | ( ~n33527 & 1'b0 ) ;
  assign n33540 = ( n33147 & n33196 ) | ( n33147 & n33528 ) | ( n33196 & n33528 ) ;
  assign n33539 = n33147 | n33528 ;
  assign n33541 = ( n33538 & ~n33540 ) | ( n33538 & n33539 ) | ( ~n33540 & n33539 ) ;
  assign n33545 = n33047 &  n33195 ;
  assign n33546 = n33194 &  n33545 ;
  assign n33534 = x77 | n33047 ;
  assign n33535 = x77 &  n33047 ;
  assign n33536 = ( n33534 & ~n33535 ) | ( n33534 & 1'b0 ) | ( ~n33535 & 1'b0 ) ;
  assign n33548 = ( n33146 & n33196 ) | ( n33146 & n33536 ) | ( n33196 & n33536 ) ;
  assign n33547 = n33146 | n33536 ;
  assign n33549 = ( n33546 & ~n33548 ) | ( n33546 & n33547 ) | ( ~n33548 & n33547 ) ;
  assign n33553 = n33055 &  n33195 ;
  assign n33554 = n33194 &  n33553 ;
  assign n33542 = x76 | n33055 ;
  assign n33543 = x76 &  n33055 ;
  assign n33544 = ( n33542 & ~n33543 ) | ( n33542 & 1'b0 ) | ( ~n33543 & 1'b0 ) ;
  assign n33556 = ( n33145 & n33196 ) | ( n33145 & n33544 ) | ( n33196 & n33544 ) ;
  assign n33555 = n33145 | n33544 ;
  assign n33557 = ( n33554 & ~n33556 ) | ( n33554 & n33555 ) | ( ~n33556 & n33555 ) ;
  assign n33561 = n33063 &  n33195 ;
  assign n33562 = n33194 &  n33561 ;
  assign n33550 = x75 | n33063 ;
  assign n33551 = x75 &  n33063 ;
  assign n33552 = ( n33550 & ~n33551 ) | ( n33550 & 1'b0 ) | ( ~n33551 & 1'b0 ) ;
  assign n33564 = ( n33144 & n33196 ) | ( n33144 & n33552 ) | ( n33196 & n33552 ) ;
  assign n33563 = n33144 | n33552 ;
  assign n33565 = ( n33562 & ~n33564 ) | ( n33562 & n33563 ) | ( ~n33564 & n33563 ) ;
  assign n33569 = n33071 &  n33195 ;
  assign n33570 = n33194 &  n33569 ;
  assign n33558 = x74 | n33071 ;
  assign n33559 = x74 &  n33071 ;
  assign n33560 = ( n33558 & ~n33559 ) | ( n33558 & 1'b0 ) | ( ~n33559 & 1'b0 ) ;
  assign n33572 = ( n33143 & n33196 ) | ( n33143 & n33560 ) | ( n33196 & n33560 ) ;
  assign n33571 = n33143 | n33560 ;
  assign n33573 = ( n33570 & ~n33572 ) | ( n33570 & n33571 ) | ( ~n33572 & n33571 ) ;
  assign n33577 = n33079 &  n33195 ;
  assign n33578 = n33194 &  n33577 ;
  assign n33566 = x73 | n33079 ;
  assign n33567 = x73 &  n33079 ;
  assign n33568 = ( n33566 & ~n33567 ) | ( n33566 & 1'b0 ) | ( ~n33567 & 1'b0 ) ;
  assign n33580 = ( n33142 & n33196 ) | ( n33142 & n33568 ) | ( n33196 & n33568 ) ;
  assign n33579 = n33142 | n33568 ;
  assign n33581 = ( n33578 & ~n33580 ) | ( n33578 & n33579 ) | ( ~n33580 & n33579 ) ;
  assign n33585 = n33087 &  n33195 ;
  assign n33586 = n33194 &  n33585 ;
  assign n33574 = x72 | n33087 ;
  assign n33575 = x72 &  n33087 ;
  assign n33576 = ( n33574 & ~n33575 ) | ( n33574 & 1'b0 ) | ( ~n33575 & 1'b0 ) ;
  assign n33588 = ( n33141 & n33196 ) | ( n33141 & n33576 ) | ( n33196 & n33576 ) ;
  assign n33587 = n33141 | n33576 ;
  assign n33589 = ( n33586 & ~n33588 ) | ( n33586 & n33587 ) | ( ~n33588 & n33587 ) ;
  assign n33593 = n33095 &  n33195 ;
  assign n33594 = n33194 &  n33593 ;
  assign n33582 = x71 | n33095 ;
  assign n33583 = x71 &  n33095 ;
  assign n33584 = ( n33582 & ~n33583 ) | ( n33582 & 1'b0 ) | ( ~n33583 & 1'b0 ) ;
  assign n33596 = ( n33140 & n33196 ) | ( n33140 & n33584 ) | ( n33196 & n33584 ) ;
  assign n33595 = n33140 | n33584 ;
  assign n33597 = ( n33594 & ~n33596 ) | ( n33594 & n33595 ) | ( ~n33596 & n33595 ) ;
  assign n33601 = n33103 &  n33195 ;
  assign n33602 = n33194 &  n33601 ;
  assign n33590 = x70 | n33103 ;
  assign n33591 = x70 &  n33103 ;
  assign n33592 = ( n33590 & ~n33591 ) | ( n33590 & 1'b0 ) | ( ~n33591 & 1'b0 ) ;
  assign n33604 = ( n33139 & n33196 ) | ( n33139 & n33592 ) | ( n33196 & n33592 ) ;
  assign n33603 = n33139 | n33592 ;
  assign n33605 = ( n33602 & ~n33604 ) | ( n33602 & n33603 ) | ( ~n33604 & n33603 ) ;
  assign n33609 = n33111 &  n33195 ;
  assign n33610 = n33194 &  n33609 ;
  assign n33598 = x69 | n33111 ;
  assign n33599 = x69 &  n33111 ;
  assign n33600 = ( n33598 & ~n33599 ) | ( n33598 & 1'b0 ) | ( ~n33599 & 1'b0 ) ;
  assign n33612 = ( n33138 & n33196 ) | ( n33138 & n33600 ) | ( n33196 & n33600 ) ;
  assign n33611 = n33138 | n33600 ;
  assign n33613 = ( n33610 & ~n33612 ) | ( n33610 & n33611 ) | ( ~n33612 & n33611 ) ;
  assign n33617 = n33119 &  n33195 ;
  assign n33618 = n33194 &  n33617 ;
  assign n33606 = x68 | n33119 ;
  assign n33607 = x68 &  n33119 ;
  assign n33608 = ( n33606 & ~n33607 ) | ( n33606 & 1'b0 ) | ( ~n33607 & 1'b0 ) ;
  assign n33620 = ( n33137 & n33196 ) | ( n33137 & n33608 ) | ( n33196 & n33608 ) ;
  assign n33619 = n33137 | n33608 ;
  assign n33621 = ( n33618 & ~n33620 ) | ( n33618 & n33619 ) | ( ~n33620 & n33619 ) ;
  assign n33625 = n33124 &  n33195 ;
  assign n33626 = n33194 &  n33625 ;
  assign n33614 = x67 | n33124 ;
  assign n33615 = x67 &  n33124 ;
  assign n33616 = ( n33614 & ~n33615 ) | ( n33614 & 1'b0 ) | ( ~n33615 & 1'b0 ) ;
  assign n33628 = ( n33136 & n33196 ) | ( n33136 & n33616 ) | ( n33196 & n33616 ) ;
  assign n33627 = n33136 | n33616 ;
  assign n33629 = ( n33626 & ~n33628 ) | ( n33626 & n33627 ) | ( ~n33628 & n33627 ) ;
  assign n33630 = n33130 &  n33195 ;
  assign n33631 = n33194 &  n33630 ;
  assign n33622 = x66 | n33130 ;
  assign n33623 = x66 &  n33130 ;
  assign n33624 = ( n33622 & ~n33623 ) | ( n33622 & 1'b0 ) | ( ~n33623 & 1'b0 ) ;
  assign n33632 = n33135 &  n33624 ;
  assign n33633 = ( n33135 & ~n33196 ) | ( n33135 & n33624 ) | ( ~n33196 & n33624 ) ;
  assign n33634 = ( n33631 & ~n33632 ) | ( n33631 & n33633 ) | ( ~n33632 & n33633 ) ;
  assign n33635 = ( x65 & ~n14798 ) | ( x65 & n33134 ) | ( ~n14798 & n33134 ) ;
  assign n33636 = ( n33135 & ~x65 ) | ( n33135 & n33635 ) | ( ~x65 & n33635 ) ;
  assign n33637 = ~n33196 & n33636 ;
  assign n33638 = n33134 &  n33195 ;
  assign n33639 = n33194 &  n33638 ;
  assign n33640 = n33637 | n33639 ;
  assign n33641 = ( x64 & ~n33196 ) | ( x64 & 1'b0 ) | ( ~n33196 & 1'b0 ) ;
  assign n33642 = ( x7 & ~n33641 ) | ( x7 & 1'b0 ) | ( ~n33641 & 1'b0 ) ;
  assign n33643 = ( n14798 & ~n33196 ) | ( n14798 & 1'b0 ) | ( ~n33196 & 1'b0 ) ;
  assign n33644 = n33642 | n33643 ;
  assign n33645 = ( x65 & ~n33644 ) | ( x65 & n15357 ) | ( ~n33644 & n15357 ) ;
  assign n33646 = ( x66 & ~n33640 ) | ( x66 & n33645 ) | ( ~n33640 & n33645 ) ;
  assign n33647 = ( x67 & ~n33634 ) | ( x67 & n33646 ) | ( ~n33634 & n33646 ) ;
  assign n33648 = ( x68 & ~n33629 ) | ( x68 & n33647 ) | ( ~n33629 & n33647 ) ;
  assign n33649 = ( x69 & ~n33621 ) | ( x69 & n33648 ) | ( ~n33621 & n33648 ) ;
  assign n33650 = ( x70 & ~n33613 ) | ( x70 & n33649 ) | ( ~n33613 & n33649 ) ;
  assign n33651 = ( x71 & ~n33605 ) | ( x71 & n33650 ) | ( ~n33605 & n33650 ) ;
  assign n33652 = ( x72 & ~n33597 ) | ( x72 & n33651 ) | ( ~n33597 & n33651 ) ;
  assign n33653 = ( x73 & ~n33589 ) | ( x73 & n33652 ) | ( ~n33589 & n33652 ) ;
  assign n33654 = ( x74 & ~n33581 ) | ( x74 & n33653 ) | ( ~n33581 & n33653 ) ;
  assign n33655 = ( x75 & ~n33573 ) | ( x75 & n33654 ) | ( ~n33573 & n33654 ) ;
  assign n33656 = ( x76 & ~n33565 ) | ( x76 & n33655 ) | ( ~n33565 & n33655 ) ;
  assign n33657 = ( x77 & ~n33557 ) | ( x77 & n33656 ) | ( ~n33557 & n33656 ) ;
  assign n33658 = ( x78 & ~n33549 ) | ( x78 & n33657 ) | ( ~n33549 & n33657 ) ;
  assign n33659 = ( x79 & ~n33541 ) | ( x79 & n33658 ) | ( ~n33541 & n33658 ) ;
  assign n33660 = ( x80 & ~n33533 ) | ( x80 & n33659 ) | ( ~n33533 & n33659 ) ;
  assign n33661 = ( x81 & ~n33525 ) | ( x81 & n33660 ) | ( ~n33525 & n33660 ) ;
  assign n33662 = ( x82 & ~n33517 ) | ( x82 & n33661 ) | ( ~n33517 & n33661 ) ;
  assign n33663 = ( x83 & ~n33509 ) | ( x83 & n33662 ) | ( ~n33509 & n33662 ) ;
  assign n33664 = ( x84 & ~n33501 ) | ( x84 & n33663 ) | ( ~n33501 & n33663 ) ;
  assign n33665 = ( x85 & ~n33493 ) | ( x85 & n33664 ) | ( ~n33493 & n33664 ) ;
  assign n33666 = ( x86 & ~n33485 ) | ( x86 & n33665 ) | ( ~n33485 & n33665 ) ;
  assign n33667 = ( x87 & ~n33477 ) | ( x87 & n33666 ) | ( ~n33477 & n33666 ) ;
  assign n33668 = ( x88 & ~n33469 ) | ( x88 & n33667 ) | ( ~n33469 & n33667 ) ;
  assign n33669 = ( x89 & ~n33461 ) | ( x89 & n33668 ) | ( ~n33461 & n33668 ) ;
  assign n33670 = ( x90 & ~n33453 ) | ( x90 & n33669 ) | ( ~n33453 & n33669 ) ;
  assign n33671 = ( x91 & ~n33445 ) | ( x91 & n33670 ) | ( ~n33445 & n33670 ) ;
  assign n33672 = ( x92 & ~n33437 ) | ( x92 & n33671 ) | ( ~n33437 & n33671 ) ;
  assign n33673 = ( x93 & ~n33429 ) | ( x93 & n33672 ) | ( ~n33429 & n33672 ) ;
  assign n33674 = ( x94 & ~n33421 ) | ( x94 & n33673 ) | ( ~n33421 & n33673 ) ;
  assign n33675 = ( x95 & ~n33413 ) | ( x95 & n33674 ) | ( ~n33413 & n33674 ) ;
  assign n33676 = ( x96 & ~n33405 ) | ( x96 & n33675 ) | ( ~n33405 & n33675 ) ;
  assign n33677 = ( x97 & ~n33397 ) | ( x97 & n33676 ) | ( ~n33397 & n33676 ) ;
  assign n33678 = ( x98 & ~n33389 ) | ( x98 & n33677 ) | ( ~n33389 & n33677 ) ;
  assign n33679 = ( x99 & ~n33381 ) | ( x99 & n33678 ) | ( ~n33381 & n33678 ) ;
  assign n33680 = ( x100 & ~n33373 ) | ( x100 & n33679 ) | ( ~n33373 & n33679 ) ;
  assign n33681 = ( x101 & ~n33365 ) | ( x101 & n33680 ) | ( ~n33365 & n33680 ) ;
  assign n33682 = ( x102 & ~n33357 ) | ( x102 & n33681 ) | ( ~n33357 & n33681 ) ;
  assign n33683 = ( x103 & ~n33349 ) | ( x103 & n33682 ) | ( ~n33349 & n33682 ) ;
  assign n33684 = ( x104 & ~n33341 ) | ( x104 & n33683 ) | ( ~n33341 & n33683 ) ;
  assign n33685 = ( x105 & ~n33333 ) | ( x105 & n33684 ) | ( ~n33333 & n33684 ) ;
  assign n33686 = ( x106 & ~n33325 ) | ( x106 & n33685 ) | ( ~n33325 & n33685 ) ;
  assign n33687 = ( x107 & ~n33317 ) | ( x107 & n33686 ) | ( ~n33317 & n33686 ) ;
  assign n33688 = ( x108 & ~n33309 ) | ( x108 & n33687 ) | ( ~n33309 & n33687 ) ;
  assign n33689 = ( x109 & ~n33301 ) | ( x109 & n33688 ) | ( ~n33301 & n33688 ) ;
  assign n33690 = ( x110 & ~n33293 ) | ( x110 & n33689 ) | ( ~n33293 & n33689 ) ;
  assign n33691 = ( x111 & ~n33285 ) | ( x111 & n33690 ) | ( ~n33285 & n33690 ) ;
  assign n33692 = ( x112 & ~n33277 ) | ( x112 & n33691 ) | ( ~n33277 & n33691 ) ;
  assign n33693 = ( x113 & ~n33269 ) | ( x113 & n33692 ) | ( ~n33269 & n33692 ) ;
  assign n33694 = ( x114 & ~n33261 ) | ( x114 & n33693 ) | ( ~n33261 & n33693 ) ;
  assign n33695 = ( x115 & ~n33253 ) | ( x115 & n33694 ) | ( ~n33253 & n33694 ) ;
  assign n33696 = ( x116 & ~n33245 ) | ( x116 & n33695 ) | ( ~n33245 & n33695 ) ;
  assign n33697 = ( x117 & ~n33237 ) | ( x117 & n33696 ) | ( ~n33237 & n33696 ) ;
  assign n33698 = ( x118 & ~n33229 ) | ( x118 & n33697 ) | ( ~n33229 & n33697 ) ;
  assign n33699 = ( x119 & ~n33221 ) | ( x119 & n33698 ) | ( ~n33221 & n33698 ) ;
  assign n33700 = ( x120 & ~n33213 ) | ( x120 & n33699 ) | ( ~n33213 & n33699 ) ;
  assign n33701 = ( x121 & ~n33205 ) | ( x121 & n33700 ) | ( ~n33205 & n33700 ) ;
  assign n33702 = n15415 | n33701 ;
  assign n33703 = n33205 &  n33702 ;
  assign n33707 = ( n15415 & n33205 ) | ( n15415 & n33700 ) | ( n33205 & n33700 ) ;
  assign n33708 = ( x121 & ~n33707 ) | ( x121 & n33205 ) | ( ~n33707 & n33205 ) ;
  assign n33709 = ~x121 & n33708 ;
  assign n33710 = n33703 | n33709 ;
  assign n33711 = ~x122 & n33710 ;
  assign n33712 = n33213 &  n33702 ;
  assign n33704 = x120 | n33213 ;
  assign n33705 = x120 &  n33213 ;
  assign n33706 = ( n33704 & ~n33705 ) | ( n33704 & 1'b0 ) | ( ~n33705 & 1'b0 ) ;
  assign n33716 = ( n15415 & n33699 ) | ( n15415 & n33706 ) | ( n33699 & n33706 ) ;
  assign n33717 = ( n33699 & ~n33701 ) | ( n33699 & n33706 ) | ( ~n33701 & n33706 ) ;
  assign n33718 = ~n33716 & n33717 ;
  assign n33719 = n33712 | n33718 ;
  assign n33720 = n33221 &  n33702 ;
  assign n33713 = x119 | n33221 ;
  assign n33714 = x119 &  n33221 ;
  assign n33715 = ( n33713 & ~n33714 ) | ( n33713 & 1'b0 ) | ( ~n33714 & 1'b0 ) ;
  assign n33724 = ( n15415 & n33698 ) | ( n15415 & n33715 ) | ( n33698 & n33715 ) ;
  assign n33725 = ( n33698 & ~n33701 ) | ( n33698 & n33715 ) | ( ~n33701 & n33715 ) ;
  assign n33726 = ~n33724 & n33725 ;
  assign n33727 = n33720 | n33726 ;
  assign n33728 = n33229 &  n33702 ;
  assign n33721 = x118 | n33229 ;
  assign n33722 = x118 &  n33229 ;
  assign n33723 = ( n33721 & ~n33722 ) | ( n33721 & 1'b0 ) | ( ~n33722 & 1'b0 ) ;
  assign n33732 = ( n15415 & n33697 ) | ( n15415 & n33723 ) | ( n33697 & n33723 ) ;
  assign n33733 = ( n33697 & ~n33701 ) | ( n33697 & n33723 ) | ( ~n33701 & n33723 ) ;
  assign n33734 = ~n33732 & n33733 ;
  assign n33735 = n33728 | n33734 ;
  assign n33736 = n33237 &  n33702 ;
  assign n33729 = x117 | n33237 ;
  assign n33730 = x117 &  n33237 ;
  assign n33731 = ( n33729 & ~n33730 ) | ( n33729 & 1'b0 ) | ( ~n33730 & 1'b0 ) ;
  assign n33740 = ( n15415 & n33696 ) | ( n15415 & n33731 ) | ( n33696 & n33731 ) ;
  assign n33741 = ( n33696 & ~n33701 ) | ( n33696 & n33731 ) | ( ~n33701 & n33731 ) ;
  assign n33742 = ~n33740 & n33741 ;
  assign n33743 = n33736 | n33742 ;
  assign n33744 = n33245 &  n33702 ;
  assign n33737 = x116 | n33245 ;
  assign n33738 = x116 &  n33245 ;
  assign n33739 = ( n33737 & ~n33738 ) | ( n33737 & 1'b0 ) | ( ~n33738 & 1'b0 ) ;
  assign n33748 = ( n15415 & n33695 ) | ( n15415 & n33739 ) | ( n33695 & n33739 ) ;
  assign n33749 = ( n33695 & ~n33701 ) | ( n33695 & n33739 ) | ( ~n33701 & n33739 ) ;
  assign n33750 = ~n33748 & n33749 ;
  assign n33751 = n33744 | n33750 ;
  assign n33752 = n33253 &  n33702 ;
  assign n33745 = x115 | n33253 ;
  assign n33746 = x115 &  n33253 ;
  assign n33747 = ( n33745 & ~n33746 ) | ( n33745 & 1'b0 ) | ( ~n33746 & 1'b0 ) ;
  assign n33756 = ( n15415 & n33694 ) | ( n15415 & n33747 ) | ( n33694 & n33747 ) ;
  assign n33757 = ( n33694 & ~n33701 ) | ( n33694 & n33747 ) | ( ~n33701 & n33747 ) ;
  assign n33758 = ~n33756 & n33757 ;
  assign n33759 = n33752 | n33758 ;
  assign n33760 = n33261 &  n33702 ;
  assign n33753 = x114 | n33261 ;
  assign n33754 = x114 &  n33261 ;
  assign n33755 = ( n33753 & ~n33754 ) | ( n33753 & 1'b0 ) | ( ~n33754 & 1'b0 ) ;
  assign n33764 = ( n15415 & n33693 ) | ( n15415 & n33755 ) | ( n33693 & n33755 ) ;
  assign n33765 = ( n33693 & ~n33701 ) | ( n33693 & n33755 ) | ( ~n33701 & n33755 ) ;
  assign n33766 = ~n33764 & n33765 ;
  assign n33767 = n33760 | n33766 ;
  assign n33768 = n33269 &  n33702 ;
  assign n33761 = x113 | n33269 ;
  assign n33762 = x113 &  n33269 ;
  assign n33763 = ( n33761 & ~n33762 ) | ( n33761 & 1'b0 ) | ( ~n33762 & 1'b0 ) ;
  assign n33772 = ( n15415 & n33692 ) | ( n15415 & n33763 ) | ( n33692 & n33763 ) ;
  assign n33773 = ( n33692 & ~n33701 ) | ( n33692 & n33763 ) | ( ~n33701 & n33763 ) ;
  assign n33774 = ~n33772 & n33773 ;
  assign n33775 = n33768 | n33774 ;
  assign n33776 = n33277 &  n33702 ;
  assign n33769 = x112 | n33277 ;
  assign n33770 = x112 &  n33277 ;
  assign n33771 = ( n33769 & ~n33770 ) | ( n33769 & 1'b0 ) | ( ~n33770 & 1'b0 ) ;
  assign n33780 = ( n15415 & n33691 ) | ( n15415 & n33771 ) | ( n33691 & n33771 ) ;
  assign n33781 = ( n33691 & ~n33701 ) | ( n33691 & n33771 ) | ( ~n33701 & n33771 ) ;
  assign n33782 = ~n33780 & n33781 ;
  assign n33783 = n33776 | n33782 ;
  assign n33784 = n33285 &  n33702 ;
  assign n33777 = x111 | n33285 ;
  assign n33778 = x111 &  n33285 ;
  assign n33779 = ( n33777 & ~n33778 ) | ( n33777 & 1'b0 ) | ( ~n33778 & 1'b0 ) ;
  assign n33788 = ( n15415 & n33690 ) | ( n15415 & n33779 ) | ( n33690 & n33779 ) ;
  assign n33789 = ( n33690 & ~n33701 ) | ( n33690 & n33779 ) | ( ~n33701 & n33779 ) ;
  assign n33790 = ~n33788 & n33789 ;
  assign n33791 = n33784 | n33790 ;
  assign n33792 = n33293 &  n33702 ;
  assign n33785 = x110 | n33293 ;
  assign n33786 = x110 &  n33293 ;
  assign n33787 = ( n33785 & ~n33786 ) | ( n33785 & 1'b0 ) | ( ~n33786 & 1'b0 ) ;
  assign n33796 = ( n15415 & n33689 ) | ( n15415 & n33787 ) | ( n33689 & n33787 ) ;
  assign n33797 = ( n33689 & ~n33701 ) | ( n33689 & n33787 ) | ( ~n33701 & n33787 ) ;
  assign n33798 = ~n33796 & n33797 ;
  assign n33799 = n33792 | n33798 ;
  assign n33800 = n33301 &  n33702 ;
  assign n33793 = x109 | n33301 ;
  assign n33794 = x109 &  n33301 ;
  assign n33795 = ( n33793 & ~n33794 ) | ( n33793 & 1'b0 ) | ( ~n33794 & 1'b0 ) ;
  assign n33804 = ( n15415 & n33688 ) | ( n15415 & n33795 ) | ( n33688 & n33795 ) ;
  assign n33805 = ( n33688 & ~n33701 ) | ( n33688 & n33795 ) | ( ~n33701 & n33795 ) ;
  assign n33806 = ~n33804 & n33805 ;
  assign n33807 = n33800 | n33806 ;
  assign n33808 = n33309 &  n33702 ;
  assign n33801 = x108 | n33309 ;
  assign n33802 = x108 &  n33309 ;
  assign n33803 = ( n33801 & ~n33802 ) | ( n33801 & 1'b0 ) | ( ~n33802 & 1'b0 ) ;
  assign n33812 = ( n15415 & n33687 ) | ( n15415 & n33803 ) | ( n33687 & n33803 ) ;
  assign n33813 = ( n33687 & ~n33701 ) | ( n33687 & n33803 ) | ( ~n33701 & n33803 ) ;
  assign n33814 = ~n33812 & n33813 ;
  assign n33815 = n33808 | n33814 ;
  assign n33816 = n33317 &  n33702 ;
  assign n33809 = x107 | n33317 ;
  assign n33810 = x107 &  n33317 ;
  assign n33811 = ( n33809 & ~n33810 ) | ( n33809 & 1'b0 ) | ( ~n33810 & 1'b0 ) ;
  assign n33820 = ( n15415 & n33686 ) | ( n15415 & n33811 ) | ( n33686 & n33811 ) ;
  assign n33821 = ( n33686 & ~n33701 ) | ( n33686 & n33811 ) | ( ~n33701 & n33811 ) ;
  assign n33822 = ~n33820 & n33821 ;
  assign n33823 = n33816 | n33822 ;
  assign n33824 = n33325 &  n33702 ;
  assign n33817 = x106 | n33325 ;
  assign n33818 = x106 &  n33325 ;
  assign n33819 = ( n33817 & ~n33818 ) | ( n33817 & 1'b0 ) | ( ~n33818 & 1'b0 ) ;
  assign n33828 = ( n15415 & n33685 ) | ( n15415 & n33819 ) | ( n33685 & n33819 ) ;
  assign n33829 = ( n33685 & ~n33701 ) | ( n33685 & n33819 ) | ( ~n33701 & n33819 ) ;
  assign n33830 = ~n33828 & n33829 ;
  assign n33831 = n33824 | n33830 ;
  assign n33832 = n33333 &  n33702 ;
  assign n33825 = x105 | n33333 ;
  assign n33826 = x105 &  n33333 ;
  assign n33827 = ( n33825 & ~n33826 ) | ( n33825 & 1'b0 ) | ( ~n33826 & 1'b0 ) ;
  assign n33836 = ( n15415 & n33684 ) | ( n15415 & n33827 ) | ( n33684 & n33827 ) ;
  assign n33837 = ( n33684 & ~n33701 ) | ( n33684 & n33827 ) | ( ~n33701 & n33827 ) ;
  assign n33838 = ~n33836 & n33837 ;
  assign n33839 = n33832 | n33838 ;
  assign n33840 = n33341 &  n33702 ;
  assign n33833 = x104 | n33341 ;
  assign n33834 = x104 &  n33341 ;
  assign n33835 = ( n33833 & ~n33834 ) | ( n33833 & 1'b0 ) | ( ~n33834 & 1'b0 ) ;
  assign n33844 = ( n15415 & n33683 ) | ( n15415 & n33835 ) | ( n33683 & n33835 ) ;
  assign n33845 = ( n33683 & ~n33701 ) | ( n33683 & n33835 ) | ( ~n33701 & n33835 ) ;
  assign n33846 = ~n33844 & n33845 ;
  assign n33847 = n33840 | n33846 ;
  assign n33848 = n33349 &  n33702 ;
  assign n33841 = x103 | n33349 ;
  assign n33842 = x103 &  n33349 ;
  assign n33843 = ( n33841 & ~n33842 ) | ( n33841 & 1'b0 ) | ( ~n33842 & 1'b0 ) ;
  assign n33852 = ( n15415 & n33682 ) | ( n15415 & n33843 ) | ( n33682 & n33843 ) ;
  assign n33853 = ( n33682 & ~n33701 ) | ( n33682 & n33843 ) | ( ~n33701 & n33843 ) ;
  assign n33854 = ~n33852 & n33853 ;
  assign n33855 = n33848 | n33854 ;
  assign n33856 = n33357 &  n33702 ;
  assign n33849 = x102 | n33357 ;
  assign n33850 = x102 &  n33357 ;
  assign n33851 = ( n33849 & ~n33850 ) | ( n33849 & 1'b0 ) | ( ~n33850 & 1'b0 ) ;
  assign n33860 = ( n15415 & n33681 ) | ( n15415 & n33851 ) | ( n33681 & n33851 ) ;
  assign n33861 = ( n33681 & ~n33701 ) | ( n33681 & n33851 ) | ( ~n33701 & n33851 ) ;
  assign n33862 = ~n33860 & n33861 ;
  assign n33863 = n33856 | n33862 ;
  assign n33864 = n33365 &  n33702 ;
  assign n33857 = x101 | n33365 ;
  assign n33858 = x101 &  n33365 ;
  assign n33859 = ( n33857 & ~n33858 ) | ( n33857 & 1'b0 ) | ( ~n33858 & 1'b0 ) ;
  assign n33868 = ( n15415 & n33680 ) | ( n15415 & n33859 ) | ( n33680 & n33859 ) ;
  assign n33869 = ( n33680 & ~n33701 ) | ( n33680 & n33859 ) | ( ~n33701 & n33859 ) ;
  assign n33870 = ~n33868 & n33869 ;
  assign n33871 = n33864 | n33870 ;
  assign n33872 = n33373 &  n33702 ;
  assign n33865 = x100 | n33373 ;
  assign n33866 = x100 &  n33373 ;
  assign n33867 = ( n33865 & ~n33866 ) | ( n33865 & 1'b0 ) | ( ~n33866 & 1'b0 ) ;
  assign n33876 = ( n15415 & n33679 ) | ( n15415 & n33867 ) | ( n33679 & n33867 ) ;
  assign n33877 = ( n33679 & ~n33701 ) | ( n33679 & n33867 ) | ( ~n33701 & n33867 ) ;
  assign n33878 = ~n33876 & n33877 ;
  assign n33879 = n33872 | n33878 ;
  assign n33880 = n33381 &  n33702 ;
  assign n33873 = x99 | n33381 ;
  assign n33874 = x99 &  n33381 ;
  assign n33875 = ( n33873 & ~n33874 ) | ( n33873 & 1'b0 ) | ( ~n33874 & 1'b0 ) ;
  assign n33884 = ( n15415 & n33678 ) | ( n15415 & n33875 ) | ( n33678 & n33875 ) ;
  assign n33885 = ( n33678 & ~n33701 ) | ( n33678 & n33875 ) | ( ~n33701 & n33875 ) ;
  assign n33886 = ~n33884 & n33885 ;
  assign n33887 = n33880 | n33886 ;
  assign n33888 = n33389 &  n33702 ;
  assign n33881 = x98 | n33389 ;
  assign n33882 = x98 &  n33389 ;
  assign n33883 = ( n33881 & ~n33882 ) | ( n33881 & 1'b0 ) | ( ~n33882 & 1'b0 ) ;
  assign n33892 = ( n15415 & n33677 ) | ( n15415 & n33883 ) | ( n33677 & n33883 ) ;
  assign n33893 = ( n33677 & ~n33701 ) | ( n33677 & n33883 ) | ( ~n33701 & n33883 ) ;
  assign n33894 = ~n33892 & n33893 ;
  assign n33895 = n33888 | n33894 ;
  assign n33896 = n33397 &  n33702 ;
  assign n33889 = x97 | n33397 ;
  assign n33890 = x97 &  n33397 ;
  assign n33891 = ( n33889 & ~n33890 ) | ( n33889 & 1'b0 ) | ( ~n33890 & 1'b0 ) ;
  assign n33900 = ( n15415 & n33676 ) | ( n15415 & n33891 ) | ( n33676 & n33891 ) ;
  assign n33901 = ( n33676 & ~n33701 ) | ( n33676 & n33891 ) | ( ~n33701 & n33891 ) ;
  assign n33902 = ~n33900 & n33901 ;
  assign n33903 = n33896 | n33902 ;
  assign n33904 = n33405 &  n33702 ;
  assign n33897 = x96 | n33405 ;
  assign n33898 = x96 &  n33405 ;
  assign n33899 = ( n33897 & ~n33898 ) | ( n33897 & 1'b0 ) | ( ~n33898 & 1'b0 ) ;
  assign n33908 = ( n15415 & n33675 ) | ( n15415 & n33899 ) | ( n33675 & n33899 ) ;
  assign n33909 = ( n33675 & ~n33701 ) | ( n33675 & n33899 ) | ( ~n33701 & n33899 ) ;
  assign n33910 = ~n33908 & n33909 ;
  assign n33911 = n33904 | n33910 ;
  assign n33912 = n33413 &  n33702 ;
  assign n33905 = x95 | n33413 ;
  assign n33906 = x95 &  n33413 ;
  assign n33907 = ( n33905 & ~n33906 ) | ( n33905 & 1'b0 ) | ( ~n33906 & 1'b0 ) ;
  assign n33916 = ( n15415 & n33674 ) | ( n15415 & n33907 ) | ( n33674 & n33907 ) ;
  assign n33917 = ( n33674 & ~n33701 ) | ( n33674 & n33907 ) | ( ~n33701 & n33907 ) ;
  assign n33918 = ~n33916 & n33917 ;
  assign n33919 = n33912 | n33918 ;
  assign n33920 = n33421 &  n33702 ;
  assign n33913 = x94 | n33421 ;
  assign n33914 = x94 &  n33421 ;
  assign n33915 = ( n33913 & ~n33914 ) | ( n33913 & 1'b0 ) | ( ~n33914 & 1'b0 ) ;
  assign n33924 = ( n15415 & n33673 ) | ( n15415 & n33915 ) | ( n33673 & n33915 ) ;
  assign n33925 = ( n33673 & ~n33701 ) | ( n33673 & n33915 ) | ( ~n33701 & n33915 ) ;
  assign n33926 = ~n33924 & n33925 ;
  assign n33927 = n33920 | n33926 ;
  assign n33928 = n33429 &  n33702 ;
  assign n33921 = x93 | n33429 ;
  assign n33922 = x93 &  n33429 ;
  assign n33923 = ( n33921 & ~n33922 ) | ( n33921 & 1'b0 ) | ( ~n33922 & 1'b0 ) ;
  assign n33932 = ( n15415 & n33672 ) | ( n15415 & n33923 ) | ( n33672 & n33923 ) ;
  assign n33933 = ( n33672 & ~n33701 ) | ( n33672 & n33923 ) | ( ~n33701 & n33923 ) ;
  assign n33934 = ~n33932 & n33933 ;
  assign n33935 = n33928 | n33934 ;
  assign n33936 = n33437 &  n33702 ;
  assign n33929 = x92 | n33437 ;
  assign n33930 = x92 &  n33437 ;
  assign n33931 = ( n33929 & ~n33930 ) | ( n33929 & 1'b0 ) | ( ~n33930 & 1'b0 ) ;
  assign n33940 = ( n15415 & n33671 ) | ( n15415 & n33931 ) | ( n33671 & n33931 ) ;
  assign n33941 = ( n33671 & ~n33701 ) | ( n33671 & n33931 ) | ( ~n33701 & n33931 ) ;
  assign n33942 = ~n33940 & n33941 ;
  assign n33943 = n33936 | n33942 ;
  assign n33944 = n33445 &  n33702 ;
  assign n33937 = x91 | n33445 ;
  assign n33938 = x91 &  n33445 ;
  assign n33939 = ( n33937 & ~n33938 ) | ( n33937 & 1'b0 ) | ( ~n33938 & 1'b0 ) ;
  assign n33948 = ( n15415 & n33670 ) | ( n15415 & n33939 ) | ( n33670 & n33939 ) ;
  assign n33949 = ( n33670 & ~n33701 ) | ( n33670 & n33939 ) | ( ~n33701 & n33939 ) ;
  assign n33950 = ~n33948 & n33949 ;
  assign n33951 = n33944 | n33950 ;
  assign n33952 = n33453 &  n33702 ;
  assign n33945 = x90 | n33453 ;
  assign n33946 = x90 &  n33453 ;
  assign n33947 = ( n33945 & ~n33946 ) | ( n33945 & 1'b0 ) | ( ~n33946 & 1'b0 ) ;
  assign n33956 = ( n15415 & n33669 ) | ( n15415 & n33947 ) | ( n33669 & n33947 ) ;
  assign n33957 = ( n33669 & ~n33701 ) | ( n33669 & n33947 ) | ( ~n33701 & n33947 ) ;
  assign n33958 = ~n33956 & n33957 ;
  assign n33959 = n33952 | n33958 ;
  assign n33960 = n33461 &  n33702 ;
  assign n33953 = x89 | n33461 ;
  assign n33954 = x89 &  n33461 ;
  assign n33955 = ( n33953 & ~n33954 ) | ( n33953 & 1'b0 ) | ( ~n33954 & 1'b0 ) ;
  assign n33964 = ( n15415 & n33668 ) | ( n15415 & n33955 ) | ( n33668 & n33955 ) ;
  assign n33965 = ( n33668 & ~n33701 ) | ( n33668 & n33955 ) | ( ~n33701 & n33955 ) ;
  assign n33966 = ~n33964 & n33965 ;
  assign n33967 = n33960 | n33966 ;
  assign n33968 = n33469 &  n33702 ;
  assign n33961 = x88 | n33469 ;
  assign n33962 = x88 &  n33469 ;
  assign n33963 = ( n33961 & ~n33962 ) | ( n33961 & 1'b0 ) | ( ~n33962 & 1'b0 ) ;
  assign n33972 = ( n15415 & n33667 ) | ( n15415 & n33963 ) | ( n33667 & n33963 ) ;
  assign n33973 = ( n33667 & ~n33701 ) | ( n33667 & n33963 ) | ( ~n33701 & n33963 ) ;
  assign n33974 = ~n33972 & n33973 ;
  assign n33975 = n33968 | n33974 ;
  assign n33976 = n33477 &  n33702 ;
  assign n33969 = x87 | n33477 ;
  assign n33970 = x87 &  n33477 ;
  assign n33971 = ( n33969 & ~n33970 ) | ( n33969 & 1'b0 ) | ( ~n33970 & 1'b0 ) ;
  assign n33980 = ( n15415 & n33666 ) | ( n15415 & n33971 ) | ( n33666 & n33971 ) ;
  assign n33981 = ( n33666 & ~n33701 ) | ( n33666 & n33971 ) | ( ~n33701 & n33971 ) ;
  assign n33982 = ~n33980 & n33981 ;
  assign n33983 = n33976 | n33982 ;
  assign n33984 = n33485 &  n33702 ;
  assign n33977 = x86 | n33485 ;
  assign n33978 = x86 &  n33485 ;
  assign n33979 = ( n33977 & ~n33978 ) | ( n33977 & 1'b0 ) | ( ~n33978 & 1'b0 ) ;
  assign n33988 = ( n15415 & n33665 ) | ( n15415 & n33979 ) | ( n33665 & n33979 ) ;
  assign n33989 = ( n33665 & ~n33701 ) | ( n33665 & n33979 ) | ( ~n33701 & n33979 ) ;
  assign n33990 = ~n33988 & n33989 ;
  assign n33991 = n33984 | n33990 ;
  assign n33992 = n33493 &  n33702 ;
  assign n33985 = x85 | n33493 ;
  assign n33986 = x85 &  n33493 ;
  assign n33987 = ( n33985 & ~n33986 ) | ( n33985 & 1'b0 ) | ( ~n33986 & 1'b0 ) ;
  assign n33996 = ( n15415 & n33664 ) | ( n15415 & n33987 ) | ( n33664 & n33987 ) ;
  assign n33997 = ( n33664 & ~n33701 ) | ( n33664 & n33987 ) | ( ~n33701 & n33987 ) ;
  assign n33998 = ~n33996 & n33997 ;
  assign n33999 = n33992 | n33998 ;
  assign n34000 = n33501 &  n33702 ;
  assign n33993 = x84 | n33501 ;
  assign n33994 = x84 &  n33501 ;
  assign n33995 = ( n33993 & ~n33994 ) | ( n33993 & 1'b0 ) | ( ~n33994 & 1'b0 ) ;
  assign n34004 = ( n15415 & n33663 ) | ( n15415 & n33995 ) | ( n33663 & n33995 ) ;
  assign n34005 = ( n33663 & ~n33701 ) | ( n33663 & n33995 ) | ( ~n33701 & n33995 ) ;
  assign n34006 = ~n34004 & n34005 ;
  assign n34007 = n34000 | n34006 ;
  assign n34008 = n33509 &  n33702 ;
  assign n34001 = x83 | n33509 ;
  assign n34002 = x83 &  n33509 ;
  assign n34003 = ( n34001 & ~n34002 ) | ( n34001 & 1'b0 ) | ( ~n34002 & 1'b0 ) ;
  assign n34012 = ( n15415 & n33662 ) | ( n15415 & n34003 ) | ( n33662 & n34003 ) ;
  assign n34013 = ( n33662 & ~n33701 ) | ( n33662 & n34003 ) | ( ~n33701 & n34003 ) ;
  assign n34014 = ~n34012 & n34013 ;
  assign n34015 = n34008 | n34014 ;
  assign n34016 = n33517 &  n33702 ;
  assign n34009 = x82 | n33517 ;
  assign n34010 = x82 &  n33517 ;
  assign n34011 = ( n34009 & ~n34010 ) | ( n34009 & 1'b0 ) | ( ~n34010 & 1'b0 ) ;
  assign n34020 = ( n15415 & n33661 ) | ( n15415 & n34011 ) | ( n33661 & n34011 ) ;
  assign n34021 = ( n33661 & ~n33701 ) | ( n33661 & n34011 ) | ( ~n33701 & n34011 ) ;
  assign n34022 = ~n34020 & n34021 ;
  assign n34023 = n34016 | n34022 ;
  assign n34024 = n33525 &  n33702 ;
  assign n34017 = x81 | n33525 ;
  assign n34018 = x81 &  n33525 ;
  assign n34019 = ( n34017 & ~n34018 ) | ( n34017 & 1'b0 ) | ( ~n34018 & 1'b0 ) ;
  assign n34028 = ( n15415 & n33660 ) | ( n15415 & n34019 ) | ( n33660 & n34019 ) ;
  assign n34029 = ( n33660 & ~n33701 ) | ( n33660 & n34019 ) | ( ~n33701 & n34019 ) ;
  assign n34030 = ~n34028 & n34029 ;
  assign n34031 = n34024 | n34030 ;
  assign n34032 = n33533 &  n33702 ;
  assign n34025 = x80 | n33533 ;
  assign n34026 = x80 &  n33533 ;
  assign n34027 = ( n34025 & ~n34026 ) | ( n34025 & 1'b0 ) | ( ~n34026 & 1'b0 ) ;
  assign n34036 = ( n15415 & n33659 ) | ( n15415 & n34027 ) | ( n33659 & n34027 ) ;
  assign n34037 = ( n33659 & ~n33701 ) | ( n33659 & n34027 ) | ( ~n33701 & n34027 ) ;
  assign n34038 = ~n34036 & n34037 ;
  assign n34039 = n34032 | n34038 ;
  assign n34040 = n33541 &  n33702 ;
  assign n34033 = x79 | n33541 ;
  assign n34034 = x79 &  n33541 ;
  assign n34035 = ( n34033 & ~n34034 ) | ( n34033 & 1'b0 ) | ( ~n34034 & 1'b0 ) ;
  assign n34044 = ( n15415 & n33658 ) | ( n15415 & n34035 ) | ( n33658 & n34035 ) ;
  assign n34045 = ( n33658 & ~n33701 ) | ( n33658 & n34035 ) | ( ~n33701 & n34035 ) ;
  assign n34046 = ~n34044 & n34045 ;
  assign n34047 = n34040 | n34046 ;
  assign n34048 = n33549 &  n33702 ;
  assign n34041 = x78 | n33549 ;
  assign n34042 = x78 &  n33549 ;
  assign n34043 = ( n34041 & ~n34042 ) | ( n34041 & 1'b0 ) | ( ~n34042 & 1'b0 ) ;
  assign n34052 = ( n15415 & n33657 ) | ( n15415 & n34043 ) | ( n33657 & n34043 ) ;
  assign n34053 = ( n33657 & ~n33701 ) | ( n33657 & n34043 ) | ( ~n33701 & n34043 ) ;
  assign n34054 = ~n34052 & n34053 ;
  assign n34055 = n34048 | n34054 ;
  assign n34056 = n33557 &  n33702 ;
  assign n34049 = x77 | n33557 ;
  assign n34050 = x77 &  n33557 ;
  assign n34051 = ( n34049 & ~n34050 ) | ( n34049 & 1'b0 ) | ( ~n34050 & 1'b0 ) ;
  assign n34060 = ( n15415 & n33656 ) | ( n15415 & n34051 ) | ( n33656 & n34051 ) ;
  assign n34061 = ( n33656 & ~n33701 ) | ( n33656 & n34051 ) | ( ~n33701 & n34051 ) ;
  assign n34062 = ~n34060 & n34061 ;
  assign n34063 = n34056 | n34062 ;
  assign n34064 = n33565 &  n33702 ;
  assign n34057 = x76 | n33565 ;
  assign n34058 = x76 &  n33565 ;
  assign n34059 = ( n34057 & ~n34058 ) | ( n34057 & 1'b0 ) | ( ~n34058 & 1'b0 ) ;
  assign n34068 = ( n15415 & n33655 ) | ( n15415 & n34059 ) | ( n33655 & n34059 ) ;
  assign n34069 = ( n33655 & ~n33701 ) | ( n33655 & n34059 ) | ( ~n33701 & n34059 ) ;
  assign n34070 = ~n34068 & n34069 ;
  assign n34071 = n34064 | n34070 ;
  assign n34072 = n33573 &  n33702 ;
  assign n34065 = x75 | n33573 ;
  assign n34066 = x75 &  n33573 ;
  assign n34067 = ( n34065 & ~n34066 ) | ( n34065 & 1'b0 ) | ( ~n34066 & 1'b0 ) ;
  assign n34076 = ( n15415 & n33654 ) | ( n15415 & n34067 ) | ( n33654 & n34067 ) ;
  assign n34077 = ( n33654 & ~n33701 ) | ( n33654 & n34067 ) | ( ~n33701 & n34067 ) ;
  assign n34078 = ~n34076 & n34077 ;
  assign n34079 = n34072 | n34078 ;
  assign n34080 = n33581 &  n33702 ;
  assign n34073 = x74 | n33581 ;
  assign n34074 = x74 &  n33581 ;
  assign n34075 = ( n34073 & ~n34074 ) | ( n34073 & 1'b0 ) | ( ~n34074 & 1'b0 ) ;
  assign n34084 = ( n15415 & n33653 ) | ( n15415 & n34075 ) | ( n33653 & n34075 ) ;
  assign n34085 = ( n33653 & ~n33701 ) | ( n33653 & n34075 ) | ( ~n33701 & n34075 ) ;
  assign n34086 = ~n34084 & n34085 ;
  assign n34087 = n34080 | n34086 ;
  assign n34088 = n33589 &  n33702 ;
  assign n34081 = x73 | n33589 ;
  assign n34082 = x73 &  n33589 ;
  assign n34083 = ( n34081 & ~n34082 ) | ( n34081 & 1'b0 ) | ( ~n34082 & 1'b0 ) ;
  assign n34092 = ( n15415 & n33652 ) | ( n15415 & n34083 ) | ( n33652 & n34083 ) ;
  assign n34093 = ( n33652 & ~n33701 ) | ( n33652 & n34083 ) | ( ~n33701 & n34083 ) ;
  assign n34094 = ~n34092 & n34093 ;
  assign n34095 = n34088 | n34094 ;
  assign n34096 = n33597 &  n33702 ;
  assign n34089 = x72 | n33597 ;
  assign n34090 = x72 &  n33597 ;
  assign n34091 = ( n34089 & ~n34090 ) | ( n34089 & 1'b0 ) | ( ~n34090 & 1'b0 ) ;
  assign n34100 = ( n15415 & n33651 ) | ( n15415 & n34091 ) | ( n33651 & n34091 ) ;
  assign n34101 = ( n33651 & ~n33701 ) | ( n33651 & n34091 ) | ( ~n33701 & n34091 ) ;
  assign n34102 = ~n34100 & n34101 ;
  assign n34103 = n34096 | n34102 ;
  assign n34104 = n33605 &  n33702 ;
  assign n34097 = x71 | n33605 ;
  assign n34098 = x71 &  n33605 ;
  assign n34099 = ( n34097 & ~n34098 ) | ( n34097 & 1'b0 ) | ( ~n34098 & 1'b0 ) ;
  assign n34108 = ( n15415 & n33650 ) | ( n15415 & n34099 ) | ( n33650 & n34099 ) ;
  assign n34109 = ( n33650 & ~n33701 ) | ( n33650 & n34099 ) | ( ~n33701 & n34099 ) ;
  assign n34110 = ~n34108 & n34109 ;
  assign n34111 = n34104 | n34110 ;
  assign n34112 = n33613 &  n33702 ;
  assign n34105 = x70 | n33613 ;
  assign n34106 = x70 &  n33613 ;
  assign n34107 = ( n34105 & ~n34106 ) | ( n34105 & 1'b0 ) | ( ~n34106 & 1'b0 ) ;
  assign n34116 = ( n15415 & n33649 ) | ( n15415 & n34107 ) | ( n33649 & n34107 ) ;
  assign n34117 = ( n33649 & ~n33701 ) | ( n33649 & n34107 ) | ( ~n33701 & n34107 ) ;
  assign n34118 = ~n34116 & n34117 ;
  assign n34119 = n34112 | n34118 ;
  assign n34120 = n33621 &  n33702 ;
  assign n34113 = x69 | n33621 ;
  assign n34114 = x69 &  n33621 ;
  assign n34115 = ( n34113 & ~n34114 ) | ( n34113 & 1'b0 ) | ( ~n34114 & 1'b0 ) ;
  assign n34124 = ( n15415 & n33648 ) | ( n15415 & n34115 ) | ( n33648 & n34115 ) ;
  assign n34125 = ( n33648 & ~n33701 ) | ( n33648 & n34115 ) | ( ~n33701 & n34115 ) ;
  assign n34126 = ~n34124 & n34125 ;
  assign n34127 = n34120 | n34126 ;
  assign n34128 = n33629 &  n33702 ;
  assign n34121 = x68 | n33629 ;
  assign n34122 = x68 &  n33629 ;
  assign n34123 = ( n34121 & ~n34122 ) | ( n34121 & 1'b0 ) | ( ~n34122 & 1'b0 ) ;
  assign n34132 = ( n15415 & n33647 ) | ( n15415 & n34123 ) | ( n33647 & n34123 ) ;
  assign n34133 = ( n33647 & ~n33701 ) | ( n33647 & n34123 ) | ( ~n33701 & n34123 ) ;
  assign n34134 = ~n34132 & n34133 ;
  assign n34135 = n34128 | n34134 ;
  assign n34136 = n33634 &  n33702 ;
  assign n34129 = x67 | n33634 ;
  assign n34130 = x67 &  n33634 ;
  assign n34131 = ( n34129 & ~n34130 ) | ( n34129 & 1'b0 ) | ( ~n34130 & 1'b0 ) ;
  assign n34140 = ( n15415 & n33646 ) | ( n15415 & n34131 ) | ( n33646 & n34131 ) ;
  assign n34141 = ( n33646 & ~n33701 ) | ( n33646 & n34131 ) | ( ~n33701 & n34131 ) ;
  assign n34142 = ~n34140 & n34141 ;
  assign n34143 = n34136 | n34142 ;
  assign n34144 = n33640 &  n33702 ;
  assign n34137 = x66 | n33640 ;
  assign n34138 = x66 &  n33640 ;
  assign n34139 = ( n34137 & ~n34138 ) | ( n34137 & 1'b0 ) | ( ~n34138 & 1'b0 ) ;
  assign n34145 = ( n15415 & n33645 ) | ( n15415 & n34139 ) | ( n33645 & n34139 ) ;
  assign n34146 = ( n33645 & ~n33701 ) | ( n33645 & n34139 ) | ( ~n33701 & n34139 ) ;
  assign n34147 = ~n34145 & n34146 ;
  assign n34148 = n34144 | n34147 ;
  assign n34149 = n33644 &  n33702 ;
  assign n34150 = ( x65 & ~x7 ) | ( x65 & n33641 ) | ( ~x7 & n33641 ) ;
  assign n34151 = ( x7 & ~n33641 ) | ( x7 & x65 ) | ( ~n33641 & x65 ) ;
  assign n34152 = ( n34150 & ~x65 ) | ( n34150 & n34151 ) | ( ~x65 & n34151 ) ;
  assign n34153 = ( n15357 & ~n15415 ) | ( n15357 & n34152 ) | ( ~n15415 & n34152 ) ;
  assign n34154 = ( n15357 & n33701 ) | ( n15357 & n34152 ) | ( n33701 & n34152 ) ;
  assign n34155 = ( n34153 & ~n34154 ) | ( n34153 & 1'b0 ) | ( ~n34154 & 1'b0 ) ;
  assign n34156 = n34149 | n34155 ;
  assign n34157 = ( n15837 & ~n33701 ) | ( n15837 & 1'b0 ) | ( ~n33701 & 1'b0 ) ;
  assign n34158 = ( x6 & ~n34157 ) | ( x6 & 1'b0 ) | ( ~n34157 & 1'b0 ) ;
  assign n34159 = ( n15841 & ~n33701 ) | ( n15841 & 1'b0 ) | ( ~n33701 & 1'b0 ) ;
  assign n34160 = n34158 | n34159 ;
  assign n34161 = ( x65 & ~n34160 ) | ( x65 & n15844 ) | ( ~n34160 & n15844 ) ;
  assign n34162 = ( x66 & ~n34156 ) | ( x66 & n34161 ) | ( ~n34156 & n34161 ) ;
  assign n34163 = ( x67 & ~n34148 ) | ( x67 & n34162 ) | ( ~n34148 & n34162 ) ;
  assign n34164 = ( x68 & ~n34143 ) | ( x68 & n34163 ) | ( ~n34143 & n34163 ) ;
  assign n34165 = ( x69 & ~n34135 ) | ( x69 & n34164 ) | ( ~n34135 & n34164 ) ;
  assign n34166 = ( x70 & ~n34127 ) | ( x70 & n34165 ) | ( ~n34127 & n34165 ) ;
  assign n34167 = ( x71 & ~n34119 ) | ( x71 & n34166 ) | ( ~n34119 & n34166 ) ;
  assign n34168 = ( x72 & ~n34111 ) | ( x72 & n34167 ) | ( ~n34111 & n34167 ) ;
  assign n34169 = ( x73 & ~n34103 ) | ( x73 & n34168 ) | ( ~n34103 & n34168 ) ;
  assign n34170 = ( x74 & ~n34095 ) | ( x74 & n34169 ) | ( ~n34095 & n34169 ) ;
  assign n34171 = ( x75 & ~n34087 ) | ( x75 & n34170 ) | ( ~n34087 & n34170 ) ;
  assign n34172 = ( x76 & ~n34079 ) | ( x76 & n34171 ) | ( ~n34079 & n34171 ) ;
  assign n34173 = ( x77 & ~n34071 ) | ( x77 & n34172 ) | ( ~n34071 & n34172 ) ;
  assign n34174 = ( x78 & ~n34063 ) | ( x78 & n34173 ) | ( ~n34063 & n34173 ) ;
  assign n34175 = ( x79 & ~n34055 ) | ( x79 & n34174 ) | ( ~n34055 & n34174 ) ;
  assign n34176 = ( x80 & ~n34047 ) | ( x80 & n34175 ) | ( ~n34047 & n34175 ) ;
  assign n34177 = ( x81 & ~n34039 ) | ( x81 & n34176 ) | ( ~n34039 & n34176 ) ;
  assign n34178 = ( x82 & ~n34031 ) | ( x82 & n34177 ) | ( ~n34031 & n34177 ) ;
  assign n34179 = ( x83 & ~n34023 ) | ( x83 & n34178 ) | ( ~n34023 & n34178 ) ;
  assign n34180 = ( x84 & ~n34015 ) | ( x84 & n34179 ) | ( ~n34015 & n34179 ) ;
  assign n34181 = ( x85 & ~n34007 ) | ( x85 & n34180 ) | ( ~n34007 & n34180 ) ;
  assign n34182 = ( x86 & ~n33999 ) | ( x86 & n34181 ) | ( ~n33999 & n34181 ) ;
  assign n34183 = ( x87 & ~n33991 ) | ( x87 & n34182 ) | ( ~n33991 & n34182 ) ;
  assign n34184 = ( x88 & ~n33983 ) | ( x88 & n34183 ) | ( ~n33983 & n34183 ) ;
  assign n34185 = ( x89 & ~n33975 ) | ( x89 & n34184 ) | ( ~n33975 & n34184 ) ;
  assign n34186 = ( x90 & ~n33967 ) | ( x90 & n34185 ) | ( ~n33967 & n34185 ) ;
  assign n34187 = ( x91 & ~n33959 ) | ( x91 & n34186 ) | ( ~n33959 & n34186 ) ;
  assign n34188 = ( x92 & ~n33951 ) | ( x92 & n34187 ) | ( ~n33951 & n34187 ) ;
  assign n34189 = ( x93 & ~n33943 ) | ( x93 & n34188 ) | ( ~n33943 & n34188 ) ;
  assign n34190 = ( x94 & ~n33935 ) | ( x94 & n34189 ) | ( ~n33935 & n34189 ) ;
  assign n34191 = ( x95 & ~n33927 ) | ( x95 & n34190 ) | ( ~n33927 & n34190 ) ;
  assign n34192 = ( x96 & ~n33919 ) | ( x96 & n34191 ) | ( ~n33919 & n34191 ) ;
  assign n34193 = ( x97 & ~n33911 ) | ( x97 & n34192 ) | ( ~n33911 & n34192 ) ;
  assign n34194 = ( x98 & ~n33903 ) | ( x98 & n34193 ) | ( ~n33903 & n34193 ) ;
  assign n34195 = ( x99 & ~n33895 ) | ( x99 & n34194 ) | ( ~n33895 & n34194 ) ;
  assign n34196 = ( x100 & ~n33887 ) | ( x100 & n34195 ) | ( ~n33887 & n34195 ) ;
  assign n34197 = ( x101 & ~n33879 ) | ( x101 & n34196 ) | ( ~n33879 & n34196 ) ;
  assign n34198 = ( x102 & ~n33871 ) | ( x102 & n34197 ) | ( ~n33871 & n34197 ) ;
  assign n34199 = ( x103 & ~n33863 ) | ( x103 & n34198 ) | ( ~n33863 & n34198 ) ;
  assign n34200 = ( x104 & ~n33855 ) | ( x104 & n34199 ) | ( ~n33855 & n34199 ) ;
  assign n34201 = ( x105 & ~n33847 ) | ( x105 & n34200 ) | ( ~n33847 & n34200 ) ;
  assign n34202 = ( x106 & ~n33839 ) | ( x106 & n34201 ) | ( ~n33839 & n34201 ) ;
  assign n34203 = ( x107 & ~n33831 ) | ( x107 & n34202 ) | ( ~n33831 & n34202 ) ;
  assign n34204 = ( x108 & ~n33823 ) | ( x108 & n34203 ) | ( ~n33823 & n34203 ) ;
  assign n34205 = ( x109 & ~n33815 ) | ( x109 & n34204 ) | ( ~n33815 & n34204 ) ;
  assign n34206 = ( x110 & ~n33807 ) | ( x110 & n34205 ) | ( ~n33807 & n34205 ) ;
  assign n34207 = ( x111 & ~n33799 ) | ( x111 & n34206 ) | ( ~n33799 & n34206 ) ;
  assign n34208 = ( x112 & ~n33791 ) | ( x112 & n34207 ) | ( ~n33791 & n34207 ) ;
  assign n34209 = ( x113 & ~n33783 ) | ( x113 & n34208 ) | ( ~n33783 & n34208 ) ;
  assign n34210 = ( x114 & ~n33775 ) | ( x114 & n34209 ) | ( ~n33775 & n34209 ) ;
  assign n34211 = ( x115 & ~n33767 ) | ( x115 & n34210 ) | ( ~n33767 & n34210 ) ;
  assign n34212 = ( x116 & ~n33759 ) | ( x116 & n34211 ) | ( ~n33759 & n34211 ) ;
  assign n34213 = ( x117 & ~n33751 ) | ( x117 & n34212 ) | ( ~n33751 & n34212 ) ;
  assign n34214 = ( x118 & ~n33743 ) | ( x118 & n34213 ) | ( ~n33743 & n34213 ) ;
  assign n34215 = ( x119 & ~n33735 ) | ( x119 & n34214 ) | ( ~n33735 & n34214 ) ;
  assign n34216 = ( x120 & ~n33727 ) | ( x120 & n34215 ) | ( ~n33727 & n34215 ) ;
  assign n34217 = ( x121 & ~n33719 ) | ( x121 & n34216 ) | ( ~n33719 & n34216 ) ;
  assign n34218 = ( x122 & ~n33703 ) | ( x122 & 1'b0 ) | ( ~n33703 & 1'b0 ) ;
  assign n34219 = ~n33709 & n34218 ;
  assign n34220 = ( n34217 & ~n33711 ) | ( n34217 & n34219 ) | ( ~n33711 & n34219 ) ;
  assign n34221 = ( n33711 & ~n15943 ) | ( n33711 & n34220 ) | ( ~n15943 & n34220 ) ;
  assign n34222 = n15943 | n34221 ;
  assign n34223 = ~n33710 |  n15415 ;
  assign n34239 = n33719 &  n34223 ;
  assign n34240 = n34222 &  n34239 ;
  assign n34224 = n34222 &  n34223 ;
  assign n34225 = x121 | n33719 ;
  assign n34226 = x121 &  n33719 ;
  assign n34227 = ( n34225 & ~n34226 ) | ( n34225 & 1'b0 ) | ( ~n34226 & 1'b0 ) ;
  assign n34242 = ( n34216 & n34224 ) | ( n34216 & n34227 ) | ( n34224 & n34227 ) ;
  assign n34241 = n34216 | n34227 ;
  assign n34243 = ( n34240 & ~n34242 ) | ( n34240 & n34241 ) | ( ~n34242 & n34241 ) ;
  assign n34247 = n33727 &  n34223 ;
  assign n34248 = n34222 &  n34247 ;
  assign n34236 = x120 | n33727 ;
  assign n34237 = x120 &  n33727 ;
  assign n34238 = ( n34236 & ~n34237 ) | ( n34236 & 1'b0 ) | ( ~n34237 & 1'b0 ) ;
  assign n34250 = ( n34215 & n34224 ) | ( n34215 & n34238 ) | ( n34224 & n34238 ) ;
  assign n34249 = n34215 | n34238 ;
  assign n34251 = ( n34248 & ~n34250 ) | ( n34248 & n34249 ) | ( ~n34250 & n34249 ) ;
  assign n34255 = n33735 &  n34223 ;
  assign n34256 = n34222 &  n34255 ;
  assign n34244 = x119 | n33735 ;
  assign n34245 = x119 &  n33735 ;
  assign n34246 = ( n34244 & ~n34245 ) | ( n34244 & 1'b0 ) | ( ~n34245 & 1'b0 ) ;
  assign n34258 = ( n34214 & n34224 ) | ( n34214 & n34246 ) | ( n34224 & n34246 ) ;
  assign n34257 = n34214 | n34246 ;
  assign n34259 = ( n34256 & ~n34258 ) | ( n34256 & n34257 ) | ( ~n34258 & n34257 ) ;
  assign n34263 = n33743 &  n34223 ;
  assign n34264 = n34222 &  n34263 ;
  assign n34252 = x118 | n33743 ;
  assign n34253 = x118 &  n33743 ;
  assign n34254 = ( n34252 & ~n34253 ) | ( n34252 & 1'b0 ) | ( ~n34253 & 1'b0 ) ;
  assign n34266 = ( n34213 & n34224 ) | ( n34213 & n34254 ) | ( n34224 & n34254 ) ;
  assign n34265 = n34213 | n34254 ;
  assign n34267 = ( n34264 & ~n34266 ) | ( n34264 & n34265 ) | ( ~n34266 & n34265 ) ;
  assign n34271 = n33751 &  n34223 ;
  assign n34272 = n34222 &  n34271 ;
  assign n34260 = x117 | n33751 ;
  assign n34261 = x117 &  n33751 ;
  assign n34262 = ( n34260 & ~n34261 ) | ( n34260 & 1'b0 ) | ( ~n34261 & 1'b0 ) ;
  assign n34274 = ( n34212 & n34224 ) | ( n34212 & n34262 ) | ( n34224 & n34262 ) ;
  assign n34273 = n34212 | n34262 ;
  assign n34275 = ( n34272 & ~n34274 ) | ( n34272 & n34273 ) | ( ~n34274 & n34273 ) ;
  assign n34279 = n33759 &  n34223 ;
  assign n34280 = n34222 &  n34279 ;
  assign n34268 = x116 | n33759 ;
  assign n34269 = x116 &  n33759 ;
  assign n34270 = ( n34268 & ~n34269 ) | ( n34268 & 1'b0 ) | ( ~n34269 & 1'b0 ) ;
  assign n34282 = ( n34211 & n34224 ) | ( n34211 & n34270 ) | ( n34224 & n34270 ) ;
  assign n34281 = n34211 | n34270 ;
  assign n34283 = ( n34280 & ~n34282 ) | ( n34280 & n34281 ) | ( ~n34282 & n34281 ) ;
  assign n34287 = n33767 &  n34223 ;
  assign n34288 = n34222 &  n34287 ;
  assign n34276 = x115 | n33767 ;
  assign n34277 = x115 &  n33767 ;
  assign n34278 = ( n34276 & ~n34277 ) | ( n34276 & 1'b0 ) | ( ~n34277 & 1'b0 ) ;
  assign n34290 = ( n34210 & n34224 ) | ( n34210 & n34278 ) | ( n34224 & n34278 ) ;
  assign n34289 = n34210 | n34278 ;
  assign n34291 = ( n34288 & ~n34290 ) | ( n34288 & n34289 ) | ( ~n34290 & n34289 ) ;
  assign n34295 = n33775 &  n34223 ;
  assign n34296 = n34222 &  n34295 ;
  assign n34284 = x114 | n33775 ;
  assign n34285 = x114 &  n33775 ;
  assign n34286 = ( n34284 & ~n34285 ) | ( n34284 & 1'b0 ) | ( ~n34285 & 1'b0 ) ;
  assign n34298 = ( n34209 & n34224 ) | ( n34209 & n34286 ) | ( n34224 & n34286 ) ;
  assign n34297 = n34209 | n34286 ;
  assign n34299 = ( n34296 & ~n34298 ) | ( n34296 & n34297 ) | ( ~n34298 & n34297 ) ;
  assign n34303 = n33783 &  n34223 ;
  assign n34304 = n34222 &  n34303 ;
  assign n34292 = x113 | n33783 ;
  assign n34293 = x113 &  n33783 ;
  assign n34294 = ( n34292 & ~n34293 ) | ( n34292 & 1'b0 ) | ( ~n34293 & 1'b0 ) ;
  assign n34306 = ( n34208 & n34224 ) | ( n34208 & n34294 ) | ( n34224 & n34294 ) ;
  assign n34305 = n34208 | n34294 ;
  assign n34307 = ( n34304 & ~n34306 ) | ( n34304 & n34305 ) | ( ~n34306 & n34305 ) ;
  assign n34311 = n33791 &  n34223 ;
  assign n34312 = n34222 &  n34311 ;
  assign n34300 = x112 | n33791 ;
  assign n34301 = x112 &  n33791 ;
  assign n34302 = ( n34300 & ~n34301 ) | ( n34300 & 1'b0 ) | ( ~n34301 & 1'b0 ) ;
  assign n34314 = ( n34207 & n34224 ) | ( n34207 & n34302 ) | ( n34224 & n34302 ) ;
  assign n34313 = n34207 | n34302 ;
  assign n34315 = ( n34312 & ~n34314 ) | ( n34312 & n34313 ) | ( ~n34314 & n34313 ) ;
  assign n34319 = n33799 &  n34223 ;
  assign n34320 = n34222 &  n34319 ;
  assign n34308 = x111 | n33799 ;
  assign n34309 = x111 &  n33799 ;
  assign n34310 = ( n34308 & ~n34309 ) | ( n34308 & 1'b0 ) | ( ~n34309 & 1'b0 ) ;
  assign n34322 = ( n34206 & n34224 ) | ( n34206 & n34310 ) | ( n34224 & n34310 ) ;
  assign n34321 = n34206 | n34310 ;
  assign n34323 = ( n34320 & ~n34322 ) | ( n34320 & n34321 ) | ( ~n34322 & n34321 ) ;
  assign n34327 = n33807 &  n34223 ;
  assign n34328 = n34222 &  n34327 ;
  assign n34316 = x110 | n33807 ;
  assign n34317 = x110 &  n33807 ;
  assign n34318 = ( n34316 & ~n34317 ) | ( n34316 & 1'b0 ) | ( ~n34317 & 1'b0 ) ;
  assign n34330 = ( n34205 & n34224 ) | ( n34205 & n34318 ) | ( n34224 & n34318 ) ;
  assign n34329 = n34205 | n34318 ;
  assign n34331 = ( n34328 & ~n34330 ) | ( n34328 & n34329 ) | ( ~n34330 & n34329 ) ;
  assign n34335 = n33815 &  n34223 ;
  assign n34336 = n34222 &  n34335 ;
  assign n34324 = x109 | n33815 ;
  assign n34325 = x109 &  n33815 ;
  assign n34326 = ( n34324 & ~n34325 ) | ( n34324 & 1'b0 ) | ( ~n34325 & 1'b0 ) ;
  assign n34338 = ( n34204 & n34224 ) | ( n34204 & n34326 ) | ( n34224 & n34326 ) ;
  assign n34337 = n34204 | n34326 ;
  assign n34339 = ( n34336 & ~n34338 ) | ( n34336 & n34337 ) | ( ~n34338 & n34337 ) ;
  assign n34343 = n33823 &  n34223 ;
  assign n34344 = n34222 &  n34343 ;
  assign n34332 = x108 | n33823 ;
  assign n34333 = x108 &  n33823 ;
  assign n34334 = ( n34332 & ~n34333 ) | ( n34332 & 1'b0 ) | ( ~n34333 & 1'b0 ) ;
  assign n34346 = ( n34203 & n34224 ) | ( n34203 & n34334 ) | ( n34224 & n34334 ) ;
  assign n34345 = n34203 | n34334 ;
  assign n34347 = ( n34344 & ~n34346 ) | ( n34344 & n34345 ) | ( ~n34346 & n34345 ) ;
  assign n34351 = n33831 &  n34223 ;
  assign n34352 = n34222 &  n34351 ;
  assign n34340 = x107 | n33831 ;
  assign n34341 = x107 &  n33831 ;
  assign n34342 = ( n34340 & ~n34341 ) | ( n34340 & 1'b0 ) | ( ~n34341 & 1'b0 ) ;
  assign n34354 = ( n34202 & n34224 ) | ( n34202 & n34342 ) | ( n34224 & n34342 ) ;
  assign n34353 = n34202 | n34342 ;
  assign n34355 = ( n34352 & ~n34354 ) | ( n34352 & n34353 ) | ( ~n34354 & n34353 ) ;
  assign n34359 = n33839 &  n34223 ;
  assign n34360 = n34222 &  n34359 ;
  assign n34348 = x106 | n33839 ;
  assign n34349 = x106 &  n33839 ;
  assign n34350 = ( n34348 & ~n34349 ) | ( n34348 & 1'b0 ) | ( ~n34349 & 1'b0 ) ;
  assign n34362 = ( n34201 & n34224 ) | ( n34201 & n34350 ) | ( n34224 & n34350 ) ;
  assign n34361 = n34201 | n34350 ;
  assign n34363 = ( n34360 & ~n34362 ) | ( n34360 & n34361 ) | ( ~n34362 & n34361 ) ;
  assign n34367 = n33847 &  n34223 ;
  assign n34368 = n34222 &  n34367 ;
  assign n34356 = x105 | n33847 ;
  assign n34357 = x105 &  n33847 ;
  assign n34358 = ( n34356 & ~n34357 ) | ( n34356 & 1'b0 ) | ( ~n34357 & 1'b0 ) ;
  assign n34370 = ( n34200 & n34224 ) | ( n34200 & n34358 ) | ( n34224 & n34358 ) ;
  assign n34369 = n34200 | n34358 ;
  assign n34371 = ( n34368 & ~n34370 ) | ( n34368 & n34369 ) | ( ~n34370 & n34369 ) ;
  assign n34375 = n33855 &  n34223 ;
  assign n34376 = n34222 &  n34375 ;
  assign n34364 = x104 | n33855 ;
  assign n34365 = x104 &  n33855 ;
  assign n34366 = ( n34364 & ~n34365 ) | ( n34364 & 1'b0 ) | ( ~n34365 & 1'b0 ) ;
  assign n34378 = ( n34199 & n34224 ) | ( n34199 & n34366 ) | ( n34224 & n34366 ) ;
  assign n34377 = n34199 | n34366 ;
  assign n34379 = ( n34376 & ~n34378 ) | ( n34376 & n34377 ) | ( ~n34378 & n34377 ) ;
  assign n34383 = n33863 &  n34223 ;
  assign n34384 = n34222 &  n34383 ;
  assign n34372 = x103 | n33863 ;
  assign n34373 = x103 &  n33863 ;
  assign n34374 = ( n34372 & ~n34373 ) | ( n34372 & 1'b0 ) | ( ~n34373 & 1'b0 ) ;
  assign n34386 = ( n34198 & n34224 ) | ( n34198 & n34374 ) | ( n34224 & n34374 ) ;
  assign n34385 = n34198 | n34374 ;
  assign n34387 = ( n34384 & ~n34386 ) | ( n34384 & n34385 ) | ( ~n34386 & n34385 ) ;
  assign n34391 = n33871 &  n34223 ;
  assign n34392 = n34222 &  n34391 ;
  assign n34380 = x102 | n33871 ;
  assign n34381 = x102 &  n33871 ;
  assign n34382 = ( n34380 & ~n34381 ) | ( n34380 & 1'b0 ) | ( ~n34381 & 1'b0 ) ;
  assign n34394 = ( n34197 & n34224 ) | ( n34197 & n34382 ) | ( n34224 & n34382 ) ;
  assign n34393 = n34197 | n34382 ;
  assign n34395 = ( n34392 & ~n34394 ) | ( n34392 & n34393 ) | ( ~n34394 & n34393 ) ;
  assign n34399 = n33879 &  n34223 ;
  assign n34400 = n34222 &  n34399 ;
  assign n34388 = x101 | n33879 ;
  assign n34389 = x101 &  n33879 ;
  assign n34390 = ( n34388 & ~n34389 ) | ( n34388 & 1'b0 ) | ( ~n34389 & 1'b0 ) ;
  assign n34402 = ( n34196 & n34224 ) | ( n34196 & n34390 ) | ( n34224 & n34390 ) ;
  assign n34401 = n34196 | n34390 ;
  assign n34403 = ( n34400 & ~n34402 ) | ( n34400 & n34401 ) | ( ~n34402 & n34401 ) ;
  assign n34407 = n33887 &  n34223 ;
  assign n34408 = n34222 &  n34407 ;
  assign n34396 = x100 | n33887 ;
  assign n34397 = x100 &  n33887 ;
  assign n34398 = ( n34396 & ~n34397 ) | ( n34396 & 1'b0 ) | ( ~n34397 & 1'b0 ) ;
  assign n34410 = ( n34195 & n34224 ) | ( n34195 & n34398 ) | ( n34224 & n34398 ) ;
  assign n34409 = n34195 | n34398 ;
  assign n34411 = ( n34408 & ~n34410 ) | ( n34408 & n34409 ) | ( ~n34410 & n34409 ) ;
  assign n34415 = n33895 &  n34223 ;
  assign n34416 = n34222 &  n34415 ;
  assign n34404 = x99 | n33895 ;
  assign n34405 = x99 &  n33895 ;
  assign n34406 = ( n34404 & ~n34405 ) | ( n34404 & 1'b0 ) | ( ~n34405 & 1'b0 ) ;
  assign n34418 = ( n34194 & n34224 ) | ( n34194 & n34406 ) | ( n34224 & n34406 ) ;
  assign n34417 = n34194 | n34406 ;
  assign n34419 = ( n34416 & ~n34418 ) | ( n34416 & n34417 ) | ( ~n34418 & n34417 ) ;
  assign n34423 = n33903 &  n34223 ;
  assign n34424 = n34222 &  n34423 ;
  assign n34412 = x98 | n33903 ;
  assign n34413 = x98 &  n33903 ;
  assign n34414 = ( n34412 & ~n34413 ) | ( n34412 & 1'b0 ) | ( ~n34413 & 1'b0 ) ;
  assign n34426 = ( n34193 & n34224 ) | ( n34193 & n34414 ) | ( n34224 & n34414 ) ;
  assign n34425 = n34193 | n34414 ;
  assign n34427 = ( n34424 & ~n34426 ) | ( n34424 & n34425 ) | ( ~n34426 & n34425 ) ;
  assign n34431 = n33911 &  n34223 ;
  assign n34432 = n34222 &  n34431 ;
  assign n34420 = x97 | n33911 ;
  assign n34421 = x97 &  n33911 ;
  assign n34422 = ( n34420 & ~n34421 ) | ( n34420 & 1'b0 ) | ( ~n34421 & 1'b0 ) ;
  assign n34434 = ( n34192 & n34224 ) | ( n34192 & n34422 ) | ( n34224 & n34422 ) ;
  assign n34433 = n34192 | n34422 ;
  assign n34435 = ( n34432 & ~n34434 ) | ( n34432 & n34433 ) | ( ~n34434 & n34433 ) ;
  assign n34439 = n33919 &  n34223 ;
  assign n34440 = n34222 &  n34439 ;
  assign n34428 = x96 | n33919 ;
  assign n34429 = x96 &  n33919 ;
  assign n34430 = ( n34428 & ~n34429 ) | ( n34428 & 1'b0 ) | ( ~n34429 & 1'b0 ) ;
  assign n34442 = ( n34191 & n34224 ) | ( n34191 & n34430 ) | ( n34224 & n34430 ) ;
  assign n34441 = n34191 | n34430 ;
  assign n34443 = ( n34440 & ~n34442 ) | ( n34440 & n34441 ) | ( ~n34442 & n34441 ) ;
  assign n34447 = n33927 &  n34223 ;
  assign n34448 = n34222 &  n34447 ;
  assign n34436 = x95 | n33927 ;
  assign n34437 = x95 &  n33927 ;
  assign n34438 = ( n34436 & ~n34437 ) | ( n34436 & 1'b0 ) | ( ~n34437 & 1'b0 ) ;
  assign n34450 = ( n34190 & n34224 ) | ( n34190 & n34438 ) | ( n34224 & n34438 ) ;
  assign n34449 = n34190 | n34438 ;
  assign n34451 = ( n34448 & ~n34450 ) | ( n34448 & n34449 ) | ( ~n34450 & n34449 ) ;
  assign n34455 = n33935 &  n34223 ;
  assign n34456 = n34222 &  n34455 ;
  assign n34444 = x94 | n33935 ;
  assign n34445 = x94 &  n33935 ;
  assign n34446 = ( n34444 & ~n34445 ) | ( n34444 & 1'b0 ) | ( ~n34445 & 1'b0 ) ;
  assign n34458 = ( n34189 & n34224 ) | ( n34189 & n34446 ) | ( n34224 & n34446 ) ;
  assign n34457 = n34189 | n34446 ;
  assign n34459 = ( n34456 & ~n34458 ) | ( n34456 & n34457 ) | ( ~n34458 & n34457 ) ;
  assign n34463 = n33943 &  n34223 ;
  assign n34464 = n34222 &  n34463 ;
  assign n34452 = x93 | n33943 ;
  assign n34453 = x93 &  n33943 ;
  assign n34454 = ( n34452 & ~n34453 ) | ( n34452 & 1'b0 ) | ( ~n34453 & 1'b0 ) ;
  assign n34466 = ( n34188 & n34224 ) | ( n34188 & n34454 ) | ( n34224 & n34454 ) ;
  assign n34465 = n34188 | n34454 ;
  assign n34467 = ( n34464 & ~n34466 ) | ( n34464 & n34465 ) | ( ~n34466 & n34465 ) ;
  assign n34471 = n33951 &  n34223 ;
  assign n34472 = n34222 &  n34471 ;
  assign n34460 = x92 | n33951 ;
  assign n34461 = x92 &  n33951 ;
  assign n34462 = ( n34460 & ~n34461 ) | ( n34460 & 1'b0 ) | ( ~n34461 & 1'b0 ) ;
  assign n34474 = ( n34187 & n34224 ) | ( n34187 & n34462 ) | ( n34224 & n34462 ) ;
  assign n34473 = n34187 | n34462 ;
  assign n34475 = ( n34472 & ~n34474 ) | ( n34472 & n34473 ) | ( ~n34474 & n34473 ) ;
  assign n34479 = n33959 &  n34223 ;
  assign n34480 = n34222 &  n34479 ;
  assign n34468 = x91 | n33959 ;
  assign n34469 = x91 &  n33959 ;
  assign n34470 = ( n34468 & ~n34469 ) | ( n34468 & 1'b0 ) | ( ~n34469 & 1'b0 ) ;
  assign n34482 = ( n34186 & n34224 ) | ( n34186 & n34470 ) | ( n34224 & n34470 ) ;
  assign n34481 = n34186 | n34470 ;
  assign n34483 = ( n34480 & ~n34482 ) | ( n34480 & n34481 ) | ( ~n34482 & n34481 ) ;
  assign n34487 = n33967 &  n34223 ;
  assign n34488 = n34222 &  n34487 ;
  assign n34476 = x90 | n33967 ;
  assign n34477 = x90 &  n33967 ;
  assign n34478 = ( n34476 & ~n34477 ) | ( n34476 & 1'b0 ) | ( ~n34477 & 1'b0 ) ;
  assign n34490 = ( n34185 & n34224 ) | ( n34185 & n34478 ) | ( n34224 & n34478 ) ;
  assign n34489 = n34185 | n34478 ;
  assign n34491 = ( n34488 & ~n34490 ) | ( n34488 & n34489 ) | ( ~n34490 & n34489 ) ;
  assign n34495 = n33975 &  n34223 ;
  assign n34496 = n34222 &  n34495 ;
  assign n34484 = x89 | n33975 ;
  assign n34485 = x89 &  n33975 ;
  assign n34486 = ( n34484 & ~n34485 ) | ( n34484 & 1'b0 ) | ( ~n34485 & 1'b0 ) ;
  assign n34498 = ( n34184 & n34224 ) | ( n34184 & n34486 ) | ( n34224 & n34486 ) ;
  assign n34497 = n34184 | n34486 ;
  assign n34499 = ( n34496 & ~n34498 ) | ( n34496 & n34497 ) | ( ~n34498 & n34497 ) ;
  assign n34503 = n33983 &  n34223 ;
  assign n34504 = n34222 &  n34503 ;
  assign n34492 = x88 | n33983 ;
  assign n34493 = x88 &  n33983 ;
  assign n34494 = ( n34492 & ~n34493 ) | ( n34492 & 1'b0 ) | ( ~n34493 & 1'b0 ) ;
  assign n34506 = ( n34183 & n34224 ) | ( n34183 & n34494 ) | ( n34224 & n34494 ) ;
  assign n34505 = n34183 | n34494 ;
  assign n34507 = ( n34504 & ~n34506 ) | ( n34504 & n34505 ) | ( ~n34506 & n34505 ) ;
  assign n34511 = n33991 &  n34223 ;
  assign n34512 = n34222 &  n34511 ;
  assign n34500 = x87 | n33991 ;
  assign n34501 = x87 &  n33991 ;
  assign n34502 = ( n34500 & ~n34501 ) | ( n34500 & 1'b0 ) | ( ~n34501 & 1'b0 ) ;
  assign n34514 = ( n34182 & n34224 ) | ( n34182 & n34502 ) | ( n34224 & n34502 ) ;
  assign n34513 = n34182 | n34502 ;
  assign n34515 = ( n34512 & ~n34514 ) | ( n34512 & n34513 ) | ( ~n34514 & n34513 ) ;
  assign n34519 = n33999 &  n34223 ;
  assign n34520 = n34222 &  n34519 ;
  assign n34508 = x86 | n33999 ;
  assign n34509 = x86 &  n33999 ;
  assign n34510 = ( n34508 & ~n34509 ) | ( n34508 & 1'b0 ) | ( ~n34509 & 1'b0 ) ;
  assign n34522 = ( n34181 & n34224 ) | ( n34181 & n34510 ) | ( n34224 & n34510 ) ;
  assign n34521 = n34181 | n34510 ;
  assign n34523 = ( n34520 & ~n34522 ) | ( n34520 & n34521 ) | ( ~n34522 & n34521 ) ;
  assign n34527 = n34007 &  n34223 ;
  assign n34528 = n34222 &  n34527 ;
  assign n34516 = x85 | n34007 ;
  assign n34517 = x85 &  n34007 ;
  assign n34518 = ( n34516 & ~n34517 ) | ( n34516 & 1'b0 ) | ( ~n34517 & 1'b0 ) ;
  assign n34530 = ( n34180 & n34224 ) | ( n34180 & n34518 ) | ( n34224 & n34518 ) ;
  assign n34529 = n34180 | n34518 ;
  assign n34531 = ( n34528 & ~n34530 ) | ( n34528 & n34529 ) | ( ~n34530 & n34529 ) ;
  assign n34535 = n34015 &  n34223 ;
  assign n34536 = n34222 &  n34535 ;
  assign n34524 = x84 | n34015 ;
  assign n34525 = x84 &  n34015 ;
  assign n34526 = ( n34524 & ~n34525 ) | ( n34524 & 1'b0 ) | ( ~n34525 & 1'b0 ) ;
  assign n34538 = ( n34179 & n34224 ) | ( n34179 & n34526 ) | ( n34224 & n34526 ) ;
  assign n34537 = n34179 | n34526 ;
  assign n34539 = ( n34536 & ~n34538 ) | ( n34536 & n34537 ) | ( ~n34538 & n34537 ) ;
  assign n34543 = n34023 &  n34223 ;
  assign n34544 = n34222 &  n34543 ;
  assign n34532 = x83 | n34023 ;
  assign n34533 = x83 &  n34023 ;
  assign n34534 = ( n34532 & ~n34533 ) | ( n34532 & 1'b0 ) | ( ~n34533 & 1'b0 ) ;
  assign n34546 = ( n34178 & n34224 ) | ( n34178 & n34534 ) | ( n34224 & n34534 ) ;
  assign n34545 = n34178 | n34534 ;
  assign n34547 = ( n34544 & ~n34546 ) | ( n34544 & n34545 ) | ( ~n34546 & n34545 ) ;
  assign n34551 = n34031 &  n34223 ;
  assign n34552 = n34222 &  n34551 ;
  assign n34540 = x82 | n34031 ;
  assign n34541 = x82 &  n34031 ;
  assign n34542 = ( n34540 & ~n34541 ) | ( n34540 & 1'b0 ) | ( ~n34541 & 1'b0 ) ;
  assign n34554 = ( n34177 & n34224 ) | ( n34177 & n34542 ) | ( n34224 & n34542 ) ;
  assign n34553 = n34177 | n34542 ;
  assign n34555 = ( n34552 & ~n34554 ) | ( n34552 & n34553 ) | ( ~n34554 & n34553 ) ;
  assign n34559 = n34039 &  n34223 ;
  assign n34560 = n34222 &  n34559 ;
  assign n34548 = x81 | n34039 ;
  assign n34549 = x81 &  n34039 ;
  assign n34550 = ( n34548 & ~n34549 ) | ( n34548 & 1'b0 ) | ( ~n34549 & 1'b0 ) ;
  assign n34562 = ( n34176 & n34224 ) | ( n34176 & n34550 ) | ( n34224 & n34550 ) ;
  assign n34561 = n34176 | n34550 ;
  assign n34563 = ( n34560 & ~n34562 ) | ( n34560 & n34561 ) | ( ~n34562 & n34561 ) ;
  assign n34567 = n34047 &  n34223 ;
  assign n34568 = n34222 &  n34567 ;
  assign n34556 = x80 | n34047 ;
  assign n34557 = x80 &  n34047 ;
  assign n34558 = ( n34556 & ~n34557 ) | ( n34556 & 1'b0 ) | ( ~n34557 & 1'b0 ) ;
  assign n34570 = ( n34175 & n34224 ) | ( n34175 & n34558 ) | ( n34224 & n34558 ) ;
  assign n34569 = n34175 | n34558 ;
  assign n34571 = ( n34568 & ~n34570 ) | ( n34568 & n34569 ) | ( ~n34570 & n34569 ) ;
  assign n34575 = n34055 &  n34223 ;
  assign n34576 = n34222 &  n34575 ;
  assign n34564 = x79 | n34055 ;
  assign n34565 = x79 &  n34055 ;
  assign n34566 = ( n34564 & ~n34565 ) | ( n34564 & 1'b0 ) | ( ~n34565 & 1'b0 ) ;
  assign n34578 = ( n34174 & n34224 ) | ( n34174 & n34566 ) | ( n34224 & n34566 ) ;
  assign n34577 = n34174 | n34566 ;
  assign n34579 = ( n34576 & ~n34578 ) | ( n34576 & n34577 ) | ( ~n34578 & n34577 ) ;
  assign n34583 = n34063 &  n34223 ;
  assign n34584 = n34222 &  n34583 ;
  assign n34572 = x78 | n34063 ;
  assign n34573 = x78 &  n34063 ;
  assign n34574 = ( n34572 & ~n34573 ) | ( n34572 & 1'b0 ) | ( ~n34573 & 1'b0 ) ;
  assign n34586 = ( n34173 & n34224 ) | ( n34173 & n34574 ) | ( n34224 & n34574 ) ;
  assign n34585 = n34173 | n34574 ;
  assign n34587 = ( n34584 & ~n34586 ) | ( n34584 & n34585 ) | ( ~n34586 & n34585 ) ;
  assign n34591 = n34071 &  n34223 ;
  assign n34592 = n34222 &  n34591 ;
  assign n34580 = x77 | n34071 ;
  assign n34581 = x77 &  n34071 ;
  assign n34582 = ( n34580 & ~n34581 ) | ( n34580 & 1'b0 ) | ( ~n34581 & 1'b0 ) ;
  assign n34594 = ( n34172 & n34224 ) | ( n34172 & n34582 ) | ( n34224 & n34582 ) ;
  assign n34593 = n34172 | n34582 ;
  assign n34595 = ( n34592 & ~n34594 ) | ( n34592 & n34593 ) | ( ~n34594 & n34593 ) ;
  assign n34599 = n34079 &  n34223 ;
  assign n34600 = n34222 &  n34599 ;
  assign n34588 = x76 | n34079 ;
  assign n34589 = x76 &  n34079 ;
  assign n34590 = ( n34588 & ~n34589 ) | ( n34588 & 1'b0 ) | ( ~n34589 & 1'b0 ) ;
  assign n34602 = ( n34171 & n34224 ) | ( n34171 & n34590 ) | ( n34224 & n34590 ) ;
  assign n34601 = n34171 | n34590 ;
  assign n34603 = ( n34600 & ~n34602 ) | ( n34600 & n34601 ) | ( ~n34602 & n34601 ) ;
  assign n34607 = n34087 &  n34223 ;
  assign n34608 = n34222 &  n34607 ;
  assign n34596 = x75 | n34087 ;
  assign n34597 = x75 &  n34087 ;
  assign n34598 = ( n34596 & ~n34597 ) | ( n34596 & 1'b0 ) | ( ~n34597 & 1'b0 ) ;
  assign n34610 = ( n34170 & n34224 ) | ( n34170 & n34598 ) | ( n34224 & n34598 ) ;
  assign n34609 = n34170 | n34598 ;
  assign n34611 = ( n34608 & ~n34610 ) | ( n34608 & n34609 ) | ( ~n34610 & n34609 ) ;
  assign n34615 = n34095 &  n34223 ;
  assign n34616 = n34222 &  n34615 ;
  assign n34604 = x74 | n34095 ;
  assign n34605 = x74 &  n34095 ;
  assign n34606 = ( n34604 & ~n34605 ) | ( n34604 & 1'b0 ) | ( ~n34605 & 1'b0 ) ;
  assign n34618 = ( n34169 & n34224 ) | ( n34169 & n34606 ) | ( n34224 & n34606 ) ;
  assign n34617 = n34169 | n34606 ;
  assign n34619 = ( n34616 & ~n34618 ) | ( n34616 & n34617 ) | ( ~n34618 & n34617 ) ;
  assign n34623 = n34103 &  n34223 ;
  assign n34624 = n34222 &  n34623 ;
  assign n34612 = x73 | n34103 ;
  assign n34613 = x73 &  n34103 ;
  assign n34614 = ( n34612 & ~n34613 ) | ( n34612 & 1'b0 ) | ( ~n34613 & 1'b0 ) ;
  assign n34626 = ( n34168 & n34224 ) | ( n34168 & n34614 ) | ( n34224 & n34614 ) ;
  assign n34625 = n34168 | n34614 ;
  assign n34627 = ( n34624 & ~n34626 ) | ( n34624 & n34625 ) | ( ~n34626 & n34625 ) ;
  assign n34631 = n34111 &  n34223 ;
  assign n34632 = n34222 &  n34631 ;
  assign n34620 = x72 | n34111 ;
  assign n34621 = x72 &  n34111 ;
  assign n34622 = ( n34620 & ~n34621 ) | ( n34620 & 1'b0 ) | ( ~n34621 & 1'b0 ) ;
  assign n34634 = ( n34167 & n34224 ) | ( n34167 & n34622 ) | ( n34224 & n34622 ) ;
  assign n34633 = n34167 | n34622 ;
  assign n34635 = ( n34632 & ~n34634 ) | ( n34632 & n34633 ) | ( ~n34634 & n34633 ) ;
  assign n34639 = n34119 &  n34223 ;
  assign n34640 = n34222 &  n34639 ;
  assign n34628 = x71 | n34119 ;
  assign n34629 = x71 &  n34119 ;
  assign n34630 = ( n34628 & ~n34629 ) | ( n34628 & 1'b0 ) | ( ~n34629 & 1'b0 ) ;
  assign n34642 = ( n34166 & n34224 ) | ( n34166 & n34630 ) | ( n34224 & n34630 ) ;
  assign n34641 = n34166 | n34630 ;
  assign n34643 = ( n34640 & ~n34642 ) | ( n34640 & n34641 ) | ( ~n34642 & n34641 ) ;
  assign n34647 = n34127 &  n34223 ;
  assign n34648 = n34222 &  n34647 ;
  assign n34636 = x70 | n34127 ;
  assign n34637 = x70 &  n34127 ;
  assign n34638 = ( n34636 & ~n34637 ) | ( n34636 & 1'b0 ) | ( ~n34637 & 1'b0 ) ;
  assign n34650 = ( n34165 & n34224 ) | ( n34165 & n34638 ) | ( n34224 & n34638 ) ;
  assign n34649 = n34165 | n34638 ;
  assign n34651 = ( n34648 & ~n34650 ) | ( n34648 & n34649 ) | ( ~n34650 & n34649 ) ;
  assign n34655 = n34135 &  n34223 ;
  assign n34656 = n34222 &  n34655 ;
  assign n34644 = x69 | n34135 ;
  assign n34645 = x69 &  n34135 ;
  assign n34646 = ( n34644 & ~n34645 ) | ( n34644 & 1'b0 ) | ( ~n34645 & 1'b0 ) ;
  assign n34658 = ( n34164 & n34224 ) | ( n34164 & n34646 ) | ( n34224 & n34646 ) ;
  assign n34657 = n34164 | n34646 ;
  assign n34659 = ( n34656 & ~n34658 ) | ( n34656 & n34657 ) | ( ~n34658 & n34657 ) ;
  assign n34663 = n34143 &  n34223 ;
  assign n34664 = n34222 &  n34663 ;
  assign n34652 = x68 | n34143 ;
  assign n34653 = x68 &  n34143 ;
  assign n34654 = ( n34652 & ~n34653 ) | ( n34652 & 1'b0 ) | ( ~n34653 & 1'b0 ) ;
  assign n34666 = ( n34163 & n34224 ) | ( n34163 & n34654 ) | ( n34224 & n34654 ) ;
  assign n34665 = n34163 | n34654 ;
  assign n34667 = ( n34664 & ~n34666 ) | ( n34664 & n34665 ) | ( ~n34666 & n34665 ) ;
  assign n34671 = n34148 &  n34223 ;
  assign n34672 = n34222 &  n34671 ;
  assign n34660 = x67 | n34148 ;
  assign n34661 = x67 &  n34148 ;
  assign n34662 = ( n34660 & ~n34661 ) | ( n34660 & 1'b0 ) | ( ~n34661 & 1'b0 ) ;
  assign n34674 = ( n34162 & n34224 ) | ( n34162 & n34662 ) | ( n34224 & n34662 ) ;
  assign n34673 = n34162 | n34662 ;
  assign n34675 = ( n34672 & ~n34674 ) | ( n34672 & n34673 ) | ( ~n34674 & n34673 ) ;
  assign n34676 = n34156 &  n34223 ;
  assign n34677 = n34222 &  n34676 ;
  assign n34668 = x66 | n34156 ;
  assign n34669 = x66 &  n34156 ;
  assign n34670 = ( n34668 & ~n34669 ) | ( n34668 & 1'b0 ) | ( ~n34669 & 1'b0 ) ;
  assign n34679 = ( n34161 & n34224 ) | ( n34161 & n34670 ) | ( n34224 & n34670 ) ;
  assign n34678 = n34161 | n34670 ;
  assign n34680 = ( n34677 & ~n34679 ) | ( n34677 & n34678 ) | ( ~n34679 & n34678 ) ;
  assign n34681 = ( x65 & ~n15844 ) | ( x65 & n34160 ) | ( ~n15844 & n34160 ) ;
  assign n34682 = ( n34161 & ~x65 ) | ( n34161 & n34681 ) | ( ~x65 & n34681 ) ;
  assign n34683 = ~n34224 & n34682 ;
  assign n34684 = n34160 &  n34223 ;
  assign n34685 = n34222 &  n34684 ;
  assign n34686 = n34683 | n34685 ;
  assign n34687 = ( x64 & ~n34224 ) | ( x64 & 1'b0 ) | ( ~n34224 & 1'b0 ) ;
  assign n34688 = ( x5 & ~n34687 ) | ( x5 & 1'b0 ) | ( ~n34687 & 1'b0 ) ;
  assign n34689 = ( n15844 & ~n34224 ) | ( n15844 & 1'b0 ) | ( ~n34224 & 1'b0 ) ;
  assign n34690 = n34688 | n34689 ;
  assign n34691 = ( x65 & ~n34690 ) | ( x65 & n16378 ) | ( ~n34690 & n16378 ) ;
  assign n34692 = ( x66 & ~n34686 ) | ( x66 & n34691 ) | ( ~n34686 & n34691 ) ;
  assign n34693 = ( x67 & ~n34680 ) | ( x67 & n34692 ) | ( ~n34680 & n34692 ) ;
  assign n34694 = ( x68 & ~n34675 ) | ( x68 & n34693 ) | ( ~n34675 & n34693 ) ;
  assign n34695 = ( x69 & ~n34667 ) | ( x69 & n34694 ) | ( ~n34667 & n34694 ) ;
  assign n34696 = ( x70 & ~n34659 ) | ( x70 & n34695 ) | ( ~n34659 & n34695 ) ;
  assign n34697 = ( x71 & ~n34651 ) | ( x71 & n34696 ) | ( ~n34651 & n34696 ) ;
  assign n34698 = ( x72 & ~n34643 ) | ( x72 & n34697 ) | ( ~n34643 & n34697 ) ;
  assign n34699 = ( x73 & ~n34635 ) | ( x73 & n34698 ) | ( ~n34635 & n34698 ) ;
  assign n34700 = ( x74 & ~n34627 ) | ( x74 & n34699 ) | ( ~n34627 & n34699 ) ;
  assign n34701 = ( x75 & ~n34619 ) | ( x75 & n34700 ) | ( ~n34619 & n34700 ) ;
  assign n34702 = ( x76 & ~n34611 ) | ( x76 & n34701 ) | ( ~n34611 & n34701 ) ;
  assign n34703 = ( x77 & ~n34603 ) | ( x77 & n34702 ) | ( ~n34603 & n34702 ) ;
  assign n34704 = ( x78 & ~n34595 ) | ( x78 & n34703 ) | ( ~n34595 & n34703 ) ;
  assign n34705 = ( x79 & ~n34587 ) | ( x79 & n34704 ) | ( ~n34587 & n34704 ) ;
  assign n34706 = ( x80 & ~n34579 ) | ( x80 & n34705 ) | ( ~n34579 & n34705 ) ;
  assign n34707 = ( x81 & ~n34571 ) | ( x81 & n34706 ) | ( ~n34571 & n34706 ) ;
  assign n34708 = ( x82 & ~n34563 ) | ( x82 & n34707 ) | ( ~n34563 & n34707 ) ;
  assign n34709 = ( x83 & ~n34555 ) | ( x83 & n34708 ) | ( ~n34555 & n34708 ) ;
  assign n34710 = ( x84 & ~n34547 ) | ( x84 & n34709 ) | ( ~n34547 & n34709 ) ;
  assign n34711 = ( x85 & ~n34539 ) | ( x85 & n34710 ) | ( ~n34539 & n34710 ) ;
  assign n34712 = ( x86 & ~n34531 ) | ( x86 & n34711 ) | ( ~n34531 & n34711 ) ;
  assign n34713 = ( x87 & ~n34523 ) | ( x87 & n34712 ) | ( ~n34523 & n34712 ) ;
  assign n34714 = ( x88 & ~n34515 ) | ( x88 & n34713 ) | ( ~n34515 & n34713 ) ;
  assign n34715 = ( x89 & ~n34507 ) | ( x89 & n34714 ) | ( ~n34507 & n34714 ) ;
  assign n34716 = ( x90 & ~n34499 ) | ( x90 & n34715 ) | ( ~n34499 & n34715 ) ;
  assign n34717 = ( x91 & ~n34491 ) | ( x91 & n34716 ) | ( ~n34491 & n34716 ) ;
  assign n34718 = ( x92 & ~n34483 ) | ( x92 & n34717 ) | ( ~n34483 & n34717 ) ;
  assign n34719 = ( x93 & ~n34475 ) | ( x93 & n34718 ) | ( ~n34475 & n34718 ) ;
  assign n34720 = ( x94 & ~n34467 ) | ( x94 & n34719 ) | ( ~n34467 & n34719 ) ;
  assign n34721 = ( x95 & ~n34459 ) | ( x95 & n34720 ) | ( ~n34459 & n34720 ) ;
  assign n34722 = ( x96 & ~n34451 ) | ( x96 & n34721 ) | ( ~n34451 & n34721 ) ;
  assign n34723 = ( x97 & ~n34443 ) | ( x97 & n34722 ) | ( ~n34443 & n34722 ) ;
  assign n34724 = ( x98 & ~n34435 ) | ( x98 & n34723 ) | ( ~n34435 & n34723 ) ;
  assign n34725 = ( x99 & ~n34427 ) | ( x99 & n34724 ) | ( ~n34427 & n34724 ) ;
  assign n34726 = ( x100 & ~n34419 ) | ( x100 & n34725 ) | ( ~n34419 & n34725 ) ;
  assign n34727 = ( x101 & ~n34411 ) | ( x101 & n34726 ) | ( ~n34411 & n34726 ) ;
  assign n34728 = ( x102 & ~n34403 ) | ( x102 & n34727 ) | ( ~n34403 & n34727 ) ;
  assign n34729 = ( x103 & ~n34395 ) | ( x103 & n34728 ) | ( ~n34395 & n34728 ) ;
  assign n34730 = ( x104 & ~n34387 ) | ( x104 & n34729 ) | ( ~n34387 & n34729 ) ;
  assign n34731 = ( x105 & ~n34379 ) | ( x105 & n34730 ) | ( ~n34379 & n34730 ) ;
  assign n34732 = ( x106 & ~n34371 ) | ( x106 & n34731 ) | ( ~n34371 & n34731 ) ;
  assign n34733 = ( x107 & ~n34363 ) | ( x107 & n34732 ) | ( ~n34363 & n34732 ) ;
  assign n34734 = ( x108 & ~n34355 ) | ( x108 & n34733 ) | ( ~n34355 & n34733 ) ;
  assign n34735 = ( x109 & ~n34347 ) | ( x109 & n34734 ) | ( ~n34347 & n34734 ) ;
  assign n34736 = ( x110 & ~n34339 ) | ( x110 & n34735 ) | ( ~n34339 & n34735 ) ;
  assign n34737 = ( x111 & ~n34331 ) | ( x111 & n34736 ) | ( ~n34331 & n34736 ) ;
  assign n34738 = ( x112 & ~n34323 ) | ( x112 & n34737 ) | ( ~n34323 & n34737 ) ;
  assign n34739 = ( x113 & ~n34315 ) | ( x113 & n34738 ) | ( ~n34315 & n34738 ) ;
  assign n34740 = ( x114 & ~n34307 ) | ( x114 & n34739 ) | ( ~n34307 & n34739 ) ;
  assign n34741 = ( x115 & ~n34299 ) | ( x115 & n34740 ) | ( ~n34299 & n34740 ) ;
  assign n34742 = ( x116 & ~n34291 ) | ( x116 & n34741 ) | ( ~n34291 & n34741 ) ;
  assign n34743 = ( x117 & ~n34283 ) | ( x117 & n34742 ) | ( ~n34283 & n34742 ) ;
  assign n34744 = ( x118 & ~n34275 ) | ( x118 & n34743 ) | ( ~n34275 & n34743 ) ;
  assign n34745 = ( x119 & ~n34267 ) | ( x119 & n34744 ) | ( ~n34267 & n34744 ) ;
  assign n34746 = ( x120 & ~n34259 ) | ( x120 & n34745 ) | ( ~n34259 & n34745 ) ;
  assign n34747 = ( x121 & ~n34251 ) | ( x121 & n34746 ) | ( ~n34251 & n34746 ) ;
  assign n34748 = ( x122 & ~n34243 ) | ( x122 & n34747 ) | ( ~n34243 & n34747 ) ;
  assign n34228 = n33711 | n34219 ;
  assign n34229 = ( n34217 & ~n34228 ) | ( n34217 & 1'b0 ) | ( ~n34228 & 1'b0 ) ;
  assign n34230 = ~n34217 & n34228 ;
  assign n34231 = ( n34229 & ~n34224 ) | ( n34229 & n34230 ) | ( ~n34224 & n34230 ) ;
  assign n34232 = n15415 &  n33205 ;
  assign n34233 = n34222 &  n34232 ;
  assign n34234 = n34231 | n34233 ;
  assign n34235 = ~x123 & n34234 ;
  assign n34749 = ( x123 & ~n34233 ) | ( x123 & 1'b0 ) | ( ~n34233 & 1'b0 ) ;
  assign n34750 = ~n34231 & n34749 ;
  assign n34759 = n34235 | n34750 ;
  assign n34760 = ( n34748 & ~n34759 ) | ( n34748 & 1'b0 ) | ( ~n34759 & 1'b0 ) ;
  assign n34751 = ( n34748 & ~n34235 ) | ( n34748 & n34750 ) | ( ~n34235 & n34750 ) ;
  assign n34752 = ( n34235 & ~n152 ) | ( n34235 & n34751 ) | ( ~n152 & n34751 ) ;
  assign n34753 = n152 | n34752 ;
  assign n34754 = ~n34234 |  n15943 ;
  assign n34755 = n34753 &  n34754 ;
  assign n34761 = ~n34748 & n34759 ;
  assign n34762 = ( n34760 & ~n34755 ) | ( n34760 & n34761 ) | ( ~n34755 & n34761 ) ;
  assign n34763 = n15943 &  n34234 ;
  assign n34764 = n34753 &  n34763 ;
  assign n34765 = n34762 | n34764 ;
  assign n34766 = ~x124 & n34765 ;
  assign n34770 = n34243 &  n34754 ;
  assign n34771 = n34753 &  n34770 ;
  assign n34756 = x122 | n34243 ;
  assign n34757 = x122 &  n34243 ;
  assign n34758 = ( n34756 & ~n34757 ) | ( n34756 & 1'b0 ) | ( ~n34757 & 1'b0 ) ;
  assign n34773 = ( n34747 & n34755 ) | ( n34747 & n34758 ) | ( n34755 & n34758 ) ;
  assign n34772 = n34747 | n34758 ;
  assign n34774 = ( n34771 & ~n34773 ) | ( n34771 & n34772 ) | ( ~n34773 & n34772 ) ;
  assign n34778 = n34251 &  n34754 ;
  assign n34779 = n34753 &  n34778 ;
  assign n34767 = x121 | n34251 ;
  assign n34768 = x121 &  n34251 ;
  assign n34769 = ( n34767 & ~n34768 ) | ( n34767 & 1'b0 ) | ( ~n34768 & 1'b0 ) ;
  assign n34781 = ( n34746 & n34755 ) | ( n34746 & n34769 ) | ( n34755 & n34769 ) ;
  assign n34780 = n34746 | n34769 ;
  assign n34782 = ( n34779 & ~n34781 ) | ( n34779 & n34780 ) | ( ~n34781 & n34780 ) ;
  assign n34786 = n34259 &  n34754 ;
  assign n34787 = n34753 &  n34786 ;
  assign n34775 = x120 | n34259 ;
  assign n34776 = x120 &  n34259 ;
  assign n34777 = ( n34775 & ~n34776 ) | ( n34775 & 1'b0 ) | ( ~n34776 & 1'b0 ) ;
  assign n34789 = ( n34745 & n34755 ) | ( n34745 & n34777 ) | ( n34755 & n34777 ) ;
  assign n34788 = n34745 | n34777 ;
  assign n34790 = ( n34787 & ~n34789 ) | ( n34787 & n34788 ) | ( ~n34789 & n34788 ) ;
  assign n34794 = n34267 &  n34754 ;
  assign n34795 = n34753 &  n34794 ;
  assign n34783 = x119 | n34267 ;
  assign n34784 = x119 &  n34267 ;
  assign n34785 = ( n34783 & ~n34784 ) | ( n34783 & 1'b0 ) | ( ~n34784 & 1'b0 ) ;
  assign n34797 = ( n34744 & n34755 ) | ( n34744 & n34785 ) | ( n34755 & n34785 ) ;
  assign n34796 = n34744 | n34785 ;
  assign n34798 = ( n34795 & ~n34797 ) | ( n34795 & n34796 ) | ( ~n34797 & n34796 ) ;
  assign n34802 = n34275 &  n34754 ;
  assign n34803 = n34753 &  n34802 ;
  assign n34791 = x118 | n34275 ;
  assign n34792 = x118 &  n34275 ;
  assign n34793 = ( n34791 & ~n34792 ) | ( n34791 & 1'b0 ) | ( ~n34792 & 1'b0 ) ;
  assign n34805 = ( n34743 & n34755 ) | ( n34743 & n34793 ) | ( n34755 & n34793 ) ;
  assign n34804 = n34743 | n34793 ;
  assign n34806 = ( n34803 & ~n34805 ) | ( n34803 & n34804 ) | ( ~n34805 & n34804 ) ;
  assign n34810 = n34283 &  n34754 ;
  assign n34811 = n34753 &  n34810 ;
  assign n34799 = x117 | n34283 ;
  assign n34800 = x117 &  n34283 ;
  assign n34801 = ( n34799 & ~n34800 ) | ( n34799 & 1'b0 ) | ( ~n34800 & 1'b0 ) ;
  assign n34813 = ( n34742 & n34755 ) | ( n34742 & n34801 ) | ( n34755 & n34801 ) ;
  assign n34812 = n34742 | n34801 ;
  assign n34814 = ( n34811 & ~n34813 ) | ( n34811 & n34812 ) | ( ~n34813 & n34812 ) ;
  assign n34818 = n34291 &  n34754 ;
  assign n34819 = n34753 &  n34818 ;
  assign n34807 = x116 | n34291 ;
  assign n34808 = x116 &  n34291 ;
  assign n34809 = ( n34807 & ~n34808 ) | ( n34807 & 1'b0 ) | ( ~n34808 & 1'b0 ) ;
  assign n34821 = ( n34741 & n34755 ) | ( n34741 & n34809 ) | ( n34755 & n34809 ) ;
  assign n34820 = n34741 | n34809 ;
  assign n34822 = ( n34819 & ~n34821 ) | ( n34819 & n34820 ) | ( ~n34821 & n34820 ) ;
  assign n34826 = n34299 &  n34754 ;
  assign n34827 = n34753 &  n34826 ;
  assign n34815 = x115 | n34299 ;
  assign n34816 = x115 &  n34299 ;
  assign n34817 = ( n34815 & ~n34816 ) | ( n34815 & 1'b0 ) | ( ~n34816 & 1'b0 ) ;
  assign n34829 = ( n34740 & n34755 ) | ( n34740 & n34817 ) | ( n34755 & n34817 ) ;
  assign n34828 = n34740 | n34817 ;
  assign n34830 = ( n34827 & ~n34829 ) | ( n34827 & n34828 ) | ( ~n34829 & n34828 ) ;
  assign n34834 = n34307 &  n34754 ;
  assign n34835 = n34753 &  n34834 ;
  assign n34823 = x114 | n34307 ;
  assign n34824 = x114 &  n34307 ;
  assign n34825 = ( n34823 & ~n34824 ) | ( n34823 & 1'b0 ) | ( ~n34824 & 1'b0 ) ;
  assign n34837 = ( n34739 & n34755 ) | ( n34739 & n34825 ) | ( n34755 & n34825 ) ;
  assign n34836 = n34739 | n34825 ;
  assign n34838 = ( n34835 & ~n34837 ) | ( n34835 & n34836 ) | ( ~n34837 & n34836 ) ;
  assign n34842 = n34315 &  n34754 ;
  assign n34843 = n34753 &  n34842 ;
  assign n34831 = x113 | n34315 ;
  assign n34832 = x113 &  n34315 ;
  assign n34833 = ( n34831 & ~n34832 ) | ( n34831 & 1'b0 ) | ( ~n34832 & 1'b0 ) ;
  assign n34845 = ( n34738 & n34755 ) | ( n34738 & n34833 ) | ( n34755 & n34833 ) ;
  assign n34844 = n34738 | n34833 ;
  assign n34846 = ( n34843 & ~n34845 ) | ( n34843 & n34844 ) | ( ~n34845 & n34844 ) ;
  assign n34850 = n34323 &  n34754 ;
  assign n34851 = n34753 &  n34850 ;
  assign n34839 = x112 | n34323 ;
  assign n34840 = x112 &  n34323 ;
  assign n34841 = ( n34839 & ~n34840 ) | ( n34839 & 1'b0 ) | ( ~n34840 & 1'b0 ) ;
  assign n34853 = ( n34737 & n34755 ) | ( n34737 & n34841 ) | ( n34755 & n34841 ) ;
  assign n34852 = n34737 | n34841 ;
  assign n34854 = ( n34851 & ~n34853 ) | ( n34851 & n34852 ) | ( ~n34853 & n34852 ) ;
  assign n34858 = n34331 &  n34754 ;
  assign n34859 = n34753 &  n34858 ;
  assign n34847 = x111 | n34331 ;
  assign n34848 = x111 &  n34331 ;
  assign n34849 = ( n34847 & ~n34848 ) | ( n34847 & 1'b0 ) | ( ~n34848 & 1'b0 ) ;
  assign n34861 = ( n34736 & n34755 ) | ( n34736 & n34849 ) | ( n34755 & n34849 ) ;
  assign n34860 = n34736 | n34849 ;
  assign n34862 = ( n34859 & ~n34861 ) | ( n34859 & n34860 ) | ( ~n34861 & n34860 ) ;
  assign n34866 = n34339 &  n34754 ;
  assign n34867 = n34753 &  n34866 ;
  assign n34855 = x110 | n34339 ;
  assign n34856 = x110 &  n34339 ;
  assign n34857 = ( n34855 & ~n34856 ) | ( n34855 & 1'b0 ) | ( ~n34856 & 1'b0 ) ;
  assign n34869 = ( n34735 & n34755 ) | ( n34735 & n34857 ) | ( n34755 & n34857 ) ;
  assign n34868 = n34735 | n34857 ;
  assign n34870 = ( n34867 & ~n34869 ) | ( n34867 & n34868 ) | ( ~n34869 & n34868 ) ;
  assign n34874 = n34347 &  n34754 ;
  assign n34875 = n34753 &  n34874 ;
  assign n34863 = x109 | n34347 ;
  assign n34864 = x109 &  n34347 ;
  assign n34865 = ( n34863 & ~n34864 ) | ( n34863 & 1'b0 ) | ( ~n34864 & 1'b0 ) ;
  assign n34877 = ( n34734 & n34755 ) | ( n34734 & n34865 ) | ( n34755 & n34865 ) ;
  assign n34876 = n34734 | n34865 ;
  assign n34878 = ( n34875 & ~n34877 ) | ( n34875 & n34876 ) | ( ~n34877 & n34876 ) ;
  assign n34882 = n34355 &  n34754 ;
  assign n34883 = n34753 &  n34882 ;
  assign n34871 = x108 | n34355 ;
  assign n34872 = x108 &  n34355 ;
  assign n34873 = ( n34871 & ~n34872 ) | ( n34871 & 1'b0 ) | ( ~n34872 & 1'b0 ) ;
  assign n34885 = ( n34733 & n34755 ) | ( n34733 & n34873 ) | ( n34755 & n34873 ) ;
  assign n34884 = n34733 | n34873 ;
  assign n34886 = ( n34883 & ~n34885 ) | ( n34883 & n34884 ) | ( ~n34885 & n34884 ) ;
  assign n34890 = n34363 &  n34754 ;
  assign n34891 = n34753 &  n34890 ;
  assign n34879 = x107 | n34363 ;
  assign n34880 = x107 &  n34363 ;
  assign n34881 = ( n34879 & ~n34880 ) | ( n34879 & 1'b0 ) | ( ~n34880 & 1'b0 ) ;
  assign n34893 = ( n34732 & n34755 ) | ( n34732 & n34881 ) | ( n34755 & n34881 ) ;
  assign n34892 = n34732 | n34881 ;
  assign n34894 = ( n34891 & ~n34893 ) | ( n34891 & n34892 ) | ( ~n34893 & n34892 ) ;
  assign n34898 = n34371 &  n34754 ;
  assign n34899 = n34753 &  n34898 ;
  assign n34887 = x106 | n34371 ;
  assign n34888 = x106 &  n34371 ;
  assign n34889 = ( n34887 & ~n34888 ) | ( n34887 & 1'b0 ) | ( ~n34888 & 1'b0 ) ;
  assign n34901 = ( n34731 & n34755 ) | ( n34731 & n34889 ) | ( n34755 & n34889 ) ;
  assign n34900 = n34731 | n34889 ;
  assign n34902 = ( n34899 & ~n34901 ) | ( n34899 & n34900 ) | ( ~n34901 & n34900 ) ;
  assign n34906 = n34379 &  n34754 ;
  assign n34907 = n34753 &  n34906 ;
  assign n34895 = x105 | n34379 ;
  assign n34896 = x105 &  n34379 ;
  assign n34897 = ( n34895 & ~n34896 ) | ( n34895 & 1'b0 ) | ( ~n34896 & 1'b0 ) ;
  assign n34909 = ( n34730 & n34755 ) | ( n34730 & n34897 ) | ( n34755 & n34897 ) ;
  assign n34908 = n34730 | n34897 ;
  assign n34910 = ( n34907 & ~n34909 ) | ( n34907 & n34908 ) | ( ~n34909 & n34908 ) ;
  assign n34914 = n34387 &  n34754 ;
  assign n34915 = n34753 &  n34914 ;
  assign n34903 = x104 | n34387 ;
  assign n34904 = x104 &  n34387 ;
  assign n34905 = ( n34903 & ~n34904 ) | ( n34903 & 1'b0 ) | ( ~n34904 & 1'b0 ) ;
  assign n34917 = ( n34729 & n34755 ) | ( n34729 & n34905 ) | ( n34755 & n34905 ) ;
  assign n34916 = n34729 | n34905 ;
  assign n34918 = ( n34915 & ~n34917 ) | ( n34915 & n34916 ) | ( ~n34917 & n34916 ) ;
  assign n34922 = n34395 &  n34754 ;
  assign n34923 = n34753 &  n34922 ;
  assign n34911 = x103 | n34395 ;
  assign n34912 = x103 &  n34395 ;
  assign n34913 = ( n34911 & ~n34912 ) | ( n34911 & 1'b0 ) | ( ~n34912 & 1'b0 ) ;
  assign n34925 = ( n34728 & n34755 ) | ( n34728 & n34913 ) | ( n34755 & n34913 ) ;
  assign n34924 = n34728 | n34913 ;
  assign n34926 = ( n34923 & ~n34925 ) | ( n34923 & n34924 ) | ( ~n34925 & n34924 ) ;
  assign n34930 = n34403 &  n34754 ;
  assign n34931 = n34753 &  n34930 ;
  assign n34919 = x102 | n34403 ;
  assign n34920 = x102 &  n34403 ;
  assign n34921 = ( n34919 & ~n34920 ) | ( n34919 & 1'b0 ) | ( ~n34920 & 1'b0 ) ;
  assign n34933 = ( n34727 & n34755 ) | ( n34727 & n34921 ) | ( n34755 & n34921 ) ;
  assign n34932 = n34727 | n34921 ;
  assign n34934 = ( n34931 & ~n34933 ) | ( n34931 & n34932 ) | ( ~n34933 & n34932 ) ;
  assign n34938 = n34411 &  n34754 ;
  assign n34939 = n34753 &  n34938 ;
  assign n34927 = x101 | n34411 ;
  assign n34928 = x101 &  n34411 ;
  assign n34929 = ( n34927 & ~n34928 ) | ( n34927 & 1'b0 ) | ( ~n34928 & 1'b0 ) ;
  assign n34941 = ( n34726 & n34755 ) | ( n34726 & n34929 ) | ( n34755 & n34929 ) ;
  assign n34940 = n34726 | n34929 ;
  assign n34942 = ( n34939 & ~n34941 ) | ( n34939 & n34940 ) | ( ~n34941 & n34940 ) ;
  assign n34946 = n34419 &  n34754 ;
  assign n34947 = n34753 &  n34946 ;
  assign n34935 = x100 | n34419 ;
  assign n34936 = x100 &  n34419 ;
  assign n34937 = ( n34935 & ~n34936 ) | ( n34935 & 1'b0 ) | ( ~n34936 & 1'b0 ) ;
  assign n34949 = ( n34725 & n34755 ) | ( n34725 & n34937 ) | ( n34755 & n34937 ) ;
  assign n34948 = n34725 | n34937 ;
  assign n34950 = ( n34947 & ~n34949 ) | ( n34947 & n34948 ) | ( ~n34949 & n34948 ) ;
  assign n34954 = n34427 &  n34754 ;
  assign n34955 = n34753 &  n34954 ;
  assign n34943 = x99 | n34427 ;
  assign n34944 = x99 &  n34427 ;
  assign n34945 = ( n34943 & ~n34944 ) | ( n34943 & 1'b0 ) | ( ~n34944 & 1'b0 ) ;
  assign n34957 = ( n34724 & n34755 ) | ( n34724 & n34945 ) | ( n34755 & n34945 ) ;
  assign n34956 = n34724 | n34945 ;
  assign n34958 = ( n34955 & ~n34957 ) | ( n34955 & n34956 ) | ( ~n34957 & n34956 ) ;
  assign n34962 = n34435 &  n34754 ;
  assign n34963 = n34753 &  n34962 ;
  assign n34951 = x98 | n34435 ;
  assign n34952 = x98 &  n34435 ;
  assign n34953 = ( n34951 & ~n34952 ) | ( n34951 & 1'b0 ) | ( ~n34952 & 1'b0 ) ;
  assign n34965 = ( n34723 & n34755 ) | ( n34723 & n34953 ) | ( n34755 & n34953 ) ;
  assign n34964 = n34723 | n34953 ;
  assign n34966 = ( n34963 & ~n34965 ) | ( n34963 & n34964 ) | ( ~n34965 & n34964 ) ;
  assign n34970 = n34443 &  n34754 ;
  assign n34971 = n34753 &  n34970 ;
  assign n34959 = x97 | n34443 ;
  assign n34960 = x97 &  n34443 ;
  assign n34961 = ( n34959 & ~n34960 ) | ( n34959 & 1'b0 ) | ( ~n34960 & 1'b0 ) ;
  assign n34973 = ( n34722 & n34755 ) | ( n34722 & n34961 ) | ( n34755 & n34961 ) ;
  assign n34972 = n34722 | n34961 ;
  assign n34974 = ( n34971 & ~n34973 ) | ( n34971 & n34972 ) | ( ~n34973 & n34972 ) ;
  assign n34978 = n34451 &  n34754 ;
  assign n34979 = n34753 &  n34978 ;
  assign n34967 = x96 | n34451 ;
  assign n34968 = x96 &  n34451 ;
  assign n34969 = ( n34967 & ~n34968 ) | ( n34967 & 1'b0 ) | ( ~n34968 & 1'b0 ) ;
  assign n34981 = ( n34721 & n34755 ) | ( n34721 & n34969 ) | ( n34755 & n34969 ) ;
  assign n34980 = n34721 | n34969 ;
  assign n34982 = ( n34979 & ~n34981 ) | ( n34979 & n34980 ) | ( ~n34981 & n34980 ) ;
  assign n34986 = n34459 &  n34754 ;
  assign n34987 = n34753 &  n34986 ;
  assign n34975 = x95 | n34459 ;
  assign n34976 = x95 &  n34459 ;
  assign n34977 = ( n34975 & ~n34976 ) | ( n34975 & 1'b0 ) | ( ~n34976 & 1'b0 ) ;
  assign n34989 = ( n34720 & n34755 ) | ( n34720 & n34977 ) | ( n34755 & n34977 ) ;
  assign n34988 = n34720 | n34977 ;
  assign n34990 = ( n34987 & ~n34989 ) | ( n34987 & n34988 ) | ( ~n34989 & n34988 ) ;
  assign n34994 = n34467 &  n34754 ;
  assign n34995 = n34753 &  n34994 ;
  assign n34983 = x94 | n34467 ;
  assign n34984 = x94 &  n34467 ;
  assign n34985 = ( n34983 & ~n34984 ) | ( n34983 & 1'b0 ) | ( ~n34984 & 1'b0 ) ;
  assign n34997 = ( n34719 & n34755 ) | ( n34719 & n34985 ) | ( n34755 & n34985 ) ;
  assign n34996 = n34719 | n34985 ;
  assign n34998 = ( n34995 & ~n34997 ) | ( n34995 & n34996 ) | ( ~n34997 & n34996 ) ;
  assign n35002 = n34475 &  n34754 ;
  assign n35003 = n34753 &  n35002 ;
  assign n34991 = x93 | n34475 ;
  assign n34992 = x93 &  n34475 ;
  assign n34993 = ( n34991 & ~n34992 ) | ( n34991 & 1'b0 ) | ( ~n34992 & 1'b0 ) ;
  assign n35005 = ( n34718 & n34755 ) | ( n34718 & n34993 ) | ( n34755 & n34993 ) ;
  assign n35004 = n34718 | n34993 ;
  assign n35006 = ( n35003 & ~n35005 ) | ( n35003 & n35004 ) | ( ~n35005 & n35004 ) ;
  assign n35010 = n34483 &  n34754 ;
  assign n35011 = n34753 &  n35010 ;
  assign n34999 = x92 | n34483 ;
  assign n35000 = x92 &  n34483 ;
  assign n35001 = ( n34999 & ~n35000 ) | ( n34999 & 1'b0 ) | ( ~n35000 & 1'b0 ) ;
  assign n35013 = ( n34717 & n34755 ) | ( n34717 & n35001 ) | ( n34755 & n35001 ) ;
  assign n35012 = n34717 | n35001 ;
  assign n35014 = ( n35011 & ~n35013 ) | ( n35011 & n35012 ) | ( ~n35013 & n35012 ) ;
  assign n35018 = n34491 &  n34754 ;
  assign n35019 = n34753 &  n35018 ;
  assign n35007 = x91 | n34491 ;
  assign n35008 = x91 &  n34491 ;
  assign n35009 = ( n35007 & ~n35008 ) | ( n35007 & 1'b0 ) | ( ~n35008 & 1'b0 ) ;
  assign n35021 = ( n34716 & n34755 ) | ( n34716 & n35009 ) | ( n34755 & n35009 ) ;
  assign n35020 = n34716 | n35009 ;
  assign n35022 = ( n35019 & ~n35021 ) | ( n35019 & n35020 ) | ( ~n35021 & n35020 ) ;
  assign n35026 = n34499 &  n34754 ;
  assign n35027 = n34753 &  n35026 ;
  assign n35015 = x90 | n34499 ;
  assign n35016 = x90 &  n34499 ;
  assign n35017 = ( n35015 & ~n35016 ) | ( n35015 & 1'b0 ) | ( ~n35016 & 1'b0 ) ;
  assign n35029 = ( n34715 & n34755 ) | ( n34715 & n35017 ) | ( n34755 & n35017 ) ;
  assign n35028 = n34715 | n35017 ;
  assign n35030 = ( n35027 & ~n35029 ) | ( n35027 & n35028 ) | ( ~n35029 & n35028 ) ;
  assign n35034 = n34507 &  n34754 ;
  assign n35035 = n34753 &  n35034 ;
  assign n35023 = x89 | n34507 ;
  assign n35024 = x89 &  n34507 ;
  assign n35025 = ( n35023 & ~n35024 ) | ( n35023 & 1'b0 ) | ( ~n35024 & 1'b0 ) ;
  assign n35037 = ( n34714 & n34755 ) | ( n34714 & n35025 ) | ( n34755 & n35025 ) ;
  assign n35036 = n34714 | n35025 ;
  assign n35038 = ( n35035 & ~n35037 ) | ( n35035 & n35036 ) | ( ~n35037 & n35036 ) ;
  assign n35042 = n34515 &  n34754 ;
  assign n35043 = n34753 &  n35042 ;
  assign n35031 = x88 | n34515 ;
  assign n35032 = x88 &  n34515 ;
  assign n35033 = ( n35031 & ~n35032 ) | ( n35031 & 1'b0 ) | ( ~n35032 & 1'b0 ) ;
  assign n35045 = ( n34713 & n34755 ) | ( n34713 & n35033 ) | ( n34755 & n35033 ) ;
  assign n35044 = n34713 | n35033 ;
  assign n35046 = ( n35043 & ~n35045 ) | ( n35043 & n35044 ) | ( ~n35045 & n35044 ) ;
  assign n35050 = n34523 &  n34754 ;
  assign n35051 = n34753 &  n35050 ;
  assign n35039 = x87 | n34523 ;
  assign n35040 = x87 &  n34523 ;
  assign n35041 = ( n35039 & ~n35040 ) | ( n35039 & 1'b0 ) | ( ~n35040 & 1'b0 ) ;
  assign n35053 = ( n34712 & n34755 ) | ( n34712 & n35041 ) | ( n34755 & n35041 ) ;
  assign n35052 = n34712 | n35041 ;
  assign n35054 = ( n35051 & ~n35053 ) | ( n35051 & n35052 ) | ( ~n35053 & n35052 ) ;
  assign n35058 = n34531 &  n34754 ;
  assign n35059 = n34753 &  n35058 ;
  assign n35047 = x86 | n34531 ;
  assign n35048 = x86 &  n34531 ;
  assign n35049 = ( n35047 & ~n35048 ) | ( n35047 & 1'b0 ) | ( ~n35048 & 1'b0 ) ;
  assign n35061 = ( n34711 & n34755 ) | ( n34711 & n35049 ) | ( n34755 & n35049 ) ;
  assign n35060 = n34711 | n35049 ;
  assign n35062 = ( n35059 & ~n35061 ) | ( n35059 & n35060 ) | ( ~n35061 & n35060 ) ;
  assign n35066 = n34539 &  n34754 ;
  assign n35067 = n34753 &  n35066 ;
  assign n35055 = x85 | n34539 ;
  assign n35056 = x85 &  n34539 ;
  assign n35057 = ( n35055 & ~n35056 ) | ( n35055 & 1'b0 ) | ( ~n35056 & 1'b0 ) ;
  assign n35069 = ( n34710 & n34755 ) | ( n34710 & n35057 ) | ( n34755 & n35057 ) ;
  assign n35068 = n34710 | n35057 ;
  assign n35070 = ( n35067 & ~n35069 ) | ( n35067 & n35068 ) | ( ~n35069 & n35068 ) ;
  assign n35074 = n34547 &  n34754 ;
  assign n35075 = n34753 &  n35074 ;
  assign n35063 = x84 | n34547 ;
  assign n35064 = x84 &  n34547 ;
  assign n35065 = ( n35063 & ~n35064 ) | ( n35063 & 1'b0 ) | ( ~n35064 & 1'b0 ) ;
  assign n35077 = ( n34709 & n34755 ) | ( n34709 & n35065 ) | ( n34755 & n35065 ) ;
  assign n35076 = n34709 | n35065 ;
  assign n35078 = ( n35075 & ~n35077 ) | ( n35075 & n35076 ) | ( ~n35077 & n35076 ) ;
  assign n35082 = n34555 &  n34754 ;
  assign n35083 = n34753 &  n35082 ;
  assign n35071 = x83 | n34555 ;
  assign n35072 = x83 &  n34555 ;
  assign n35073 = ( n35071 & ~n35072 ) | ( n35071 & 1'b0 ) | ( ~n35072 & 1'b0 ) ;
  assign n35085 = ( n34708 & n34755 ) | ( n34708 & n35073 ) | ( n34755 & n35073 ) ;
  assign n35084 = n34708 | n35073 ;
  assign n35086 = ( n35083 & ~n35085 ) | ( n35083 & n35084 ) | ( ~n35085 & n35084 ) ;
  assign n35090 = n34563 &  n34754 ;
  assign n35091 = n34753 &  n35090 ;
  assign n35079 = x82 | n34563 ;
  assign n35080 = x82 &  n34563 ;
  assign n35081 = ( n35079 & ~n35080 ) | ( n35079 & 1'b0 ) | ( ~n35080 & 1'b0 ) ;
  assign n35093 = ( n34707 & n34755 ) | ( n34707 & n35081 ) | ( n34755 & n35081 ) ;
  assign n35092 = n34707 | n35081 ;
  assign n35094 = ( n35091 & ~n35093 ) | ( n35091 & n35092 ) | ( ~n35093 & n35092 ) ;
  assign n35098 = n34571 &  n34754 ;
  assign n35099 = n34753 &  n35098 ;
  assign n35087 = x81 | n34571 ;
  assign n35088 = x81 &  n34571 ;
  assign n35089 = ( n35087 & ~n35088 ) | ( n35087 & 1'b0 ) | ( ~n35088 & 1'b0 ) ;
  assign n35101 = ( n34706 & n34755 ) | ( n34706 & n35089 ) | ( n34755 & n35089 ) ;
  assign n35100 = n34706 | n35089 ;
  assign n35102 = ( n35099 & ~n35101 ) | ( n35099 & n35100 ) | ( ~n35101 & n35100 ) ;
  assign n35106 = n34579 &  n34754 ;
  assign n35107 = n34753 &  n35106 ;
  assign n35095 = x80 | n34579 ;
  assign n35096 = x80 &  n34579 ;
  assign n35097 = ( n35095 & ~n35096 ) | ( n35095 & 1'b0 ) | ( ~n35096 & 1'b0 ) ;
  assign n35109 = ( n34705 & n34755 ) | ( n34705 & n35097 ) | ( n34755 & n35097 ) ;
  assign n35108 = n34705 | n35097 ;
  assign n35110 = ( n35107 & ~n35109 ) | ( n35107 & n35108 ) | ( ~n35109 & n35108 ) ;
  assign n35114 = n34587 &  n34754 ;
  assign n35115 = n34753 &  n35114 ;
  assign n35103 = x79 | n34587 ;
  assign n35104 = x79 &  n34587 ;
  assign n35105 = ( n35103 & ~n35104 ) | ( n35103 & 1'b0 ) | ( ~n35104 & 1'b0 ) ;
  assign n35117 = ( n34704 & n34755 ) | ( n34704 & n35105 ) | ( n34755 & n35105 ) ;
  assign n35116 = n34704 | n35105 ;
  assign n35118 = ( n35115 & ~n35117 ) | ( n35115 & n35116 ) | ( ~n35117 & n35116 ) ;
  assign n35122 = n34595 &  n34754 ;
  assign n35123 = n34753 &  n35122 ;
  assign n35111 = x78 | n34595 ;
  assign n35112 = x78 &  n34595 ;
  assign n35113 = ( n35111 & ~n35112 ) | ( n35111 & 1'b0 ) | ( ~n35112 & 1'b0 ) ;
  assign n35125 = ( n34703 & n34755 ) | ( n34703 & n35113 ) | ( n34755 & n35113 ) ;
  assign n35124 = n34703 | n35113 ;
  assign n35126 = ( n35123 & ~n35125 ) | ( n35123 & n35124 ) | ( ~n35125 & n35124 ) ;
  assign n35130 = n34603 &  n34754 ;
  assign n35131 = n34753 &  n35130 ;
  assign n35119 = x77 | n34603 ;
  assign n35120 = x77 &  n34603 ;
  assign n35121 = ( n35119 & ~n35120 ) | ( n35119 & 1'b0 ) | ( ~n35120 & 1'b0 ) ;
  assign n35133 = ( n34702 & n34755 ) | ( n34702 & n35121 ) | ( n34755 & n35121 ) ;
  assign n35132 = n34702 | n35121 ;
  assign n35134 = ( n35131 & ~n35133 ) | ( n35131 & n35132 ) | ( ~n35133 & n35132 ) ;
  assign n35138 = n34611 &  n34754 ;
  assign n35139 = n34753 &  n35138 ;
  assign n35127 = x76 | n34611 ;
  assign n35128 = x76 &  n34611 ;
  assign n35129 = ( n35127 & ~n35128 ) | ( n35127 & 1'b0 ) | ( ~n35128 & 1'b0 ) ;
  assign n35141 = ( n34701 & n34755 ) | ( n34701 & n35129 ) | ( n34755 & n35129 ) ;
  assign n35140 = n34701 | n35129 ;
  assign n35142 = ( n35139 & ~n35141 ) | ( n35139 & n35140 ) | ( ~n35141 & n35140 ) ;
  assign n35146 = n34619 &  n34754 ;
  assign n35147 = n34753 &  n35146 ;
  assign n35135 = x75 | n34619 ;
  assign n35136 = x75 &  n34619 ;
  assign n35137 = ( n35135 & ~n35136 ) | ( n35135 & 1'b0 ) | ( ~n35136 & 1'b0 ) ;
  assign n35149 = ( n34700 & n34755 ) | ( n34700 & n35137 ) | ( n34755 & n35137 ) ;
  assign n35148 = n34700 | n35137 ;
  assign n35150 = ( n35147 & ~n35149 ) | ( n35147 & n35148 ) | ( ~n35149 & n35148 ) ;
  assign n35154 = n34627 &  n34754 ;
  assign n35155 = n34753 &  n35154 ;
  assign n35143 = x74 | n34627 ;
  assign n35144 = x74 &  n34627 ;
  assign n35145 = ( n35143 & ~n35144 ) | ( n35143 & 1'b0 ) | ( ~n35144 & 1'b0 ) ;
  assign n35157 = ( n34699 & n34755 ) | ( n34699 & n35145 ) | ( n34755 & n35145 ) ;
  assign n35156 = n34699 | n35145 ;
  assign n35158 = ( n35155 & ~n35157 ) | ( n35155 & n35156 ) | ( ~n35157 & n35156 ) ;
  assign n35162 = n34635 &  n34754 ;
  assign n35163 = n34753 &  n35162 ;
  assign n35151 = x73 | n34635 ;
  assign n35152 = x73 &  n34635 ;
  assign n35153 = ( n35151 & ~n35152 ) | ( n35151 & 1'b0 ) | ( ~n35152 & 1'b0 ) ;
  assign n35165 = ( n34698 & n34755 ) | ( n34698 & n35153 ) | ( n34755 & n35153 ) ;
  assign n35164 = n34698 | n35153 ;
  assign n35166 = ( n35163 & ~n35165 ) | ( n35163 & n35164 ) | ( ~n35165 & n35164 ) ;
  assign n35170 = n34643 &  n34754 ;
  assign n35171 = n34753 &  n35170 ;
  assign n35159 = x72 | n34643 ;
  assign n35160 = x72 &  n34643 ;
  assign n35161 = ( n35159 & ~n35160 ) | ( n35159 & 1'b0 ) | ( ~n35160 & 1'b0 ) ;
  assign n35173 = ( n34697 & n34755 ) | ( n34697 & n35161 ) | ( n34755 & n35161 ) ;
  assign n35172 = n34697 | n35161 ;
  assign n35174 = ( n35171 & ~n35173 ) | ( n35171 & n35172 ) | ( ~n35173 & n35172 ) ;
  assign n35178 = n34651 &  n34754 ;
  assign n35179 = n34753 &  n35178 ;
  assign n35167 = x71 | n34651 ;
  assign n35168 = x71 &  n34651 ;
  assign n35169 = ( n35167 & ~n35168 ) | ( n35167 & 1'b0 ) | ( ~n35168 & 1'b0 ) ;
  assign n35181 = ( n34696 & n34755 ) | ( n34696 & n35169 ) | ( n34755 & n35169 ) ;
  assign n35180 = n34696 | n35169 ;
  assign n35182 = ( n35179 & ~n35181 ) | ( n35179 & n35180 ) | ( ~n35181 & n35180 ) ;
  assign n35186 = n34659 &  n34754 ;
  assign n35187 = n34753 &  n35186 ;
  assign n35175 = x70 | n34659 ;
  assign n35176 = x70 &  n34659 ;
  assign n35177 = ( n35175 & ~n35176 ) | ( n35175 & 1'b0 ) | ( ~n35176 & 1'b0 ) ;
  assign n35189 = ( n34695 & n34755 ) | ( n34695 & n35177 ) | ( n34755 & n35177 ) ;
  assign n35188 = n34695 | n35177 ;
  assign n35190 = ( n35187 & ~n35189 ) | ( n35187 & n35188 ) | ( ~n35189 & n35188 ) ;
  assign n35194 = n34667 &  n34754 ;
  assign n35195 = n34753 &  n35194 ;
  assign n35183 = x69 | n34667 ;
  assign n35184 = x69 &  n34667 ;
  assign n35185 = ( n35183 & ~n35184 ) | ( n35183 & 1'b0 ) | ( ~n35184 & 1'b0 ) ;
  assign n35197 = ( n34694 & n34755 ) | ( n34694 & n35185 ) | ( n34755 & n35185 ) ;
  assign n35196 = n34694 | n35185 ;
  assign n35198 = ( n35195 & ~n35197 ) | ( n35195 & n35196 ) | ( ~n35197 & n35196 ) ;
  assign n35202 = n34675 &  n34754 ;
  assign n35203 = n34753 &  n35202 ;
  assign n35191 = x68 | n34675 ;
  assign n35192 = x68 &  n34675 ;
  assign n35193 = ( n35191 & ~n35192 ) | ( n35191 & 1'b0 ) | ( ~n35192 & 1'b0 ) ;
  assign n35205 = ( n34693 & n34755 ) | ( n34693 & n35193 ) | ( n34755 & n35193 ) ;
  assign n35204 = n34693 | n35193 ;
  assign n35206 = ( n35203 & ~n35205 ) | ( n35203 & n35204 ) | ( ~n35205 & n35204 ) ;
  assign n35210 = n34680 &  n34754 ;
  assign n35211 = n34753 &  n35210 ;
  assign n35199 = x67 | n34680 ;
  assign n35200 = x67 &  n34680 ;
  assign n35201 = ( n35199 & ~n35200 ) | ( n35199 & 1'b0 ) | ( ~n35200 & 1'b0 ) ;
  assign n35213 = ( n34692 & n34755 ) | ( n34692 & n35201 ) | ( n34755 & n35201 ) ;
  assign n35212 = n34692 | n35201 ;
  assign n35214 = ( n35211 & ~n35213 ) | ( n35211 & n35212 ) | ( ~n35213 & n35212 ) ;
  assign n35215 = n34686 &  n34754 ;
  assign n35216 = n34753 &  n35215 ;
  assign n35207 = x66 | n34686 ;
  assign n35208 = x66 &  n34686 ;
  assign n35209 = ( n35207 & ~n35208 ) | ( n35207 & 1'b0 ) | ( ~n35208 & 1'b0 ) ;
  assign n35217 = n34691 &  n35209 ;
  assign n35218 = ( n34691 & ~n34755 ) | ( n34691 & n35209 ) | ( ~n34755 & n35209 ) ;
  assign n35219 = ( n35216 & ~n35217 ) | ( n35216 & n35218 ) | ( ~n35217 & n35218 ) ;
  assign n35220 = ( x65 & ~n16378 ) | ( x65 & n34690 ) | ( ~n16378 & n34690 ) ;
  assign n35221 = ( n34691 & ~x65 ) | ( n34691 & n35220 ) | ( ~x65 & n35220 ) ;
  assign n35222 = ~n34755 & n35221 ;
  assign n35223 = n34690 &  n34754 ;
  assign n35224 = n34753 &  n35223 ;
  assign n35225 = n35222 | n35224 ;
  assign n35226 = ( x64 & ~n34755 ) | ( x64 & 1'b0 ) | ( ~n34755 & 1'b0 ) ;
  assign n35227 = ( x4 & ~n35226 ) | ( x4 & 1'b0 ) | ( ~n35226 & 1'b0 ) ;
  assign n35228 = ( n16378 & ~n34755 ) | ( n16378 & 1'b0 ) | ( ~n34755 & 1'b0 ) ;
  assign n35229 = n35227 | n35228 ;
  assign n35230 = ( x65 & ~n35229 ) | ( x65 & n16926 ) | ( ~n35229 & n16926 ) ;
  assign n35231 = ( x66 & ~n35225 ) | ( x66 & n35230 ) | ( ~n35225 & n35230 ) ;
  assign n35232 = ( x67 & ~n35219 ) | ( x67 & n35231 ) | ( ~n35219 & n35231 ) ;
  assign n35233 = ( x68 & ~n35214 ) | ( x68 & n35232 ) | ( ~n35214 & n35232 ) ;
  assign n35234 = ( x69 & ~n35206 ) | ( x69 & n35233 ) | ( ~n35206 & n35233 ) ;
  assign n35235 = ( x70 & ~n35198 ) | ( x70 & n35234 ) | ( ~n35198 & n35234 ) ;
  assign n35236 = ( x71 & ~n35190 ) | ( x71 & n35235 ) | ( ~n35190 & n35235 ) ;
  assign n35237 = ( x72 & ~n35182 ) | ( x72 & n35236 ) | ( ~n35182 & n35236 ) ;
  assign n35238 = ( x73 & ~n35174 ) | ( x73 & n35237 ) | ( ~n35174 & n35237 ) ;
  assign n35239 = ( x74 & ~n35166 ) | ( x74 & n35238 ) | ( ~n35166 & n35238 ) ;
  assign n35240 = ( x75 & ~n35158 ) | ( x75 & n35239 ) | ( ~n35158 & n35239 ) ;
  assign n35241 = ( x76 & ~n35150 ) | ( x76 & n35240 ) | ( ~n35150 & n35240 ) ;
  assign n35242 = ( x77 & ~n35142 ) | ( x77 & n35241 ) | ( ~n35142 & n35241 ) ;
  assign n35243 = ( x78 & ~n35134 ) | ( x78 & n35242 ) | ( ~n35134 & n35242 ) ;
  assign n35244 = ( x79 & ~n35126 ) | ( x79 & n35243 ) | ( ~n35126 & n35243 ) ;
  assign n35245 = ( x80 & ~n35118 ) | ( x80 & n35244 ) | ( ~n35118 & n35244 ) ;
  assign n35246 = ( x81 & ~n35110 ) | ( x81 & n35245 ) | ( ~n35110 & n35245 ) ;
  assign n35247 = ( x82 & ~n35102 ) | ( x82 & n35246 ) | ( ~n35102 & n35246 ) ;
  assign n35248 = ( x83 & ~n35094 ) | ( x83 & n35247 ) | ( ~n35094 & n35247 ) ;
  assign n35249 = ( x84 & ~n35086 ) | ( x84 & n35248 ) | ( ~n35086 & n35248 ) ;
  assign n35250 = ( x85 & ~n35078 ) | ( x85 & n35249 ) | ( ~n35078 & n35249 ) ;
  assign n35251 = ( x86 & ~n35070 ) | ( x86 & n35250 ) | ( ~n35070 & n35250 ) ;
  assign n35252 = ( x87 & ~n35062 ) | ( x87 & n35251 ) | ( ~n35062 & n35251 ) ;
  assign n35253 = ( x88 & ~n35054 ) | ( x88 & n35252 ) | ( ~n35054 & n35252 ) ;
  assign n35254 = ( x89 & ~n35046 ) | ( x89 & n35253 ) | ( ~n35046 & n35253 ) ;
  assign n35255 = ( x90 & ~n35038 ) | ( x90 & n35254 ) | ( ~n35038 & n35254 ) ;
  assign n35256 = ( x91 & ~n35030 ) | ( x91 & n35255 ) | ( ~n35030 & n35255 ) ;
  assign n35257 = ( x92 & ~n35022 ) | ( x92 & n35256 ) | ( ~n35022 & n35256 ) ;
  assign n35258 = ( x93 & ~n35014 ) | ( x93 & n35257 ) | ( ~n35014 & n35257 ) ;
  assign n35259 = ( x94 & ~n35006 ) | ( x94 & n35258 ) | ( ~n35006 & n35258 ) ;
  assign n35260 = ( x95 & ~n34998 ) | ( x95 & n35259 ) | ( ~n34998 & n35259 ) ;
  assign n35261 = ( x96 & ~n34990 ) | ( x96 & n35260 ) | ( ~n34990 & n35260 ) ;
  assign n35262 = ( x97 & ~n34982 ) | ( x97 & n35261 ) | ( ~n34982 & n35261 ) ;
  assign n35263 = ( x98 & ~n34974 ) | ( x98 & n35262 ) | ( ~n34974 & n35262 ) ;
  assign n35264 = ( x99 & ~n34966 ) | ( x99 & n35263 ) | ( ~n34966 & n35263 ) ;
  assign n35265 = ( x100 & ~n34958 ) | ( x100 & n35264 ) | ( ~n34958 & n35264 ) ;
  assign n35266 = ( x101 & ~n34950 ) | ( x101 & n35265 ) | ( ~n34950 & n35265 ) ;
  assign n35267 = ( x102 & ~n34942 ) | ( x102 & n35266 ) | ( ~n34942 & n35266 ) ;
  assign n35268 = ( x103 & ~n34934 ) | ( x103 & n35267 ) | ( ~n34934 & n35267 ) ;
  assign n35269 = ( x104 & ~n34926 ) | ( x104 & n35268 ) | ( ~n34926 & n35268 ) ;
  assign n35270 = ( x105 & ~n34918 ) | ( x105 & n35269 ) | ( ~n34918 & n35269 ) ;
  assign n35271 = ( x106 & ~n34910 ) | ( x106 & n35270 ) | ( ~n34910 & n35270 ) ;
  assign n35272 = ( x107 & ~n34902 ) | ( x107 & n35271 ) | ( ~n34902 & n35271 ) ;
  assign n35273 = ( x108 & ~n34894 ) | ( x108 & n35272 ) | ( ~n34894 & n35272 ) ;
  assign n35274 = ( x109 & ~n34886 ) | ( x109 & n35273 ) | ( ~n34886 & n35273 ) ;
  assign n35275 = ( x110 & ~n34878 ) | ( x110 & n35274 ) | ( ~n34878 & n35274 ) ;
  assign n35276 = ( x111 & ~n34870 ) | ( x111 & n35275 ) | ( ~n34870 & n35275 ) ;
  assign n35277 = ( x112 & ~n34862 ) | ( x112 & n35276 ) | ( ~n34862 & n35276 ) ;
  assign n35278 = ( x113 & ~n34854 ) | ( x113 & n35277 ) | ( ~n34854 & n35277 ) ;
  assign n35279 = ( x114 & ~n34846 ) | ( x114 & n35278 ) | ( ~n34846 & n35278 ) ;
  assign n35280 = ( x115 & ~n34838 ) | ( x115 & n35279 ) | ( ~n34838 & n35279 ) ;
  assign n35281 = ( x116 & ~n34830 ) | ( x116 & n35280 ) | ( ~n34830 & n35280 ) ;
  assign n35282 = ( x117 & ~n34822 ) | ( x117 & n35281 ) | ( ~n34822 & n35281 ) ;
  assign n35283 = ( x118 & ~n34814 ) | ( x118 & n35282 ) | ( ~n34814 & n35282 ) ;
  assign n35284 = ( x119 & ~n34806 ) | ( x119 & n35283 ) | ( ~n34806 & n35283 ) ;
  assign n35285 = ( x120 & ~n34798 ) | ( x120 & n35284 ) | ( ~n34798 & n35284 ) ;
  assign n35286 = ( x121 & ~n34790 ) | ( x121 & n35285 ) | ( ~n34790 & n35285 ) ;
  assign n35287 = ( x122 & ~n34782 ) | ( x122 & n35286 ) | ( ~n34782 & n35286 ) ;
  assign n35288 = ( x123 & ~n34774 ) | ( x123 & n35287 ) | ( ~n34774 & n35287 ) ;
  assign n35289 = ( x124 & ~n34764 ) | ( x124 & 1'b0 ) | ( ~n34764 & 1'b0 ) ;
  assign n35290 = ~n34762 & n35289 ;
  assign n35291 = ( n35288 & ~n34766 ) | ( n35288 & n35290 ) | ( ~n34766 & n35290 ) ;
  assign n35292 = ( n34766 & ~n235 ) | ( n34766 & n35291 ) | ( ~n235 & n35291 ) ;
  assign n35293 = n235 | n35292 ;
  assign n35294 = ~n34765 |  n152 ;
  assign n35310 = n34774 &  n35294 ;
  assign n35311 = n35293 &  n35310 ;
  assign n35295 = n35293 &  n35294 ;
  assign n35296 = x123 | n34774 ;
  assign n35297 = x123 &  n34774 ;
  assign n35298 = ( n35296 & ~n35297 ) | ( n35296 & 1'b0 ) | ( ~n35297 & 1'b0 ) ;
  assign n35313 = ( n35287 & n35295 ) | ( n35287 & n35298 ) | ( n35295 & n35298 ) ;
  assign n35312 = n35287 | n35298 ;
  assign n35314 = ( n35311 & ~n35313 ) | ( n35311 & n35312 ) | ( ~n35313 & n35312 ) ;
  assign n35318 = n34782 &  n35294 ;
  assign n35319 = n35293 &  n35318 ;
  assign n35307 = x122 | n34782 ;
  assign n35308 = x122 &  n34782 ;
  assign n35309 = ( n35307 & ~n35308 ) | ( n35307 & 1'b0 ) | ( ~n35308 & 1'b0 ) ;
  assign n35321 = ( n35286 & n35295 ) | ( n35286 & n35309 ) | ( n35295 & n35309 ) ;
  assign n35320 = n35286 | n35309 ;
  assign n35322 = ( n35319 & ~n35321 ) | ( n35319 & n35320 ) | ( ~n35321 & n35320 ) ;
  assign n35326 = n34790 &  n35294 ;
  assign n35327 = n35293 &  n35326 ;
  assign n35315 = x121 | n34790 ;
  assign n35316 = x121 &  n34790 ;
  assign n35317 = ( n35315 & ~n35316 ) | ( n35315 & 1'b0 ) | ( ~n35316 & 1'b0 ) ;
  assign n35329 = ( n35285 & n35295 ) | ( n35285 & n35317 ) | ( n35295 & n35317 ) ;
  assign n35328 = n35285 | n35317 ;
  assign n35330 = ( n35327 & ~n35329 ) | ( n35327 & n35328 ) | ( ~n35329 & n35328 ) ;
  assign n35334 = n34798 &  n35294 ;
  assign n35335 = n35293 &  n35334 ;
  assign n35323 = x120 | n34798 ;
  assign n35324 = x120 &  n34798 ;
  assign n35325 = ( n35323 & ~n35324 ) | ( n35323 & 1'b0 ) | ( ~n35324 & 1'b0 ) ;
  assign n35337 = ( n35284 & n35295 ) | ( n35284 & n35325 ) | ( n35295 & n35325 ) ;
  assign n35336 = n35284 | n35325 ;
  assign n35338 = ( n35335 & ~n35337 ) | ( n35335 & n35336 ) | ( ~n35337 & n35336 ) ;
  assign n35342 = n34806 &  n35294 ;
  assign n35343 = n35293 &  n35342 ;
  assign n35331 = x119 | n34806 ;
  assign n35332 = x119 &  n34806 ;
  assign n35333 = ( n35331 & ~n35332 ) | ( n35331 & 1'b0 ) | ( ~n35332 & 1'b0 ) ;
  assign n35345 = ( n35283 & n35295 ) | ( n35283 & n35333 ) | ( n35295 & n35333 ) ;
  assign n35344 = n35283 | n35333 ;
  assign n35346 = ( n35343 & ~n35345 ) | ( n35343 & n35344 ) | ( ~n35345 & n35344 ) ;
  assign n35350 = n34814 &  n35294 ;
  assign n35351 = n35293 &  n35350 ;
  assign n35339 = x118 | n34814 ;
  assign n35340 = x118 &  n34814 ;
  assign n35341 = ( n35339 & ~n35340 ) | ( n35339 & 1'b0 ) | ( ~n35340 & 1'b0 ) ;
  assign n35353 = ( n35282 & n35295 ) | ( n35282 & n35341 ) | ( n35295 & n35341 ) ;
  assign n35352 = n35282 | n35341 ;
  assign n35354 = ( n35351 & ~n35353 ) | ( n35351 & n35352 ) | ( ~n35353 & n35352 ) ;
  assign n35358 = n34822 &  n35294 ;
  assign n35359 = n35293 &  n35358 ;
  assign n35347 = x117 | n34822 ;
  assign n35348 = x117 &  n34822 ;
  assign n35349 = ( n35347 & ~n35348 ) | ( n35347 & 1'b0 ) | ( ~n35348 & 1'b0 ) ;
  assign n35361 = ( n35281 & n35295 ) | ( n35281 & n35349 ) | ( n35295 & n35349 ) ;
  assign n35360 = n35281 | n35349 ;
  assign n35362 = ( n35359 & ~n35361 ) | ( n35359 & n35360 ) | ( ~n35361 & n35360 ) ;
  assign n35366 = n34830 &  n35294 ;
  assign n35367 = n35293 &  n35366 ;
  assign n35355 = x116 | n34830 ;
  assign n35356 = x116 &  n34830 ;
  assign n35357 = ( n35355 & ~n35356 ) | ( n35355 & 1'b0 ) | ( ~n35356 & 1'b0 ) ;
  assign n35369 = ( n35280 & n35295 ) | ( n35280 & n35357 ) | ( n35295 & n35357 ) ;
  assign n35368 = n35280 | n35357 ;
  assign n35370 = ( n35367 & ~n35369 ) | ( n35367 & n35368 ) | ( ~n35369 & n35368 ) ;
  assign n35374 = n34838 &  n35294 ;
  assign n35375 = n35293 &  n35374 ;
  assign n35363 = x115 | n34838 ;
  assign n35364 = x115 &  n34838 ;
  assign n35365 = ( n35363 & ~n35364 ) | ( n35363 & 1'b0 ) | ( ~n35364 & 1'b0 ) ;
  assign n35377 = ( n35279 & n35295 ) | ( n35279 & n35365 ) | ( n35295 & n35365 ) ;
  assign n35376 = n35279 | n35365 ;
  assign n35378 = ( n35375 & ~n35377 ) | ( n35375 & n35376 ) | ( ~n35377 & n35376 ) ;
  assign n35382 = n34846 &  n35294 ;
  assign n35383 = n35293 &  n35382 ;
  assign n35371 = x114 | n34846 ;
  assign n35372 = x114 &  n34846 ;
  assign n35373 = ( n35371 & ~n35372 ) | ( n35371 & 1'b0 ) | ( ~n35372 & 1'b0 ) ;
  assign n35385 = ( n35278 & n35295 ) | ( n35278 & n35373 ) | ( n35295 & n35373 ) ;
  assign n35384 = n35278 | n35373 ;
  assign n35386 = ( n35383 & ~n35385 ) | ( n35383 & n35384 ) | ( ~n35385 & n35384 ) ;
  assign n35390 = n34854 &  n35294 ;
  assign n35391 = n35293 &  n35390 ;
  assign n35379 = x113 | n34854 ;
  assign n35380 = x113 &  n34854 ;
  assign n35381 = ( n35379 & ~n35380 ) | ( n35379 & 1'b0 ) | ( ~n35380 & 1'b0 ) ;
  assign n35393 = ( n35277 & n35295 ) | ( n35277 & n35381 ) | ( n35295 & n35381 ) ;
  assign n35392 = n35277 | n35381 ;
  assign n35394 = ( n35391 & ~n35393 ) | ( n35391 & n35392 ) | ( ~n35393 & n35392 ) ;
  assign n35398 = n34862 &  n35294 ;
  assign n35399 = n35293 &  n35398 ;
  assign n35387 = x112 | n34862 ;
  assign n35388 = x112 &  n34862 ;
  assign n35389 = ( n35387 & ~n35388 ) | ( n35387 & 1'b0 ) | ( ~n35388 & 1'b0 ) ;
  assign n35401 = ( n35276 & n35295 ) | ( n35276 & n35389 ) | ( n35295 & n35389 ) ;
  assign n35400 = n35276 | n35389 ;
  assign n35402 = ( n35399 & ~n35401 ) | ( n35399 & n35400 ) | ( ~n35401 & n35400 ) ;
  assign n35406 = n34870 &  n35294 ;
  assign n35407 = n35293 &  n35406 ;
  assign n35395 = x111 | n34870 ;
  assign n35396 = x111 &  n34870 ;
  assign n35397 = ( n35395 & ~n35396 ) | ( n35395 & 1'b0 ) | ( ~n35396 & 1'b0 ) ;
  assign n35409 = ( n35275 & n35295 ) | ( n35275 & n35397 ) | ( n35295 & n35397 ) ;
  assign n35408 = n35275 | n35397 ;
  assign n35410 = ( n35407 & ~n35409 ) | ( n35407 & n35408 ) | ( ~n35409 & n35408 ) ;
  assign n35414 = n34878 &  n35294 ;
  assign n35415 = n35293 &  n35414 ;
  assign n35403 = x110 | n34878 ;
  assign n35404 = x110 &  n34878 ;
  assign n35405 = ( n35403 & ~n35404 ) | ( n35403 & 1'b0 ) | ( ~n35404 & 1'b0 ) ;
  assign n35417 = ( n35274 & n35295 ) | ( n35274 & n35405 ) | ( n35295 & n35405 ) ;
  assign n35416 = n35274 | n35405 ;
  assign n35418 = ( n35415 & ~n35417 ) | ( n35415 & n35416 ) | ( ~n35417 & n35416 ) ;
  assign n35422 = n34886 &  n35294 ;
  assign n35423 = n35293 &  n35422 ;
  assign n35411 = x109 | n34886 ;
  assign n35412 = x109 &  n34886 ;
  assign n35413 = ( n35411 & ~n35412 ) | ( n35411 & 1'b0 ) | ( ~n35412 & 1'b0 ) ;
  assign n35425 = ( n35273 & n35295 ) | ( n35273 & n35413 ) | ( n35295 & n35413 ) ;
  assign n35424 = n35273 | n35413 ;
  assign n35426 = ( n35423 & ~n35425 ) | ( n35423 & n35424 ) | ( ~n35425 & n35424 ) ;
  assign n35430 = n34894 &  n35294 ;
  assign n35431 = n35293 &  n35430 ;
  assign n35419 = x108 | n34894 ;
  assign n35420 = x108 &  n34894 ;
  assign n35421 = ( n35419 & ~n35420 ) | ( n35419 & 1'b0 ) | ( ~n35420 & 1'b0 ) ;
  assign n35433 = ( n35272 & n35295 ) | ( n35272 & n35421 ) | ( n35295 & n35421 ) ;
  assign n35432 = n35272 | n35421 ;
  assign n35434 = ( n35431 & ~n35433 ) | ( n35431 & n35432 ) | ( ~n35433 & n35432 ) ;
  assign n35438 = n34902 &  n35294 ;
  assign n35439 = n35293 &  n35438 ;
  assign n35427 = x107 | n34902 ;
  assign n35428 = x107 &  n34902 ;
  assign n35429 = ( n35427 & ~n35428 ) | ( n35427 & 1'b0 ) | ( ~n35428 & 1'b0 ) ;
  assign n35441 = ( n35271 & n35295 ) | ( n35271 & n35429 ) | ( n35295 & n35429 ) ;
  assign n35440 = n35271 | n35429 ;
  assign n35442 = ( n35439 & ~n35441 ) | ( n35439 & n35440 ) | ( ~n35441 & n35440 ) ;
  assign n35446 = n34910 &  n35294 ;
  assign n35447 = n35293 &  n35446 ;
  assign n35435 = x106 | n34910 ;
  assign n35436 = x106 &  n34910 ;
  assign n35437 = ( n35435 & ~n35436 ) | ( n35435 & 1'b0 ) | ( ~n35436 & 1'b0 ) ;
  assign n35449 = ( n35270 & n35295 ) | ( n35270 & n35437 ) | ( n35295 & n35437 ) ;
  assign n35448 = n35270 | n35437 ;
  assign n35450 = ( n35447 & ~n35449 ) | ( n35447 & n35448 ) | ( ~n35449 & n35448 ) ;
  assign n35454 = n34918 &  n35294 ;
  assign n35455 = n35293 &  n35454 ;
  assign n35443 = x105 | n34918 ;
  assign n35444 = x105 &  n34918 ;
  assign n35445 = ( n35443 & ~n35444 ) | ( n35443 & 1'b0 ) | ( ~n35444 & 1'b0 ) ;
  assign n35457 = ( n35269 & n35295 ) | ( n35269 & n35445 ) | ( n35295 & n35445 ) ;
  assign n35456 = n35269 | n35445 ;
  assign n35458 = ( n35455 & ~n35457 ) | ( n35455 & n35456 ) | ( ~n35457 & n35456 ) ;
  assign n35462 = n34926 &  n35294 ;
  assign n35463 = n35293 &  n35462 ;
  assign n35451 = x104 | n34926 ;
  assign n35452 = x104 &  n34926 ;
  assign n35453 = ( n35451 & ~n35452 ) | ( n35451 & 1'b0 ) | ( ~n35452 & 1'b0 ) ;
  assign n35465 = ( n35268 & n35295 ) | ( n35268 & n35453 ) | ( n35295 & n35453 ) ;
  assign n35464 = n35268 | n35453 ;
  assign n35466 = ( n35463 & ~n35465 ) | ( n35463 & n35464 ) | ( ~n35465 & n35464 ) ;
  assign n35470 = n34934 &  n35294 ;
  assign n35471 = n35293 &  n35470 ;
  assign n35459 = x103 | n34934 ;
  assign n35460 = x103 &  n34934 ;
  assign n35461 = ( n35459 & ~n35460 ) | ( n35459 & 1'b0 ) | ( ~n35460 & 1'b0 ) ;
  assign n35473 = ( n35267 & n35295 ) | ( n35267 & n35461 ) | ( n35295 & n35461 ) ;
  assign n35472 = n35267 | n35461 ;
  assign n35474 = ( n35471 & ~n35473 ) | ( n35471 & n35472 ) | ( ~n35473 & n35472 ) ;
  assign n35478 = n34942 &  n35294 ;
  assign n35479 = n35293 &  n35478 ;
  assign n35467 = x102 | n34942 ;
  assign n35468 = x102 &  n34942 ;
  assign n35469 = ( n35467 & ~n35468 ) | ( n35467 & 1'b0 ) | ( ~n35468 & 1'b0 ) ;
  assign n35481 = ( n35266 & n35295 ) | ( n35266 & n35469 ) | ( n35295 & n35469 ) ;
  assign n35480 = n35266 | n35469 ;
  assign n35482 = ( n35479 & ~n35481 ) | ( n35479 & n35480 ) | ( ~n35481 & n35480 ) ;
  assign n35486 = n34950 &  n35294 ;
  assign n35487 = n35293 &  n35486 ;
  assign n35475 = x101 | n34950 ;
  assign n35476 = x101 &  n34950 ;
  assign n35477 = ( n35475 & ~n35476 ) | ( n35475 & 1'b0 ) | ( ~n35476 & 1'b0 ) ;
  assign n35489 = ( n35265 & n35295 ) | ( n35265 & n35477 ) | ( n35295 & n35477 ) ;
  assign n35488 = n35265 | n35477 ;
  assign n35490 = ( n35487 & ~n35489 ) | ( n35487 & n35488 ) | ( ~n35489 & n35488 ) ;
  assign n35494 = n34958 &  n35294 ;
  assign n35495 = n35293 &  n35494 ;
  assign n35483 = x100 | n34958 ;
  assign n35484 = x100 &  n34958 ;
  assign n35485 = ( n35483 & ~n35484 ) | ( n35483 & 1'b0 ) | ( ~n35484 & 1'b0 ) ;
  assign n35497 = ( n35264 & n35295 ) | ( n35264 & n35485 ) | ( n35295 & n35485 ) ;
  assign n35496 = n35264 | n35485 ;
  assign n35498 = ( n35495 & ~n35497 ) | ( n35495 & n35496 ) | ( ~n35497 & n35496 ) ;
  assign n35502 = n34966 &  n35294 ;
  assign n35503 = n35293 &  n35502 ;
  assign n35491 = x99 | n34966 ;
  assign n35492 = x99 &  n34966 ;
  assign n35493 = ( n35491 & ~n35492 ) | ( n35491 & 1'b0 ) | ( ~n35492 & 1'b0 ) ;
  assign n35505 = ( n35263 & n35295 ) | ( n35263 & n35493 ) | ( n35295 & n35493 ) ;
  assign n35504 = n35263 | n35493 ;
  assign n35506 = ( n35503 & ~n35505 ) | ( n35503 & n35504 ) | ( ~n35505 & n35504 ) ;
  assign n35510 = n34974 &  n35294 ;
  assign n35511 = n35293 &  n35510 ;
  assign n35499 = x98 | n34974 ;
  assign n35500 = x98 &  n34974 ;
  assign n35501 = ( n35499 & ~n35500 ) | ( n35499 & 1'b0 ) | ( ~n35500 & 1'b0 ) ;
  assign n35513 = ( n35262 & n35295 ) | ( n35262 & n35501 ) | ( n35295 & n35501 ) ;
  assign n35512 = n35262 | n35501 ;
  assign n35514 = ( n35511 & ~n35513 ) | ( n35511 & n35512 ) | ( ~n35513 & n35512 ) ;
  assign n35518 = n34982 &  n35294 ;
  assign n35519 = n35293 &  n35518 ;
  assign n35507 = x97 | n34982 ;
  assign n35508 = x97 &  n34982 ;
  assign n35509 = ( n35507 & ~n35508 ) | ( n35507 & 1'b0 ) | ( ~n35508 & 1'b0 ) ;
  assign n35521 = ( n35261 & n35295 ) | ( n35261 & n35509 ) | ( n35295 & n35509 ) ;
  assign n35520 = n35261 | n35509 ;
  assign n35522 = ( n35519 & ~n35521 ) | ( n35519 & n35520 ) | ( ~n35521 & n35520 ) ;
  assign n35526 = n34990 &  n35294 ;
  assign n35527 = n35293 &  n35526 ;
  assign n35515 = x96 | n34990 ;
  assign n35516 = x96 &  n34990 ;
  assign n35517 = ( n35515 & ~n35516 ) | ( n35515 & 1'b0 ) | ( ~n35516 & 1'b0 ) ;
  assign n35529 = ( n35260 & n35295 ) | ( n35260 & n35517 ) | ( n35295 & n35517 ) ;
  assign n35528 = n35260 | n35517 ;
  assign n35530 = ( n35527 & ~n35529 ) | ( n35527 & n35528 ) | ( ~n35529 & n35528 ) ;
  assign n35534 = n34998 &  n35294 ;
  assign n35535 = n35293 &  n35534 ;
  assign n35523 = x95 | n34998 ;
  assign n35524 = x95 &  n34998 ;
  assign n35525 = ( n35523 & ~n35524 ) | ( n35523 & 1'b0 ) | ( ~n35524 & 1'b0 ) ;
  assign n35537 = ( n35259 & n35295 ) | ( n35259 & n35525 ) | ( n35295 & n35525 ) ;
  assign n35536 = n35259 | n35525 ;
  assign n35538 = ( n35535 & ~n35537 ) | ( n35535 & n35536 ) | ( ~n35537 & n35536 ) ;
  assign n35542 = n35006 &  n35294 ;
  assign n35543 = n35293 &  n35542 ;
  assign n35531 = x94 | n35006 ;
  assign n35532 = x94 &  n35006 ;
  assign n35533 = ( n35531 & ~n35532 ) | ( n35531 & 1'b0 ) | ( ~n35532 & 1'b0 ) ;
  assign n35545 = ( n35258 & n35295 ) | ( n35258 & n35533 ) | ( n35295 & n35533 ) ;
  assign n35544 = n35258 | n35533 ;
  assign n35546 = ( n35543 & ~n35545 ) | ( n35543 & n35544 ) | ( ~n35545 & n35544 ) ;
  assign n35550 = n35014 &  n35294 ;
  assign n35551 = n35293 &  n35550 ;
  assign n35539 = x93 | n35014 ;
  assign n35540 = x93 &  n35014 ;
  assign n35541 = ( n35539 & ~n35540 ) | ( n35539 & 1'b0 ) | ( ~n35540 & 1'b0 ) ;
  assign n35553 = ( n35257 & n35295 ) | ( n35257 & n35541 ) | ( n35295 & n35541 ) ;
  assign n35552 = n35257 | n35541 ;
  assign n35554 = ( n35551 & ~n35553 ) | ( n35551 & n35552 ) | ( ~n35553 & n35552 ) ;
  assign n35558 = n35022 &  n35294 ;
  assign n35559 = n35293 &  n35558 ;
  assign n35547 = x92 | n35022 ;
  assign n35548 = x92 &  n35022 ;
  assign n35549 = ( n35547 & ~n35548 ) | ( n35547 & 1'b0 ) | ( ~n35548 & 1'b0 ) ;
  assign n35561 = ( n35256 & n35295 ) | ( n35256 & n35549 ) | ( n35295 & n35549 ) ;
  assign n35560 = n35256 | n35549 ;
  assign n35562 = ( n35559 & ~n35561 ) | ( n35559 & n35560 ) | ( ~n35561 & n35560 ) ;
  assign n35566 = n35030 &  n35294 ;
  assign n35567 = n35293 &  n35566 ;
  assign n35555 = x91 | n35030 ;
  assign n35556 = x91 &  n35030 ;
  assign n35557 = ( n35555 & ~n35556 ) | ( n35555 & 1'b0 ) | ( ~n35556 & 1'b0 ) ;
  assign n35569 = ( n35255 & n35295 ) | ( n35255 & n35557 ) | ( n35295 & n35557 ) ;
  assign n35568 = n35255 | n35557 ;
  assign n35570 = ( n35567 & ~n35569 ) | ( n35567 & n35568 ) | ( ~n35569 & n35568 ) ;
  assign n35574 = n35038 &  n35294 ;
  assign n35575 = n35293 &  n35574 ;
  assign n35563 = x90 | n35038 ;
  assign n35564 = x90 &  n35038 ;
  assign n35565 = ( n35563 & ~n35564 ) | ( n35563 & 1'b0 ) | ( ~n35564 & 1'b0 ) ;
  assign n35577 = ( n35254 & n35295 ) | ( n35254 & n35565 ) | ( n35295 & n35565 ) ;
  assign n35576 = n35254 | n35565 ;
  assign n35578 = ( n35575 & ~n35577 ) | ( n35575 & n35576 ) | ( ~n35577 & n35576 ) ;
  assign n35582 = n35046 &  n35294 ;
  assign n35583 = n35293 &  n35582 ;
  assign n35571 = x89 | n35046 ;
  assign n35572 = x89 &  n35046 ;
  assign n35573 = ( n35571 & ~n35572 ) | ( n35571 & 1'b0 ) | ( ~n35572 & 1'b0 ) ;
  assign n35585 = ( n35253 & n35295 ) | ( n35253 & n35573 ) | ( n35295 & n35573 ) ;
  assign n35584 = n35253 | n35573 ;
  assign n35586 = ( n35583 & ~n35585 ) | ( n35583 & n35584 ) | ( ~n35585 & n35584 ) ;
  assign n35590 = n35054 &  n35294 ;
  assign n35591 = n35293 &  n35590 ;
  assign n35579 = x88 | n35054 ;
  assign n35580 = x88 &  n35054 ;
  assign n35581 = ( n35579 & ~n35580 ) | ( n35579 & 1'b0 ) | ( ~n35580 & 1'b0 ) ;
  assign n35593 = ( n35252 & n35295 ) | ( n35252 & n35581 ) | ( n35295 & n35581 ) ;
  assign n35592 = n35252 | n35581 ;
  assign n35594 = ( n35591 & ~n35593 ) | ( n35591 & n35592 ) | ( ~n35593 & n35592 ) ;
  assign n35598 = n35062 &  n35294 ;
  assign n35599 = n35293 &  n35598 ;
  assign n35587 = x87 | n35062 ;
  assign n35588 = x87 &  n35062 ;
  assign n35589 = ( n35587 & ~n35588 ) | ( n35587 & 1'b0 ) | ( ~n35588 & 1'b0 ) ;
  assign n35601 = ( n35251 & n35295 ) | ( n35251 & n35589 ) | ( n35295 & n35589 ) ;
  assign n35600 = n35251 | n35589 ;
  assign n35602 = ( n35599 & ~n35601 ) | ( n35599 & n35600 ) | ( ~n35601 & n35600 ) ;
  assign n35606 = n35070 &  n35294 ;
  assign n35607 = n35293 &  n35606 ;
  assign n35595 = x86 | n35070 ;
  assign n35596 = x86 &  n35070 ;
  assign n35597 = ( n35595 & ~n35596 ) | ( n35595 & 1'b0 ) | ( ~n35596 & 1'b0 ) ;
  assign n35609 = ( n35250 & n35295 ) | ( n35250 & n35597 ) | ( n35295 & n35597 ) ;
  assign n35608 = n35250 | n35597 ;
  assign n35610 = ( n35607 & ~n35609 ) | ( n35607 & n35608 ) | ( ~n35609 & n35608 ) ;
  assign n35614 = n35078 &  n35294 ;
  assign n35615 = n35293 &  n35614 ;
  assign n35603 = x85 | n35078 ;
  assign n35604 = x85 &  n35078 ;
  assign n35605 = ( n35603 & ~n35604 ) | ( n35603 & 1'b0 ) | ( ~n35604 & 1'b0 ) ;
  assign n35617 = ( n35249 & n35295 ) | ( n35249 & n35605 ) | ( n35295 & n35605 ) ;
  assign n35616 = n35249 | n35605 ;
  assign n35618 = ( n35615 & ~n35617 ) | ( n35615 & n35616 ) | ( ~n35617 & n35616 ) ;
  assign n35622 = n35086 &  n35294 ;
  assign n35623 = n35293 &  n35622 ;
  assign n35611 = x84 | n35086 ;
  assign n35612 = x84 &  n35086 ;
  assign n35613 = ( n35611 & ~n35612 ) | ( n35611 & 1'b0 ) | ( ~n35612 & 1'b0 ) ;
  assign n35625 = ( n35248 & n35295 ) | ( n35248 & n35613 ) | ( n35295 & n35613 ) ;
  assign n35624 = n35248 | n35613 ;
  assign n35626 = ( n35623 & ~n35625 ) | ( n35623 & n35624 ) | ( ~n35625 & n35624 ) ;
  assign n35630 = n35094 &  n35294 ;
  assign n35631 = n35293 &  n35630 ;
  assign n35619 = x83 | n35094 ;
  assign n35620 = x83 &  n35094 ;
  assign n35621 = ( n35619 & ~n35620 ) | ( n35619 & 1'b0 ) | ( ~n35620 & 1'b0 ) ;
  assign n35633 = ( n35247 & n35295 ) | ( n35247 & n35621 ) | ( n35295 & n35621 ) ;
  assign n35632 = n35247 | n35621 ;
  assign n35634 = ( n35631 & ~n35633 ) | ( n35631 & n35632 ) | ( ~n35633 & n35632 ) ;
  assign n35638 = n35102 &  n35294 ;
  assign n35639 = n35293 &  n35638 ;
  assign n35627 = x82 | n35102 ;
  assign n35628 = x82 &  n35102 ;
  assign n35629 = ( n35627 & ~n35628 ) | ( n35627 & 1'b0 ) | ( ~n35628 & 1'b0 ) ;
  assign n35641 = ( n35246 & n35295 ) | ( n35246 & n35629 ) | ( n35295 & n35629 ) ;
  assign n35640 = n35246 | n35629 ;
  assign n35642 = ( n35639 & ~n35641 ) | ( n35639 & n35640 ) | ( ~n35641 & n35640 ) ;
  assign n35646 = n35110 &  n35294 ;
  assign n35647 = n35293 &  n35646 ;
  assign n35635 = x81 | n35110 ;
  assign n35636 = x81 &  n35110 ;
  assign n35637 = ( n35635 & ~n35636 ) | ( n35635 & 1'b0 ) | ( ~n35636 & 1'b0 ) ;
  assign n35649 = ( n35245 & n35295 ) | ( n35245 & n35637 ) | ( n35295 & n35637 ) ;
  assign n35648 = n35245 | n35637 ;
  assign n35650 = ( n35647 & ~n35649 ) | ( n35647 & n35648 ) | ( ~n35649 & n35648 ) ;
  assign n35654 = n35118 &  n35294 ;
  assign n35655 = n35293 &  n35654 ;
  assign n35643 = x80 | n35118 ;
  assign n35644 = x80 &  n35118 ;
  assign n35645 = ( n35643 & ~n35644 ) | ( n35643 & 1'b0 ) | ( ~n35644 & 1'b0 ) ;
  assign n35657 = ( n35244 & n35295 ) | ( n35244 & n35645 ) | ( n35295 & n35645 ) ;
  assign n35656 = n35244 | n35645 ;
  assign n35658 = ( n35655 & ~n35657 ) | ( n35655 & n35656 ) | ( ~n35657 & n35656 ) ;
  assign n35662 = n35126 &  n35294 ;
  assign n35663 = n35293 &  n35662 ;
  assign n35651 = x79 | n35126 ;
  assign n35652 = x79 &  n35126 ;
  assign n35653 = ( n35651 & ~n35652 ) | ( n35651 & 1'b0 ) | ( ~n35652 & 1'b0 ) ;
  assign n35665 = ( n35243 & n35295 ) | ( n35243 & n35653 ) | ( n35295 & n35653 ) ;
  assign n35664 = n35243 | n35653 ;
  assign n35666 = ( n35663 & ~n35665 ) | ( n35663 & n35664 ) | ( ~n35665 & n35664 ) ;
  assign n35670 = n35134 &  n35294 ;
  assign n35671 = n35293 &  n35670 ;
  assign n35659 = x78 | n35134 ;
  assign n35660 = x78 &  n35134 ;
  assign n35661 = ( n35659 & ~n35660 ) | ( n35659 & 1'b0 ) | ( ~n35660 & 1'b0 ) ;
  assign n35673 = ( n35242 & n35295 ) | ( n35242 & n35661 ) | ( n35295 & n35661 ) ;
  assign n35672 = n35242 | n35661 ;
  assign n35674 = ( n35671 & ~n35673 ) | ( n35671 & n35672 ) | ( ~n35673 & n35672 ) ;
  assign n35678 = n35142 &  n35294 ;
  assign n35679 = n35293 &  n35678 ;
  assign n35667 = x77 | n35142 ;
  assign n35668 = x77 &  n35142 ;
  assign n35669 = ( n35667 & ~n35668 ) | ( n35667 & 1'b0 ) | ( ~n35668 & 1'b0 ) ;
  assign n35681 = ( n35241 & n35295 ) | ( n35241 & n35669 ) | ( n35295 & n35669 ) ;
  assign n35680 = n35241 | n35669 ;
  assign n35682 = ( n35679 & ~n35681 ) | ( n35679 & n35680 ) | ( ~n35681 & n35680 ) ;
  assign n35686 = n35150 &  n35294 ;
  assign n35687 = n35293 &  n35686 ;
  assign n35675 = x76 | n35150 ;
  assign n35676 = x76 &  n35150 ;
  assign n35677 = ( n35675 & ~n35676 ) | ( n35675 & 1'b0 ) | ( ~n35676 & 1'b0 ) ;
  assign n35689 = ( n35240 & n35295 ) | ( n35240 & n35677 ) | ( n35295 & n35677 ) ;
  assign n35688 = n35240 | n35677 ;
  assign n35690 = ( n35687 & ~n35689 ) | ( n35687 & n35688 ) | ( ~n35689 & n35688 ) ;
  assign n35694 = n35158 &  n35294 ;
  assign n35695 = n35293 &  n35694 ;
  assign n35683 = x75 | n35158 ;
  assign n35684 = x75 &  n35158 ;
  assign n35685 = ( n35683 & ~n35684 ) | ( n35683 & 1'b0 ) | ( ~n35684 & 1'b0 ) ;
  assign n35697 = ( n35239 & n35295 ) | ( n35239 & n35685 ) | ( n35295 & n35685 ) ;
  assign n35696 = n35239 | n35685 ;
  assign n35698 = ( n35695 & ~n35697 ) | ( n35695 & n35696 ) | ( ~n35697 & n35696 ) ;
  assign n35702 = n35166 &  n35294 ;
  assign n35703 = n35293 &  n35702 ;
  assign n35691 = x74 | n35166 ;
  assign n35692 = x74 &  n35166 ;
  assign n35693 = ( n35691 & ~n35692 ) | ( n35691 & 1'b0 ) | ( ~n35692 & 1'b0 ) ;
  assign n35705 = ( n35238 & n35295 ) | ( n35238 & n35693 ) | ( n35295 & n35693 ) ;
  assign n35704 = n35238 | n35693 ;
  assign n35706 = ( n35703 & ~n35705 ) | ( n35703 & n35704 ) | ( ~n35705 & n35704 ) ;
  assign n35710 = n35174 &  n35294 ;
  assign n35711 = n35293 &  n35710 ;
  assign n35699 = x73 | n35174 ;
  assign n35700 = x73 &  n35174 ;
  assign n35701 = ( n35699 & ~n35700 ) | ( n35699 & 1'b0 ) | ( ~n35700 & 1'b0 ) ;
  assign n35713 = ( n35237 & n35295 ) | ( n35237 & n35701 ) | ( n35295 & n35701 ) ;
  assign n35712 = n35237 | n35701 ;
  assign n35714 = ( n35711 & ~n35713 ) | ( n35711 & n35712 ) | ( ~n35713 & n35712 ) ;
  assign n35718 = n35182 &  n35294 ;
  assign n35719 = n35293 &  n35718 ;
  assign n35707 = x72 | n35182 ;
  assign n35708 = x72 &  n35182 ;
  assign n35709 = ( n35707 & ~n35708 ) | ( n35707 & 1'b0 ) | ( ~n35708 & 1'b0 ) ;
  assign n35721 = ( n35236 & n35295 ) | ( n35236 & n35709 ) | ( n35295 & n35709 ) ;
  assign n35720 = n35236 | n35709 ;
  assign n35722 = ( n35719 & ~n35721 ) | ( n35719 & n35720 ) | ( ~n35721 & n35720 ) ;
  assign n35726 = n35190 &  n35294 ;
  assign n35727 = n35293 &  n35726 ;
  assign n35715 = x71 | n35190 ;
  assign n35716 = x71 &  n35190 ;
  assign n35717 = ( n35715 & ~n35716 ) | ( n35715 & 1'b0 ) | ( ~n35716 & 1'b0 ) ;
  assign n35729 = ( n35235 & n35295 ) | ( n35235 & n35717 ) | ( n35295 & n35717 ) ;
  assign n35728 = n35235 | n35717 ;
  assign n35730 = ( n35727 & ~n35729 ) | ( n35727 & n35728 ) | ( ~n35729 & n35728 ) ;
  assign n35734 = n35198 &  n35294 ;
  assign n35735 = n35293 &  n35734 ;
  assign n35723 = x70 | n35198 ;
  assign n35724 = x70 &  n35198 ;
  assign n35725 = ( n35723 & ~n35724 ) | ( n35723 & 1'b0 ) | ( ~n35724 & 1'b0 ) ;
  assign n35737 = ( n35234 & n35295 ) | ( n35234 & n35725 ) | ( n35295 & n35725 ) ;
  assign n35736 = n35234 | n35725 ;
  assign n35738 = ( n35735 & ~n35737 ) | ( n35735 & n35736 ) | ( ~n35737 & n35736 ) ;
  assign n35742 = n35206 &  n35294 ;
  assign n35743 = n35293 &  n35742 ;
  assign n35731 = x69 | n35206 ;
  assign n35732 = x69 &  n35206 ;
  assign n35733 = ( n35731 & ~n35732 ) | ( n35731 & 1'b0 ) | ( ~n35732 & 1'b0 ) ;
  assign n35745 = ( n35233 & n35295 ) | ( n35233 & n35733 ) | ( n35295 & n35733 ) ;
  assign n35744 = n35233 | n35733 ;
  assign n35746 = ( n35743 & ~n35745 ) | ( n35743 & n35744 ) | ( ~n35745 & n35744 ) ;
  assign n35750 = n35214 &  n35294 ;
  assign n35751 = n35293 &  n35750 ;
  assign n35739 = x68 | n35214 ;
  assign n35740 = x68 &  n35214 ;
  assign n35741 = ( n35739 & ~n35740 ) | ( n35739 & 1'b0 ) | ( ~n35740 & 1'b0 ) ;
  assign n35753 = ( n35232 & n35295 ) | ( n35232 & n35741 ) | ( n35295 & n35741 ) ;
  assign n35752 = n35232 | n35741 ;
  assign n35754 = ( n35751 & ~n35753 ) | ( n35751 & n35752 ) | ( ~n35753 & n35752 ) ;
  assign n35758 = n35219 &  n35294 ;
  assign n35759 = n35293 &  n35758 ;
  assign n35747 = x67 | n35219 ;
  assign n35748 = x67 &  n35219 ;
  assign n35749 = ( n35747 & ~n35748 ) | ( n35747 & 1'b0 ) | ( ~n35748 & 1'b0 ) ;
  assign n35761 = ( n35231 & n35295 ) | ( n35231 & n35749 ) | ( n35295 & n35749 ) ;
  assign n35760 = n35231 | n35749 ;
  assign n35762 = ( n35759 & ~n35761 ) | ( n35759 & n35760 ) | ( ~n35761 & n35760 ) ;
  assign n35763 = n35225 &  n35294 ;
  assign n35764 = n35293 &  n35763 ;
  assign n35755 = x66 | n35225 ;
  assign n35756 = x66 &  n35225 ;
  assign n35757 = ( n35755 & ~n35756 ) | ( n35755 & 1'b0 ) | ( ~n35756 & 1'b0 ) ;
  assign n35765 = n35230 &  n35757 ;
  assign n35766 = ( n35230 & ~n35295 ) | ( n35230 & n35757 ) | ( ~n35295 & n35757 ) ;
  assign n35767 = ( n35764 & ~n35765 ) | ( n35764 & n35766 ) | ( ~n35765 & n35766 ) ;
  assign n35768 = ( x65 & ~n16926 ) | ( x65 & n35229 ) | ( ~n16926 & n35229 ) ;
  assign n35769 = ( n35230 & ~x65 ) | ( n35230 & n35768 ) | ( ~x65 & n35768 ) ;
  assign n35770 = ~n35295 & n35769 ;
  assign n35771 = n35229 &  n35294 ;
  assign n35772 = n35293 &  n35771 ;
  assign n35773 = n35770 | n35772 ;
  assign n35774 = ( x64 & ~n35295 ) | ( x64 & 1'b0 ) | ( ~n35295 & 1'b0 ) ;
  assign n35775 = ( x3 & ~n35774 ) | ( x3 & 1'b0 ) | ( ~n35774 & 1'b0 ) ;
  assign n35776 = ( n16926 & ~n35295 ) | ( n16926 & 1'b0 ) | ( ~n35295 & 1'b0 ) ;
  assign n35777 = n35775 | n35776 ;
  assign n35778 = ( x65 & ~n35777 ) | ( x65 & n17483 ) | ( ~n35777 & n17483 ) ;
  assign n35779 = ( x66 & ~n35773 ) | ( x66 & n35778 ) | ( ~n35773 & n35778 ) ;
  assign n35780 = ( x67 & ~n35767 ) | ( x67 & n35779 ) | ( ~n35767 & n35779 ) ;
  assign n35781 = ( x68 & ~n35762 ) | ( x68 & n35780 ) | ( ~n35762 & n35780 ) ;
  assign n35782 = ( x69 & ~n35754 ) | ( x69 & n35781 ) | ( ~n35754 & n35781 ) ;
  assign n35783 = ( x70 & ~n35746 ) | ( x70 & n35782 ) | ( ~n35746 & n35782 ) ;
  assign n35784 = ( x71 & ~n35738 ) | ( x71 & n35783 ) | ( ~n35738 & n35783 ) ;
  assign n35785 = ( x72 & ~n35730 ) | ( x72 & n35784 ) | ( ~n35730 & n35784 ) ;
  assign n35786 = ( x73 & ~n35722 ) | ( x73 & n35785 ) | ( ~n35722 & n35785 ) ;
  assign n35787 = ( x74 & ~n35714 ) | ( x74 & n35786 ) | ( ~n35714 & n35786 ) ;
  assign n35788 = ( x75 & ~n35706 ) | ( x75 & n35787 ) | ( ~n35706 & n35787 ) ;
  assign n35789 = ( x76 & ~n35698 ) | ( x76 & n35788 ) | ( ~n35698 & n35788 ) ;
  assign n35790 = ( x77 & ~n35690 ) | ( x77 & n35789 ) | ( ~n35690 & n35789 ) ;
  assign n35791 = ( x78 & ~n35682 ) | ( x78 & n35790 ) | ( ~n35682 & n35790 ) ;
  assign n35792 = ( x79 & ~n35674 ) | ( x79 & n35791 ) | ( ~n35674 & n35791 ) ;
  assign n35793 = ( x80 & ~n35666 ) | ( x80 & n35792 ) | ( ~n35666 & n35792 ) ;
  assign n35794 = ( x81 & ~n35658 ) | ( x81 & n35793 ) | ( ~n35658 & n35793 ) ;
  assign n35795 = ( x82 & ~n35650 ) | ( x82 & n35794 ) | ( ~n35650 & n35794 ) ;
  assign n35796 = ( x83 & ~n35642 ) | ( x83 & n35795 ) | ( ~n35642 & n35795 ) ;
  assign n35797 = ( x84 & ~n35634 ) | ( x84 & n35796 ) | ( ~n35634 & n35796 ) ;
  assign n35798 = ( x85 & ~n35626 ) | ( x85 & n35797 ) | ( ~n35626 & n35797 ) ;
  assign n35799 = ( x86 & ~n35618 ) | ( x86 & n35798 ) | ( ~n35618 & n35798 ) ;
  assign n35800 = ( x87 & ~n35610 ) | ( x87 & n35799 ) | ( ~n35610 & n35799 ) ;
  assign n35801 = ( x88 & ~n35602 ) | ( x88 & n35800 ) | ( ~n35602 & n35800 ) ;
  assign n35802 = ( x89 & ~n35594 ) | ( x89 & n35801 ) | ( ~n35594 & n35801 ) ;
  assign n35803 = ( x90 & ~n35586 ) | ( x90 & n35802 ) | ( ~n35586 & n35802 ) ;
  assign n35804 = ( x91 & ~n35578 ) | ( x91 & n35803 ) | ( ~n35578 & n35803 ) ;
  assign n35805 = ( x92 & ~n35570 ) | ( x92 & n35804 ) | ( ~n35570 & n35804 ) ;
  assign n35806 = ( x93 & ~n35562 ) | ( x93 & n35805 ) | ( ~n35562 & n35805 ) ;
  assign n35807 = ( x94 & ~n35554 ) | ( x94 & n35806 ) | ( ~n35554 & n35806 ) ;
  assign n35808 = ( x95 & ~n35546 ) | ( x95 & n35807 ) | ( ~n35546 & n35807 ) ;
  assign n35809 = ( x96 & ~n35538 ) | ( x96 & n35808 ) | ( ~n35538 & n35808 ) ;
  assign n35810 = ( x97 & ~n35530 ) | ( x97 & n35809 ) | ( ~n35530 & n35809 ) ;
  assign n35811 = ( x98 & ~n35522 ) | ( x98 & n35810 ) | ( ~n35522 & n35810 ) ;
  assign n35812 = ( x99 & ~n35514 ) | ( x99 & n35811 ) | ( ~n35514 & n35811 ) ;
  assign n35813 = ( x100 & ~n35506 ) | ( x100 & n35812 ) | ( ~n35506 & n35812 ) ;
  assign n35814 = ( x101 & ~n35498 ) | ( x101 & n35813 ) | ( ~n35498 & n35813 ) ;
  assign n35815 = ( x102 & ~n35490 ) | ( x102 & n35814 ) | ( ~n35490 & n35814 ) ;
  assign n35816 = ( x103 & ~n35482 ) | ( x103 & n35815 ) | ( ~n35482 & n35815 ) ;
  assign n35817 = ( x104 & ~n35474 ) | ( x104 & n35816 ) | ( ~n35474 & n35816 ) ;
  assign n35818 = ( x105 & ~n35466 ) | ( x105 & n35817 ) | ( ~n35466 & n35817 ) ;
  assign n35819 = ( x106 & ~n35458 ) | ( x106 & n35818 ) | ( ~n35458 & n35818 ) ;
  assign n35820 = ( x107 & ~n35450 ) | ( x107 & n35819 ) | ( ~n35450 & n35819 ) ;
  assign n35821 = ( x108 & ~n35442 ) | ( x108 & n35820 ) | ( ~n35442 & n35820 ) ;
  assign n35822 = ( x109 & ~n35434 ) | ( x109 & n35821 ) | ( ~n35434 & n35821 ) ;
  assign n35823 = ( x110 & ~n35426 ) | ( x110 & n35822 ) | ( ~n35426 & n35822 ) ;
  assign n35824 = ( x111 & ~n35418 ) | ( x111 & n35823 ) | ( ~n35418 & n35823 ) ;
  assign n35825 = ( x112 & ~n35410 ) | ( x112 & n35824 ) | ( ~n35410 & n35824 ) ;
  assign n35826 = ( x113 & ~n35402 ) | ( x113 & n35825 ) | ( ~n35402 & n35825 ) ;
  assign n35827 = ( x114 & ~n35394 ) | ( x114 & n35826 ) | ( ~n35394 & n35826 ) ;
  assign n35828 = ( x115 & ~n35386 ) | ( x115 & n35827 ) | ( ~n35386 & n35827 ) ;
  assign n35829 = ( x116 & ~n35378 ) | ( x116 & n35828 ) | ( ~n35378 & n35828 ) ;
  assign n35830 = ( x117 & ~n35370 ) | ( x117 & n35829 ) | ( ~n35370 & n35829 ) ;
  assign n35831 = ( x118 & ~n35362 ) | ( x118 & n35830 ) | ( ~n35362 & n35830 ) ;
  assign n35832 = ( x119 & ~n35354 ) | ( x119 & n35831 ) | ( ~n35354 & n35831 ) ;
  assign n35833 = ( x120 & ~n35346 ) | ( x120 & n35832 ) | ( ~n35346 & n35832 ) ;
  assign n35834 = ( x121 & ~n35338 ) | ( x121 & n35833 ) | ( ~n35338 & n35833 ) ;
  assign n35835 = ( x122 & ~n35330 ) | ( x122 & n35834 ) | ( ~n35330 & n35834 ) ;
  assign n35836 = ( x123 & ~n35322 ) | ( x123 & n35835 ) | ( ~n35322 & n35835 ) ;
  assign n35837 = ( x124 & ~n35314 ) | ( x124 & n35836 ) | ( ~n35314 & n35836 ) ;
  assign n35299 = n34766 | n35290 ;
  assign n35300 = ( n35288 & ~n35299 ) | ( n35288 & 1'b0 ) | ( ~n35299 & 1'b0 ) ;
  assign n35301 = ~n35288 & n35299 ;
  assign n35302 = ( n35300 & ~n35295 ) | ( n35300 & n35301 ) | ( ~n35295 & n35301 ) ;
  assign n35303 = n152 &  n34765 ;
  assign n35304 = n35293 &  n35303 ;
  assign n35305 = n35302 | n35304 ;
  assign n35306 = ~x125 & n35305 ;
  assign n35838 = ( x125 & ~n35304 ) | ( x125 & 1'b0 ) | ( ~n35304 & 1'b0 ) ;
  assign n35839 = ~n35302 & n35838 ;
  assign n35848 = n35306 | n35839 ;
  assign n35849 = ( n35837 & ~n35848 ) | ( n35837 & 1'b0 ) | ( ~n35848 & 1'b0 ) ;
  assign n35840 = ( n35837 & ~n35306 ) | ( n35837 & n35839 ) | ( ~n35306 & n35839 ) ;
  assign n35841 = ( n35306 & ~n151 ) | ( n35306 & n35840 ) | ( ~n151 & n35840 ) ;
  assign n35842 = n151 | n35841 ;
  assign n35843 = ~n35305 |  n235 ;
  assign n35844 = n35842 &  n35843 ;
  assign n35850 = ~n35837 & n35848 ;
  assign n35851 = ( n35849 & ~n35844 ) | ( n35849 & n35850 ) | ( ~n35844 & n35850 ) ;
  assign n35852 = n235 &  n35305 ;
  assign n35853 = n35842 &  n35852 ;
  assign n35854 = n35851 | n35853 ;
  assign n35855 = ~x126 & n35854 ;
  assign n35859 = n35314 &  n35843 ;
  assign n35860 = n35842 &  n35859 ;
  assign n35845 = x124 | n35314 ;
  assign n35846 = x124 &  n35314 ;
  assign n35847 = ( n35845 & ~n35846 ) | ( n35845 & 1'b0 ) | ( ~n35846 & 1'b0 ) ;
  assign n35862 = ( n35836 & n35844 ) | ( n35836 & n35847 ) | ( n35844 & n35847 ) ;
  assign n35861 = n35836 | n35847 ;
  assign n35863 = ( n35860 & ~n35862 ) | ( n35860 & n35861 ) | ( ~n35862 & n35861 ) ;
  assign n35867 = n35322 &  n35843 ;
  assign n35868 = n35842 &  n35867 ;
  assign n35856 = x123 | n35322 ;
  assign n35857 = x123 &  n35322 ;
  assign n35858 = ( n35856 & ~n35857 ) | ( n35856 & 1'b0 ) | ( ~n35857 & 1'b0 ) ;
  assign n35870 = ( n35835 & n35844 ) | ( n35835 & n35858 ) | ( n35844 & n35858 ) ;
  assign n35869 = n35835 | n35858 ;
  assign n35871 = ( n35868 & ~n35870 ) | ( n35868 & n35869 ) | ( ~n35870 & n35869 ) ;
  assign n35875 = n35330 &  n35843 ;
  assign n35876 = n35842 &  n35875 ;
  assign n35864 = x122 | n35330 ;
  assign n35865 = x122 &  n35330 ;
  assign n35866 = ( n35864 & ~n35865 ) | ( n35864 & 1'b0 ) | ( ~n35865 & 1'b0 ) ;
  assign n35878 = ( n35834 & n35844 ) | ( n35834 & n35866 ) | ( n35844 & n35866 ) ;
  assign n35877 = n35834 | n35866 ;
  assign n35879 = ( n35876 & ~n35878 ) | ( n35876 & n35877 ) | ( ~n35878 & n35877 ) ;
  assign n35883 = n35338 &  n35843 ;
  assign n35884 = n35842 &  n35883 ;
  assign n35872 = x121 | n35338 ;
  assign n35873 = x121 &  n35338 ;
  assign n35874 = ( n35872 & ~n35873 ) | ( n35872 & 1'b0 ) | ( ~n35873 & 1'b0 ) ;
  assign n35886 = ( n35833 & n35844 ) | ( n35833 & n35874 ) | ( n35844 & n35874 ) ;
  assign n35885 = n35833 | n35874 ;
  assign n35887 = ( n35884 & ~n35886 ) | ( n35884 & n35885 ) | ( ~n35886 & n35885 ) ;
  assign n35891 = n35346 &  n35843 ;
  assign n35892 = n35842 &  n35891 ;
  assign n35880 = x120 | n35346 ;
  assign n35881 = x120 &  n35346 ;
  assign n35882 = ( n35880 & ~n35881 ) | ( n35880 & 1'b0 ) | ( ~n35881 & 1'b0 ) ;
  assign n35894 = ( n35832 & n35844 ) | ( n35832 & n35882 ) | ( n35844 & n35882 ) ;
  assign n35893 = n35832 | n35882 ;
  assign n35895 = ( n35892 & ~n35894 ) | ( n35892 & n35893 ) | ( ~n35894 & n35893 ) ;
  assign n35899 = n35354 &  n35843 ;
  assign n35900 = n35842 &  n35899 ;
  assign n35888 = x119 | n35354 ;
  assign n35889 = x119 &  n35354 ;
  assign n35890 = ( n35888 & ~n35889 ) | ( n35888 & 1'b0 ) | ( ~n35889 & 1'b0 ) ;
  assign n35902 = ( n35831 & n35844 ) | ( n35831 & n35890 ) | ( n35844 & n35890 ) ;
  assign n35901 = n35831 | n35890 ;
  assign n35903 = ( n35900 & ~n35902 ) | ( n35900 & n35901 ) | ( ~n35902 & n35901 ) ;
  assign n35907 = n35362 &  n35843 ;
  assign n35908 = n35842 &  n35907 ;
  assign n35896 = x118 | n35362 ;
  assign n35897 = x118 &  n35362 ;
  assign n35898 = ( n35896 & ~n35897 ) | ( n35896 & 1'b0 ) | ( ~n35897 & 1'b0 ) ;
  assign n35910 = ( n35830 & n35844 ) | ( n35830 & n35898 ) | ( n35844 & n35898 ) ;
  assign n35909 = n35830 | n35898 ;
  assign n35911 = ( n35908 & ~n35910 ) | ( n35908 & n35909 ) | ( ~n35910 & n35909 ) ;
  assign n35915 = n35370 &  n35843 ;
  assign n35916 = n35842 &  n35915 ;
  assign n35904 = x117 | n35370 ;
  assign n35905 = x117 &  n35370 ;
  assign n35906 = ( n35904 & ~n35905 ) | ( n35904 & 1'b0 ) | ( ~n35905 & 1'b0 ) ;
  assign n35918 = ( n35829 & n35844 ) | ( n35829 & n35906 ) | ( n35844 & n35906 ) ;
  assign n35917 = n35829 | n35906 ;
  assign n35919 = ( n35916 & ~n35918 ) | ( n35916 & n35917 ) | ( ~n35918 & n35917 ) ;
  assign n35923 = n35378 &  n35843 ;
  assign n35924 = n35842 &  n35923 ;
  assign n35912 = x116 | n35378 ;
  assign n35913 = x116 &  n35378 ;
  assign n35914 = ( n35912 & ~n35913 ) | ( n35912 & 1'b0 ) | ( ~n35913 & 1'b0 ) ;
  assign n35926 = ( n35828 & n35844 ) | ( n35828 & n35914 ) | ( n35844 & n35914 ) ;
  assign n35925 = n35828 | n35914 ;
  assign n35927 = ( n35924 & ~n35926 ) | ( n35924 & n35925 ) | ( ~n35926 & n35925 ) ;
  assign n35931 = n35386 &  n35843 ;
  assign n35932 = n35842 &  n35931 ;
  assign n35920 = x115 | n35386 ;
  assign n35921 = x115 &  n35386 ;
  assign n35922 = ( n35920 & ~n35921 ) | ( n35920 & 1'b0 ) | ( ~n35921 & 1'b0 ) ;
  assign n35934 = ( n35827 & n35844 ) | ( n35827 & n35922 ) | ( n35844 & n35922 ) ;
  assign n35933 = n35827 | n35922 ;
  assign n35935 = ( n35932 & ~n35934 ) | ( n35932 & n35933 ) | ( ~n35934 & n35933 ) ;
  assign n35939 = n35394 &  n35843 ;
  assign n35940 = n35842 &  n35939 ;
  assign n35928 = x114 | n35394 ;
  assign n35929 = x114 &  n35394 ;
  assign n35930 = ( n35928 & ~n35929 ) | ( n35928 & 1'b0 ) | ( ~n35929 & 1'b0 ) ;
  assign n35942 = ( n35826 & n35844 ) | ( n35826 & n35930 ) | ( n35844 & n35930 ) ;
  assign n35941 = n35826 | n35930 ;
  assign n35943 = ( n35940 & ~n35942 ) | ( n35940 & n35941 ) | ( ~n35942 & n35941 ) ;
  assign n35947 = n35402 &  n35843 ;
  assign n35948 = n35842 &  n35947 ;
  assign n35936 = x113 | n35402 ;
  assign n35937 = x113 &  n35402 ;
  assign n35938 = ( n35936 & ~n35937 ) | ( n35936 & 1'b0 ) | ( ~n35937 & 1'b0 ) ;
  assign n35950 = ( n35825 & n35844 ) | ( n35825 & n35938 ) | ( n35844 & n35938 ) ;
  assign n35949 = n35825 | n35938 ;
  assign n35951 = ( n35948 & ~n35950 ) | ( n35948 & n35949 ) | ( ~n35950 & n35949 ) ;
  assign n35955 = n35410 &  n35843 ;
  assign n35956 = n35842 &  n35955 ;
  assign n35944 = x112 | n35410 ;
  assign n35945 = x112 &  n35410 ;
  assign n35946 = ( n35944 & ~n35945 ) | ( n35944 & 1'b0 ) | ( ~n35945 & 1'b0 ) ;
  assign n35958 = ( n35824 & n35844 ) | ( n35824 & n35946 ) | ( n35844 & n35946 ) ;
  assign n35957 = n35824 | n35946 ;
  assign n35959 = ( n35956 & ~n35958 ) | ( n35956 & n35957 ) | ( ~n35958 & n35957 ) ;
  assign n35963 = n35418 &  n35843 ;
  assign n35964 = n35842 &  n35963 ;
  assign n35952 = x111 | n35418 ;
  assign n35953 = x111 &  n35418 ;
  assign n35954 = ( n35952 & ~n35953 ) | ( n35952 & 1'b0 ) | ( ~n35953 & 1'b0 ) ;
  assign n35966 = ( n35823 & n35844 ) | ( n35823 & n35954 ) | ( n35844 & n35954 ) ;
  assign n35965 = n35823 | n35954 ;
  assign n35967 = ( n35964 & ~n35966 ) | ( n35964 & n35965 ) | ( ~n35966 & n35965 ) ;
  assign n35971 = n35426 &  n35843 ;
  assign n35972 = n35842 &  n35971 ;
  assign n35960 = x110 | n35426 ;
  assign n35961 = x110 &  n35426 ;
  assign n35962 = ( n35960 & ~n35961 ) | ( n35960 & 1'b0 ) | ( ~n35961 & 1'b0 ) ;
  assign n35974 = ( n35822 & n35844 ) | ( n35822 & n35962 ) | ( n35844 & n35962 ) ;
  assign n35973 = n35822 | n35962 ;
  assign n35975 = ( n35972 & ~n35974 ) | ( n35972 & n35973 ) | ( ~n35974 & n35973 ) ;
  assign n35979 = n35434 &  n35843 ;
  assign n35980 = n35842 &  n35979 ;
  assign n35968 = x109 | n35434 ;
  assign n35969 = x109 &  n35434 ;
  assign n35970 = ( n35968 & ~n35969 ) | ( n35968 & 1'b0 ) | ( ~n35969 & 1'b0 ) ;
  assign n35982 = ( n35821 & n35844 ) | ( n35821 & n35970 ) | ( n35844 & n35970 ) ;
  assign n35981 = n35821 | n35970 ;
  assign n35983 = ( n35980 & ~n35982 ) | ( n35980 & n35981 ) | ( ~n35982 & n35981 ) ;
  assign n35987 = n35442 &  n35843 ;
  assign n35988 = n35842 &  n35987 ;
  assign n35976 = x108 | n35442 ;
  assign n35977 = x108 &  n35442 ;
  assign n35978 = ( n35976 & ~n35977 ) | ( n35976 & 1'b0 ) | ( ~n35977 & 1'b0 ) ;
  assign n35990 = ( n35820 & n35844 ) | ( n35820 & n35978 ) | ( n35844 & n35978 ) ;
  assign n35989 = n35820 | n35978 ;
  assign n35991 = ( n35988 & ~n35990 ) | ( n35988 & n35989 ) | ( ~n35990 & n35989 ) ;
  assign n35995 = n35450 &  n35843 ;
  assign n35996 = n35842 &  n35995 ;
  assign n35984 = x107 | n35450 ;
  assign n35985 = x107 &  n35450 ;
  assign n35986 = ( n35984 & ~n35985 ) | ( n35984 & 1'b0 ) | ( ~n35985 & 1'b0 ) ;
  assign n35998 = ( n35819 & n35844 ) | ( n35819 & n35986 ) | ( n35844 & n35986 ) ;
  assign n35997 = n35819 | n35986 ;
  assign n35999 = ( n35996 & ~n35998 ) | ( n35996 & n35997 ) | ( ~n35998 & n35997 ) ;
  assign n36003 = n35458 &  n35843 ;
  assign n36004 = n35842 &  n36003 ;
  assign n35992 = x106 | n35458 ;
  assign n35993 = x106 &  n35458 ;
  assign n35994 = ( n35992 & ~n35993 ) | ( n35992 & 1'b0 ) | ( ~n35993 & 1'b0 ) ;
  assign n36006 = ( n35818 & n35844 ) | ( n35818 & n35994 ) | ( n35844 & n35994 ) ;
  assign n36005 = n35818 | n35994 ;
  assign n36007 = ( n36004 & ~n36006 ) | ( n36004 & n36005 ) | ( ~n36006 & n36005 ) ;
  assign n36011 = n35466 &  n35843 ;
  assign n36012 = n35842 &  n36011 ;
  assign n36000 = x105 | n35466 ;
  assign n36001 = x105 &  n35466 ;
  assign n36002 = ( n36000 & ~n36001 ) | ( n36000 & 1'b0 ) | ( ~n36001 & 1'b0 ) ;
  assign n36014 = ( n35817 & n35844 ) | ( n35817 & n36002 ) | ( n35844 & n36002 ) ;
  assign n36013 = n35817 | n36002 ;
  assign n36015 = ( n36012 & ~n36014 ) | ( n36012 & n36013 ) | ( ~n36014 & n36013 ) ;
  assign n36019 = n35474 &  n35843 ;
  assign n36020 = n35842 &  n36019 ;
  assign n36008 = x104 | n35474 ;
  assign n36009 = x104 &  n35474 ;
  assign n36010 = ( n36008 & ~n36009 ) | ( n36008 & 1'b0 ) | ( ~n36009 & 1'b0 ) ;
  assign n36022 = ( n35816 & n35844 ) | ( n35816 & n36010 ) | ( n35844 & n36010 ) ;
  assign n36021 = n35816 | n36010 ;
  assign n36023 = ( n36020 & ~n36022 ) | ( n36020 & n36021 ) | ( ~n36022 & n36021 ) ;
  assign n36027 = n35482 &  n35843 ;
  assign n36028 = n35842 &  n36027 ;
  assign n36016 = x103 | n35482 ;
  assign n36017 = x103 &  n35482 ;
  assign n36018 = ( n36016 & ~n36017 ) | ( n36016 & 1'b0 ) | ( ~n36017 & 1'b0 ) ;
  assign n36030 = ( n35815 & n35844 ) | ( n35815 & n36018 ) | ( n35844 & n36018 ) ;
  assign n36029 = n35815 | n36018 ;
  assign n36031 = ( n36028 & ~n36030 ) | ( n36028 & n36029 ) | ( ~n36030 & n36029 ) ;
  assign n36035 = n35490 &  n35843 ;
  assign n36036 = n35842 &  n36035 ;
  assign n36024 = x102 | n35490 ;
  assign n36025 = x102 &  n35490 ;
  assign n36026 = ( n36024 & ~n36025 ) | ( n36024 & 1'b0 ) | ( ~n36025 & 1'b0 ) ;
  assign n36038 = ( n35814 & n35844 ) | ( n35814 & n36026 ) | ( n35844 & n36026 ) ;
  assign n36037 = n35814 | n36026 ;
  assign n36039 = ( n36036 & ~n36038 ) | ( n36036 & n36037 ) | ( ~n36038 & n36037 ) ;
  assign n36043 = n35498 &  n35843 ;
  assign n36044 = n35842 &  n36043 ;
  assign n36032 = x101 | n35498 ;
  assign n36033 = x101 &  n35498 ;
  assign n36034 = ( n36032 & ~n36033 ) | ( n36032 & 1'b0 ) | ( ~n36033 & 1'b0 ) ;
  assign n36046 = ( n35813 & n35844 ) | ( n35813 & n36034 ) | ( n35844 & n36034 ) ;
  assign n36045 = n35813 | n36034 ;
  assign n36047 = ( n36044 & ~n36046 ) | ( n36044 & n36045 ) | ( ~n36046 & n36045 ) ;
  assign n36051 = n35506 &  n35843 ;
  assign n36052 = n35842 &  n36051 ;
  assign n36040 = x100 | n35506 ;
  assign n36041 = x100 &  n35506 ;
  assign n36042 = ( n36040 & ~n36041 ) | ( n36040 & 1'b0 ) | ( ~n36041 & 1'b0 ) ;
  assign n36054 = ( n35812 & n35844 ) | ( n35812 & n36042 ) | ( n35844 & n36042 ) ;
  assign n36053 = n35812 | n36042 ;
  assign n36055 = ( n36052 & ~n36054 ) | ( n36052 & n36053 ) | ( ~n36054 & n36053 ) ;
  assign n36059 = n35514 &  n35843 ;
  assign n36060 = n35842 &  n36059 ;
  assign n36048 = x99 | n35514 ;
  assign n36049 = x99 &  n35514 ;
  assign n36050 = ( n36048 & ~n36049 ) | ( n36048 & 1'b0 ) | ( ~n36049 & 1'b0 ) ;
  assign n36062 = ( n35811 & n35844 ) | ( n35811 & n36050 ) | ( n35844 & n36050 ) ;
  assign n36061 = n35811 | n36050 ;
  assign n36063 = ( n36060 & ~n36062 ) | ( n36060 & n36061 ) | ( ~n36062 & n36061 ) ;
  assign n36067 = n35522 &  n35843 ;
  assign n36068 = n35842 &  n36067 ;
  assign n36056 = x98 | n35522 ;
  assign n36057 = x98 &  n35522 ;
  assign n36058 = ( n36056 & ~n36057 ) | ( n36056 & 1'b0 ) | ( ~n36057 & 1'b0 ) ;
  assign n36070 = ( n35810 & n35844 ) | ( n35810 & n36058 ) | ( n35844 & n36058 ) ;
  assign n36069 = n35810 | n36058 ;
  assign n36071 = ( n36068 & ~n36070 ) | ( n36068 & n36069 ) | ( ~n36070 & n36069 ) ;
  assign n36075 = n35530 &  n35843 ;
  assign n36076 = n35842 &  n36075 ;
  assign n36064 = x97 | n35530 ;
  assign n36065 = x97 &  n35530 ;
  assign n36066 = ( n36064 & ~n36065 ) | ( n36064 & 1'b0 ) | ( ~n36065 & 1'b0 ) ;
  assign n36078 = ( n35809 & n35844 ) | ( n35809 & n36066 ) | ( n35844 & n36066 ) ;
  assign n36077 = n35809 | n36066 ;
  assign n36079 = ( n36076 & ~n36078 ) | ( n36076 & n36077 ) | ( ~n36078 & n36077 ) ;
  assign n36083 = n35538 &  n35843 ;
  assign n36084 = n35842 &  n36083 ;
  assign n36072 = x96 | n35538 ;
  assign n36073 = x96 &  n35538 ;
  assign n36074 = ( n36072 & ~n36073 ) | ( n36072 & 1'b0 ) | ( ~n36073 & 1'b0 ) ;
  assign n36086 = ( n35808 & n35844 ) | ( n35808 & n36074 ) | ( n35844 & n36074 ) ;
  assign n36085 = n35808 | n36074 ;
  assign n36087 = ( n36084 & ~n36086 ) | ( n36084 & n36085 ) | ( ~n36086 & n36085 ) ;
  assign n36091 = n35546 &  n35843 ;
  assign n36092 = n35842 &  n36091 ;
  assign n36080 = x95 | n35546 ;
  assign n36081 = x95 &  n35546 ;
  assign n36082 = ( n36080 & ~n36081 ) | ( n36080 & 1'b0 ) | ( ~n36081 & 1'b0 ) ;
  assign n36094 = ( n35807 & n35844 ) | ( n35807 & n36082 ) | ( n35844 & n36082 ) ;
  assign n36093 = n35807 | n36082 ;
  assign n36095 = ( n36092 & ~n36094 ) | ( n36092 & n36093 ) | ( ~n36094 & n36093 ) ;
  assign n36099 = n35554 &  n35843 ;
  assign n36100 = n35842 &  n36099 ;
  assign n36088 = x94 | n35554 ;
  assign n36089 = x94 &  n35554 ;
  assign n36090 = ( n36088 & ~n36089 ) | ( n36088 & 1'b0 ) | ( ~n36089 & 1'b0 ) ;
  assign n36102 = ( n35806 & n35844 ) | ( n35806 & n36090 ) | ( n35844 & n36090 ) ;
  assign n36101 = n35806 | n36090 ;
  assign n36103 = ( n36100 & ~n36102 ) | ( n36100 & n36101 ) | ( ~n36102 & n36101 ) ;
  assign n36107 = n35562 &  n35843 ;
  assign n36108 = n35842 &  n36107 ;
  assign n36096 = x93 | n35562 ;
  assign n36097 = x93 &  n35562 ;
  assign n36098 = ( n36096 & ~n36097 ) | ( n36096 & 1'b0 ) | ( ~n36097 & 1'b0 ) ;
  assign n36110 = ( n35805 & n35844 ) | ( n35805 & n36098 ) | ( n35844 & n36098 ) ;
  assign n36109 = n35805 | n36098 ;
  assign n36111 = ( n36108 & ~n36110 ) | ( n36108 & n36109 ) | ( ~n36110 & n36109 ) ;
  assign n36115 = n35570 &  n35843 ;
  assign n36116 = n35842 &  n36115 ;
  assign n36104 = x92 | n35570 ;
  assign n36105 = x92 &  n35570 ;
  assign n36106 = ( n36104 & ~n36105 ) | ( n36104 & 1'b0 ) | ( ~n36105 & 1'b0 ) ;
  assign n36118 = ( n35804 & n35844 ) | ( n35804 & n36106 ) | ( n35844 & n36106 ) ;
  assign n36117 = n35804 | n36106 ;
  assign n36119 = ( n36116 & ~n36118 ) | ( n36116 & n36117 ) | ( ~n36118 & n36117 ) ;
  assign n36123 = n35578 &  n35843 ;
  assign n36124 = n35842 &  n36123 ;
  assign n36112 = x91 | n35578 ;
  assign n36113 = x91 &  n35578 ;
  assign n36114 = ( n36112 & ~n36113 ) | ( n36112 & 1'b0 ) | ( ~n36113 & 1'b0 ) ;
  assign n36126 = ( n35803 & n35844 ) | ( n35803 & n36114 ) | ( n35844 & n36114 ) ;
  assign n36125 = n35803 | n36114 ;
  assign n36127 = ( n36124 & ~n36126 ) | ( n36124 & n36125 ) | ( ~n36126 & n36125 ) ;
  assign n36131 = n35586 &  n35843 ;
  assign n36132 = n35842 &  n36131 ;
  assign n36120 = x90 | n35586 ;
  assign n36121 = x90 &  n35586 ;
  assign n36122 = ( n36120 & ~n36121 ) | ( n36120 & 1'b0 ) | ( ~n36121 & 1'b0 ) ;
  assign n36134 = ( n35802 & n35844 ) | ( n35802 & n36122 ) | ( n35844 & n36122 ) ;
  assign n36133 = n35802 | n36122 ;
  assign n36135 = ( n36132 & ~n36134 ) | ( n36132 & n36133 ) | ( ~n36134 & n36133 ) ;
  assign n36139 = n35594 &  n35843 ;
  assign n36140 = n35842 &  n36139 ;
  assign n36128 = x89 | n35594 ;
  assign n36129 = x89 &  n35594 ;
  assign n36130 = ( n36128 & ~n36129 ) | ( n36128 & 1'b0 ) | ( ~n36129 & 1'b0 ) ;
  assign n36142 = ( n35801 & n35844 ) | ( n35801 & n36130 ) | ( n35844 & n36130 ) ;
  assign n36141 = n35801 | n36130 ;
  assign n36143 = ( n36140 & ~n36142 ) | ( n36140 & n36141 ) | ( ~n36142 & n36141 ) ;
  assign n36147 = n35602 &  n35843 ;
  assign n36148 = n35842 &  n36147 ;
  assign n36136 = x88 | n35602 ;
  assign n36137 = x88 &  n35602 ;
  assign n36138 = ( n36136 & ~n36137 ) | ( n36136 & 1'b0 ) | ( ~n36137 & 1'b0 ) ;
  assign n36150 = ( n35800 & n35844 ) | ( n35800 & n36138 ) | ( n35844 & n36138 ) ;
  assign n36149 = n35800 | n36138 ;
  assign n36151 = ( n36148 & ~n36150 ) | ( n36148 & n36149 ) | ( ~n36150 & n36149 ) ;
  assign n36155 = n35610 &  n35843 ;
  assign n36156 = n35842 &  n36155 ;
  assign n36144 = x87 | n35610 ;
  assign n36145 = x87 &  n35610 ;
  assign n36146 = ( n36144 & ~n36145 ) | ( n36144 & 1'b0 ) | ( ~n36145 & 1'b0 ) ;
  assign n36158 = ( n35799 & n35844 ) | ( n35799 & n36146 ) | ( n35844 & n36146 ) ;
  assign n36157 = n35799 | n36146 ;
  assign n36159 = ( n36156 & ~n36158 ) | ( n36156 & n36157 ) | ( ~n36158 & n36157 ) ;
  assign n36163 = n35618 &  n35843 ;
  assign n36164 = n35842 &  n36163 ;
  assign n36152 = x86 | n35618 ;
  assign n36153 = x86 &  n35618 ;
  assign n36154 = ( n36152 & ~n36153 ) | ( n36152 & 1'b0 ) | ( ~n36153 & 1'b0 ) ;
  assign n36166 = ( n35798 & n35844 ) | ( n35798 & n36154 ) | ( n35844 & n36154 ) ;
  assign n36165 = n35798 | n36154 ;
  assign n36167 = ( n36164 & ~n36166 ) | ( n36164 & n36165 ) | ( ~n36166 & n36165 ) ;
  assign n36171 = n35626 &  n35843 ;
  assign n36172 = n35842 &  n36171 ;
  assign n36160 = x85 | n35626 ;
  assign n36161 = x85 &  n35626 ;
  assign n36162 = ( n36160 & ~n36161 ) | ( n36160 & 1'b0 ) | ( ~n36161 & 1'b0 ) ;
  assign n36174 = ( n35797 & n35844 ) | ( n35797 & n36162 ) | ( n35844 & n36162 ) ;
  assign n36173 = n35797 | n36162 ;
  assign n36175 = ( n36172 & ~n36174 ) | ( n36172 & n36173 ) | ( ~n36174 & n36173 ) ;
  assign n36179 = n35634 &  n35843 ;
  assign n36180 = n35842 &  n36179 ;
  assign n36168 = x84 | n35634 ;
  assign n36169 = x84 &  n35634 ;
  assign n36170 = ( n36168 & ~n36169 ) | ( n36168 & 1'b0 ) | ( ~n36169 & 1'b0 ) ;
  assign n36182 = ( n35796 & n35844 ) | ( n35796 & n36170 ) | ( n35844 & n36170 ) ;
  assign n36181 = n35796 | n36170 ;
  assign n36183 = ( n36180 & ~n36182 ) | ( n36180 & n36181 ) | ( ~n36182 & n36181 ) ;
  assign n36187 = n35642 &  n35843 ;
  assign n36188 = n35842 &  n36187 ;
  assign n36176 = x83 | n35642 ;
  assign n36177 = x83 &  n35642 ;
  assign n36178 = ( n36176 & ~n36177 ) | ( n36176 & 1'b0 ) | ( ~n36177 & 1'b0 ) ;
  assign n36190 = ( n35795 & n35844 ) | ( n35795 & n36178 ) | ( n35844 & n36178 ) ;
  assign n36189 = n35795 | n36178 ;
  assign n36191 = ( n36188 & ~n36190 ) | ( n36188 & n36189 ) | ( ~n36190 & n36189 ) ;
  assign n36195 = n35650 &  n35843 ;
  assign n36196 = n35842 &  n36195 ;
  assign n36184 = x82 | n35650 ;
  assign n36185 = x82 &  n35650 ;
  assign n36186 = ( n36184 & ~n36185 ) | ( n36184 & 1'b0 ) | ( ~n36185 & 1'b0 ) ;
  assign n36198 = ( n35794 & n35844 ) | ( n35794 & n36186 ) | ( n35844 & n36186 ) ;
  assign n36197 = n35794 | n36186 ;
  assign n36199 = ( n36196 & ~n36198 ) | ( n36196 & n36197 ) | ( ~n36198 & n36197 ) ;
  assign n36203 = n35658 &  n35843 ;
  assign n36204 = n35842 &  n36203 ;
  assign n36192 = x81 | n35658 ;
  assign n36193 = x81 &  n35658 ;
  assign n36194 = ( n36192 & ~n36193 ) | ( n36192 & 1'b0 ) | ( ~n36193 & 1'b0 ) ;
  assign n36206 = ( n35793 & n35844 ) | ( n35793 & n36194 ) | ( n35844 & n36194 ) ;
  assign n36205 = n35793 | n36194 ;
  assign n36207 = ( n36204 & ~n36206 ) | ( n36204 & n36205 ) | ( ~n36206 & n36205 ) ;
  assign n36211 = n35666 &  n35843 ;
  assign n36212 = n35842 &  n36211 ;
  assign n36200 = x80 | n35666 ;
  assign n36201 = x80 &  n35666 ;
  assign n36202 = ( n36200 & ~n36201 ) | ( n36200 & 1'b0 ) | ( ~n36201 & 1'b0 ) ;
  assign n36214 = ( n35792 & n35844 ) | ( n35792 & n36202 ) | ( n35844 & n36202 ) ;
  assign n36213 = n35792 | n36202 ;
  assign n36215 = ( n36212 & ~n36214 ) | ( n36212 & n36213 ) | ( ~n36214 & n36213 ) ;
  assign n36219 = n35674 &  n35843 ;
  assign n36220 = n35842 &  n36219 ;
  assign n36208 = x79 | n35674 ;
  assign n36209 = x79 &  n35674 ;
  assign n36210 = ( n36208 & ~n36209 ) | ( n36208 & 1'b0 ) | ( ~n36209 & 1'b0 ) ;
  assign n36222 = ( n35791 & n35844 ) | ( n35791 & n36210 ) | ( n35844 & n36210 ) ;
  assign n36221 = n35791 | n36210 ;
  assign n36223 = ( n36220 & ~n36222 ) | ( n36220 & n36221 ) | ( ~n36222 & n36221 ) ;
  assign n36227 = n35682 &  n35843 ;
  assign n36228 = n35842 &  n36227 ;
  assign n36216 = x78 | n35682 ;
  assign n36217 = x78 &  n35682 ;
  assign n36218 = ( n36216 & ~n36217 ) | ( n36216 & 1'b0 ) | ( ~n36217 & 1'b0 ) ;
  assign n36230 = ( n35790 & n35844 ) | ( n35790 & n36218 ) | ( n35844 & n36218 ) ;
  assign n36229 = n35790 | n36218 ;
  assign n36231 = ( n36228 & ~n36230 ) | ( n36228 & n36229 ) | ( ~n36230 & n36229 ) ;
  assign n36235 = n35690 &  n35843 ;
  assign n36236 = n35842 &  n36235 ;
  assign n36224 = x77 | n35690 ;
  assign n36225 = x77 &  n35690 ;
  assign n36226 = ( n36224 & ~n36225 ) | ( n36224 & 1'b0 ) | ( ~n36225 & 1'b0 ) ;
  assign n36238 = ( n35789 & n35844 ) | ( n35789 & n36226 ) | ( n35844 & n36226 ) ;
  assign n36237 = n35789 | n36226 ;
  assign n36239 = ( n36236 & ~n36238 ) | ( n36236 & n36237 ) | ( ~n36238 & n36237 ) ;
  assign n36243 = n35698 &  n35843 ;
  assign n36244 = n35842 &  n36243 ;
  assign n36232 = x76 | n35698 ;
  assign n36233 = x76 &  n35698 ;
  assign n36234 = ( n36232 & ~n36233 ) | ( n36232 & 1'b0 ) | ( ~n36233 & 1'b0 ) ;
  assign n36246 = ( n35788 & n35844 ) | ( n35788 & n36234 ) | ( n35844 & n36234 ) ;
  assign n36245 = n35788 | n36234 ;
  assign n36247 = ( n36244 & ~n36246 ) | ( n36244 & n36245 ) | ( ~n36246 & n36245 ) ;
  assign n36251 = n35706 &  n35843 ;
  assign n36252 = n35842 &  n36251 ;
  assign n36240 = x75 | n35706 ;
  assign n36241 = x75 &  n35706 ;
  assign n36242 = ( n36240 & ~n36241 ) | ( n36240 & 1'b0 ) | ( ~n36241 & 1'b0 ) ;
  assign n36254 = ( n35787 & n35844 ) | ( n35787 & n36242 ) | ( n35844 & n36242 ) ;
  assign n36253 = n35787 | n36242 ;
  assign n36255 = ( n36252 & ~n36254 ) | ( n36252 & n36253 ) | ( ~n36254 & n36253 ) ;
  assign n36259 = n35714 &  n35843 ;
  assign n36260 = n35842 &  n36259 ;
  assign n36248 = x74 | n35714 ;
  assign n36249 = x74 &  n35714 ;
  assign n36250 = ( n36248 & ~n36249 ) | ( n36248 & 1'b0 ) | ( ~n36249 & 1'b0 ) ;
  assign n36262 = ( n35786 & n35844 ) | ( n35786 & n36250 ) | ( n35844 & n36250 ) ;
  assign n36261 = n35786 | n36250 ;
  assign n36263 = ( n36260 & ~n36262 ) | ( n36260 & n36261 ) | ( ~n36262 & n36261 ) ;
  assign n36267 = n35722 &  n35843 ;
  assign n36268 = n35842 &  n36267 ;
  assign n36256 = x73 | n35722 ;
  assign n36257 = x73 &  n35722 ;
  assign n36258 = ( n36256 & ~n36257 ) | ( n36256 & 1'b0 ) | ( ~n36257 & 1'b0 ) ;
  assign n36270 = ( n35785 & n35844 ) | ( n35785 & n36258 ) | ( n35844 & n36258 ) ;
  assign n36269 = n35785 | n36258 ;
  assign n36271 = ( n36268 & ~n36270 ) | ( n36268 & n36269 ) | ( ~n36270 & n36269 ) ;
  assign n36275 = n35730 &  n35843 ;
  assign n36276 = n35842 &  n36275 ;
  assign n36264 = x72 | n35730 ;
  assign n36265 = x72 &  n35730 ;
  assign n36266 = ( n36264 & ~n36265 ) | ( n36264 & 1'b0 ) | ( ~n36265 & 1'b0 ) ;
  assign n36278 = ( n35784 & n35844 ) | ( n35784 & n36266 ) | ( n35844 & n36266 ) ;
  assign n36277 = n35784 | n36266 ;
  assign n36279 = ( n36276 & ~n36278 ) | ( n36276 & n36277 ) | ( ~n36278 & n36277 ) ;
  assign n36283 = n35738 &  n35843 ;
  assign n36284 = n35842 &  n36283 ;
  assign n36272 = x71 | n35738 ;
  assign n36273 = x71 &  n35738 ;
  assign n36274 = ( n36272 & ~n36273 ) | ( n36272 & 1'b0 ) | ( ~n36273 & 1'b0 ) ;
  assign n36286 = ( n35783 & n35844 ) | ( n35783 & n36274 ) | ( n35844 & n36274 ) ;
  assign n36285 = n35783 | n36274 ;
  assign n36287 = ( n36284 & ~n36286 ) | ( n36284 & n36285 ) | ( ~n36286 & n36285 ) ;
  assign n36291 = n35746 &  n35843 ;
  assign n36292 = n35842 &  n36291 ;
  assign n36280 = x70 | n35746 ;
  assign n36281 = x70 &  n35746 ;
  assign n36282 = ( n36280 & ~n36281 ) | ( n36280 & 1'b0 ) | ( ~n36281 & 1'b0 ) ;
  assign n36294 = ( n35782 & n35844 ) | ( n35782 & n36282 ) | ( n35844 & n36282 ) ;
  assign n36293 = n35782 | n36282 ;
  assign n36295 = ( n36292 & ~n36294 ) | ( n36292 & n36293 ) | ( ~n36294 & n36293 ) ;
  assign n36299 = n35754 &  n35843 ;
  assign n36300 = n35842 &  n36299 ;
  assign n36288 = x69 | n35754 ;
  assign n36289 = x69 &  n35754 ;
  assign n36290 = ( n36288 & ~n36289 ) | ( n36288 & 1'b0 ) | ( ~n36289 & 1'b0 ) ;
  assign n36302 = ( n35781 & n35844 ) | ( n35781 & n36290 ) | ( n35844 & n36290 ) ;
  assign n36301 = n35781 | n36290 ;
  assign n36303 = ( n36300 & ~n36302 ) | ( n36300 & n36301 ) | ( ~n36302 & n36301 ) ;
  assign n36307 = n35762 &  n35843 ;
  assign n36308 = n35842 &  n36307 ;
  assign n36296 = x68 | n35762 ;
  assign n36297 = x68 &  n35762 ;
  assign n36298 = ( n36296 & ~n36297 ) | ( n36296 & 1'b0 ) | ( ~n36297 & 1'b0 ) ;
  assign n36310 = ( n35780 & n35844 ) | ( n35780 & n36298 ) | ( n35844 & n36298 ) ;
  assign n36309 = n35780 | n36298 ;
  assign n36311 = ( n36308 & ~n36310 ) | ( n36308 & n36309 ) | ( ~n36310 & n36309 ) ;
  assign n36315 = n35767 &  n35843 ;
  assign n36316 = n35842 &  n36315 ;
  assign n36304 = x67 | n35767 ;
  assign n36305 = x67 &  n35767 ;
  assign n36306 = ( n36304 & ~n36305 ) | ( n36304 & 1'b0 ) | ( ~n36305 & 1'b0 ) ;
  assign n36318 = ( n35779 & n35844 ) | ( n35779 & n36306 ) | ( n35844 & n36306 ) ;
  assign n36317 = n35779 | n36306 ;
  assign n36319 = ( n36316 & ~n36318 ) | ( n36316 & n36317 ) | ( ~n36318 & n36317 ) ;
  assign n36320 = n35773 &  n35843 ;
  assign n36321 = n35842 &  n36320 ;
  assign n36312 = x66 | n35773 ;
  assign n36313 = x66 &  n35773 ;
  assign n36314 = ( n36312 & ~n36313 ) | ( n36312 & 1'b0 ) | ( ~n36313 & 1'b0 ) ;
  assign n36322 = n35778 &  n36314 ;
  assign n36323 = ( n35778 & ~n35844 ) | ( n35778 & n36314 ) | ( ~n35844 & n36314 ) ;
  assign n36324 = ( n36321 & ~n36322 ) | ( n36321 & n36323 ) | ( ~n36322 & n36323 ) ;
  assign n36325 = ( x65 & ~n17483 ) | ( x65 & n35777 ) | ( ~n17483 & n35777 ) ;
  assign n36326 = ( n35778 & ~x65 ) | ( n35778 & n36325 ) | ( ~x65 & n36325 ) ;
  assign n36327 = ~n35844 & n36326 ;
  assign n36328 = n35777 &  n35843 ;
  assign n36329 = n35842 &  n36328 ;
  assign n36330 = n36327 | n36329 ;
  assign n36331 = ( x64 & ~n35844 ) | ( x64 & 1'b0 ) | ( ~n35844 & 1'b0 ) ;
  assign n36332 = ( x2 & ~n36331 ) | ( x2 & 1'b0 ) | ( ~n36331 & 1'b0 ) ;
  assign n36333 = ( n17483 & ~n35844 ) | ( n17483 & 1'b0 ) | ( ~n35844 & 1'b0 ) ;
  assign n36334 = n36332 | n36333 ;
  assign n36335 = ( x65 & ~n36334 ) | ( x65 & n18049 ) | ( ~n36334 & n18049 ) ;
  assign n36336 = ( x66 & ~n36330 ) | ( x66 & n36335 ) | ( ~n36330 & n36335 ) ;
  assign n36337 = ( x67 & ~n36324 ) | ( x67 & n36336 ) | ( ~n36324 & n36336 ) ;
  assign n36338 = ( x68 & ~n36319 ) | ( x68 & n36337 ) | ( ~n36319 & n36337 ) ;
  assign n36339 = ( x69 & ~n36311 ) | ( x69 & n36338 ) | ( ~n36311 & n36338 ) ;
  assign n36340 = ( x70 & ~n36303 ) | ( x70 & n36339 ) | ( ~n36303 & n36339 ) ;
  assign n36341 = ( x71 & ~n36295 ) | ( x71 & n36340 ) | ( ~n36295 & n36340 ) ;
  assign n36342 = ( x72 & ~n36287 ) | ( x72 & n36341 ) | ( ~n36287 & n36341 ) ;
  assign n36343 = ( x73 & ~n36279 ) | ( x73 & n36342 ) | ( ~n36279 & n36342 ) ;
  assign n36344 = ( x74 & ~n36271 ) | ( x74 & n36343 ) | ( ~n36271 & n36343 ) ;
  assign n36345 = ( x75 & ~n36263 ) | ( x75 & n36344 ) | ( ~n36263 & n36344 ) ;
  assign n36346 = ( x76 & ~n36255 ) | ( x76 & n36345 ) | ( ~n36255 & n36345 ) ;
  assign n36347 = ( x77 & ~n36247 ) | ( x77 & n36346 ) | ( ~n36247 & n36346 ) ;
  assign n36348 = ( x78 & ~n36239 ) | ( x78 & n36347 ) | ( ~n36239 & n36347 ) ;
  assign n36349 = ( x79 & ~n36231 ) | ( x79 & n36348 ) | ( ~n36231 & n36348 ) ;
  assign n36350 = ( x80 & ~n36223 ) | ( x80 & n36349 ) | ( ~n36223 & n36349 ) ;
  assign n36351 = ( x81 & ~n36215 ) | ( x81 & n36350 ) | ( ~n36215 & n36350 ) ;
  assign n36352 = ( x82 & ~n36207 ) | ( x82 & n36351 ) | ( ~n36207 & n36351 ) ;
  assign n36353 = ( x83 & ~n36199 ) | ( x83 & n36352 ) | ( ~n36199 & n36352 ) ;
  assign n36354 = ( x84 & ~n36191 ) | ( x84 & n36353 ) | ( ~n36191 & n36353 ) ;
  assign n36355 = ( x85 & ~n36183 ) | ( x85 & n36354 ) | ( ~n36183 & n36354 ) ;
  assign n36356 = ( x86 & ~n36175 ) | ( x86 & n36355 ) | ( ~n36175 & n36355 ) ;
  assign n36357 = ( x87 & ~n36167 ) | ( x87 & n36356 ) | ( ~n36167 & n36356 ) ;
  assign n36358 = ( x88 & ~n36159 ) | ( x88 & n36357 ) | ( ~n36159 & n36357 ) ;
  assign n36359 = ( x89 & ~n36151 ) | ( x89 & n36358 ) | ( ~n36151 & n36358 ) ;
  assign n36360 = ( x90 & ~n36143 ) | ( x90 & n36359 ) | ( ~n36143 & n36359 ) ;
  assign n36361 = ( x91 & ~n36135 ) | ( x91 & n36360 ) | ( ~n36135 & n36360 ) ;
  assign n36362 = ( x92 & ~n36127 ) | ( x92 & n36361 ) | ( ~n36127 & n36361 ) ;
  assign n36363 = ( x93 & ~n36119 ) | ( x93 & n36362 ) | ( ~n36119 & n36362 ) ;
  assign n36364 = ( x94 & ~n36111 ) | ( x94 & n36363 ) | ( ~n36111 & n36363 ) ;
  assign n36365 = ( x95 & ~n36103 ) | ( x95 & n36364 ) | ( ~n36103 & n36364 ) ;
  assign n36366 = ( x96 & ~n36095 ) | ( x96 & n36365 ) | ( ~n36095 & n36365 ) ;
  assign n36367 = ( x97 & ~n36087 ) | ( x97 & n36366 ) | ( ~n36087 & n36366 ) ;
  assign n36368 = ( x98 & ~n36079 ) | ( x98 & n36367 ) | ( ~n36079 & n36367 ) ;
  assign n36369 = ( x99 & ~n36071 ) | ( x99 & n36368 ) | ( ~n36071 & n36368 ) ;
  assign n36370 = ( x100 & ~n36063 ) | ( x100 & n36369 ) | ( ~n36063 & n36369 ) ;
  assign n36371 = ( x101 & ~n36055 ) | ( x101 & n36370 ) | ( ~n36055 & n36370 ) ;
  assign n36372 = ( x102 & ~n36047 ) | ( x102 & n36371 ) | ( ~n36047 & n36371 ) ;
  assign n36373 = ( x103 & ~n36039 ) | ( x103 & n36372 ) | ( ~n36039 & n36372 ) ;
  assign n36374 = ( x104 & ~n36031 ) | ( x104 & n36373 ) | ( ~n36031 & n36373 ) ;
  assign n36375 = ( x105 & ~n36023 ) | ( x105 & n36374 ) | ( ~n36023 & n36374 ) ;
  assign n36376 = ( x106 & ~n36015 ) | ( x106 & n36375 ) | ( ~n36015 & n36375 ) ;
  assign n36377 = ( x107 & ~n36007 ) | ( x107 & n36376 ) | ( ~n36007 & n36376 ) ;
  assign n36378 = ( x108 & ~n35999 ) | ( x108 & n36377 ) | ( ~n35999 & n36377 ) ;
  assign n36379 = ( x109 & ~n35991 ) | ( x109 & n36378 ) | ( ~n35991 & n36378 ) ;
  assign n36380 = ( x110 & ~n35983 ) | ( x110 & n36379 ) | ( ~n35983 & n36379 ) ;
  assign n36381 = ( x111 & ~n35975 ) | ( x111 & n36380 ) | ( ~n35975 & n36380 ) ;
  assign n36382 = ( x112 & ~n35967 ) | ( x112 & n36381 ) | ( ~n35967 & n36381 ) ;
  assign n36383 = ( x113 & ~n35959 ) | ( x113 & n36382 ) | ( ~n35959 & n36382 ) ;
  assign n36384 = ( x114 & ~n35951 ) | ( x114 & n36383 ) | ( ~n35951 & n36383 ) ;
  assign n36385 = ( x115 & ~n35943 ) | ( x115 & n36384 ) | ( ~n35943 & n36384 ) ;
  assign n36386 = ( x116 & ~n35935 ) | ( x116 & n36385 ) | ( ~n35935 & n36385 ) ;
  assign n36387 = ( x117 & ~n35927 ) | ( x117 & n36386 ) | ( ~n35927 & n36386 ) ;
  assign n36388 = ( x118 & ~n35919 ) | ( x118 & n36387 ) | ( ~n35919 & n36387 ) ;
  assign n36389 = ( x119 & ~n35911 ) | ( x119 & n36388 ) | ( ~n35911 & n36388 ) ;
  assign n36390 = ( x120 & ~n35903 ) | ( x120 & n36389 ) | ( ~n35903 & n36389 ) ;
  assign n36391 = ( x121 & ~n35895 ) | ( x121 & n36390 ) | ( ~n35895 & n36390 ) ;
  assign n36392 = ( x122 & ~n35887 ) | ( x122 & n36391 ) | ( ~n35887 & n36391 ) ;
  assign n36393 = ( x123 & ~n35879 ) | ( x123 & n36392 ) | ( ~n35879 & n36392 ) ;
  assign n36394 = ( x124 & ~n35871 ) | ( x124 & n36393 ) | ( ~n35871 & n36393 ) ;
  assign n36395 = ( x125 & ~n35863 ) | ( x125 & n36394 ) | ( ~n35863 & n36394 ) ;
  assign n36396 = ( x126 & ~n35305 ) | ( x126 & 1'b0 ) | ( ~n35305 & 1'b0 ) ;
  assign n36397 = ~n35851 & n36396 ;
  assign n36398 = ( n36395 & ~n35855 ) | ( n36395 & n36397 ) | ( ~n35855 & n36397 ) ;
  assign n36399 = ( n35855 & ~x127 ) | ( n35855 & n36398 ) | ( ~x127 & n36398 ) ;
  assign n36400 = x127 | n36399 ;
  assign n36407 = n151 &  n35854 ;
  assign n36408 = n36400 &  n36407 ;
  assign n36401 = ~n35854 |  n151 ;
  assign n36402 = n36400 &  n36401 ;
  assign n36406 = n35855 | n36397 ;
  assign n36410 = ( n36395 & n36402 ) | ( n36395 & n36406 ) | ( n36402 & n36406 ) ;
  assign n36409 = n36395 | n36406 ;
  assign n36411 = ( n36408 & ~n36410 ) | ( n36408 & n36409 ) | ( ~n36410 & n36409 ) ;
  assign n36415 = n35863 &  n36401 ;
  assign n36416 = n36400 &  n36415 ;
  assign n36403 = x125 | n35863 ;
  assign n36404 = x125 &  n35863 ;
  assign n36405 = ( n36403 & ~n36404 ) | ( n36403 & 1'b0 ) | ( ~n36404 & 1'b0 ) ;
  assign n36418 = ( n36394 & n36402 ) | ( n36394 & n36405 ) | ( n36402 & n36405 ) ;
  assign n36417 = n36394 | n36405 ;
  assign n36419 = ( n36416 & ~n36418 ) | ( n36416 & n36417 ) | ( ~n36418 & n36417 ) ;
  assign n36423 = n35871 &  n36401 ;
  assign n36424 = n36400 &  n36423 ;
  assign n36412 = x124 | n35871 ;
  assign n36413 = x124 &  n35871 ;
  assign n36414 = ( n36412 & ~n36413 ) | ( n36412 & 1'b0 ) | ( ~n36413 & 1'b0 ) ;
  assign n36426 = ( n36393 & n36402 ) | ( n36393 & n36414 ) | ( n36402 & n36414 ) ;
  assign n36425 = n36393 | n36414 ;
  assign n36427 = ( n36424 & ~n36426 ) | ( n36424 & n36425 ) | ( ~n36426 & n36425 ) ;
  assign n36431 = n35879 &  n36401 ;
  assign n36432 = n36400 &  n36431 ;
  assign n36420 = x123 | n35879 ;
  assign n36421 = x123 &  n35879 ;
  assign n36422 = ( n36420 & ~n36421 ) | ( n36420 & 1'b0 ) | ( ~n36421 & 1'b0 ) ;
  assign n36434 = ( n36392 & n36402 ) | ( n36392 & n36422 ) | ( n36402 & n36422 ) ;
  assign n36433 = n36392 | n36422 ;
  assign n36435 = ( n36432 & ~n36434 ) | ( n36432 & n36433 ) | ( ~n36434 & n36433 ) ;
  assign n36439 = n35887 &  n36401 ;
  assign n36440 = n36400 &  n36439 ;
  assign n36428 = x122 | n35887 ;
  assign n36429 = x122 &  n35887 ;
  assign n36430 = ( n36428 & ~n36429 ) | ( n36428 & 1'b0 ) | ( ~n36429 & 1'b0 ) ;
  assign n36442 = ( n36391 & n36402 ) | ( n36391 & n36430 ) | ( n36402 & n36430 ) ;
  assign n36441 = n36391 | n36430 ;
  assign n36443 = ( n36440 & ~n36442 ) | ( n36440 & n36441 ) | ( ~n36442 & n36441 ) ;
  assign n36447 = n35895 &  n36401 ;
  assign n36448 = n36400 &  n36447 ;
  assign n36436 = x121 | n35895 ;
  assign n36437 = x121 &  n35895 ;
  assign n36438 = ( n36436 & ~n36437 ) | ( n36436 & 1'b0 ) | ( ~n36437 & 1'b0 ) ;
  assign n36450 = ( n36390 & n36402 ) | ( n36390 & n36438 ) | ( n36402 & n36438 ) ;
  assign n36449 = n36390 | n36438 ;
  assign n36451 = ( n36448 & ~n36450 ) | ( n36448 & n36449 ) | ( ~n36450 & n36449 ) ;
  assign n36455 = n35903 &  n36401 ;
  assign n36456 = n36400 &  n36455 ;
  assign n36444 = x120 | n35903 ;
  assign n36445 = x120 &  n35903 ;
  assign n36446 = ( n36444 & ~n36445 ) | ( n36444 & 1'b0 ) | ( ~n36445 & 1'b0 ) ;
  assign n36458 = ( n36389 & n36402 ) | ( n36389 & n36446 ) | ( n36402 & n36446 ) ;
  assign n36457 = n36389 | n36446 ;
  assign n36459 = ( n36456 & ~n36458 ) | ( n36456 & n36457 ) | ( ~n36458 & n36457 ) ;
  assign n36463 = n35911 &  n36401 ;
  assign n36464 = n36400 &  n36463 ;
  assign n36452 = x119 | n35911 ;
  assign n36453 = x119 &  n35911 ;
  assign n36454 = ( n36452 & ~n36453 ) | ( n36452 & 1'b0 ) | ( ~n36453 & 1'b0 ) ;
  assign n36466 = ( n36388 & n36402 ) | ( n36388 & n36454 ) | ( n36402 & n36454 ) ;
  assign n36465 = n36388 | n36454 ;
  assign n36467 = ( n36464 & ~n36466 ) | ( n36464 & n36465 ) | ( ~n36466 & n36465 ) ;
  assign n36471 = n35919 &  n36401 ;
  assign n36472 = n36400 &  n36471 ;
  assign n36460 = x118 | n35919 ;
  assign n36461 = x118 &  n35919 ;
  assign n36462 = ( n36460 & ~n36461 ) | ( n36460 & 1'b0 ) | ( ~n36461 & 1'b0 ) ;
  assign n36474 = ( n36387 & n36402 ) | ( n36387 & n36462 ) | ( n36402 & n36462 ) ;
  assign n36473 = n36387 | n36462 ;
  assign n36475 = ( n36472 & ~n36474 ) | ( n36472 & n36473 ) | ( ~n36474 & n36473 ) ;
  assign n36479 = n35927 &  n36401 ;
  assign n36480 = n36400 &  n36479 ;
  assign n36468 = x117 | n35927 ;
  assign n36469 = x117 &  n35927 ;
  assign n36470 = ( n36468 & ~n36469 ) | ( n36468 & 1'b0 ) | ( ~n36469 & 1'b0 ) ;
  assign n36482 = ( n36386 & n36402 ) | ( n36386 & n36470 ) | ( n36402 & n36470 ) ;
  assign n36481 = n36386 | n36470 ;
  assign n36483 = ( n36480 & ~n36482 ) | ( n36480 & n36481 ) | ( ~n36482 & n36481 ) ;
  assign n36487 = n35935 &  n36401 ;
  assign n36488 = n36400 &  n36487 ;
  assign n36476 = x116 | n35935 ;
  assign n36477 = x116 &  n35935 ;
  assign n36478 = ( n36476 & ~n36477 ) | ( n36476 & 1'b0 ) | ( ~n36477 & 1'b0 ) ;
  assign n36490 = ( n36385 & n36402 ) | ( n36385 & n36478 ) | ( n36402 & n36478 ) ;
  assign n36489 = n36385 | n36478 ;
  assign n36491 = ( n36488 & ~n36490 ) | ( n36488 & n36489 ) | ( ~n36490 & n36489 ) ;
  assign n36495 = n35943 &  n36401 ;
  assign n36496 = n36400 &  n36495 ;
  assign n36484 = x115 | n35943 ;
  assign n36485 = x115 &  n35943 ;
  assign n36486 = ( n36484 & ~n36485 ) | ( n36484 & 1'b0 ) | ( ~n36485 & 1'b0 ) ;
  assign n36498 = ( n36384 & n36402 ) | ( n36384 & n36486 ) | ( n36402 & n36486 ) ;
  assign n36497 = n36384 | n36486 ;
  assign n36499 = ( n36496 & ~n36498 ) | ( n36496 & n36497 ) | ( ~n36498 & n36497 ) ;
  assign n36503 = n35951 &  n36401 ;
  assign n36504 = n36400 &  n36503 ;
  assign n36492 = x114 | n35951 ;
  assign n36493 = x114 &  n35951 ;
  assign n36494 = ( n36492 & ~n36493 ) | ( n36492 & 1'b0 ) | ( ~n36493 & 1'b0 ) ;
  assign n36506 = ( n36383 & n36402 ) | ( n36383 & n36494 ) | ( n36402 & n36494 ) ;
  assign n36505 = n36383 | n36494 ;
  assign n36507 = ( n36504 & ~n36506 ) | ( n36504 & n36505 ) | ( ~n36506 & n36505 ) ;
  assign n36511 = n35959 &  n36401 ;
  assign n36512 = n36400 &  n36511 ;
  assign n36500 = x113 | n35959 ;
  assign n36501 = x113 &  n35959 ;
  assign n36502 = ( n36500 & ~n36501 ) | ( n36500 & 1'b0 ) | ( ~n36501 & 1'b0 ) ;
  assign n36514 = ( n36382 & n36402 ) | ( n36382 & n36502 ) | ( n36402 & n36502 ) ;
  assign n36513 = n36382 | n36502 ;
  assign n36515 = ( n36512 & ~n36514 ) | ( n36512 & n36513 ) | ( ~n36514 & n36513 ) ;
  assign n36519 = n35967 &  n36401 ;
  assign n36520 = n36400 &  n36519 ;
  assign n36508 = x112 | n35967 ;
  assign n36509 = x112 &  n35967 ;
  assign n36510 = ( n36508 & ~n36509 ) | ( n36508 & 1'b0 ) | ( ~n36509 & 1'b0 ) ;
  assign n36522 = ( n36381 & n36402 ) | ( n36381 & n36510 ) | ( n36402 & n36510 ) ;
  assign n36521 = n36381 | n36510 ;
  assign n36523 = ( n36520 & ~n36522 ) | ( n36520 & n36521 ) | ( ~n36522 & n36521 ) ;
  assign n36527 = n35975 &  n36401 ;
  assign n36528 = n36400 &  n36527 ;
  assign n36516 = x111 | n35975 ;
  assign n36517 = x111 &  n35975 ;
  assign n36518 = ( n36516 & ~n36517 ) | ( n36516 & 1'b0 ) | ( ~n36517 & 1'b0 ) ;
  assign n36530 = ( n36380 & n36402 ) | ( n36380 & n36518 ) | ( n36402 & n36518 ) ;
  assign n36529 = n36380 | n36518 ;
  assign n36531 = ( n36528 & ~n36530 ) | ( n36528 & n36529 ) | ( ~n36530 & n36529 ) ;
  assign n36535 = n35983 &  n36401 ;
  assign n36536 = n36400 &  n36535 ;
  assign n36524 = x110 | n35983 ;
  assign n36525 = x110 &  n35983 ;
  assign n36526 = ( n36524 & ~n36525 ) | ( n36524 & 1'b0 ) | ( ~n36525 & 1'b0 ) ;
  assign n36538 = ( n36379 & n36402 ) | ( n36379 & n36526 ) | ( n36402 & n36526 ) ;
  assign n36537 = n36379 | n36526 ;
  assign n36539 = ( n36536 & ~n36538 ) | ( n36536 & n36537 ) | ( ~n36538 & n36537 ) ;
  assign n36543 = n35991 &  n36401 ;
  assign n36544 = n36400 &  n36543 ;
  assign n36532 = x109 | n35991 ;
  assign n36533 = x109 &  n35991 ;
  assign n36534 = ( n36532 & ~n36533 ) | ( n36532 & 1'b0 ) | ( ~n36533 & 1'b0 ) ;
  assign n36546 = ( n36378 & n36402 ) | ( n36378 & n36534 ) | ( n36402 & n36534 ) ;
  assign n36545 = n36378 | n36534 ;
  assign n36547 = ( n36544 & ~n36546 ) | ( n36544 & n36545 ) | ( ~n36546 & n36545 ) ;
  assign n36551 = n35999 &  n36401 ;
  assign n36552 = n36400 &  n36551 ;
  assign n36540 = x108 | n35999 ;
  assign n36541 = x108 &  n35999 ;
  assign n36542 = ( n36540 & ~n36541 ) | ( n36540 & 1'b0 ) | ( ~n36541 & 1'b0 ) ;
  assign n36554 = ( n36377 & n36402 ) | ( n36377 & n36542 ) | ( n36402 & n36542 ) ;
  assign n36553 = n36377 | n36542 ;
  assign n36555 = ( n36552 & ~n36554 ) | ( n36552 & n36553 ) | ( ~n36554 & n36553 ) ;
  assign n36559 = n36007 &  n36401 ;
  assign n36560 = n36400 &  n36559 ;
  assign n36548 = x107 | n36007 ;
  assign n36549 = x107 &  n36007 ;
  assign n36550 = ( n36548 & ~n36549 ) | ( n36548 & 1'b0 ) | ( ~n36549 & 1'b0 ) ;
  assign n36562 = ( n36376 & n36402 ) | ( n36376 & n36550 ) | ( n36402 & n36550 ) ;
  assign n36561 = n36376 | n36550 ;
  assign n36563 = ( n36560 & ~n36562 ) | ( n36560 & n36561 ) | ( ~n36562 & n36561 ) ;
  assign n36567 = n36015 &  n36401 ;
  assign n36568 = n36400 &  n36567 ;
  assign n36556 = x106 | n36015 ;
  assign n36557 = x106 &  n36015 ;
  assign n36558 = ( n36556 & ~n36557 ) | ( n36556 & 1'b0 ) | ( ~n36557 & 1'b0 ) ;
  assign n36570 = ( n36375 & n36402 ) | ( n36375 & n36558 ) | ( n36402 & n36558 ) ;
  assign n36569 = n36375 | n36558 ;
  assign n36571 = ( n36568 & ~n36570 ) | ( n36568 & n36569 ) | ( ~n36570 & n36569 ) ;
  assign n36575 = n36023 &  n36401 ;
  assign n36576 = n36400 &  n36575 ;
  assign n36564 = x105 | n36023 ;
  assign n36565 = x105 &  n36023 ;
  assign n36566 = ( n36564 & ~n36565 ) | ( n36564 & 1'b0 ) | ( ~n36565 & 1'b0 ) ;
  assign n36578 = ( n36374 & n36402 ) | ( n36374 & n36566 ) | ( n36402 & n36566 ) ;
  assign n36577 = n36374 | n36566 ;
  assign n36579 = ( n36576 & ~n36578 ) | ( n36576 & n36577 ) | ( ~n36578 & n36577 ) ;
  assign n36583 = n36031 &  n36401 ;
  assign n36584 = n36400 &  n36583 ;
  assign n36572 = x104 | n36031 ;
  assign n36573 = x104 &  n36031 ;
  assign n36574 = ( n36572 & ~n36573 ) | ( n36572 & 1'b0 ) | ( ~n36573 & 1'b0 ) ;
  assign n36586 = ( n36373 & n36402 ) | ( n36373 & n36574 ) | ( n36402 & n36574 ) ;
  assign n36585 = n36373 | n36574 ;
  assign n36587 = ( n36584 & ~n36586 ) | ( n36584 & n36585 ) | ( ~n36586 & n36585 ) ;
  assign n36591 = n36039 &  n36401 ;
  assign n36592 = n36400 &  n36591 ;
  assign n36580 = x103 | n36039 ;
  assign n36581 = x103 &  n36039 ;
  assign n36582 = ( n36580 & ~n36581 ) | ( n36580 & 1'b0 ) | ( ~n36581 & 1'b0 ) ;
  assign n36594 = ( n36372 & n36402 ) | ( n36372 & n36582 ) | ( n36402 & n36582 ) ;
  assign n36593 = n36372 | n36582 ;
  assign n36595 = ( n36592 & ~n36594 ) | ( n36592 & n36593 ) | ( ~n36594 & n36593 ) ;
  assign n36599 = n36047 &  n36401 ;
  assign n36600 = n36400 &  n36599 ;
  assign n36588 = x102 | n36047 ;
  assign n36589 = x102 &  n36047 ;
  assign n36590 = ( n36588 & ~n36589 ) | ( n36588 & 1'b0 ) | ( ~n36589 & 1'b0 ) ;
  assign n36602 = ( n36371 & n36402 ) | ( n36371 & n36590 ) | ( n36402 & n36590 ) ;
  assign n36601 = n36371 | n36590 ;
  assign n36603 = ( n36600 & ~n36602 ) | ( n36600 & n36601 ) | ( ~n36602 & n36601 ) ;
  assign n36607 = n36055 &  n36401 ;
  assign n36608 = n36400 &  n36607 ;
  assign n36596 = x101 | n36055 ;
  assign n36597 = x101 &  n36055 ;
  assign n36598 = ( n36596 & ~n36597 ) | ( n36596 & 1'b0 ) | ( ~n36597 & 1'b0 ) ;
  assign n36610 = ( n36370 & n36402 ) | ( n36370 & n36598 ) | ( n36402 & n36598 ) ;
  assign n36609 = n36370 | n36598 ;
  assign n36611 = ( n36608 & ~n36610 ) | ( n36608 & n36609 ) | ( ~n36610 & n36609 ) ;
  assign n36615 = n36063 &  n36401 ;
  assign n36616 = n36400 &  n36615 ;
  assign n36604 = x100 | n36063 ;
  assign n36605 = x100 &  n36063 ;
  assign n36606 = ( n36604 & ~n36605 ) | ( n36604 & 1'b0 ) | ( ~n36605 & 1'b0 ) ;
  assign n36618 = ( n36369 & n36402 ) | ( n36369 & n36606 ) | ( n36402 & n36606 ) ;
  assign n36617 = n36369 | n36606 ;
  assign n36619 = ( n36616 & ~n36618 ) | ( n36616 & n36617 ) | ( ~n36618 & n36617 ) ;
  assign n36623 = n36071 &  n36401 ;
  assign n36624 = n36400 &  n36623 ;
  assign n36612 = x99 | n36071 ;
  assign n36613 = x99 &  n36071 ;
  assign n36614 = ( n36612 & ~n36613 ) | ( n36612 & 1'b0 ) | ( ~n36613 & 1'b0 ) ;
  assign n36626 = ( n36368 & n36402 ) | ( n36368 & n36614 ) | ( n36402 & n36614 ) ;
  assign n36625 = n36368 | n36614 ;
  assign n36627 = ( n36624 & ~n36626 ) | ( n36624 & n36625 ) | ( ~n36626 & n36625 ) ;
  assign n36631 = n36079 &  n36401 ;
  assign n36632 = n36400 &  n36631 ;
  assign n36620 = x98 | n36079 ;
  assign n36621 = x98 &  n36079 ;
  assign n36622 = ( n36620 & ~n36621 ) | ( n36620 & 1'b0 ) | ( ~n36621 & 1'b0 ) ;
  assign n36634 = ( n36367 & n36402 ) | ( n36367 & n36622 ) | ( n36402 & n36622 ) ;
  assign n36633 = n36367 | n36622 ;
  assign n36635 = ( n36632 & ~n36634 ) | ( n36632 & n36633 ) | ( ~n36634 & n36633 ) ;
  assign n36639 = n36087 &  n36401 ;
  assign n36640 = n36400 &  n36639 ;
  assign n36628 = x97 | n36087 ;
  assign n36629 = x97 &  n36087 ;
  assign n36630 = ( n36628 & ~n36629 ) | ( n36628 & 1'b0 ) | ( ~n36629 & 1'b0 ) ;
  assign n36642 = ( n36366 & n36402 ) | ( n36366 & n36630 ) | ( n36402 & n36630 ) ;
  assign n36641 = n36366 | n36630 ;
  assign n36643 = ( n36640 & ~n36642 ) | ( n36640 & n36641 ) | ( ~n36642 & n36641 ) ;
  assign n36647 = n36095 &  n36401 ;
  assign n36648 = n36400 &  n36647 ;
  assign n36636 = x96 | n36095 ;
  assign n36637 = x96 &  n36095 ;
  assign n36638 = ( n36636 & ~n36637 ) | ( n36636 & 1'b0 ) | ( ~n36637 & 1'b0 ) ;
  assign n36650 = ( n36365 & n36402 ) | ( n36365 & n36638 ) | ( n36402 & n36638 ) ;
  assign n36649 = n36365 | n36638 ;
  assign n36651 = ( n36648 & ~n36650 ) | ( n36648 & n36649 ) | ( ~n36650 & n36649 ) ;
  assign n36655 = n36103 &  n36401 ;
  assign n36656 = n36400 &  n36655 ;
  assign n36644 = x95 | n36103 ;
  assign n36645 = x95 &  n36103 ;
  assign n36646 = ( n36644 & ~n36645 ) | ( n36644 & 1'b0 ) | ( ~n36645 & 1'b0 ) ;
  assign n36658 = ( n36364 & n36402 ) | ( n36364 & n36646 ) | ( n36402 & n36646 ) ;
  assign n36657 = n36364 | n36646 ;
  assign n36659 = ( n36656 & ~n36658 ) | ( n36656 & n36657 ) | ( ~n36658 & n36657 ) ;
  assign n36663 = n36111 &  n36401 ;
  assign n36664 = n36400 &  n36663 ;
  assign n36652 = x94 | n36111 ;
  assign n36653 = x94 &  n36111 ;
  assign n36654 = ( n36652 & ~n36653 ) | ( n36652 & 1'b0 ) | ( ~n36653 & 1'b0 ) ;
  assign n36666 = ( n36363 & n36402 ) | ( n36363 & n36654 ) | ( n36402 & n36654 ) ;
  assign n36665 = n36363 | n36654 ;
  assign n36667 = ( n36664 & ~n36666 ) | ( n36664 & n36665 ) | ( ~n36666 & n36665 ) ;
  assign n36671 = n36119 &  n36401 ;
  assign n36672 = n36400 &  n36671 ;
  assign n36660 = x93 | n36119 ;
  assign n36661 = x93 &  n36119 ;
  assign n36662 = ( n36660 & ~n36661 ) | ( n36660 & 1'b0 ) | ( ~n36661 & 1'b0 ) ;
  assign n36674 = ( n36362 & n36402 ) | ( n36362 & n36662 ) | ( n36402 & n36662 ) ;
  assign n36673 = n36362 | n36662 ;
  assign n36675 = ( n36672 & ~n36674 ) | ( n36672 & n36673 ) | ( ~n36674 & n36673 ) ;
  assign n36679 = n36127 &  n36401 ;
  assign n36680 = n36400 &  n36679 ;
  assign n36668 = x92 | n36127 ;
  assign n36669 = x92 &  n36127 ;
  assign n36670 = ( n36668 & ~n36669 ) | ( n36668 & 1'b0 ) | ( ~n36669 & 1'b0 ) ;
  assign n36682 = ( n36361 & n36402 ) | ( n36361 & n36670 ) | ( n36402 & n36670 ) ;
  assign n36681 = n36361 | n36670 ;
  assign n36683 = ( n36680 & ~n36682 ) | ( n36680 & n36681 ) | ( ~n36682 & n36681 ) ;
  assign n36687 = n36135 &  n36401 ;
  assign n36688 = n36400 &  n36687 ;
  assign n36676 = x91 | n36135 ;
  assign n36677 = x91 &  n36135 ;
  assign n36678 = ( n36676 & ~n36677 ) | ( n36676 & 1'b0 ) | ( ~n36677 & 1'b0 ) ;
  assign n36690 = ( n36360 & n36402 ) | ( n36360 & n36678 ) | ( n36402 & n36678 ) ;
  assign n36689 = n36360 | n36678 ;
  assign n36691 = ( n36688 & ~n36690 ) | ( n36688 & n36689 ) | ( ~n36690 & n36689 ) ;
  assign n36695 = n36143 &  n36401 ;
  assign n36696 = n36400 &  n36695 ;
  assign n36684 = x90 | n36143 ;
  assign n36685 = x90 &  n36143 ;
  assign n36686 = ( n36684 & ~n36685 ) | ( n36684 & 1'b0 ) | ( ~n36685 & 1'b0 ) ;
  assign n36698 = ( n36359 & n36402 ) | ( n36359 & n36686 ) | ( n36402 & n36686 ) ;
  assign n36697 = n36359 | n36686 ;
  assign n36699 = ( n36696 & ~n36698 ) | ( n36696 & n36697 ) | ( ~n36698 & n36697 ) ;
  assign n36703 = n36151 &  n36401 ;
  assign n36704 = n36400 &  n36703 ;
  assign n36692 = x89 | n36151 ;
  assign n36693 = x89 &  n36151 ;
  assign n36694 = ( n36692 & ~n36693 ) | ( n36692 & 1'b0 ) | ( ~n36693 & 1'b0 ) ;
  assign n36706 = ( n36358 & n36402 ) | ( n36358 & n36694 ) | ( n36402 & n36694 ) ;
  assign n36705 = n36358 | n36694 ;
  assign n36707 = ( n36704 & ~n36706 ) | ( n36704 & n36705 ) | ( ~n36706 & n36705 ) ;
  assign n36711 = n36159 &  n36401 ;
  assign n36712 = n36400 &  n36711 ;
  assign n36700 = x88 | n36159 ;
  assign n36701 = x88 &  n36159 ;
  assign n36702 = ( n36700 & ~n36701 ) | ( n36700 & 1'b0 ) | ( ~n36701 & 1'b0 ) ;
  assign n36714 = ( n36357 & n36402 ) | ( n36357 & n36702 ) | ( n36402 & n36702 ) ;
  assign n36713 = n36357 | n36702 ;
  assign n36715 = ( n36712 & ~n36714 ) | ( n36712 & n36713 ) | ( ~n36714 & n36713 ) ;
  assign n36719 = n36167 &  n36401 ;
  assign n36720 = n36400 &  n36719 ;
  assign n36708 = x87 | n36167 ;
  assign n36709 = x87 &  n36167 ;
  assign n36710 = ( n36708 & ~n36709 ) | ( n36708 & 1'b0 ) | ( ~n36709 & 1'b0 ) ;
  assign n36722 = ( n36356 & n36402 ) | ( n36356 & n36710 ) | ( n36402 & n36710 ) ;
  assign n36721 = n36356 | n36710 ;
  assign n36723 = ( n36720 & ~n36722 ) | ( n36720 & n36721 ) | ( ~n36722 & n36721 ) ;
  assign n36727 = n36175 &  n36401 ;
  assign n36728 = n36400 &  n36727 ;
  assign n36716 = x86 | n36175 ;
  assign n36717 = x86 &  n36175 ;
  assign n36718 = ( n36716 & ~n36717 ) | ( n36716 & 1'b0 ) | ( ~n36717 & 1'b0 ) ;
  assign n36730 = ( n36355 & n36402 ) | ( n36355 & n36718 ) | ( n36402 & n36718 ) ;
  assign n36729 = n36355 | n36718 ;
  assign n36731 = ( n36728 & ~n36730 ) | ( n36728 & n36729 ) | ( ~n36730 & n36729 ) ;
  assign n36735 = n36183 &  n36401 ;
  assign n36736 = n36400 &  n36735 ;
  assign n36724 = x85 | n36183 ;
  assign n36725 = x85 &  n36183 ;
  assign n36726 = ( n36724 & ~n36725 ) | ( n36724 & 1'b0 ) | ( ~n36725 & 1'b0 ) ;
  assign n36738 = ( n36354 & n36402 ) | ( n36354 & n36726 ) | ( n36402 & n36726 ) ;
  assign n36737 = n36354 | n36726 ;
  assign n36739 = ( n36736 & ~n36738 ) | ( n36736 & n36737 ) | ( ~n36738 & n36737 ) ;
  assign n36743 = n36191 &  n36401 ;
  assign n36744 = n36400 &  n36743 ;
  assign n36732 = x84 | n36191 ;
  assign n36733 = x84 &  n36191 ;
  assign n36734 = ( n36732 & ~n36733 ) | ( n36732 & 1'b0 ) | ( ~n36733 & 1'b0 ) ;
  assign n36746 = ( n36353 & n36402 ) | ( n36353 & n36734 ) | ( n36402 & n36734 ) ;
  assign n36745 = n36353 | n36734 ;
  assign n36747 = ( n36744 & ~n36746 ) | ( n36744 & n36745 ) | ( ~n36746 & n36745 ) ;
  assign n36751 = n36199 &  n36401 ;
  assign n36752 = n36400 &  n36751 ;
  assign n36740 = x83 | n36199 ;
  assign n36741 = x83 &  n36199 ;
  assign n36742 = ( n36740 & ~n36741 ) | ( n36740 & 1'b0 ) | ( ~n36741 & 1'b0 ) ;
  assign n36754 = ( n36352 & n36402 ) | ( n36352 & n36742 ) | ( n36402 & n36742 ) ;
  assign n36753 = n36352 | n36742 ;
  assign n36755 = ( n36752 & ~n36754 ) | ( n36752 & n36753 ) | ( ~n36754 & n36753 ) ;
  assign n36759 = n36207 &  n36401 ;
  assign n36760 = n36400 &  n36759 ;
  assign n36748 = x82 | n36207 ;
  assign n36749 = x82 &  n36207 ;
  assign n36750 = ( n36748 & ~n36749 ) | ( n36748 & 1'b0 ) | ( ~n36749 & 1'b0 ) ;
  assign n36762 = ( n36351 & n36402 ) | ( n36351 & n36750 ) | ( n36402 & n36750 ) ;
  assign n36761 = n36351 | n36750 ;
  assign n36763 = ( n36760 & ~n36762 ) | ( n36760 & n36761 ) | ( ~n36762 & n36761 ) ;
  assign n36767 = n36215 &  n36401 ;
  assign n36768 = n36400 &  n36767 ;
  assign n36756 = x81 | n36215 ;
  assign n36757 = x81 &  n36215 ;
  assign n36758 = ( n36756 & ~n36757 ) | ( n36756 & 1'b0 ) | ( ~n36757 & 1'b0 ) ;
  assign n36770 = ( n36350 & n36402 ) | ( n36350 & n36758 ) | ( n36402 & n36758 ) ;
  assign n36769 = n36350 | n36758 ;
  assign n36771 = ( n36768 & ~n36770 ) | ( n36768 & n36769 ) | ( ~n36770 & n36769 ) ;
  assign n36775 = n36223 &  n36401 ;
  assign n36776 = n36400 &  n36775 ;
  assign n36764 = x80 | n36223 ;
  assign n36765 = x80 &  n36223 ;
  assign n36766 = ( n36764 & ~n36765 ) | ( n36764 & 1'b0 ) | ( ~n36765 & 1'b0 ) ;
  assign n36778 = ( n36349 & n36402 ) | ( n36349 & n36766 ) | ( n36402 & n36766 ) ;
  assign n36777 = n36349 | n36766 ;
  assign n36779 = ( n36776 & ~n36778 ) | ( n36776 & n36777 ) | ( ~n36778 & n36777 ) ;
  assign n36783 = n36231 &  n36401 ;
  assign n36784 = n36400 &  n36783 ;
  assign n36772 = x79 | n36231 ;
  assign n36773 = x79 &  n36231 ;
  assign n36774 = ( n36772 & ~n36773 ) | ( n36772 & 1'b0 ) | ( ~n36773 & 1'b0 ) ;
  assign n36786 = ( n36348 & n36402 ) | ( n36348 & n36774 ) | ( n36402 & n36774 ) ;
  assign n36785 = n36348 | n36774 ;
  assign n36787 = ( n36784 & ~n36786 ) | ( n36784 & n36785 ) | ( ~n36786 & n36785 ) ;
  assign n36791 = n36239 &  n36401 ;
  assign n36792 = n36400 &  n36791 ;
  assign n36780 = x78 | n36239 ;
  assign n36781 = x78 &  n36239 ;
  assign n36782 = ( n36780 & ~n36781 ) | ( n36780 & 1'b0 ) | ( ~n36781 & 1'b0 ) ;
  assign n36794 = ( n36347 & n36402 ) | ( n36347 & n36782 ) | ( n36402 & n36782 ) ;
  assign n36793 = n36347 | n36782 ;
  assign n36795 = ( n36792 & ~n36794 ) | ( n36792 & n36793 ) | ( ~n36794 & n36793 ) ;
  assign n36799 = n36247 &  n36401 ;
  assign n36800 = n36400 &  n36799 ;
  assign n36788 = x77 | n36247 ;
  assign n36789 = x77 &  n36247 ;
  assign n36790 = ( n36788 & ~n36789 ) | ( n36788 & 1'b0 ) | ( ~n36789 & 1'b0 ) ;
  assign n36802 = ( n36346 & n36402 ) | ( n36346 & n36790 ) | ( n36402 & n36790 ) ;
  assign n36801 = n36346 | n36790 ;
  assign n36803 = ( n36800 & ~n36802 ) | ( n36800 & n36801 ) | ( ~n36802 & n36801 ) ;
  assign n36807 = n36255 &  n36401 ;
  assign n36808 = n36400 &  n36807 ;
  assign n36796 = x76 | n36255 ;
  assign n36797 = x76 &  n36255 ;
  assign n36798 = ( n36796 & ~n36797 ) | ( n36796 & 1'b0 ) | ( ~n36797 & 1'b0 ) ;
  assign n36810 = ( n36345 & n36402 ) | ( n36345 & n36798 ) | ( n36402 & n36798 ) ;
  assign n36809 = n36345 | n36798 ;
  assign n36811 = ( n36808 & ~n36810 ) | ( n36808 & n36809 ) | ( ~n36810 & n36809 ) ;
  assign n36815 = n36263 &  n36401 ;
  assign n36816 = n36400 &  n36815 ;
  assign n36804 = x75 | n36263 ;
  assign n36805 = x75 &  n36263 ;
  assign n36806 = ( n36804 & ~n36805 ) | ( n36804 & 1'b0 ) | ( ~n36805 & 1'b0 ) ;
  assign n36818 = ( n36344 & n36402 ) | ( n36344 & n36806 ) | ( n36402 & n36806 ) ;
  assign n36817 = n36344 | n36806 ;
  assign n36819 = ( n36816 & ~n36818 ) | ( n36816 & n36817 ) | ( ~n36818 & n36817 ) ;
  assign n36823 = n36271 &  n36401 ;
  assign n36824 = n36400 &  n36823 ;
  assign n36812 = x74 | n36271 ;
  assign n36813 = x74 &  n36271 ;
  assign n36814 = ( n36812 & ~n36813 ) | ( n36812 & 1'b0 ) | ( ~n36813 & 1'b0 ) ;
  assign n36826 = ( n36343 & n36402 ) | ( n36343 & n36814 ) | ( n36402 & n36814 ) ;
  assign n36825 = n36343 | n36814 ;
  assign n36827 = ( n36824 & ~n36826 ) | ( n36824 & n36825 ) | ( ~n36826 & n36825 ) ;
  assign n36831 = n36279 &  n36401 ;
  assign n36832 = n36400 &  n36831 ;
  assign n36820 = x73 | n36279 ;
  assign n36821 = x73 &  n36279 ;
  assign n36822 = ( n36820 & ~n36821 ) | ( n36820 & 1'b0 ) | ( ~n36821 & 1'b0 ) ;
  assign n36834 = ( n36342 & n36402 ) | ( n36342 & n36822 ) | ( n36402 & n36822 ) ;
  assign n36833 = n36342 | n36822 ;
  assign n36835 = ( n36832 & ~n36834 ) | ( n36832 & n36833 ) | ( ~n36834 & n36833 ) ;
  assign n36839 = n36287 &  n36401 ;
  assign n36840 = n36400 &  n36839 ;
  assign n36828 = x72 | n36287 ;
  assign n36829 = x72 &  n36287 ;
  assign n36830 = ( n36828 & ~n36829 ) | ( n36828 & 1'b0 ) | ( ~n36829 & 1'b0 ) ;
  assign n36842 = ( n36341 & n36402 ) | ( n36341 & n36830 ) | ( n36402 & n36830 ) ;
  assign n36841 = n36341 | n36830 ;
  assign n36843 = ( n36840 & ~n36842 ) | ( n36840 & n36841 ) | ( ~n36842 & n36841 ) ;
  assign n36847 = n36295 &  n36401 ;
  assign n36848 = n36400 &  n36847 ;
  assign n36836 = x71 | n36295 ;
  assign n36837 = x71 &  n36295 ;
  assign n36838 = ( n36836 & ~n36837 ) | ( n36836 & 1'b0 ) | ( ~n36837 & 1'b0 ) ;
  assign n36850 = ( n36340 & n36402 ) | ( n36340 & n36838 ) | ( n36402 & n36838 ) ;
  assign n36849 = n36340 | n36838 ;
  assign n36851 = ( n36848 & ~n36850 ) | ( n36848 & n36849 ) | ( ~n36850 & n36849 ) ;
  assign n36855 = n36303 &  n36401 ;
  assign n36856 = n36400 &  n36855 ;
  assign n36844 = x70 | n36303 ;
  assign n36845 = x70 &  n36303 ;
  assign n36846 = ( n36844 & ~n36845 ) | ( n36844 & 1'b0 ) | ( ~n36845 & 1'b0 ) ;
  assign n36858 = ( n36339 & n36402 ) | ( n36339 & n36846 ) | ( n36402 & n36846 ) ;
  assign n36857 = n36339 | n36846 ;
  assign n36859 = ( n36856 & ~n36858 ) | ( n36856 & n36857 ) | ( ~n36858 & n36857 ) ;
  assign n36863 = n36311 &  n36401 ;
  assign n36864 = n36400 &  n36863 ;
  assign n36852 = x69 | n36311 ;
  assign n36853 = x69 &  n36311 ;
  assign n36854 = ( n36852 & ~n36853 ) | ( n36852 & 1'b0 ) | ( ~n36853 & 1'b0 ) ;
  assign n36866 = ( n36338 & n36402 ) | ( n36338 & n36854 ) | ( n36402 & n36854 ) ;
  assign n36865 = n36338 | n36854 ;
  assign n36867 = ( n36864 & ~n36866 ) | ( n36864 & n36865 ) | ( ~n36866 & n36865 ) ;
  assign n36871 = n36319 &  n36401 ;
  assign n36872 = n36400 &  n36871 ;
  assign n36860 = x68 | n36319 ;
  assign n36861 = x68 &  n36319 ;
  assign n36862 = ( n36860 & ~n36861 ) | ( n36860 & 1'b0 ) | ( ~n36861 & 1'b0 ) ;
  assign n36874 = ( n36337 & n36402 ) | ( n36337 & n36862 ) | ( n36402 & n36862 ) ;
  assign n36873 = n36337 | n36862 ;
  assign n36875 = ( n36872 & ~n36874 ) | ( n36872 & n36873 ) | ( ~n36874 & n36873 ) ;
  assign n36879 = n36324 &  n36401 ;
  assign n36880 = n36400 &  n36879 ;
  assign n36868 = x67 | n36324 ;
  assign n36869 = x67 &  n36324 ;
  assign n36870 = ( n36868 & ~n36869 ) | ( n36868 & 1'b0 ) | ( ~n36869 & 1'b0 ) ;
  assign n36882 = ( n36336 & n36402 ) | ( n36336 & n36870 ) | ( n36402 & n36870 ) ;
  assign n36881 = n36336 | n36870 ;
  assign n36883 = ( n36880 & ~n36882 ) | ( n36880 & n36881 ) | ( ~n36882 & n36881 ) ;
  assign n36884 = n36330 &  n36401 ;
  assign n36885 = n36400 &  n36884 ;
  assign n36876 = x66 | n36330 ;
  assign n36877 = x66 &  n36330 ;
  assign n36878 = ( n36876 & ~n36877 ) | ( n36876 & 1'b0 ) | ( ~n36877 & 1'b0 ) ;
  assign n36886 = n36335 &  n36878 ;
  assign n36887 = ( n36335 & ~n36402 ) | ( n36335 & n36878 ) | ( ~n36402 & n36878 ) ;
  assign n36888 = ( n36885 & ~n36886 ) | ( n36885 & n36887 ) | ( ~n36886 & n36887 ) ;
  assign n36889 = ( x65 & ~n18049 ) | ( x65 & n36334 ) | ( ~n18049 & n36334 ) ;
  assign n36890 = ( n36335 & ~x65 ) | ( n36335 & n36889 ) | ( ~x65 & n36889 ) ;
  assign n36891 = ~n36402 & n36890 ;
  assign n36892 = n36334 &  n36401 ;
  assign n36893 = n36400 &  n36892 ;
  assign n36894 = n36891 | n36893 ;
  assign n36895 = ( x64 & ~n36402 ) | ( x64 & 1'b0 ) | ( ~n36402 & 1'b0 ) ;
  assign n36896 = ( x1 & ~n36895 ) | ( x1 & 1'b0 ) | ( ~n36895 & 1'b0 ) ;
  assign n36897 = ( n18049 & ~n36402 ) | ( n18049 & 1'b0 ) | ( ~n36402 & 1'b0 ) ;
  assign n36898 = n36896 | n36897 ;
  assign n36899 = ( x65 & ~n36898 ) | ( x65 & n18135 ) | ( ~n36898 & n18135 ) ;
  assign n36900 = ( x66 & ~n36894 ) | ( x66 & n36899 ) | ( ~n36894 & n36899 ) ;
  assign n36901 = ( x67 & ~n36888 ) | ( x67 & n36900 ) | ( ~n36888 & n36900 ) ;
  assign n36902 = ( x68 & ~n36883 ) | ( x68 & n36901 ) | ( ~n36883 & n36901 ) ;
  assign n36903 = ( x69 & ~n36875 ) | ( x69 & n36902 ) | ( ~n36875 & n36902 ) ;
  assign n36904 = ( x70 & ~n36867 ) | ( x70 & n36903 ) | ( ~n36867 & n36903 ) ;
  assign n36905 = ( x71 & ~n36859 ) | ( x71 & n36904 ) | ( ~n36859 & n36904 ) ;
  assign n36906 = ( x72 & ~n36851 ) | ( x72 & n36905 ) | ( ~n36851 & n36905 ) ;
  assign n36907 = ( x73 & ~n36843 ) | ( x73 & n36906 ) | ( ~n36843 & n36906 ) ;
  assign n36908 = ( x74 & ~n36835 ) | ( x74 & n36907 ) | ( ~n36835 & n36907 ) ;
  assign n36909 = ( x75 & ~n36827 ) | ( x75 & n36908 ) | ( ~n36827 & n36908 ) ;
  assign n36910 = ( x76 & ~n36819 ) | ( x76 & n36909 ) | ( ~n36819 & n36909 ) ;
  assign n36911 = ( x77 & ~n36811 ) | ( x77 & n36910 ) | ( ~n36811 & n36910 ) ;
  assign n36912 = ( x78 & ~n36803 ) | ( x78 & n36911 ) | ( ~n36803 & n36911 ) ;
  assign n36913 = ( x79 & ~n36795 ) | ( x79 & n36912 ) | ( ~n36795 & n36912 ) ;
  assign n36914 = ( x80 & ~n36787 ) | ( x80 & n36913 ) | ( ~n36787 & n36913 ) ;
  assign n36915 = ( x81 & ~n36779 ) | ( x81 & n36914 ) | ( ~n36779 & n36914 ) ;
  assign n36916 = ( x82 & ~n36771 ) | ( x82 & n36915 ) | ( ~n36771 & n36915 ) ;
  assign n36917 = ( x83 & ~n36763 ) | ( x83 & n36916 ) | ( ~n36763 & n36916 ) ;
  assign n36918 = ( x84 & ~n36755 ) | ( x84 & n36917 ) | ( ~n36755 & n36917 ) ;
  assign n36919 = ( x85 & ~n36747 ) | ( x85 & n36918 ) | ( ~n36747 & n36918 ) ;
  assign n36920 = ( x86 & ~n36739 ) | ( x86 & n36919 ) | ( ~n36739 & n36919 ) ;
  assign n36921 = ( x87 & ~n36731 ) | ( x87 & n36920 ) | ( ~n36731 & n36920 ) ;
  assign n36922 = ( x88 & ~n36723 ) | ( x88 & n36921 ) | ( ~n36723 & n36921 ) ;
  assign n36923 = ( x89 & ~n36715 ) | ( x89 & n36922 ) | ( ~n36715 & n36922 ) ;
  assign n36924 = ( x90 & ~n36707 ) | ( x90 & n36923 ) | ( ~n36707 & n36923 ) ;
  assign n36925 = ( x91 & ~n36699 ) | ( x91 & n36924 ) | ( ~n36699 & n36924 ) ;
  assign n36926 = ( x92 & ~n36691 ) | ( x92 & n36925 ) | ( ~n36691 & n36925 ) ;
  assign n36927 = ( x93 & ~n36683 ) | ( x93 & n36926 ) | ( ~n36683 & n36926 ) ;
  assign n36928 = ( x94 & ~n36675 ) | ( x94 & n36927 ) | ( ~n36675 & n36927 ) ;
  assign n36929 = ( x95 & ~n36667 ) | ( x95 & n36928 ) | ( ~n36667 & n36928 ) ;
  assign n36930 = ( x96 & ~n36659 ) | ( x96 & n36929 ) | ( ~n36659 & n36929 ) ;
  assign n36931 = ( x97 & ~n36651 ) | ( x97 & n36930 ) | ( ~n36651 & n36930 ) ;
  assign n36932 = ( x98 & ~n36643 ) | ( x98 & n36931 ) | ( ~n36643 & n36931 ) ;
  assign n36933 = ( x99 & ~n36635 ) | ( x99 & n36932 ) | ( ~n36635 & n36932 ) ;
  assign n36934 = ( x100 & ~n36627 ) | ( x100 & n36933 ) | ( ~n36627 & n36933 ) ;
  assign n36935 = ( x101 & ~n36619 ) | ( x101 & n36934 ) | ( ~n36619 & n36934 ) ;
  assign n36936 = ( x102 & ~n36611 ) | ( x102 & n36935 ) | ( ~n36611 & n36935 ) ;
  assign n36937 = ( x103 & ~n36603 ) | ( x103 & n36936 ) | ( ~n36603 & n36936 ) ;
  assign n36938 = ( x104 & ~n36595 ) | ( x104 & n36937 ) | ( ~n36595 & n36937 ) ;
  assign n36939 = ( x105 & ~n36587 ) | ( x105 & n36938 ) | ( ~n36587 & n36938 ) ;
  assign n36940 = ( x106 & ~n36579 ) | ( x106 & n36939 ) | ( ~n36579 & n36939 ) ;
  assign n36941 = ( x107 & ~n36571 ) | ( x107 & n36940 ) | ( ~n36571 & n36940 ) ;
  assign n36942 = ( x108 & ~n36563 ) | ( x108 & n36941 ) | ( ~n36563 & n36941 ) ;
  assign n36943 = ( x109 & ~n36555 ) | ( x109 & n36942 ) | ( ~n36555 & n36942 ) ;
  assign n36944 = ( x110 & ~n36547 ) | ( x110 & n36943 ) | ( ~n36547 & n36943 ) ;
  assign n36945 = ( x111 & ~n36539 ) | ( x111 & n36944 ) | ( ~n36539 & n36944 ) ;
  assign n36946 = ( x112 & ~n36531 ) | ( x112 & n36945 ) | ( ~n36531 & n36945 ) ;
  assign n36947 = ( x113 & ~n36523 ) | ( x113 & n36946 ) | ( ~n36523 & n36946 ) ;
  assign n36948 = ( x114 & ~n36515 ) | ( x114 & n36947 ) | ( ~n36515 & n36947 ) ;
  assign n36949 = ( x115 & ~n36507 ) | ( x115 & n36948 ) | ( ~n36507 & n36948 ) ;
  assign n36950 = ( x116 & ~n36499 ) | ( x116 & n36949 ) | ( ~n36499 & n36949 ) ;
  assign n36951 = ( x117 & ~n36491 ) | ( x117 & n36950 ) | ( ~n36491 & n36950 ) ;
  assign n36952 = ( x118 & ~n36483 ) | ( x118 & n36951 ) | ( ~n36483 & n36951 ) ;
  assign n36953 = ( x119 & ~n36475 ) | ( x119 & n36952 ) | ( ~n36475 & n36952 ) ;
  assign n36954 = ( x120 & ~n36467 ) | ( x120 & n36953 ) | ( ~n36467 & n36953 ) ;
  assign n36955 = ( x121 & ~n36459 ) | ( x121 & n36954 ) | ( ~n36459 & n36954 ) ;
  assign n36956 = ( x122 & ~n36451 ) | ( x122 & n36955 ) | ( ~n36451 & n36955 ) ;
  assign n36957 = ( x123 & ~n36443 ) | ( x123 & n36956 ) | ( ~n36443 & n36956 ) ;
  assign n36958 = ( x124 & ~n36435 ) | ( x124 & n36957 ) | ( ~n36435 & n36957 ) ;
  assign n36959 = ( x125 & ~n36427 ) | ( x125 & n36958 ) | ( ~n36427 & n36958 ) ;
  assign n36960 = ( x126 & ~n36419 ) | ( x126 & n36959 ) | ( ~n36419 & n36959 ) ;
  assign n36961 = ( x127 & ~n36411 ) | ( x127 & n36960 ) | ( ~n36411 & n36960 ) ;
  assign n36962 = x64 | n36961 ;
  assign n36963 = ( x0 & ~n36962 ) | ( x0 & n36961 ) | ( ~n36962 & n36961 ) ;
  assign n36964 = ( n18135 & ~n36961 ) | ( n18135 & 1'b0 ) | ( ~n36961 & 1'b0 ) ;
  assign n36965 = n36963 | n36964 ;
  assign n36968 = ~x127 & n36411 ;
  assign n36966 = ( n36411 & ~x127 ) | ( n36411 & n36960 ) | ( ~x127 & n36960 ) ;
  assign n36967 = n36961 | n36966 ;
  assign n36972 = ( n36967 & ~n36898 ) | ( n36967 & n36968 ) | ( ~n36898 & n36968 ) ;
  assign n36969 = ( x65 & ~n18135 ) | ( x65 & n36898 ) | ( ~n18135 & n36898 ) ;
  assign n36970 = ( n36899 & ~x65 ) | ( n36899 & n36969 ) | ( ~x65 & n36969 ) ;
  assign n36971 = ( n36967 & ~n36968 ) | ( n36967 & n36970 ) | ( ~n36968 & n36970 ) ;
  assign n36973 = ( n36968 & ~n36972 ) | ( n36968 & n36971 ) | ( ~n36972 & n36971 ) ;
  assign n36975 = x66 | n36961 ;
  assign n36974 = n36899 | n36961 ;
  assign n36976 = ( n36894 & ~n36975 ) | ( n36894 & n36974 ) | ( ~n36975 & n36974 ) ;
  assign n36977 = ( n36974 & ~n36894 ) | ( n36974 & n36975 ) | ( ~n36894 & n36975 ) ;
  assign n36978 = ( n36976 & ~n36974 ) | ( n36976 & n36977 ) | ( ~n36974 & n36977 ) ;
  assign n36980 = x67 | n36961 ;
  assign n36979 = n36900 | n36961 ;
  assign n36981 = ( n36888 & ~n36980 ) | ( n36888 & n36979 ) | ( ~n36980 & n36979 ) ;
  assign n36982 = ( n36979 & ~n36888 ) | ( n36979 & n36980 ) | ( ~n36888 & n36980 ) ;
  assign n36983 = ( n36981 & ~n36979 ) | ( n36981 & n36982 ) | ( ~n36979 & n36982 ) ;
  assign n36985 = x68 | n36961 ;
  assign n36984 = n36901 | n36961 ;
  assign n36986 = ( n36883 & ~n36985 ) | ( n36883 & n36984 ) | ( ~n36985 & n36984 ) ;
  assign n36987 = ( n36984 & ~n36883 ) | ( n36984 & n36985 ) | ( ~n36883 & n36985 ) ;
  assign n36988 = ( n36986 & ~n36984 ) | ( n36986 & n36987 ) | ( ~n36984 & n36987 ) ;
  assign n36990 = x69 | n36961 ;
  assign n36989 = n36902 | n36961 ;
  assign n36991 = ( n36875 & ~n36990 ) | ( n36875 & n36989 ) | ( ~n36990 & n36989 ) ;
  assign n36992 = ( n36989 & ~n36875 ) | ( n36989 & n36990 ) | ( ~n36875 & n36990 ) ;
  assign n36993 = ( n36991 & ~n36989 ) | ( n36991 & n36992 ) | ( ~n36989 & n36992 ) ;
  assign n36995 = x70 | n36961 ;
  assign n36994 = n36903 | n36961 ;
  assign n36996 = ( n36867 & ~n36995 ) | ( n36867 & n36994 ) | ( ~n36995 & n36994 ) ;
  assign n36997 = ( n36994 & ~n36867 ) | ( n36994 & n36995 ) | ( ~n36867 & n36995 ) ;
  assign n36998 = ( n36996 & ~n36994 ) | ( n36996 & n36997 ) | ( ~n36994 & n36997 ) ;
  assign n37000 = x71 | n36961 ;
  assign n36999 = n36904 | n36961 ;
  assign n37001 = ( n36859 & ~n37000 ) | ( n36859 & n36999 ) | ( ~n37000 & n36999 ) ;
  assign n37002 = ( n36999 & ~n36859 ) | ( n36999 & n37000 ) | ( ~n36859 & n37000 ) ;
  assign n37003 = ( n37001 & ~n36999 ) | ( n37001 & n37002 ) | ( ~n36999 & n37002 ) ;
  assign n37005 = x72 | n36961 ;
  assign n37004 = n36905 | n36961 ;
  assign n37006 = ( n36851 & ~n37005 ) | ( n36851 & n37004 ) | ( ~n37005 & n37004 ) ;
  assign n37007 = ( n37004 & ~n36851 ) | ( n37004 & n37005 ) | ( ~n36851 & n37005 ) ;
  assign n37008 = ( n37006 & ~n37004 ) | ( n37006 & n37007 ) | ( ~n37004 & n37007 ) ;
  assign n37010 = x73 | n36961 ;
  assign n37009 = n36906 | n36961 ;
  assign n37011 = ( n36843 & ~n37010 ) | ( n36843 & n37009 ) | ( ~n37010 & n37009 ) ;
  assign n37012 = ( n37009 & ~n36843 ) | ( n37009 & n37010 ) | ( ~n36843 & n37010 ) ;
  assign n37013 = ( n37011 & ~n37009 ) | ( n37011 & n37012 ) | ( ~n37009 & n37012 ) ;
  assign n37015 = x74 | n36961 ;
  assign n37014 = n36907 | n36961 ;
  assign n37016 = ( n36835 & ~n37015 ) | ( n36835 & n37014 ) | ( ~n37015 & n37014 ) ;
  assign n37017 = ( n37014 & ~n36835 ) | ( n37014 & n37015 ) | ( ~n36835 & n37015 ) ;
  assign n37018 = ( n37016 & ~n37014 ) | ( n37016 & n37017 ) | ( ~n37014 & n37017 ) ;
  assign n37020 = x75 | n36961 ;
  assign n37019 = n36908 | n36961 ;
  assign n37021 = ( n36827 & ~n37020 ) | ( n36827 & n37019 ) | ( ~n37020 & n37019 ) ;
  assign n37022 = ( n37019 & ~n36827 ) | ( n37019 & n37020 ) | ( ~n36827 & n37020 ) ;
  assign n37023 = ( n37021 & ~n37019 ) | ( n37021 & n37022 ) | ( ~n37019 & n37022 ) ;
  assign n37025 = x76 | n36961 ;
  assign n37024 = n36909 | n36961 ;
  assign n37026 = ( n36819 & ~n37025 ) | ( n36819 & n37024 ) | ( ~n37025 & n37024 ) ;
  assign n37027 = ( n37024 & ~n36819 ) | ( n37024 & n37025 ) | ( ~n36819 & n37025 ) ;
  assign n37028 = ( n37026 & ~n37024 ) | ( n37026 & n37027 ) | ( ~n37024 & n37027 ) ;
  assign n37030 = x77 | n36961 ;
  assign n37029 = n36910 | n36961 ;
  assign n37031 = ( n36811 & ~n37030 ) | ( n36811 & n37029 ) | ( ~n37030 & n37029 ) ;
  assign n37032 = ( n37029 & ~n36811 ) | ( n37029 & n37030 ) | ( ~n36811 & n37030 ) ;
  assign n37033 = ( n37031 & ~n37029 ) | ( n37031 & n37032 ) | ( ~n37029 & n37032 ) ;
  assign n37035 = x78 | n36961 ;
  assign n37034 = n36911 | n36961 ;
  assign n37036 = ( n36803 & ~n37035 ) | ( n36803 & n37034 ) | ( ~n37035 & n37034 ) ;
  assign n37037 = ( n37034 & ~n36803 ) | ( n37034 & n37035 ) | ( ~n36803 & n37035 ) ;
  assign n37038 = ( n37036 & ~n37034 ) | ( n37036 & n37037 ) | ( ~n37034 & n37037 ) ;
  assign n37040 = x79 | n36961 ;
  assign n37039 = n36912 | n36961 ;
  assign n37041 = ( n36795 & ~n37040 ) | ( n36795 & n37039 ) | ( ~n37040 & n37039 ) ;
  assign n37042 = ( n37039 & ~n36795 ) | ( n37039 & n37040 ) | ( ~n36795 & n37040 ) ;
  assign n37043 = ( n37041 & ~n37039 ) | ( n37041 & n37042 ) | ( ~n37039 & n37042 ) ;
  assign n37045 = x80 | n36961 ;
  assign n37044 = n36913 | n36961 ;
  assign n37046 = ( n36787 & ~n37045 ) | ( n36787 & n37044 ) | ( ~n37045 & n37044 ) ;
  assign n37047 = ( n37044 & ~n36787 ) | ( n37044 & n37045 ) | ( ~n36787 & n37045 ) ;
  assign n37048 = ( n37046 & ~n37044 ) | ( n37046 & n37047 ) | ( ~n37044 & n37047 ) ;
  assign n37050 = x81 | n36961 ;
  assign n37049 = n36914 | n36961 ;
  assign n37051 = ( n36779 & ~n37050 ) | ( n36779 & n37049 ) | ( ~n37050 & n37049 ) ;
  assign n37052 = ( n37049 & ~n36779 ) | ( n37049 & n37050 ) | ( ~n36779 & n37050 ) ;
  assign n37053 = ( n37051 & ~n37049 ) | ( n37051 & n37052 ) | ( ~n37049 & n37052 ) ;
  assign n37055 = x82 | n36961 ;
  assign n37054 = n36915 | n36961 ;
  assign n37056 = ( n36771 & ~n37055 ) | ( n36771 & n37054 ) | ( ~n37055 & n37054 ) ;
  assign n37057 = ( n37054 & ~n36771 ) | ( n37054 & n37055 ) | ( ~n36771 & n37055 ) ;
  assign n37058 = ( n37056 & ~n37054 ) | ( n37056 & n37057 ) | ( ~n37054 & n37057 ) ;
  assign n37060 = x83 | n36961 ;
  assign n37059 = n36916 | n36961 ;
  assign n37061 = ( n36763 & ~n37060 ) | ( n36763 & n37059 ) | ( ~n37060 & n37059 ) ;
  assign n37062 = ( n37059 & ~n36763 ) | ( n37059 & n37060 ) | ( ~n36763 & n37060 ) ;
  assign n37063 = ( n37061 & ~n37059 ) | ( n37061 & n37062 ) | ( ~n37059 & n37062 ) ;
  assign n37065 = x84 | n36961 ;
  assign n37064 = n36917 | n36961 ;
  assign n37066 = ( n36755 & ~n37065 ) | ( n36755 & n37064 ) | ( ~n37065 & n37064 ) ;
  assign n37067 = ( n37064 & ~n36755 ) | ( n37064 & n37065 ) | ( ~n36755 & n37065 ) ;
  assign n37068 = ( n37066 & ~n37064 ) | ( n37066 & n37067 ) | ( ~n37064 & n37067 ) ;
  assign n37070 = x85 | n36961 ;
  assign n37069 = n36918 | n36961 ;
  assign n37071 = ( n36747 & ~n37070 ) | ( n36747 & n37069 ) | ( ~n37070 & n37069 ) ;
  assign n37072 = ( n37069 & ~n36747 ) | ( n37069 & n37070 ) | ( ~n36747 & n37070 ) ;
  assign n37073 = ( n37071 & ~n37069 ) | ( n37071 & n37072 ) | ( ~n37069 & n37072 ) ;
  assign n37075 = x86 | n36961 ;
  assign n37074 = n36919 | n36961 ;
  assign n37076 = ( n36739 & ~n37075 ) | ( n36739 & n37074 ) | ( ~n37075 & n37074 ) ;
  assign n37077 = ( n37074 & ~n36739 ) | ( n37074 & n37075 ) | ( ~n36739 & n37075 ) ;
  assign n37078 = ( n37076 & ~n37074 ) | ( n37076 & n37077 ) | ( ~n37074 & n37077 ) ;
  assign n37080 = x87 | n36961 ;
  assign n37079 = n36920 | n36961 ;
  assign n37081 = ( n36731 & ~n37080 ) | ( n36731 & n37079 ) | ( ~n37080 & n37079 ) ;
  assign n37082 = ( n37079 & ~n36731 ) | ( n37079 & n37080 ) | ( ~n36731 & n37080 ) ;
  assign n37083 = ( n37081 & ~n37079 ) | ( n37081 & n37082 ) | ( ~n37079 & n37082 ) ;
  assign n37085 = x88 | n36961 ;
  assign n37084 = n36921 | n36961 ;
  assign n37086 = ( n36723 & ~n37085 ) | ( n36723 & n37084 ) | ( ~n37085 & n37084 ) ;
  assign n37087 = ( n37084 & ~n36723 ) | ( n37084 & n37085 ) | ( ~n36723 & n37085 ) ;
  assign n37088 = ( n37086 & ~n37084 ) | ( n37086 & n37087 ) | ( ~n37084 & n37087 ) ;
  assign n37090 = x89 | n36961 ;
  assign n37089 = n36922 | n36961 ;
  assign n37091 = ( n36715 & ~n37090 ) | ( n36715 & n37089 ) | ( ~n37090 & n37089 ) ;
  assign n37092 = ( n37089 & ~n36715 ) | ( n37089 & n37090 ) | ( ~n36715 & n37090 ) ;
  assign n37093 = ( n37091 & ~n37089 ) | ( n37091 & n37092 ) | ( ~n37089 & n37092 ) ;
  assign n37095 = x90 | n36961 ;
  assign n37094 = n36923 | n36961 ;
  assign n37096 = ( n36707 & ~n37095 ) | ( n36707 & n37094 ) | ( ~n37095 & n37094 ) ;
  assign n37097 = ( n37094 & ~n36707 ) | ( n37094 & n37095 ) | ( ~n36707 & n37095 ) ;
  assign n37098 = ( n37096 & ~n37094 ) | ( n37096 & n37097 ) | ( ~n37094 & n37097 ) ;
  assign n37100 = x91 | n36961 ;
  assign n37099 = n36924 | n36961 ;
  assign n37101 = ( n36699 & ~n37100 ) | ( n36699 & n37099 ) | ( ~n37100 & n37099 ) ;
  assign n37102 = ( n37099 & ~n36699 ) | ( n37099 & n37100 ) | ( ~n36699 & n37100 ) ;
  assign n37103 = ( n37101 & ~n37099 ) | ( n37101 & n37102 ) | ( ~n37099 & n37102 ) ;
  assign n37105 = x92 | n36961 ;
  assign n37104 = n36925 | n36961 ;
  assign n37106 = ( n36691 & ~n37105 ) | ( n36691 & n37104 ) | ( ~n37105 & n37104 ) ;
  assign n37107 = ( n37104 & ~n36691 ) | ( n37104 & n37105 ) | ( ~n36691 & n37105 ) ;
  assign n37108 = ( n37106 & ~n37104 ) | ( n37106 & n37107 ) | ( ~n37104 & n37107 ) ;
  assign n37110 = x93 | n36961 ;
  assign n37109 = n36926 | n36961 ;
  assign n37111 = ( n36683 & ~n37110 ) | ( n36683 & n37109 ) | ( ~n37110 & n37109 ) ;
  assign n37112 = ( n37109 & ~n36683 ) | ( n37109 & n37110 ) | ( ~n36683 & n37110 ) ;
  assign n37113 = ( n37111 & ~n37109 ) | ( n37111 & n37112 ) | ( ~n37109 & n37112 ) ;
  assign n37115 = x94 | n36961 ;
  assign n37114 = n36927 | n36961 ;
  assign n37116 = ( n36675 & ~n37115 ) | ( n36675 & n37114 ) | ( ~n37115 & n37114 ) ;
  assign n37117 = ( n37114 & ~n36675 ) | ( n37114 & n37115 ) | ( ~n36675 & n37115 ) ;
  assign n37118 = ( n37116 & ~n37114 ) | ( n37116 & n37117 ) | ( ~n37114 & n37117 ) ;
  assign n37120 = x95 | n36961 ;
  assign n37119 = n36928 | n36961 ;
  assign n37121 = ( n36667 & ~n37120 ) | ( n36667 & n37119 ) | ( ~n37120 & n37119 ) ;
  assign n37122 = ( n37119 & ~n36667 ) | ( n37119 & n37120 ) | ( ~n36667 & n37120 ) ;
  assign n37123 = ( n37121 & ~n37119 ) | ( n37121 & n37122 ) | ( ~n37119 & n37122 ) ;
  assign n37125 = x96 | n36961 ;
  assign n37124 = n36929 | n36961 ;
  assign n37126 = ( n36659 & ~n37125 ) | ( n36659 & n37124 ) | ( ~n37125 & n37124 ) ;
  assign n37127 = ( n37124 & ~n36659 ) | ( n37124 & n37125 ) | ( ~n36659 & n37125 ) ;
  assign n37128 = ( n37126 & ~n37124 ) | ( n37126 & n37127 ) | ( ~n37124 & n37127 ) ;
  assign n37130 = x97 | n36961 ;
  assign n37129 = n36930 | n36961 ;
  assign n37131 = ( n36651 & ~n37130 ) | ( n36651 & n37129 ) | ( ~n37130 & n37129 ) ;
  assign n37132 = ( n37129 & ~n36651 ) | ( n37129 & n37130 ) | ( ~n36651 & n37130 ) ;
  assign n37133 = ( n37131 & ~n37129 ) | ( n37131 & n37132 ) | ( ~n37129 & n37132 ) ;
  assign n37135 = x98 | n36961 ;
  assign n37134 = n36931 | n36961 ;
  assign n37136 = ( n36643 & ~n37135 ) | ( n36643 & n37134 ) | ( ~n37135 & n37134 ) ;
  assign n37137 = ( n37134 & ~n36643 ) | ( n37134 & n37135 ) | ( ~n36643 & n37135 ) ;
  assign n37138 = ( n37136 & ~n37134 ) | ( n37136 & n37137 ) | ( ~n37134 & n37137 ) ;
  assign n37140 = x99 | n36961 ;
  assign n37139 = n36932 | n36961 ;
  assign n37141 = ( n36635 & ~n37140 ) | ( n36635 & n37139 ) | ( ~n37140 & n37139 ) ;
  assign n37142 = ( n37139 & ~n36635 ) | ( n37139 & n37140 ) | ( ~n36635 & n37140 ) ;
  assign n37143 = ( n37141 & ~n37139 ) | ( n37141 & n37142 ) | ( ~n37139 & n37142 ) ;
  assign n37145 = x100 | n36961 ;
  assign n37144 = n36933 | n36961 ;
  assign n37146 = ( n36627 & ~n37145 ) | ( n36627 & n37144 ) | ( ~n37145 & n37144 ) ;
  assign n37147 = ( n37144 & ~n36627 ) | ( n37144 & n37145 ) | ( ~n36627 & n37145 ) ;
  assign n37148 = ( n37146 & ~n37144 ) | ( n37146 & n37147 ) | ( ~n37144 & n37147 ) ;
  assign n37150 = x101 | n36961 ;
  assign n37149 = n36934 | n36961 ;
  assign n37151 = ( n36619 & ~n37150 ) | ( n36619 & n37149 ) | ( ~n37150 & n37149 ) ;
  assign n37152 = ( n37149 & ~n36619 ) | ( n37149 & n37150 ) | ( ~n36619 & n37150 ) ;
  assign n37153 = ( n37151 & ~n37149 ) | ( n37151 & n37152 ) | ( ~n37149 & n37152 ) ;
  assign n37155 = x102 | n36961 ;
  assign n37154 = n36935 | n36961 ;
  assign n37156 = ( n36611 & ~n37155 ) | ( n36611 & n37154 ) | ( ~n37155 & n37154 ) ;
  assign n37157 = ( n37154 & ~n36611 ) | ( n37154 & n37155 ) | ( ~n36611 & n37155 ) ;
  assign n37158 = ( n37156 & ~n37154 ) | ( n37156 & n37157 ) | ( ~n37154 & n37157 ) ;
  assign n37160 = x103 | n36961 ;
  assign n37159 = n36936 | n36961 ;
  assign n37161 = ( n36603 & ~n37160 ) | ( n36603 & n37159 ) | ( ~n37160 & n37159 ) ;
  assign n37162 = ( n37159 & ~n36603 ) | ( n37159 & n37160 ) | ( ~n36603 & n37160 ) ;
  assign n37163 = ( n37161 & ~n37159 ) | ( n37161 & n37162 ) | ( ~n37159 & n37162 ) ;
  assign n37165 = x104 | n36961 ;
  assign n37164 = n36937 | n36961 ;
  assign n37166 = ( n36595 & ~n37165 ) | ( n36595 & n37164 ) | ( ~n37165 & n37164 ) ;
  assign n37167 = ( n37164 & ~n36595 ) | ( n37164 & n37165 ) | ( ~n36595 & n37165 ) ;
  assign n37168 = ( n37166 & ~n37164 ) | ( n37166 & n37167 ) | ( ~n37164 & n37167 ) ;
  assign n37170 = x105 | n36961 ;
  assign n37169 = n36938 | n36961 ;
  assign n37171 = ( n36587 & ~n37170 ) | ( n36587 & n37169 ) | ( ~n37170 & n37169 ) ;
  assign n37172 = ( n37169 & ~n36587 ) | ( n37169 & n37170 ) | ( ~n36587 & n37170 ) ;
  assign n37173 = ( n37171 & ~n37169 ) | ( n37171 & n37172 ) | ( ~n37169 & n37172 ) ;
  assign n37175 = x106 | n36961 ;
  assign n37174 = n36939 | n36961 ;
  assign n37176 = ( n36579 & ~n37175 ) | ( n36579 & n37174 ) | ( ~n37175 & n37174 ) ;
  assign n37177 = ( n37174 & ~n36579 ) | ( n37174 & n37175 ) | ( ~n36579 & n37175 ) ;
  assign n37178 = ( n37176 & ~n37174 ) | ( n37176 & n37177 ) | ( ~n37174 & n37177 ) ;
  assign n37180 = x107 | n36961 ;
  assign n37179 = n36940 | n36961 ;
  assign n37181 = ( n36571 & ~n37180 ) | ( n36571 & n37179 ) | ( ~n37180 & n37179 ) ;
  assign n37182 = ( n37179 & ~n36571 ) | ( n37179 & n37180 ) | ( ~n36571 & n37180 ) ;
  assign n37183 = ( n37181 & ~n37179 ) | ( n37181 & n37182 ) | ( ~n37179 & n37182 ) ;
  assign n37185 = x108 | n36961 ;
  assign n37184 = n36941 | n36961 ;
  assign n37186 = ( n36563 & ~n37185 ) | ( n36563 & n37184 ) | ( ~n37185 & n37184 ) ;
  assign n37187 = ( n37184 & ~n36563 ) | ( n37184 & n37185 ) | ( ~n36563 & n37185 ) ;
  assign n37188 = ( n37186 & ~n37184 ) | ( n37186 & n37187 ) | ( ~n37184 & n37187 ) ;
  assign n37190 = x109 | n36961 ;
  assign n37189 = n36942 | n36961 ;
  assign n37191 = ( n36555 & ~n37190 ) | ( n36555 & n37189 ) | ( ~n37190 & n37189 ) ;
  assign n37192 = ( n37189 & ~n36555 ) | ( n37189 & n37190 ) | ( ~n36555 & n37190 ) ;
  assign n37193 = ( n37191 & ~n37189 ) | ( n37191 & n37192 ) | ( ~n37189 & n37192 ) ;
  assign n37195 = x110 | n36961 ;
  assign n37194 = n36943 | n36961 ;
  assign n37196 = ( n36547 & ~n37195 ) | ( n36547 & n37194 ) | ( ~n37195 & n37194 ) ;
  assign n37197 = ( n37194 & ~n36547 ) | ( n37194 & n37195 ) | ( ~n36547 & n37195 ) ;
  assign n37198 = ( n37196 & ~n37194 ) | ( n37196 & n37197 ) | ( ~n37194 & n37197 ) ;
  assign n37200 = x111 | n36961 ;
  assign n37199 = n36944 | n36961 ;
  assign n37201 = ( n36539 & ~n37200 ) | ( n36539 & n37199 ) | ( ~n37200 & n37199 ) ;
  assign n37202 = ( n37199 & ~n36539 ) | ( n37199 & n37200 ) | ( ~n36539 & n37200 ) ;
  assign n37203 = ( n37201 & ~n37199 ) | ( n37201 & n37202 ) | ( ~n37199 & n37202 ) ;
  assign n37205 = x112 | n36961 ;
  assign n37204 = n36945 | n36961 ;
  assign n37206 = ( n36531 & ~n37205 ) | ( n36531 & n37204 ) | ( ~n37205 & n37204 ) ;
  assign n37207 = ( n37204 & ~n36531 ) | ( n37204 & n37205 ) | ( ~n36531 & n37205 ) ;
  assign n37208 = ( n37206 & ~n37204 ) | ( n37206 & n37207 ) | ( ~n37204 & n37207 ) ;
  assign n37210 = x113 | n36961 ;
  assign n37209 = n36946 | n36961 ;
  assign n37211 = ( n36523 & ~n37210 ) | ( n36523 & n37209 ) | ( ~n37210 & n37209 ) ;
  assign n37212 = ( n37209 & ~n36523 ) | ( n37209 & n37210 ) | ( ~n36523 & n37210 ) ;
  assign n37213 = ( n37211 & ~n37209 ) | ( n37211 & n37212 ) | ( ~n37209 & n37212 ) ;
  assign n37215 = x114 | n36961 ;
  assign n37214 = n36947 | n36961 ;
  assign n37216 = ( n36515 & ~n37215 ) | ( n36515 & n37214 ) | ( ~n37215 & n37214 ) ;
  assign n37217 = ( n37214 & ~n36515 ) | ( n37214 & n37215 ) | ( ~n36515 & n37215 ) ;
  assign n37218 = ( n37216 & ~n37214 ) | ( n37216 & n37217 ) | ( ~n37214 & n37217 ) ;
  assign n37220 = x115 | n36961 ;
  assign n37219 = n36948 | n36961 ;
  assign n37221 = ( n36507 & ~n37220 ) | ( n36507 & n37219 ) | ( ~n37220 & n37219 ) ;
  assign n37222 = ( n37219 & ~n36507 ) | ( n37219 & n37220 ) | ( ~n36507 & n37220 ) ;
  assign n37223 = ( n37221 & ~n37219 ) | ( n37221 & n37222 ) | ( ~n37219 & n37222 ) ;
  assign n37225 = x116 | n36961 ;
  assign n37224 = n36949 | n36961 ;
  assign n37226 = ( n36499 & ~n37225 ) | ( n36499 & n37224 ) | ( ~n37225 & n37224 ) ;
  assign n37227 = ( n37224 & ~n36499 ) | ( n37224 & n37225 ) | ( ~n36499 & n37225 ) ;
  assign n37228 = ( n37226 & ~n37224 ) | ( n37226 & n37227 ) | ( ~n37224 & n37227 ) ;
  assign n37230 = x117 | n36961 ;
  assign n37229 = n36950 | n36961 ;
  assign n37231 = ( n36491 & ~n37230 ) | ( n36491 & n37229 ) | ( ~n37230 & n37229 ) ;
  assign n37232 = ( n37229 & ~n36491 ) | ( n37229 & n37230 ) | ( ~n36491 & n37230 ) ;
  assign n37233 = ( n37231 & ~n37229 ) | ( n37231 & n37232 ) | ( ~n37229 & n37232 ) ;
  assign n37235 = x118 | n36961 ;
  assign n37234 = n36951 | n36961 ;
  assign n37236 = ( n36483 & ~n37235 ) | ( n36483 & n37234 ) | ( ~n37235 & n37234 ) ;
  assign n37237 = ( n37234 & ~n36483 ) | ( n37234 & n37235 ) | ( ~n36483 & n37235 ) ;
  assign n37238 = ( n37236 & ~n37234 ) | ( n37236 & n37237 ) | ( ~n37234 & n37237 ) ;
  assign n37240 = x119 | n36961 ;
  assign n37239 = n36952 | n36961 ;
  assign n37241 = ( n36475 & ~n37240 ) | ( n36475 & n37239 ) | ( ~n37240 & n37239 ) ;
  assign n37242 = ( n37239 & ~n36475 ) | ( n37239 & n37240 ) | ( ~n36475 & n37240 ) ;
  assign n37243 = ( n37241 & ~n37239 ) | ( n37241 & n37242 ) | ( ~n37239 & n37242 ) ;
  assign n37245 = x120 | n36961 ;
  assign n37244 = n36953 | n36961 ;
  assign n37246 = ( n36467 & ~n37245 ) | ( n36467 & n37244 ) | ( ~n37245 & n37244 ) ;
  assign n37247 = ( n37244 & ~n36467 ) | ( n37244 & n37245 ) | ( ~n36467 & n37245 ) ;
  assign n37248 = ( n37246 & ~n37244 ) | ( n37246 & n37247 ) | ( ~n37244 & n37247 ) ;
  assign n37250 = x121 | n36961 ;
  assign n37249 = n36954 | n36961 ;
  assign n37251 = ( n36459 & ~n37250 ) | ( n36459 & n37249 ) | ( ~n37250 & n37249 ) ;
  assign n37252 = ( n37249 & ~n36459 ) | ( n37249 & n37250 ) | ( ~n36459 & n37250 ) ;
  assign n37253 = ( n37251 & ~n37249 ) | ( n37251 & n37252 ) | ( ~n37249 & n37252 ) ;
  assign n37255 = x122 | n36961 ;
  assign n37254 = n36955 | n36961 ;
  assign n37256 = ( n36451 & ~n37255 ) | ( n36451 & n37254 ) | ( ~n37255 & n37254 ) ;
  assign n37257 = ( n37254 & ~n36451 ) | ( n37254 & n37255 ) | ( ~n36451 & n37255 ) ;
  assign n37258 = ( n37256 & ~n37254 ) | ( n37256 & n37257 ) | ( ~n37254 & n37257 ) ;
  assign n37260 = x123 | n36961 ;
  assign n37259 = n36956 | n36961 ;
  assign n37261 = ( n36443 & ~n37260 ) | ( n36443 & n37259 ) | ( ~n37260 & n37259 ) ;
  assign n37262 = ( n37259 & ~n36443 ) | ( n37259 & n37260 ) | ( ~n36443 & n37260 ) ;
  assign n37263 = ( n37261 & ~n37259 ) | ( n37261 & n37262 ) | ( ~n37259 & n37262 ) ;
  assign n37265 = x124 | n36961 ;
  assign n37264 = n36957 | n36961 ;
  assign n37266 = ( n36435 & ~n37265 ) | ( n36435 & n37264 ) | ( ~n37265 & n37264 ) ;
  assign n37267 = ( n37264 & ~n36435 ) | ( n37264 & n37265 ) | ( ~n36435 & n37265 ) ;
  assign n37268 = ( n37266 & ~n37264 ) | ( n37266 & n37267 ) | ( ~n37264 & n37267 ) ;
  assign n37269 = n36958 | n36961 ;
  assign n37270 = x125 | n36961 ;
  assign n37271 = ( n36427 & ~n37269 ) | ( n36427 & n37270 ) | ( ~n37269 & n37270 ) ;
  assign n37272 = ( n37269 & n36427 ) | ( n37269 & n37270 ) | ( n36427 & n37270 ) ;
  assign n37273 = ( n37271 & ~n37272 ) | ( n37271 & n37269 ) | ( ~n37272 & n37269 ) ;
  assign n37274 = n36959 | n36961 ;
  assign n37275 = x126 | n36961 ;
  assign n37276 = ( n36419 & ~n37274 ) | ( n36419 & n37275 ) | ( ~n37274 & n37275 ) ;
  assign n37277 = ( n37274 & n36419 ) | ( n37274 & n37275 ) | ( n36419 & n37275 ) ;
  assign n37278 = ( n37276 & ~n37277 ) | ( n37276 & n37274 ) | ( ~n37277 & n37274 ) ;
  assign n37279 = ( x127 & ~n36960 ) | ( x127 & n36411 ) | ( ~n36960 & n36411 ) ;
  assign n37280 = n36966 &  n37279 ;
  assign y0 = ~n19024 ;
  assign y1 = ~n18125 ;
  assign y2 = ~n17572 ;
  assign y3 = ~n17022 ;
  assign y4 = ~n16481 ;
  assign y5 = ~n15949 ;
  assign y6 = ~n15416 ;
  assign y7 = ~n14914 ;
  assign y8 = ~n14409 ;
  assign y9 = ~n13899 ;
  assign y10 = ~n13422 ;
  assign y11 = ~n12945 ;
  assign y12 = ~n12465 ;
  assign y13 = ~n12017 ;
  assign y14 = ~n11566 ;
  assign y15 = ~n11114 ;
  assign y16 = ~n10694 ;
  assign y17 = ~n10270 ;
  assign y18 = ~n9842 ;
  assign y19 = ~n9446 ;
  assign y20 = ~n9050 ;
  assign y21 = ~n8651 ;
  assign y22 = ~n8282 ;
  assign y23 = ~n7899 ;
  assign y24 = ~n7536 ;
  assign y25 = ~n7195 ;
  assign y26 = ~n6836 ;
  assign y27 = ~n6499 ;
  assign y28 = ~n6187 ;
  assign y29 = ~n5855 ;
  assign y30 = ~n5542 ;
  assign y31 = ~n5254 ;
  assign y32 = ~n4951 ;
  assign y33 = ~n4669 ;
  assign y34 = ~n4407 ;
  assign y35 = ~n4130 ;
  assign y36 = ~n3874 ;
  assign y37 = ~n3640 ;
  assign y38 = ~n3389 ;
  assign y39 = ~n3157 ;
  assign y40 = ~n2947 ;
  assign y41 = ~n2742 ;
  assign y42 = ~n2518 ;
  assign y43 = ~n2331 ;
  assign y44 = ~n2140 ;
  assign y45 = ~n1964 ;
  assign y46 = ~n1809 ;
  assign y47 = ~n1639 ;
  assign y48 = ~n1495 ;
  assign y49 = ~n1371 ;
  assign y50 = ~n1228 ;
  assign y51 = ~n1105 ;
  assign y52 = ~n1006 ;
  assign y53 = ~n892 ;
  assign y54 = ~n795 ;
  assign y55 = ~n722 ;
  assign y56 = ~n634 ;
  assign y57 = ~n564 ;
  assign y58 = ~n513 ;
  assign y59 = ~n435 ;
  assign y60 = ~n362 ;
  assign y61 = ~n346 ;
  assign y62 = ~n19027 ;
  assign y63 = ~n19032 ;
  assign y64 = n36965 ;
  assign y65 = n36973 ;
  assign y66 = n36978 ;
  assign y67 = n36983 ;
  assign y68 = n36988 ;
  assign y69 = n36993 ;
  assign y70 = n36998 ;
  assign y71 = n37003 ;
  assign y72 = n37008 ;
  assign y73 = n37013 ;
  assign y74 = n37018 ;
  assign y75 = n37023 ;
  assign y76 = n37028 ;
  assign y77 = n37033 ;
  assign y78 = n37038 ;
  assign y79 = n37043 ;
  assign y80 = n37048 ;
  assign y81 = n37053 ;
  assign y82 = n37058 ;
  assign y83 = n37063 ;
  assign y84 = n37068 ;
  assign y85 = n37073 ;
  assign y86 = n37078 ;
  assign y87 = n37083 ;
  assign y88 = n37088 ;
  assign y89 = n37093 ;
  assign y90 = n37098 ;
  assign y91 = n37103 ;
  assign y92 = n37108 ;
  assign y93 = n37113 ;
  assign y94 = n37118 ;
  assign y95 = n37123 ;
  assign y96 = n37128 ;
  assign y97 = n37133 ;
  assign y98 = n37138 ;
  assign y99 = n37143 ;
  assign y100 = n37148 ;
  assign y101 = n37153 ;
  assign y102 = n37158 ;
  assign y103 = n37163 ;
  assign y104 = n37168 ;
  assign y105 = n37173 ;
  assign y106 = n37178 ;
  assign y107 = n37183 ;
  assign y108 = n37188 ;
  assign y109 = n37193 ;
  assign y110 = n37198 ;
  assign y111 = n37203 ;
  assign y112 = n37208 ;
  assign y113 = n37213 ;
  assign y114 = n37218 ;
  assign y115 = n37223 ;
  assign y116 = n37228 ;
  assign y117 = n37233 ;
  assign y118 = n37238 ;
  assign y119 = n37243 ;
  assign y120 = n37248 ;
  assign y121 = n37253 ;
  assign y122 = n37258 ;
  assign y123 = n37263 ;
  assign y124 = n37268 ;
  assign y125 = n37273 ;
  assign y126 = n37278 ;
  assign y127 = n37280 ;
endmodule
