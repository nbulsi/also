module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 ;
  assign n133 = x126 | x127 ;
  assign n397 = x110 | x111 ;
  assign n135 = x126 &  x127 ;
  assign n129 = x124 | x125 ;
  assign n149 = ~x126 & n129 ;
  assign n150 = n135 | n149 ;
  assign n134 = x122 | x123 ;
  assign n130 = ( x126 & ~n129 ) | ( x126 & x127 ) | ( ~n129 & x127 ) ;
  assign n131 = ( x127 & ~x126 ) | ( x127 & n129 ) | ( ~x126 & n129 ) ;
  assign n132 = n130 &  n131 ;
  assign n136 = ( x124 & ~x126 ) | ( x124 & n135 ) | ( ~x126 & n135 ) ;
  assign n137 = ~x124 & n134 ;
  assign n138 = ( x124 & ~n136 ) | ( x124 & n137 ) | ( ~n136 & n137 ) ;
  assign n139 = ( x125 & ~x126 ) | ( x125 & x127 ) | ( ~x126 & x127 ) ;
  assign n140 = x124 | n139 ;
  assign n141 = x125 &  x127 ;
  assign n142 = ( x124 & ~n141 ) | ( x124 & x127 ) | ( ~n141 & x127 ) ;
  assign n143 = ( x125 & ~n140 ) | ( x125 & n142 ) | ( ~n140 & n142 ) ;
  assign n144 = ( n138 & ~n133 ) | ( n138 & n143 ) | ( ~n133 & n143 ) ;
  assign n145 = ~n132 &  ~n144 ;
  assign n148 = n134 | n145 ;
  assign n151 = ~n132 & n150 ;
  assign n152 = ~n144 & n151 ;
  assign n153 = n148 | n152 ;
  assign n154 = ( x124 & ~n153 ) | ( x124 & n152 ) | ( ~n153 & n152 ) ;
  assign n157 = x120 | x121 ;
  assign n158 = x122 | n157 ;
  assign n159 = ( x122 & ~n145 ) | ( x122 & 1'b0 ) | ( ~n145 & 1'b0 ) ;
  assign n160 = ( n150 & ~n158 ) | ( n150 & n159 ) | ( ~n158 & n159 ) ;
  assign n162 = ~x122 & n157 ;
  assign n163 = ( x122 & ~n150 ) | ( x122 & n162 ) | ( ~n150 & n162 ) ;
  assign n164 = ( x123 & ~n163 ) | ( x123 & n145 ) | ( ~n163 & n145 ) ;
  assign n161 = ( x122 & x123 ) | ( x122 & n145 ) | ( x123 & n145 ) ;
  assign n165 = ( x122 & ~x123 ) | ( x122 & 1'b0 ) | ( ~x123 & 1'b0 ) ;
  assign n166 = ( n164 & ~n161 ) | ( n164 & n165 ) | ( ~n161 & n165 ) ;
  assign n167 = n160 | n166 ;
  assign n170 = ( n138 & ~n143 ) | ( n138 & 1'b0 ) | ( ~n143 & 1'b0 ) ;
  assign n168 = ( n132 & n138 ) | ( n132 & n143 ) | ( n138 & n143 ) ;
  assign n169 = ( n132 & ~n168 ) | ( n132 & 1'b0 ) | ( ~n168 & 1'b0 ) ;
  assign n171 = ( n138 & ~n170 ) | ( n138 & n169 ) | ( ~n170 & n169 ) ;
  assign n172 = ( n167 & ~n171 ) | ( n167 & 1'b0 ) | ( ~n171 & 1'b0 ) ;
  assign n155 = x124 | n152 ;
  assign n156 = ( n148 & ~n155 ) | ( n148 & 1'b0 ) | ( ~n155 & 1'b0 ) ;
  assign n173 = ~n154 & n156 ;
  assign n174 = ( n154 & n172 ) | ( n154 & n173 ) | ( n172 & n173 ) ;
  assign n175 = n133 | n174 ;
  assign n176 = n154 | n156 ;
  assign n177 = n167 | n176 ;
  assign n178 = ~n143 & n168 ;
  assign n179 = ( n143 & ~n144 ) | ( n143 & n178 ) | ( ~n144 & n178 ) ;
  assign n180 = ( n177 & ~n179 ) | ( n177 & 1'b0 ) | ( ~n179 & 1'b0 ) ;
  assign n181 = ~n175 | ~n180 ;
  assign n184 = ( x120 & ~n181 ) | ( x120 & x121 ) | ( ~n181 & x121 ) ;
  assign n189 = ( x120 & ~x121 ) | ( x120 & 1'b0 ) | ( ~x121 & 1'b0 ) ;
  assign n146 = x118 | x119 ;
  assign n185 = ~x120 & n146 ;
  assign n186 = ( x120 & ~n132 ) | ( x120 & n185 ) | ( ~n132 & n185 ) ;
  assign n187 = ~n144 & n186 ;
  assign n188 = ( n181 & ~x121 ) | ( n181 & n187 ) | ( ~x121 & n187 ) ;
  assign n190 = ( n184 & ~n189 ) | ( n184 & n188 ) | ( ~n189 & n188 ) ;
  assign n182 = x120 &  n181 ;
  assign n147 = x120 | n146 ;
  assign n183 = ( n145 & ~n182 ) | ( n145 & n147 ) | ( ~n182 & n147 ) ;
  assign n222 = ~n183 & n190 ;
  assign n223 = ( n150 & ~n190 ) | ( n150 & n222 ) | ( ~n190 & n222 ) ;
  assign n191 = n183 &  n190 ;
  assign n192 = n145 | n179 ;
  assign n193 = ( n177 & ~n192 ) | ( n177 & 1'b0 ) | ( ~n192 & 1'b0 ) ;
  assign n194 = ~n133 & n174 ;
  assign n195 = ( n133 & n193 ) | ( n133 & n194 ) | ( n193 & n194 ) ;
  assign n196 = ( n157 & n181 ) | ( n157 & n195 ) | ( n181 & n195 ) ;
  assign n197 = ( n181 & ~n196 ) | ( n181 & 1'b0 ) | ( ~n196 & 1'b0 ) ;
  assign n198 = ( n195 & ~x122 ) | ( n195 & n197 ) | ( ~x122 & n197 ) ;
  assign n199 = ( x122 & ~n195 ) | ( x122 & n197 ) | ( ~n195 & n197 ) ;
  assign n200 = ( n198 & ~n197 ) | ( n198 & n199 ) | ( ~n197 & n199 ) ;
  assign n201 = ( n191 & ~n150 ) | ( n191 & n200 ) | ( ~n150 & n200 ) ;
  assign n202 = x122 | n145 ;
  assign n203 = x123 | n202 ;
  assign n204 = x123 &  n202 ;
  assign n205 = ( n203 & ~n204 ) | ( n203 & 1'b0 ) | ( ~n204 & 1'b0 ) ;
  assign n206 = ( x122 & ~n163 ) | ( x122 & n145 ) | ( ~n163 & n145 ) ;
  assign n207 = ( x122 & ~n206 ) | ( x122 & 1'b0 ) | ( ~n206 & 1'b0 ) ;
  assign n208 = ( n160 & ~n207 ) | ( n160 & n163 ) | ( ~n207 & n163 ) ;
  assign n209 = ( n181 & ~n208 ) | ( n181 & n205 ) | ( ~n208 & n205 ) ;
  assign n210 = ~n205 & n209 ;
  assign n211 = ( n181 & ~n208 ) | ( n181 & 1'b0 ) | ( ~n208 & 1'b0 ) ;
  assign n212 = ( n205 & ~n211 ) | ( n205 & 1'b0 ) | ( ~n211 & 1'b0 ) ;
  assign n213 = n210 | n212 ;
  assign n214 = n167 &  n176 ;
  assign n215 = ~n181 & n214 ;
  assign n216 = ( n177 & ~n214 ) | ( n177 & n215 ) | ( ~n214 & n215 ) ;
  assign n217 = n213 &  n216 ;
  assign n218 = n201 &  n217 ;
  assign n219 = ( n133 & ~n218 ) | ( n133 & n217 ) | ( ~n218 & n217 ) ;
  assign n224 = n213 | n223 ;
  assign n220 = ~n150 & n183 ;
  assign n221 = n190 &  n220 ;
  assign n225 = ~n200 & n221 ;
  assign n226 = ( n200 & ~n224 ) | ( n200 & n225 ) | ( ~n224 & n225 ) ;
  assign n228 = ( n133 & n167 ) | ( n133 & n176 ) | ( n167 & n176 ) ;
  assign n227 = ( n167 & ~n179 ) | ( n167 & n176 ) | ( ~n179 & n176 ) ;
  assign n229 = ( n176 & ~n227 ) | ( n176 & 1'b0 ) | ( ~n227 & 1'b0 ) ;
  assign n230 = ( n228 & ~n176 ) | ( n228 & n229 ) | ( ~n176 & n229 ) ;
  assign n231 = ~n132 & n143 ;
  assign n232 = ~n144 & n231 ;
  assign n233 = ( n156 & ~n154 ) | ( n156 & n232 ) | ( ~n154 & n232 ) ;
  assign n234 = n154 | n233 ;
  assign n235 = ( n177 & n179 ) | ( n177 & n234 ) | ( n179 & n234 ) ;
  assign n236 = ( n177 & ~n235 ) | ( n177 & 1'b0 ) | ( ~n235 & 1'b0 ) ;
  assign n237 = n175 &  n236 ;
  assign n238 = n230 | n237 ;
  assign n239 = n226 | n238 ;
  assign n240 = ~n219 |  n239 ;
  assign n283 = ( n200 & ~n221 ) | ( n200 & 1'b0 ) | ( ~n221 & 1'b0 ) ;
  assign n284 = ( n223 & n240 ) | ( n223 & n283 ) | ( n240 & n283 ) ;
  assign n285 = ~n223 & n284 ;
  assign n286 = n221 | n223 ;
  assign n287 = n240 | n286 ;
  assign n288 = ( n200 & ~n286 ) | ( n200 & n287 ) | ( ~n286 & n287 ) ;
  assign n289 = ~n285 & n288 ;
  assign n290 = ~n201 & n213 ;
  assign n291 = ~n240 & n290 ;
  assign n292 = ( n226 & ~n291 ) | ( n226 & n290 ) | ( ~n291 & n290 ) ;
  assign n293 = n289 | n292 ;
  assign n243 = x116 | x117 ;
  assign n244 = x118 | n243 ;
  assign n245 = x118 &  n240 ;
  assign n246 = ( n181 & ~n244 ) | ( n181 & n245 ) | ( ~n244 & n245 ) ;
  assign n247 = ( x118 & ~n240 ) | ( x118 & x119 ) | ( ~n240 & x119 ) ;
  assign n254 = ( x118 & ~x119 ) | ( x118 & 1'b0 ) | ( ~x119 & 1'b0 ) ;
  assign n248 = ~x118 & n243 ;
  assign n249 = ( x118 & ~n232 ) | ( x118 & n248 ) | ( ~n232 & n248 ) ;
  assign n250 = ( n177 & ~n249 ) | ( n177 & n179 ) | ( ~n249 & n179 ) ;
  assign n251 = ( n177 & ~n250 ) | ( n177 & 1'b0 ) | ( ~n250 & 1'b0 ) ;
  assign n252 = n175 &  n251 ;
  assign n253 = ( n240 & ~x119 ) | ( n240 & n252 ) | ( ~x119 & n252 ) ;
  assign n255 = ( n247 & ~n254 ) | ( n247 & n253 ) | ( ~n254 & n253 ) ;
  assign n256 = n246 &  n255 ;
  assign n257 = ( n145 & ~n256 ) | ( n145 & n255 ) | ( ~n256 & n255 ) ;
  assign n258 = ( n145 & ~n246 ) | ( n145 & 1'b0 ) | ( ~n246 & 1'b0 ) ;
  assign n259 = n255 &  n258 ;
  assign n261 = ( n181 & ~n237 ) | ( n181 & 1'b0 ) | ( ~n237 & 1'b0 ) ;
  assign n262 = ( n226 & ~n230 ) | ( n226 & n261 ) | ( ~n230 & n261 ) ;
  assign n263 = ~n226 & n262 ;
  assign n264 = n219 &  n263 ;
  assign n260 = ~n146 & n240 ;
  assign n265 = ( n260 & ~n264 ) | ( n260 & 1'b0 ) | ( ~n264 & 1'b0 ) ;
  assign n266 = ( x120 & n264 ) | ( x120 & n265 ) | ( n264 & n265 ) ;
  assign n267 = x120 | n264 ;
  assign n268 = n260 | n267 ;
  assign n269 = ~n266 & n268 ;
  assign n270 = n259 | n269 ;
  assign n271 = n257 &  n270 ;
  assign n272 = ~x120 & n181 ;
  assign n273 = ~x121 & n272 ;
  assign n274 = ( x121 & ~n272 ) | ( x121 & 1'b0 ) | ( ~n272 & 1'b0 ) ;
  assign n275 = n273 | n274 ;
  assign n277 = ( n183 & ~n240 ) | ( n183 & 1'b0 ) | ( ~n240 & 1'b0 ) ;
  assign n276 = ~n182 & n187 ;
  assign n278 = ( n183 & n275 ) | ( n183 & n276 ) | ( n275 & n276 ) ;
  assign n279 = ( n277 & ~n276 ) | ( n277 & n278 ) | ( ~n276 & n278 ) ;
  assign n280 = ( n183 & ~n278 ) | ( n183 & n277 ) | ( ~n278 & n277 ) ;
  assign n281 = ( n275 & ~n279 ) | ( n275 & n280 ) | ( ~n279 & n280 ) ;
  assign n282 = ( n271 & ~n150 ) | ( n271 & n281 ) | ( ~n150 & n281 ) ;
  assign n294 = ~n293 & n282 ;
  assign n295 = ( n294 & ~n133 ) | ( n294 & n293 ) | ( ~n133 & n293 ) ;
  assign n298 = ~n246 & n255 ;
  assign n299 = ( n145 & n269 ) | ( n145 & n298 ) | ( n269 & n298 ) ;
  assign n300 = ( n150 & ~n299 ) | ( n150 & 1'b0 ) | ( ~n299 & 1'b0 ) ;
  assign n301 = ( n289 & ~n300 ) | ( n289 & 1'b0 ) | ( ~n300 & 1'b0 ) ;
  assign n296 = ~n150 & n257 ;
  assign n297 = n270 &  n296 ;
  assign n302 = ~n281 & n297 ;
  assign n303 = ( n281 & n301 ) | ( n281 & n302 ) | ( n301 & n302 ) ;
  assign n305 = ( n133 & ~n226 ) | ( n133 & 1'b0 ) | ( ~n226 & 1'b0 ) ;
  assign n304 = n201 &  n240 ;
  assign n306 = n213 &  n304 ;
  assign n307 = ( n305 & ~n213 ) | ( n305 & n306 ) | ( ~n213 & n306 ) ;
  assign n308 = n210 | n237 ;
  assign n309 = ( n230 & ~n212 ) | ( n230 & n308 ) | ( ~n212 & n308 ) ;
  assign n310 = n212 | n309 ;
  assign n311 = ( n219 & n226 ) | ( n219 & n310 ) | ( n226 & n310 ) ;
  assign n312 = ( n219 & ~n311 ) | ( n219 & 1'b0 ) | ( ~n311 & 1'b0 ) ;
  assign n328 = ( n240 & ~n312 ) | ( n240 & 1'b0 ) | ( ~n312 & 1'b0 ) ;
  assign n329 = ( n303 & ~n307 ) | ( n303 & n328 ) | ( ~n307 & n328 ) ;
  assign n330 = ~n303 & n329 ;
  assign n331 = ~n295 & n330 ;
  assign n313 = n307 | n312 ;
  assign n314 = n303 | n313 ;
  assign n315 = n295 | n314 ;
  assign n327 = ~n243 & n315 ;
  assign n332 = ~n331 & n327 ;
  assign n333 = ( x118 & n332 ) | ( x118 & n331 ) | ( n332 & n331 ) ;
  assign n334 = x118 | n331 ;
  assign n335 = n327 | n334 ;
  assign n336 = ~n333 & n335 ;
  assign n318 = ( x116 & ~n315 ) | ( x116 & x117 ) | ( ~n315 & x117 ) ;
  assign n324 = ( x116 & ~x117 ) | ( x116 & 1'b0 ) | ( ~x117 & 1'b0 ) ;
  assign n241 = x114 | x115 ;
  assign n319 = ~x116 & n241 ;
  assign n320 = ( x116 & ~n238 ) | ( x116 & n319 ) | ( ~n238 & n319 ) ;
  assign n321 = ( n219 & ~n320 ) | ( n219 & n226 ) | ( ~n320 & n226 ) ;
  assign n322 = ( n219 & ~n321 ) | ( n219 & 1'b0 ) | ( ~n321 & 1'b0 ) ;
  assign n323 = ( n315 & ~x117 ) | ( n315 & n322 ) | ( ~x117 & n322 ) ;
  assign n325 = ( n318 & ~n324 ) | ( n318 & n323 ) | ( ~n324 & n323 ) ;
  assign n242 = x116 | n241 ;
  assign n316 = x116 &  n315 ;
  assign n317 = ( n240 & ~n242 ) | ( n240 & n316 ) | ( ~n242 & n316 ) ;
  assign n349 = n181 | n317 ;
  assign n350 = ( n325 & ~n349 ) | ( n325 & 1'b0 ) | ( ~n349 & 1'b0 ) ;
  assign n364 = ( n281 & ~n300 ) | ( n281 & 1'b0 ) | ( ~n300 & 1'b0 ) ;
  assign n365 = ( n297 & n315 ) | ( n297 & n364 ) | ( n315 & n364 ) ;
  assign n366 = ~n297 & n365 ;
  assign n367 = n297 | n300 ;
  assign n368 = n315 | n367 ;
  assign n369 = ( n281 & ~n367 ) | ( n281 & n368 ) | ( ~n367 & n368 ) ;
  assign n370 = ~n366 & n369 ;
  assign n371 = n282 | n289 ;
  assign n372 = n315 | n371 ;
  assign n373 = ( n303 & ~n371 ) | ( n303 & n372 ) | ( ~n371 & n372 ) ;
  assign n374 = n370 | n373 ;
  assign n326 = ~n317 & n325 ;
  assign n337 = ( n326 & ~n181 ) | ( n326 & n336 ) | ( ~n181 & n336 ) ;
  assign n338 = n145 | n337 ;
  assign n342 = ~x118 & n240 ;
  assign n343 = ( x119 & ~n342 ) | ( x119 & 1'b0 ) | ( ~n342 & 1'b0 ) ;
  assign n344 = n260 | n343 ;
  assign n339 = ( n240 & ~x118 ) | ( n240 & n252 ) | ( ~x118 & n252 ) ;
  assign n340 = x118 &  n339 ;
  assign n341 = ( n246 & ~n340 ) | ( n246 & n252 ) | ( ~n340 & n252 ) ;
  assign n345 = ( n315 & ~n344 ) | ( n315 & n341 ) | ( ~n344 & n341 ) ;
  assign n347 = ( n315 & ~n345 ) | ( n315 & 1'b0 ) | ( ~n345 & 1'b0 ) ;
  assign n346 = ~n341 & n345 ;
  assign n348 = ( n344 & ~n347 ) | ( n344 & n346 ) | ( ~n347 & n346 ) ;
  assign n351 = n336 | n350 ;
  assign n352 = n317 &  n325 ;
  assign n353 = ( n181 & ~n325 ) | ( n181 & n352 ) | ( ~n325 & n352 ) ;
  assign n354 = ( n145 & ~n353 ) | ( n145 & 1'b0 ) | ( ~n353 & 1'b0 ) ;
  assign n355 = n351 &  n354 ;
  assign n356 = n348 | n355 ;
  assign n357 = n338 &  n356 ;
  assign n358 = n257 | n259 ;
  assign n359 = ( n259 & n269 ) | ( n259 & n358 ) | ( n269 & n358 ) ;
  assign n361 = ( n315 & ~n358 ) | ( n315 & n359 ) | ( ~n358 & n359 ) ;
  assign n360 = ( n259 & ~n359 ) | ( n259 & n315 ) | ( ~n359 & n315 ) ;
  assign n362 = ( n269 & ~n361 ) | ( n269 & n360 ) | ( ~n361 & n360 ) ;
  assign n363 = ( n357 & ~n150 ) | ( n357 & n362 ) | ( ~n150 & n362 ) ;
  assign n375 = ~n374 & n363 ;
  assign n376 = ( n375 & ~n133 ) | ( n375 & n374 ) | ( ~n133 & n374 ) ;
  assign n379 = ( n351 & ~n353 ) | ( n351 & 1'b0 ) | ( ~n353 & 1'b0 ) ;
  assign n380 = ( n145 & n348 ) | ( n145 & n379 ) | ( n348 & n379 ) ;
  assign n381 = ( n150 & ~n380 ) | ( n150 & 1'b0 ) | ( ~n380 & 1'b0 ) ;
  assign n382 = ( n370 & ~n381 ) | ( n370 & 1'b0 ) | ( ~n381 & 1'b0 ) ;
  assign n377 = ~n150 & n338 ;
  assign n378 = n356 &  n377 ;
  assign n383 = ~n362 & n378 ;
  assign n384 = ( n362 & n382 ) | ( n362 & n383 ) | ( n382 & n383 ) ;
  assign n386 = ( n282 & ~n133 ) | ( n282 & n289 ) | ( ~n133 & n289 ) ;
  assign n385 = ( n282 & n289 ) | ( n282 & n315 ) | ( n289 & n315 ) ;
  assign n387 = ~n289 & n385 ;
  assign n388 = ( n289 & ~n386 ) | ( n289 & n387 ) | ( ~n386 & n387 ) ;
  assign n389 = n285 | n312 ;
  assign n390 = ( n288 & n307 ) | ( n288 & n389 ) | ( n307 & n389 ) ;
  assign n391 = ( n288 & ~n390 ) | ( n288 & 1'b0 ) | ( ~n390 & 1'b0 ) ;
  assign n392 = ( n295 & ~n303 ) | ( n295 & n391 ) | ( ~n303 & n391 ) ;
  assign n393 = ~n295 & n392 ;
  assign n394 = n388 | n393 ;
  assign n395 = n384 | n394 ;
  assign n396 = n376 | n395 ;
  assign n439 = ~n350 & n353 ;
  assign n440 = ( n336 & ~n350 ) | ( n336 & n439 ) | ( ~n350 & n439 ) ;
  assign n442 = ( n350 & n396 ) | ( n350 & n440 ) | ( n396 & n440 ) ;
  assign n441 = ( n396 & ~n440 ) | ( n396 & n439 ) | ( ~n440 & n439 ) ;
  assign n443 = ( n336 & ~n442 ) | ( n336 & n441 ) | ( ~n442 & n441 ) ;
  assign n430 = ~x116 & n315 ;
  assign n431 = ( x117 & ~n430 ) | ( x117 & 1'b0 ) | ( ~n430 & 1'b0 ) ;
  assign n432 = n327 | n431 ;
  assign n427 = ( n315 & ~x116 ) | ( n315 & n322 ) | ( ~x116 & n322 ) ;
  assign n428 = x116 &  n427 ;
  assign n429 = ( n317 & ~n428 ) | ( n317 & n322 ) | ( ~n428 & n322 ) ;
  assign n433 = ( n396 & ~n432 ) | ( n396 & n429 ) | ( ~n432 & n429 ) ;
  assign n435 = ( n396 & ~n433 ) | ( n396 & 1'b0 ) | ( ~n433 & 1'b0 ) ;
  assign n434 = ~n429 & n433 ;
  assign n436 = ( n432 & ~n435 ) | ( n432 & n434 ) | ( ~n435 & n434 ) ;
  assign n403 = ( x114 & ~n396 ) | ( x114 & x115 ) | ( ~n396 & x115 ) ;
  assign n409 = ( x114 & ~x115 ) | ( x114 & 1'b0 ) | ( ~x115 & 1'b0 ) ;
  assign n399 = x112 | x113 ;
  assign n404 = ~x114 & n399 ;
  assign n405 = ( x114 & ~n313 ) | ( x114 & n404 ) | ( ~n313 & n404 ) ;
  assign n406 = ( n295 & ~n303 ) | ( n295 & n405 ) | ( ~n303 & n405 ) ;
  assign n407 = ~n295 & n406 ;
  assign n408 = ( n396 & ~x115 ) | ( n396 & n407 ) | ( ~x115 & n407 ) ;
  assign n410 = ( n403 & ~n409 ) | ( n403 & n408 ) | ( ~n409 & n408 ) ;
  assign n400 = x114 | n399 ;
  assign n401 = x114 &  n396 ;
  assign n402 = ( n315 & ~n400 ) | ( n315 & n401 ) | ( ~n400 & n401 ) ;
  assign n413 = n240 | n402 ;
  assign n414 = ( n410 & ~n413 ) | ( n410 & 1'b0 ) | ( ~n413 & 1'b0 ) ;
  assign n416 = ( n315 & ~n393 ) | ( n315 & 1'b0 ) | ( ~n393 & 1'b0 ) ;
  assign n417 = ( n384 & ~n388 ) | ( n384 & n416 ) | ( ~n388 & n416 ) ;
  assign n418 = ~n384 & n417 ;
  assign n419 = ~n376 & n418 ;
  assign n415 = ~n241 & n396 ;
  assign n420 = ( n415 & ~n419 ) | ( n415 & 1'b0 ) | ( ~n419 & 1'b0 ) ;
  assign n421 = ( x116 & n419 ) | ( x116 & n420 ) | ( n419 & n420 ) ;
  assign n422 = x116 | n419 ;
  assign n423 = n415 | n422 ;
  assign n424 = ~n421 & n423 ;
  assign n425 = n414 | n424 ;
  assign n411 = n402 &  n410 ;
  assign n412 = ( n240 & ~n410 ) | ( n240 & n411 ) | ( ~n410 & n411 ) ;
  assign n444 = n181 | n412 ;
  assign n445 = ( n425 & ~n444 ) | ( n425 & 1'b0 ) | ( ~n444 & 1'b0 ) ;
  assign n446 = n436 | n445 ;
  assign n447 = ~n402 & n410 ;
  assign n448 = ( n424 & ~n240 ) | ( n424 & n447 ) | ( ~n240 & n447 ) ;
  assign n449 = ( n181 & ~n448 ) | ( n181 & 1'b0 ) | ( ~n448 & 1'b0 ) ;
  assign n450 = ( n145 & ~n449 ) | ( n145 & 1'b0 ) | ( ~n449 & 1'b0 ) ;
  assign n451 = n446 &  n450 ;
  assign n452 = n443 | n451 ;
  assign n426 = ~n412 & n425 ;
  assign n437 = ( n426 & ~n181 ) | ( n426 & n436 ) | ( ~n181 & n436 ) ;
  assign n438 = n145 | n437 ;
  assign n473 = ~n150 & n438 ;
  assign n474 = n452 &  n473 ;
  assign n460 = ( n362 & ~n378 ) | ( n362 & 1'b0 ) | ( ~n378 & 1'b0 ) ;
  assign n461 = ( n381 & n396 ) | ( n381 & n460 ) | ( n396 & n460 ) ;
  assign n462 = ~n381 & n461 ;
  assign n463 = n378 | n381 ;
  assign n464 = n396 | n463 ;
  assign n465 = ( n362 & ~n463 ) | ( n362 & n464 ) | ( ~n463 & n464 ) ;
  assign n466 = ~n462 & n465 ;
  assign n467 = n363 | n370 ;
  assign n468 = n396 | n467 ;
  assign n469 = ( n384 & ~n467 ) | ( n384 & n468 ) | ( ~n467 & n468 ) ;
  assign n470 = n466 | n469 ;
  assign n453 = n438 &  n452 ;
  assign n455 = ( n338 & ~n348 ) | ( n338 & n355 ) | ( ~n348 & n355 ) ;
  assign n454 = ( n338 & ~n396 ) | ( n338 & 1'b0 ) | ( ~n396 & 1'b0 ) ;
  assign n457 = ( n338 & ~n455 ) | ( n338 & n454 ) | ( ~n455 & n454 ) ;
  assign n456 = ( n454 & ~n355 ) | ( n454 & n455 ) | ( ~n355 & n455 ) ;
  assign n458 = ( n348 & ~n457 ) | ( n348 & n456 ) | ( ~n457 & n456 ) ;
  assign n459 = ( n453 & ~n150 ) | ( n453 & n458 ) | ( ~n150 & n458 ) ;
  assign n471 = ~n470 & n459 ;
  assign n472 = ( n471 & ~n133 ) | ( n471 & n470 ) | ( ~n133 & n470 ) ;
  assign n475 = ( n446 & ~n449 ) | ( n446 & 1'b0 ) | ( ~n449 & 1'b0 ) ;
  assign n476 = ( n145 & n443 ) | ( n145 & n475 ) | ( n443 & n475 ) ;
  assign n477 = ( n150 & ~n476 ) | ( n150 & 1'b0 ) | ( ~n476 & 1'b0 ) ;
  assign n478 = ( n466 & ~n477 ) | ( n466 & 1'b0 ) | ( ~n477 & 1'b0 ) ;
  assign n479 = ~n458 & n474 ;
  assign n480 = ( n458 & n478 ) | ( n458 & n479 ) | ( n478 & n479 ) ;
  assign n482 = ( n363 & ~n133 ) | ( n363 & n370 ) | ( ~n133 & n370 ) ;
  assign n481 = ( n363 & n370 ) | ( n363 & n396 ) | ( n370 & n396 ) ;
  assign n483 = ~n370 & n481 ;
  assign n484 = ( n370 & ~n482 ) | ( n370 & n483 ) | ( ~n482 & n483 ) ;
  assign n485 = n366 | n393 ;
  assign n486 = ( n369 & n388 ) | ( n369 & n485 ) | ( n388 & n485 ) ;
  assign n487 = ( n369 & ~n486 ) | ( n369 & 1'b0 ) | ( ~n486 & 1'b0 ) ;
  assign n488 = ( n376 & ~n384 ) | ( n376 & n487 ) | ( ~n384 & n487 ) ;
  assign n489 = ~n376 & n488 ;
  assign n490 = n484 | n489 ;
  assign n491 = n480 | n490 ;
  assign n492 = n472 | n491 ;
  assign n563 = ( n458 & ~n477 ) | ( n458 & 1'b0 ) | ( ~n477 & 1'b0 ) ;
  assign n564 = ( n474 & n492 ) | ( n474 & n563 ) | ( n492 & n563 ) ;
  assign n565 = ~n474 & n564 ;
  assign n566 = n474 | n477 ;
  assign n567 = n492 | n566 ;
  assign n568 = ( n458 & ~n566 ) | ( n458 & n567 ) | ( ~n566 & n567 ) ;
  assign n569 = ~n565 & n568 ;
  assign n570 = n459 | n466 ;
  assign n571 = n492 | n570 ;
  assign n572 = ( n480 & ~n570 ) | ( n480 & n571 ) | ( ~n570 & n571 ) ;
  assign n573 = n569 | n572 ;
  assign n398 = x112 | n397 ;
  assign n493 = x112 &  n492 ;
  assign n494 = ( n396 & ~n398 ) | ( n396 & n493 ) | ( ~n398 & n493 ) ;
  assign n495 = ( x112 & ~n492 ) | ( x112 & x113 ) | ( ~n492 & x113 ) ;
  assign n501 = ( x112 & ~x113 ) | ( x112 & 1'b0 ) | ( ~x113 & 1'b0 ) ;
  assign n496 = ~x112 & n397 ;
  assign n497 = ( x112 & ~n394 ) | ( x112 & n496 ) | ( ~n394 & n496 ) ;
  assign n498 = ( n376 & ~n384 ) | ( n376 & n497 ) | ( ~n384 & n497 ) ;
  assign n499 = ~n376 & n498 ;
  assign n500 = ( n492 & ~x113 ) | ( n492 & n499 ) | ( ~x113 & n499 ) ;
  assign n502 = ( n495 & ~n501 ) | ( n495 & n500 ) | ( ~n501 & n500 ) ;
  assign n503 = ~n494 & n502 ;
  assign n505 = ( n396 & ~n489 ) | ( n396 & 1'b0 ) | ( ~n489 & 1'b0 ) ;
  assign n506 = ( n480 & ~n484 ) | ( n480 & n505 ) | ( ~n484 & n505 ) ;
  assign n507 = ~n480 & n506 ;
  assign n508 = ~n472 & n507 ;
  assign n504 = ~n399 & n492 ;
  assign n509 = ( n504 & ~n508 ) | ( n504 & 1'b0 ) | ( ~n508 & 1'b0 ) ;
  assign n510 = ( x114 & n508 ) | ( x114 & n509 ) | ( n508 & n509 ) ;
  assign n511 = x114 | n508 ;
  assign n512 = n504 | n511 ;
  assign n513 = ~n510 & n512 ;
  assign n514 = ( n503 & ~n315 ) | ( n503 & n513 ) | ( ~n315 & n513 ) ;
  assign n515 = ( n240 & ~n514 ) | ( n240 & 1'b0 ) | ( ~n514 & 1'b0 ) ;
  assign n519 = ~x114 & n396 ;
  assign n520 = ( x115 & ~n519 ) | ( x115 & 1'b0 ) | ( ~n519 & 1'b0 ) ;
  assign n521 = n415 | n520 ;
  assign n516 = ( n396 & ~x114 ) | ( n396 & n407 ) | ( ~x114 & n407 ) ;
  assign n517 = x114 &  n516 ;
  assign n518 = ( n402 & ~n517 ) | ( n402 & n407 ) | ( ~n517 & n407 ) ;
  assign n522 = ( n492 & ~n521 ) | ( n492 & n518 ) | ( ~n521 & n518 ) ;
  assign n524 = ( n492 & ~n522 ) | ( n492 & 1'b0 ) | ( ~n522 & 1'b0 ) ;
  assign n523 = ~n518 & n522 ;
  assign n525 = ( n521 & ~n524 ) | ( n521 & n523 ) | ( ~n524 & n523 ) ;
  assign n526 = n315 | n494 ;
  assign n527 = ( n502 & ~n526 ) | ( n502 & 1'b0 ) | ( ~n526 & 1'b0 ) ;
  assign n528 = n513 | n527 ;
  assign n529 = n494 &  n502 ;
  assign n530 = ( n315 & ~n502 ) | ( n315 & n529 ) | ( ~n502 & n529 ) ;
  assign n531 = n240 | n530 ;
  assign n532 = ( n528 & ~n531 ) | ( n528 & 1'b0 ) | ( ~n531 & 1'b0 ) ;
  assign n533 = n525 | n532 ;
  assign n534 = ~n515 & n533 ;
  assign n535 = ( n412 & ~n414 ) | ( n412 & 1'b0 ) | ( ~n414 & 1'b0 ) ;
  assign n536 = ( n414 & ~n535 ) | ( n414 & n424 ) | ( ~n535 & n424 ) ;
  assign n538 = ( n492 & n535 ) | ( n492 & n536 ) | ( n535 & n536 ) ;
  assign n537 = ( n414 & ~n536 ) | ( n414 & n492 ) | ( ~n536 & n492 ) ;
  assign n539 = ( n424 & ~n538 ) | ( n424 & n537 ) | ( ~n538 & n537 ) ;
  assign n540 = ( n534 & ~n181 ) | ( n534 & n539 ) | ( ~n181 & n539 ) ;
  assign n541 = n145 | n540 ;
  assign n542 = n449 | n492 ;
  assign n543 = ( n436 & ~n445 ) | ( n436 & n449 ) | ( ~n445 & n449 ) ;
  assign n544 = ( n445 & n542 ) | ( n445 & n543 ) | ( n542 & n543 ) ;
  assign n545 = ( n449 & ~n543 ) | ( n449 & n542 ) | ( ~n543 & n542 ) ;
  assign n546 = ( n436 & ~n544 ) | ( n436 & n545 ) | ( ~n544 & n545 ) ;
  assign n547 = n181 | n515 ;
  assign n548 = ( n533 & ~n547 ) | ( n533 & 1'b0 ) | ( ~n547 & 1'b0 ) ;
  assign n549 = n539 | n548 ;
  assign n550 = ( n528 & ~n530 ) | ( n528 & 1'b0 ) | ( ~n530 & 1'b0 ) ;
  assign n551 = ( n525 & ~n240 ) | ( n525 & n550 ) | ( ~n240 & n550 ) ;
  assign n552 = ( n181 & ~n551 ) | ( n181 & 1'b0 ) | ( ~n551 & 1'b0 ) ;
  assign n553 = ( n145 & ~n552 ) | ( n145 & 1'b0 ) | ( ~n552 & 1'b0 ) ;
  assign n554 = n549 &  n553 ;
  assign n555 = n546 | n554 ;
  assign n556 = n541 &  n555 ;
  assign n557 = n451 &  n492 ;
  assign n558 = ( n438 & ~n492 ) | ( n438 & n557 ) | ( ~n492 & n557 ) ;
  assign n559 = ( n438 & ~n558 ) | ( n438 & n443 ) | ( ~n558 & n443 ) ;
  assign n560 = ( n443 & ~n438 ) | ( n443 & n558 ) | ( ~n438 & n558 ) ;
  assign n561 = ( n559 & ~n443 ) | ( n559 & n560 ) | ( ~n443 & n560 ) ;
  assign n562 = ( n556 & ~n150 ) | ( n556 & n561 ) | ( ~n150 & n561 ) ;
  assign n574 = ~n573 & n562 ;
  assign n575 = ( n574 & ~n133 ) | ( n574 & n573 ) | ( ~n133 & n573 ) ;
  assign n578 = ( n549 & ~n552 ) | ( n549 & 1'b0 ) | ( ~n552 & 1'b0 ) ;
  assign n579 = ( n145 & n546 ) | ( n145 & n578 ) | ( n546 & n578 ) ;
  assign n580 = ( n150 & ~n579 ) | ( n150 & 1'b0 ) | ( ~n579 & 1'b0 ) ;
  assign n581 = ( n569 & ~n580 ) | ( n569 & 1'b0 ) | ( ~n580 & 1'b0 ) ;
  assign n576 = ~n150 & n541 ;
  assign n577 = n555 &  n576 ;
  assign n582 = ~n561 & n577 ;
  assign n583 = ( n561 & n581 ) | ( n561 & n582 ) | ( n581 & n582 ) ;
  assign n585 = ( n459 & ~n133 ) | ( n459 & n466 ) | ( ~n133 & n466 ) ;
  assign n584 = ( n459 & n466 ) | ( n459 & n492 ) | ( n466 & n492 ) ;
  assign n586 = ~n466 & n584 ;
  assign n587 = ( n466 & ~n585 ) | ( n466 & n586 ) | ( ~n585 & n586 ) ;
  assign n588 = n462 | n489 ;
  assign n589 = ( n465 & n484 ) | ( n465 & n588 ) | ( n484 & n588 ) ;
  assign n590 = ( n465 & ~n589 ) | ( n465 & 1'b0 ) | ( ~n589 & 1'b0 ) ;
  assign n591 = ( n472 & ~n480 ) | ( n472 & n590 ) | ( ~n480 & n590 ) ;
  assign n592 = ~n472 & n591 ;
  assign n593 = n587 | n592 ;
  assign n594 = n583 | n593 ;
  assign n595 = n575 | n594 ;
  assign n614 = ~n397 & n595 ;
  assign n740 = ~x110 & n595 ;
  assign n741 = ( x111 & ~n740 ) | ( x111 & 1'b0 ) | ( ~n740 & 1'b0 ) ;
  assign n742 = n614 | n741 ;
  assign n681 = ( n561 & ~n577 ) | ( n561 & 1'b0 ) | ( ~n577 & 1'b0 ) ;
  assign n682 = ( n580 & n595 ) | ( n580 & n681 ) | ( n595 & n681 ) ;
  assign n683 = ~n580 & n682 ;
  assign n684 = n577 | n580 ;
  assign n685 = n595 | n684 ;
  assign n686 = ( n561 & ~n684 ) | ( n561 & n685 ) | ( ~n684 & n685 ) ;
  assign n687 = ~n683 & n686 ;
  assign n688 = n562 | n569 ;
  assign n689 = n595 | n688 ;
  assign n690 = ( n583 & ~n688 ) | ( n583 & n689 ) | ( ~n688 & n689 ) ;
  assign n691 = n687 | n690 ;
  assign n602 = ( x110 & ~n595 ) | ( x110 & x111 ) | ( ~n595 & x111 ) ;
  assign n608 = ( x110 & ~x111 ) | ( x110 & 1'b0 ) | ( ~x111 & 1'b0 ) ;
  assign n598 = x108 | x109 ;
  assign n603 = ~x110 & n598 ;
  assign n604 = ( x110 & ~n490 ) | ( x110 & n603 ) | ( ~n490 & n603 ) ;
  assign n605 = ( n472 & ~n480 ) | ( n472 & n604 ) | ( ~n480 & n604 ) ;
  assign n606 = ~n472 & n605 ;
  assign n607 = ( n595 & ~x111 ) | ( n595 & n606 ) | ( ~x111 & n606 ) ;
  assign n609 = ( n602 & ~n608 ) | ( n602 & n607 ) | ( ~n608 & n607 ) ;
  assign n599 = x110 | n598 ;
  assign n600 = x110 &  n595 ;
  assign n601 = ( n492 & ~n599 ) | ( n492 & n600 ) | ( ~n599 & n600 ) ;
  assign n610 = n601 &  n609 ;
  assign n611 = ( n396 & ~n609 ) | ( n396 & n610 ) | ( ~n609 & n610 ) ;
  assign n612 = n396 | n601 ;
  assign n613 = ( n609 & ~n612 ) | ( n609 & 1'b0 ) | ( ~n612 & 1'b0 ) ;
  assign n615 = ( n492 & ~n592 ) | ( n492 & 1'b0 ) | ( ~n592 & 1'b0 ) ;
  assign n616 = ( n583 & ~n587 ) | ( n583 & n615 ) | ( ~n587 & n615 ) ;
  assign n617 = ~n583 & n616 ;
  assign n618 = ~n575 & n617 ;
  assign n619 = ~n618 & n614 ;
  assign n620 = ( x112 & n619 ) | ( x112 & n618 ) | ( n619 & n618 ) ;
  assign n621 = x112 | n618 ;
  assign n622 = n614 | n621 ;
  assign n623 = ~n620 & n622 ;
  assign n624 = n613 | n623 ;
  assign n625 = ~n611 & n624 ;
  assign n626 = ~x112 & n492 ;
  assign n627 = ~x113 & n626 ;
  assign n628 = ( x113 & ~n626 ) | ( x113 & 1'b0 ) | ( ~n626 & 1'b0 ) ;
  assign n629 = n627 | n628 ;
  assign n630 = ~n493 & n499 ;
  assign n631 = n494 | n595 ;
  assign n632 = ( n494 & ~n630 ) | ( n494 & n629 ) | ( ~n630 & n629 ) ;
  assign n633 = ( n630 & n631 ) | ( n630 & n632 ) | ( n631 & n632 ) ;
  assign n634 = ( n494 & ~n632 ) | ( n494 & n631 ) | ( ~n632 & n631 ) ;
  assign n635 = ( n629 & ~n633 ) | ( n629 & n634 ) | ( ~n633 & n634 ) ;
  assign n636 = ( n625 & ~n315 ) | ( n625 & n635 ) | ( ~n315 & n635 ) ;
  assign n637 = ( n240 & ~n636 ) | ( n240 & 1'b0 ) | ( ~n636 & 1'b0 ) ;
  assign n638 = ~n527 & n530 ;
  assign n639 = ( n527 & ~n638 ) | ( n527 & n513 ) | ( ~n638 & n513 ) ;
  assign n640 = ( n595 & n639 ) | ( n595 & n638 ) | ( n639 & n638 ) ;
  assign n641 = ( n595 & ~n639 ) | ( n595 & n527 ) | ( ~n639 & n527 ) ;
  assign n642 = ( n513 & ~n640 ) | ( n513 & n641 ) | ( ~n640 & n641 ) ;
  assign n643 = n315 | n611 ;
  assign n644 = ( n624 & ~n643 ) | ( n624 & 1'b0 ) | ( ~n643 & 1'b0 ) ;
  assign n645 = n635 | n644 ;
  assign n646 = ~n601 & n609 ;
  assign n647 = ( n623 & ~n396 ) | ( n623 & n646 ) | ( ~n396 & n646 ) ;
  assign n648 = ( n315 & ~n647 ) | ( n315 & 1'b0 ) | ( ~n647 & 1'b0 ) ;
  assign n649 = n240 | n648 ;
  assign n650 = ( n645 & ~n649 ) | ( n645 & 1'b0 ) | ( ~n649 & 1'b0 ) ;
  assign n651 = n642 | n650 ;
  assign n652 = ~n637 & n651 ;
  assign n653 = n515 | n595 ;
  assign n654 = ( n515 & ~n532 ) | ( n515 & n525 ) | ( ~n532 & n525 ) ;
  assign n655 = ( n532 & n653 ) | ( n532 & n654 ) | ( n653 & n654 ) ;
  assign n656 = ( n515 & ~n654 ) | ( n515 & n653 ) | ( ~n654 & n653 ) ;
  assign n657 = ( n525 & ~n655 ) | ( n525 & n656 ) | ( ~n655 & n656 ) ;
  assign n658 = ( n652 & ~n181 ) | ( n652 & n657 ) | ( ~n181 & n657 ) ;
  assign n659 = n145 | n658 ;
  assign n660 = n552 | n595 ;
  assign n661 = ( n539 & ~n552 ) | ( n539 & n548 ) | ( ~n552 & n548 ) ;
  assign n663 = ( n552 & n660 ) | ( n552 & n661 ) | ( n660 & n661 ) ;
  assign n662 = ( n548 & ~n661 ) | ( n548 & n660 ) | ( ~n661 & n660 ) ;
  assign n664 = ( n539 & ~n663 ) | ( n539 & n662 ) | ( ~n663 & n662 ) ;
  assign n665 = n181 | n637 ;
  assign n666 = ( n651 & ~n665 ) | ( n651 & 1'b0 ) | ( ~n665 & 1'b0 ) ;
  assign n667 = n657 | n666 ;
  assign n668 = ( n645 & ~n648 ) | ( n645 & 1'b0 ) | ( ~n648 & 1'b0 ) ;
  assign n669 = ( n642 & ~n240 ) | ( n642 & n668 ) | ( ~n240 & n668 ) ;
  assign n670 = ( n181 & ~n669 ) | ( n181 & 1'b0 ) | ( ~n669 & 1'b0 ) ;
  assign n671 = ( n145 & ~n670 ) | ( n145 & 1'b0 ) | ( ~n670 & 1'b0 ) ;
  assign n672 = n667 &  n671 ;
  assign n673 = n664 | n672 ;
  assign n674 = n659 &  n673 ;
  assign n676 = ( n541 & ~n546 ) | ( n541 & n554 ) | ( ~n546 & n554 ) ;
  assign n675 = ( n541 & ~n595 ) | ( n541 & 1'b0 ) | ( ~n595 & 1'b0 ) ;
  assign n678 = ( n541 & ~n676 ) | ( n541 & n675 ) | ( ~n676 & n675 ) ;
  assign n677 = ( n675 & ~n554 ) | ( n675 & n676 ) | ( ~n554 & n676 ) ;
  assign n679 = ( n546 & ~n678 ) | ( n546 & n677 ) | ( ~n678 & n677 ) ;
  assign n680 = ( n674 & ~n150 ) | ( n674 & n679 ) | ( ~n150 & n679 ) ;
  assign n692 = ~n691 & n680 ;
  assign n693 = ( n692 & ~n133 ) | ( n692 & n691 ) | ( ~n133 & n691 ) ;
  assign n696 = ( n667 & ~n670 ) | ( n667 & 1'b0 ) | ( ~n670 & 1'b0 ) ;
  assign n697 = ( n145 & n664 ) | ( n145 & n696 ) | ( n664 & n696 ) ;
  assign n698 = ( n150 & ~n697 ) | ( n150 & 1'b0 ) | ( ~n697 & 1'b0 ) ;
  assign n699 = ( n687 & ~n698 ) | ( n687 & 1'b0 ) | ( ~n698 & 1'b0 ) ;
  assign n694 = ~n150 & n659 ;
  assign n695 = n673 &  n694 ;
  assign n700 = ~n679 & n695 ;
  assign n701 = ( n679 & n699 ) | ( n679 & n700 ) | ( n699 & n700 ) ;
  assign n703 = ( n562 & ~n133 ) | ( n562 & n569 ) | ( ~n133 & n569 ) ;
  assign n702 = ( n562 & n569 ) | ( n562 & n595 ) | ( n569 & n595 ) ;
  assign n704 = ~n569 & n702 ;
  assign n705 = ( n569 & ~n703 ) | ( n569 & n704 ) | ( ~n703 & n704 ) ;
  assign n706 = n565 | n592 ;
  assign n707 = ( n568 & n587 ) | ( n568 & n706 ) | ( n587 & n706 ) ;
  assign n708 = ( n568 & ~n707 ) | ( n568 & 1'b0 ) | ( ~n707 & 1'b0 ) ;
  assign n709 = ( n575 & ~n583 ) | ( n575 & n708 ) | ( ~n583 & n708 ) ;
  assign n710 = ~n575 & n709 ;
  assign n711 = n705 | n710 ;
  assign n712 = n701 | n711 ;
  assign n713 = n693 | n712 ;
  assign n737 = ( n595 & ~x110 ) | ( n595 & n606 ) | ( ~x110 & n606 ) ;
  assign n738 = x110 &  n737 ;
  assign n739 = ( n601 & ~n738 ) | ( n601 & n606 ) | ( ~n738 & n606 ) ;
  assign n743 = ( n713 & ~n742 ) | ( n713 & n739 ) | ( ~n742 & n739 ) ;
  assign n745 = ( n713 & ~n743 ) | ( n713 & 1'b0 ) | ( ~n743 & 1'b0 ) ;
  assign n744 = ~n739 & n743 ;
  assign n746 = ( n742 & ~n745 ) | ( n742 & n744 ) | ( ~n745 & n744 ) ;
  assign n726 = ( n595 & ~n710 ) | ( n595 & 1'b0 ) | ( ~n710 & 1'b0 ) ;
  assign n727 = ( n701 & ~n705 ) | ( n701 & n726 ) | ( ~n705 & n726 ) ;
  assign n728 = ~n701 & n727 ;
  assign n729 = ~n693 & n728 ;
  assign n725 = ~n598 & n713 ;
  assign n730 = ~n729 & n725 ;
  assign n731 = ( x110 & n730 ) | ( x110 & n729 ) | ( n730 & n729 ) ;
  assign n732 = x110 | n729 ;
  assign n733 = n725 | n732 ;
  assign n734 = ~n731 & n733 ;
  assign n716 = ( x108 & ~n713 ) | ( x108 & x109 ) | ( ~n713 & x109 ) ;
  assign n722 = ( x108 & ~x109 ) | ( x108 & 1'b0 ) | ( ~x109 & 1'b0 ) ;
  assign n596 = x106 | x107 ;
  assign n717 = ~x108 & n596 ;
  assign n718 = ( x108 & ~n593 ) | ( x108 & n717 ) | ( ~n593 & n717 ) ;
  assign n719 = ( n575 & ~n583 ) | ( n575 & n718 ) | ( ~n583 & n718 ) ;
  assign n720 = ~n575 & n719 ;
  assign n721 = ( n713 & ~x109 ) | ( n713 & n720 ) | ( ~x109 & n720 ) ;
  assign n723 = ( n716 & ~n722 ) | ( n716 & n721 ) | ( ~n722 & n721 ) ;
  assign n597 = x108 | n596 ;
  assign n714 = x108 &  n713 ;
  assign n715 = ( n595 & ~n597 ) | ( n595 & n714 ) | ( ~n597 & n714 ) ;
  assign n747 = n492 | n715 ;
  assign n748 = ( n723 & ~n747 ) | ( n723 & 1'b0 ) | ( ~n747 & 1'b0 ) ;
  assign n749 = n734 | n748 ;
  assign n750 = n715 &  n723 ;
  assign n751 = ( n492 & ~n723 ) | ( n492 & n750 ) | ( ~n723 & n750 ) ;
  assign n752 = n396 | n751 ;
  assign n753 = ( n749 & ~n752 ) | ( n749 & 1'b0 ) | ( ~n752 & 1'b0 ) ;
  assign n724 = ~n715 & n723 ;
  assign n735 = ( n724 & ~n492 ) | ( n724 & n734 ) | ( ~n492 & n734 ) ;
  assign n736 = ( n396 & ~n735 ) | ( n396 & 1'b0 ) | ( ~n735 & 1'b0 ) ;
  assign n805 = ( n679 & ~n698 ) | ( n679 & 1'b0 ) | ( ~n698 & 1'b0 ) ;
  assign n806 = ( n695 & n713 ) | ( n695 & n805 ) | ( n713 & n805 ) ;
  assign n807 = ~n695 & n806 ;
  assign n808 = n695 | n698 ;
  assign n809 = n713 | n808 ;
  assign n810 = ( n679 & ~n808 ) | ( n679 & n809 ) | ( ~n808 & n809 ) ;
  assign n811 = ~n807 & n810 ;
  assign n812 = n680 | n687 ;
  assign n813 = n713 | n812 ;
  assign n814 = ( n701 & ~n812 ) | ( n701 & n813 ) | ( ~n812 & n813 ) ;
  assign n815 = n811 | n814 ;
  assign n754 = n746 | n753 ;
  assign n755 = ~n736 & n754 ;
  assign n756 = ( n611 & ~n613 ) | ( n611 & 1'b0 ) | ( ~n613 & 1'b0 ) ;
  assign n757 = ( n613 & ~n756 ) | ( n613 & n623 ) | ( ~n756 & n623 ) ;
  assign n759 = ( n713 & n756 ) | ( n713 & n757 ) | ( n756 & n757 ) ;
  assign n758 = ( n613 & ~n757 ) | ( n613 & n713 ) | ( ~n757 & n713 ) ;
  assign n760 = ( n623 & ~n759 ) | ( n623 & n758 ) | ( ~n759 & n758 ) ;
  assign n761 = ( n755 & ~n315 ) | ( n755 & n760 ) | ( ~n315 & n760 ) ;
  assign n762 = ( n240 & ~n761 ) | ( n240 & 1'b0 ) | ( ~n761 & 1'b0 ) ;
  assign n763 = n315 | n736 ;
  assign n764 = ( n754 & ~n763 ) | ( n754 & 1'b0 ) | ( ~n763 & 1'b0 ) ;
  assign n765 = n760 | n764 ;
  assign n766 = ( n749 & ~n751 ) | ( n749 & 1'b0 ) | ( ~n751 & 1'b0 ) ;
  assign n767 = ( n746 & ~n396 ) | ( n746 & n766 ) | ( ~n396 & n766 ) ;
  assign n768 = ( n315 & ~n767 ) | ( n315 & 1'b0 ) | ( ~n767 & 1'b0 ) ;
  assign n769 = n240 | n768 ;
  assign n770 = ( n765 & ~n769 ) | ( n765 & 1'b0 ) | ( ~n769 & 1'b0 ) ;
  assign n771 = ( n635 & ~n648 ) | ( n635 & n644 ) | ( ~n648 & n644 ) ;
  assign n772 = ( n648 & n713 ) | ( n648 & n771 ) | ( n713 & n771 ) ;
  assign n773 = ( n644 & ~n771 ) | ( n644 & n713 ) | ( ~n771 & n713 ) ;
  assign n774 = ( n635 & ~n772 ) | ( n635 & n773 ) | ( ~n772 & n773 ) ;
  assign n775 = n770 | n774 ;
  assign n776 = ~n762 & n775 ;
  assign n777 = n650 &  n713 ;
  assign n778 = ( n637 & ~n777 ) | ( n637 & n713 ) | ( ~n777 & n713 ) ;
  assign n779 = ( n642 & ~n637 ) | ( n642 & n778 ) | ( ~n637 & n778 ) ;
  assign n780 = ( n637 & ~n778 ) | ( n637 & n642 ) | ( ~n778 & n642 ) ;
  assign n781 = ( n779 & ~n642 ) | ( n779 & n780 ) | ( ~n642 & n780 ) ;
  assign n782 = ( n776 & ~n181 ) | ( n776 & n781 ) | ( ~n181 & n781 ) ;
  assign n783 = n145 | n782 ;
  assign n784 = n670 | n713 ;
  assign n785 = ( n657 & ~n670 ) | ( n657 & n666 ) | ( ~n670 & n666 ) ;
  assign n787 = ( n670 & n784 ) | ( n670 & n785 ) | ( n784 & n785 ) ;
  assign n786 = ( n666 & ~n785 ) | ( n666 & n784 ) | ( ~n785 & n784 ) ;
  assign n788 = ( n657 & ~n787 ) | ( n657 & n786 ) | ( ~n787 & n786 ) ;
  assign n789 = n181 | n762 ;
  assign n790 = ( n775 & ~n789 ) | ( n775 & 1'b0 ) | ( ~n789 & 1'b0 ) ;
  assign n791 = n781 | n790 ;
  assign n792 = ( n765 & ~n768 ) | ( n765 & 1'b0 ) | ( ~n768 & 1'b0 ) ;
  assign n793 = ( n774 & ~n240 ) | ( n774 & n792 ) | ( ~n240 & n792 ) ;
  assign n794 = ( n181 & ~n793 ) | ( n181 & 1'b0 ) | ( ~n793 & 1'b0 ) ;
  assign n795 = ( n145 & ~n794 ) | ( n145 & 1'b0 ) | ( ~n794 & 1'b0 ) ;
  assign n796 = n791 &  n795 ;
  assign n797 = n788 | n796 ;
  assign n798 = n783 &  n797 ;
  assign n800 = ( n659 & ~n664 ) | ( n659 & n672 ) | ( ~n664 & n672 ) ;
  assign n799 = ( n659 & ~n713 ) | ( n659 & 1'b0 ) | ( ~n713 & 1'b0 ) ;
  assign n802 = ( n659 & ~n800 ) | ( n659 & n799 ) | ( ~n800 & n799 ) ;
  assign n801 = ( n799 & ~n672 ) | ( n799 & n800 ) | ( ~n672 & n800 ) ;
  assign n803 = ( n664 & ~n802 ) | ( n664 & n801 ) | ( ~n802 & n801 ) ;
  assign n804 = ( n798 & ~n150 ) | ( n798 & n803 ) | ( ~n150 & n803 ) ;
  assign n816 = ~n815 & n804 ;
  assign n817 = ( n816 & ~n133 ) | ( n816 & n815 ) | ( ~n133 & n815 ) ;
  assign n820 = ( n791 & ~n794 ) | ( n791 & 1'b0 ) | ( ~n794 & 1'b0 ) ;
  assign n821 = ( n145 & n788 ) | ( n145 & n820 ) | ( n788 & n820 ) ;
  assign n822 = ( n150 & ~n821 ) | ( n150 & 1'b0 ) | ( ~n821 & 1'b0 ) ;
  assign n823 = ( n811 & ~n822 ) | ( n811 & 1'b0 ) | ( ~n822 & 1'b0 ) ;
  assign n818 = ~n150 & n783 ;
  assign n819 = n797 &  n818 ;
  assign n824 = ~n803 & n819 ;
  assign n825 = ( n803 & n823 ) | ( n803 & n824 ) | ( n823 & n824 ) ;
  assign n827 = ( n680 & ~n133 ) | ( n680 & n687 ) | ( ~n133 & n687 ) ;
  assign n826 = ( n680 & n687 ) | ( n680 & n713 ) | ( n687 & n713 ) ;
  assign n828 = ~n687 & n826 ;
  assign n829 = ( n687 & ~n827 ) | ( n687 & n828 ) | ( ~n827 & n828 ) ;
  assign n830 = n683 | n710 ;
  assign n831 = ( n686 & n705 ) | ( n686 & n830 ) | ( n705 & n830 ) ;
  assign n832 = ( n686 & ~n831 ) | ( n686 & 1'b0 ) | ( ~n831 & 1'b0 ) ;
  assign n833 = ( n693 & ~n701 ) | ( n693 & n832 ) | ( ~n701 & n832 ) ;
  assign n834 = ~n693 & n833 ;
  assign n835 = n829 | n834 ;
  assign n836 = n825 | n835 ;
  assign n837 = n817 | n836 ;
  assign n895 = n736 | n837 ;
  assign n896 = ( n736 & ~n753 ) | ( n736 & n746 ) | ( ~n753 & n746 ) ;
  assign n897 = ( n753 & n895 ) | ( n753 & n896 ) | ( n895 & n896 ) ;
  assign n898 = ( n736 & ~n896 ) | ( n736 & n895 ) | ( ~n896 & n895 ) ;
  assign n899 = ( n746 & ~n897 ) | ( n746 & n898 ) | ( ~n897 & n898 ) ;
  assign n880 = ~n748 & n751 ;
  assign n881 = ( n734 & ~n748 ) | ( n734 & n880 ) | ( ~n748 & n880 ) ;
  assign n883 = ( n748 & n837 ) | ( n748 & n881 ) | ( n837 & n881 ) ;
  assign n882 = ( n837 & ~n881 ) | ( n837 & n880 ) | ( ~n881 & n880 ) ;
  assign n884 = ( n734 & ~n883 ) | ( n734 & n882 ) | ( ~n883 & n882 ) ;
  assign n871 = ~x108 & n713 ;
  assign n872 = ( x109 & ~n871 ) | ( x109 & 1'b0 ) | ( ~n871 & 1'b0 ) ;
  assign n873 = n725 | n872 ;
  assign n868 = ( n713 & ~x108 ) | ( n713 & n720 ) | ( ~x108 & n720 ) ;
  assign n869 = x108 &  n868 ;
  assign n870 = ( n715 & ~n869 ) | ( n715 & n720 ) | ( ~n869 & n720 ) ;
  assign n874 = ( n837 & ~n873 ) | ( n837 & n870 ) | ( ~n873 & n870 ) ;
  assign n876 = ( n837 & ~n874 ) | ( n837 & 1'b0 ) | ( ~n874 & 1'b0 ) ;
  assign n875 = ~n870 & n874 ;
  assign n877 = ( n873 & ~n876 ) | ( n873 & n875 ) | ( ~n876 & n875 ) ;
  assign n844 = ( x106 & ~n837 ) | ( x106 & x107 ) | ( ~n837 & x107 ) ;
  assign n850 = ( x106 & ~x107 ) | ( x106 & 1'b0 ) | ( ~x107 & 1'b0 ) ;
  assign n840 = x104 | x105 ;
  assign n845 = ~x106 & n840 ;
  assign n846 = ( x106 & ~n711 ) | ( x106 & n845 ) | ( ~n711 & n845 ) ;
  assign n847 = ( n693 & ~n701 ) | ( n693 & n846 ) | ( ~n701 & n846 ) ;
  assign n848 = ~n693 & n847 ;
  assign n849 = ( n837 & ~x107 ) | ( n837 & n848 ) | ( ~x107 & n848 ) ;
  assign n851 = ( n844 & ~n850 ) | ( n844 & n849 ) | ( ~n850 & n849 ) ;
  assign n841 = x106 | n840 ;
  assign n842 = x106 &  n837 ;
  assign n843 = ( n713 & ~n841 ) | ( n713 & n842 ) | ( ~n841 & n842 ) ;
  assign n854 = n595 | n843 ;
  assign n855 = ( n851 & ~n854 ) | ( n851 & 1'b0 ) | ( ~n854 & 1'b0 ) ;
  assign n857 = ( n713 & ~n834 ) | ( n713 & 1'b0 ) | ( ~n834 & 1'b0 ) ;
  assign n858 = ( n825 & ~n829 ) | ( n825 & n857 ) | ( ~n829 & n857 ) ;
  assign n859 = ~n825 & n858 ;
  assign n860 = ~n817 & n859 ;
  assign n856 = ~n596 & n837 ;
  assign n861 = ( n856 & ~n860 ) | ( n856 & 1'b0 ) | ( ~n860 & 1'b0 ) ;
  assign n862 = ( x108 & n860 ) | ( x108 & n861 ) | ( n860 & n861 ) ;
  assign n863 = x108 | n860 ;
  assign n864 = n856 | n863 ;
  assign n865 = ~n862 & n864 ;
  assign n866 = n855 | n865 ;
  assign n852 = n843 &  n851 ;
  assign n853 = ( n595 & ~n851 ) | ( n595 & n852 ) | ( ~n851 & n852 ) ;
  assign n885 = n492 | n853 ;
  assign n886 = ( n866 & ~n885 ) | ( n866 & 1'b0 ) | ( ~n885 & 1'b0 ) ;
  assign n887 = n877 | n886 ;
  assign n888 = ~n843 & n851 ;
  assign n889 = ( n865 & ~n595 ) | ( n865 & n888 ) | ( ~n595 & n888 ) ;
  assign n890 = ( n492 & ~n889 ) | ( n492 & 1'b0 ) | ( ~n889 & 1'b0 ) ;
  assign n891 = n396 | n890 ;
  assign n892 = ( n887 & ~n891 ) | ( n887 & 1'b0 ) | ( ~n891 & 1'b0 ) ;
  assign n893 = n884 | n892 ;
  assign n867 = ~n853 & n866 ;
  assign n878 = ( n867 & ~n492 ) | ( n867 & n877 ) | ( ~n492 & n877 ) ;
  assign n879 = ( n396 & ~n878 ) | ( n396 & 1'b0 ) | ( ~n878 & 1'b0 ) ;
  assign n907 = n315 | n879 ;
  assign n908 = ( n893 & ~n907 ) | ( n893 & 1'b0 ) | ( ~n907 & 1'b0 ) ;
  assign n909 = n899 | n908 ;
  assign n910 = ( n887 & ~n890 ) | ( n887 & 1'b0 ) | ( ~n890 & 1'b0 ) ;
  assign n911 = ( n884 & ~n396 ) | ( n884 & n910 ) | ( ~n396 & n910 ) ;
  assign n912 = ( n315 & ~n911 ) | ( n315 & 1'b0 ) | ( ~n911 & 1'b0 ) ;
  assign n913 = n240 | n912 ;
  assign n914 = ( n909 & ~n913 ) | ( n909 & 1'b0 ) | ( ~n913 & 1'b0 ) ;
  assign n894 = ~n879 & n893 ;
  assign n900 = ( n894 & ~n315 ) | ( n894 & n899 ) | ( ~n315 & n899 ) ;
  assign n901 = ( n240 & ~n900 ) | ( n240 & 1'b0 ) | ( ~n900 & 1'b0 ) ;
  assign n944 = ( n803 & ~n819 ) | ( n803 & 1'b0 ) | ( ~n819 & 1'b0 ) ;
  assign n945 = ( n822 & n837 ) | ( n822 & n944 ) | ( n837 & n944 ) ;
  assign n946 = ~n822 & n945 ;
  assign n947 = n819 | n822 ;
  assign n948 = n837 | n947 ;
  assign n949 = ( n803 & ~n947 ) | ( n803 & n948 ) | ( ~n947 & n948 ) ;
  assign n950 = ~n946 & n949 ;
  assign n951 = n804 | n811 ;
  assign n952 = n837 | n951 ;
  assign n953 = ( n825 & ~n951 ) | ( n825 & n952 ) | ( ~n951 & n952 ) ;
  assign n954 = n950 | n953 ;
  assign n902 = n768 | n837 ;
  assign n903 = ( n760 & ~n768 ) | ( n760 & n764 ) | ( ~n768 & n764 ) ;
  assign n905 = ( n768 & n902 ) | ( n768 & n903 ) | ( n902 & n903 ) ;
  assign n904 = ( n764 & ~n903 ) | ( n764 & n902 ) | ( ~n903 & n902 ) ;
  assign n906 = ( n760 & ~n905 ) | ( n760 & n904 ) | ( ~n905 & n904 ) ;
  assign n915 = n906 | n914 ;
  assign n916 = ~n901 & n915 ;
  assign n917 = ( n762 & ~n770 ) | ( n762 & n774 ) | ( ~n770 & n774 ) ;
  assign n918 = ( n770 & n837 ) | ( n770 & n917 ) | ( n837 & n917 ) ;
  assign n919 = ( n762 & ~n917 ) | ( n762 & n837 ) | ( ~n917 & n837 ) ;
  assign n920 = ( n774 & ~n918 ) | ( n774 & n919 ) | ( ~n918 & n919 ) ;
  assign n921 = ( n916 & ~n181 ) | ( n916 & n920 ) | ( ~n181 & n920 ) ;
  assign n922 = n145 | n921 ;
  assign n923 = n794 | n837 ;
  assign n924 = ( n781 & ~n790 ) | ( n781 & n794 ) | ( ~n790 & n794 ) ;
  assign n925 = ( n790 & n923 ) | ( n790 & n924 ) | ( n923 & n924 ) ;
  assign n926 = ( n794 & ~n924 ) | ( n794 & n923 ) | ( ~n924 & n923 ) ;
  assign n927 = ( n781 & ~n925 ) | ( n781 & n926 ) | ( ~n925 & n926 ) ;
  assign n928 = n181 | n901 ;
  assign n929 = ( n915 & ~n928 ) | ( n915 & 1'b0 ) | ( ~n928 & 1'b0 ) ;
  assign n930 = n920 | n929 ;
  assign n931 = ( n909 & ~n912 ) | ( n909 & 1'b0 ) | ( ~n912 & 1'b0 ) ;
  assign n932 = ( n906 & ~n240 ) | ( n906 & n931 ) | ( ~n240 & n931 ) ;
  assign n933 = ( n181 & ~n932 ) | ( n181 & 1'b0 ) | ( ~n932 & 1'b0 ) ;
  assign n934 = ( n145 & ~n933 ) | ( n145 & 1'b0 ) | ( ~n933 & 1'b0 ) ;
  assign n935 = n930 &  n934 ;
  assign n936 = n927 | n935 ;
  assign n937 = n922 &  n936 ;
  assign n939 = ( n783 & ~n788 ) | ( n783 & n796 ) | ( ~n788 & n796 ) ;
  assign n938 = ( n783 & ~n837 ) | ( n783 & 1'b0 ) | ( ~n837 & 1'b0 ) ;
  assign n941 = ( n783 & ~n939 ) | ( n783 & n938 ) | ( ~n939 & n938 ) ;
  assign n940 = ( n938 & ~n796 ) | ( n938 & n939 ) | ( ~n796 & n939 ) ;
  assign n942 = ( n788 & ~n941 ) | ( n788 & n940 ) | ( ~n941 & n940 ) ;
  assign n943 = ( n937 & ~n150 ) | ( n937 & n942 ) | ( ~n150 & n942 ) ;
  assign n955 = ~n954 & n943 ;
  assign n956 = ( n955 & ~n133 ) | ( n955 & n954 ) | ( ~n133 & n954 ) ;
  assign n957 = ~n150 & n922 ;
  assign n958 = n936 &  n957 ;
  assign n963 = ~n942 & n958 ;
  assign n959 = ( n930 & ~n933 ) | ( n930 & 1'b0 ) | ( ~n933 & 1'b0 ) ;
  assign n960 = ( n145 & n927 ) | ( n145 & n959 ) | ( n927 & n959 ) ;
  assign n961 = ( n150 & ~n960 ) | ( n150 & 1'b0 ) | ( ~n960 & 1'b0 ) ;
  assign n962 = ( n950 & ~n961 ) | ( n950 & 1'b0 ) | ( ~n961 & 1'b0 ) ;
  assign n964 = ( n942 & n963 ) | ( n942 & n962 ) | ( n963 & n962 ) ;
  assign n966 = ( n804 & ~n133 ) | ( n804 & n811 ) | ( ~n133 & n811 ) ;
  assign n965 = ( n804 & n811 ) | ( n804 & n837 ) | ( n811 & n837 ) ;
  assign n967 = ~n811 & n965 ;
  assign n968 = ( n811 & ~n966 ) | ( n811 & n967 ) | ( ~n966 & n967 ) ;
  assign n969 = n807 | n834 ;
  assign n970 = ( n810 & n829 ) | ( n810 & n969 ) | ( n829 & n969 ) ;
  assign n971 = ( n810 & ~n970 ) | ( n810 & 1'b0 ) | ( ~n970 & 1'b0 ) ;
  assign n972 = ( n817 & ~n825 ) | ( n817 & n971 ) | ( ~n825 & n971 ) ;
  assign n973 = ~n817 & n972 ;
  assign n974 = n968 | n973 ;
  assign n975 = n964 | n974 ;
  assign n976 = ~n956 &  ~n975 ;
  assign n1063 = ~n901 & n976 ;
  assign n1064 = ( n901 & ~n914 ) | ( n901 & n906 ) | ( ~n914 & n906 ) ;
  assign n1065 = ( n914 & ~n1063 ) | ( n914 & n1064 ) | ( ~n1063 & n1064 ) ;
  assign n1066 = ( n1063 & ~n901 ) | ( n1063 & n1064 ) | ( ~n901 & n1064 ) ;
  assign n1067 = ( n1065 & ~n906 ) | ( n1065 & n1066 ) | ( ~n906 & n1066 ) ;
  assign n1048 = ~n912 & n976 ;
  assign n1049 = ( n899 & ~n908 ) | ( n899 & n912 ) | ( ~n908 & n912 ) ;
  assign n1050 = ( n908 & ~n1048 ) | ( n908 & n1049 ) | ( ~n1048 & n1049 ) ;
  assign n1051 = ( n1048 & ~n912 ) | ( n1048 & n1049 ) | ( ~n912 & n1049 ) ;
  assign n1052 = ( n1050 & ~n899 ) | ( n1050 & n1051 ) | ( ~n899 & n1051 ) ;
  assign n1041 = ~n879 & n976 ;
  assign n1042 = ( n884 & ~n879 ) | ( n884 & n892 ) | ( ~n879 & n892 ) ;
  assign n1043 = ( n1041 & ~n892 ) | ( n1041 & n1042 ) | ( ~n892 & n1042 ) ;
  assign n1044 = ( n879 & ~n1041 ) | ( n879 & n1042 ) | ( ~n1041 & n1042 ) ;
  assign n1045 = ( n1043 & ~n884 ) | ( n1043 & n1044 ) | ( ~n884 & n1044 ) ;
  assign n1026 = ~n890 & n976 ;
  assign n1027 = ( n877 & ~n886 ) | ( n877 & n890 ) | ( ~n886 & n890 ) ;
  assign n1028 = ( n886 & ~n1026 ) | ( n886 & n1027 ) | ( ~n1026 & n1027 ) ;
  assign n1029 = ( n1026 & ~n890 ) | ( n1026 & n1027 ) | ( ~n890 & n1027 ) ;
  assign n1030 = ( n1028 & ~n877 ) | ( n1028 & n1029 ) | ( ~n877 & n1029 ) ;
  assign n1019 = ( n853 & ~n855 ) | ( n853 & 1'b0 ) | ( ~n855 & 1'b0 ) ;
  assign n1020 = ( n855 & ~n1019 ) | ( n855 & n865 ) | ( ~n1019 & n865 ) ;
  assign n1021 = ( n976 & ~n855 ) | ( n976 & n1020 ) | ( ~n855 & n1020 ) ;
  assign n1022 = ( n1019 & ~n976 ) | ( n1019 & n1020 ) | ( ~n976 & n1020 ) ;
  assign n1023 = ( n1021 & ~n865 ) | ( n1021 & n1022 ) | ( ~n865 & n1022 ) ;
  assign n1000 = ( n837 & ~x106 ) | ( n837 & n848 ) | ( ~x106 & n848 ) ;
  assign n1001 = x106 &  n1000 ;
  assign n1002 = ( n843 & ~n1001 ) | ( n843 & n848 ) | ( ~n1001 & n848 ) ;
  assign n1003 = ~x106 & n837 ;
  assign n1004 = ( x107 & ~n1003 ) | ( x107 & 1'b0 ) | ( ~n1003 & 1'b0 ) ;
  assign n1005 = n856 | n1004 ;
  assign n1006 = ( n976 & ~n1002 ) | ( n976 & n1005 ) | ( ~n1002 & n1005 ) ;
  assign n1007 = n1002 | n1006 ;
  assign n1008 = ~n976 & n1006 ;
  assign n1009 = ( n1007 & ~n1005 ) | ( n1007 & n1008 ) | ( ~n1005 & n1008 ) ;
  assign n988 = n840 | n976 ;
  assign n989 = ( n837 & ~n973 ) | ( n837 & 1'b0 ) | ( ~n973 & 1'b0 ) ;
  assign n990 = ( n964 & ~n968 ) | ( n964 & n989 ) | ( ~n968 & n989 ) ;
  assign n991 = ~n964 & n990 ;
  assign n992 = ~n956 & n991 ;
  assign n993 = n988 | n992 ;
  assign n994 = ( x106 & ~n993 ) | ( x106 & n992 ) | ( ~n993 & n992 ) ;
  assign n995 = x106 | n992 ;
  assign n996 = ( n988 & ~n995 ) | ( n988 & 1'b0 ) | ( ~n995 & 1'b0 ) ;
  assign n997 = n994 | n996 ;
  assign n838 = x102 | x103 ;
  assign n980 = ~x104 & n838 ;
  assign n981 = ( x104 & ~n835 ) | ( x104 & n980 ) | ( ~n835 & n980 ) ;
  assign n982 = ( n817 & ~n825 ) | ( n817 & n981 ) | ( ~n825 & n981 ) ;
  assign n983 = ~n817 & n982 ;
  assign n984 = ( x105 & ~n983 ) | ( x105 & n976 ) | ( ~n983 & n976 ) ;
  assign n979 = ( x104 & x105 ) | ( x104 & n976 ) | ( x105 & n976 ) ;
  assign n985 = ( x104 & ~x105 ) | ( x104 & 1'b0 ) | ( ~x105 & 1'b0 ) ;
  assign n986 = ( n984 & ~n979 ) | ( n984 & n985 ) | ( ~n979 & n985 ) ;
  assign n839 = x104 | n838 ;
  assign n977 = ( x104 & ~n976 ) | ( x104 & 1'b0 ) | ( ~n976 & 1'b0 ) ;
  assign n978 = ( n837 & ~n839 ) | ( n837 & n977 ) | ( ~n839 & n977 ) ;
  assign n1010 = n713 | n978 ;
  assign n1011 = n986 | n1010 ;
  assign n1012 = n997 &  n1011 ;
  assign n1013 = ~n986 & n978 ;
  assign n1014 = ( n713 & n1013 ) | ( n713 & n986 ) | ( n1013 & n986 ) ;
  assign n1015 = n595 | n1014 ;
  assign n1016 = n1012 | n1015 ;
  assign n1017 = n1009 &  n1016 ;
  assign n987 = n978 | n986 ;
  assign n998 = ( n713 & n987 ) | ( n713 & n997 ) | ( n987 & n997 ) ;
  assign n999 = n595 &  n998 ;
  assign n1031 = n492 | n999 ;
  assign n1032 = n1017 | n1031 ;
  assign n1033 = n1023 &  n1032 ;
  assign n1034 = n1012 | n1014 ;
  assign n1035 = ( n595 & n1009 ) | ( n595 & n1034 ) | ( n1009 & n1034 ) ;
  assign n1036 = n492 &  n1035 ;
  assign n1037 = n396 | n1036 ;
  assign n1038 = n1033 | n1037 ;
  assign n1039 = n1030 &  n1038 ;
  assign n1018 = n999 | n1017 ;
  assign n1024 = ( n492 & n1018 ) | ( n492 & n1023 ) | ( n1018 & n1023 ) ;
  assign n1025 = n396 &  n1024 ;
  assign n1053 = n315 | n1025 ;
  assign n1054 = n1039 | n1053 ;
  assign n1055 = n1045 &  n1054 ;
  assign n1056 = n1033 | n1036 ;
  assign n1057 = ( n396 & n1030 ) | ( n396 & n1056 ) | ( n1030 & n1056 ) ;
  assign n1058 = n315 &  n1057 ;
  assign n1059 = n240 | n1058 ;
  assign n1060 = n1055 | n1059 ;
  assign n1061 = n1052 &  n1060 ;
  assign n1040 = n1025 | n1039 ;
  assign n1046 = ( n315 & n1040 ) | ( n315 & n1045 ) | ( n1040 & n1045 ) ;
  assign n1047 = n240 &  n1046 ;
  assign n1070 = n181 | n1047 ;
  assign n1071 = n1061 | n1070 ;
  assign n1073 = n1055 | n1058 ;
  assign n1074 = ( n240 & n1052 ) | ( n240 & n1073 ) | ( n1052 & n1073 ) ;
  assign n1075 = n181 &  n1074 ;
  assign n1232 = ( n1071 & ~n1067 ) | ( n1071 & n1075 ) | ( ~n1067 & n1075 ) ;
  assign n1085 = ( n922 & ~n927 ) | ( n922 & n935 ) | ( ~n927 & n935 ) ;
  assign n1084 = n922 &  n976 ;
  assign n1087 = ( n922 & ~n1085 ) | ( n922 & n1084 ) | ( ~n1085 & n1084 ) ;
  assign n1086 = ( n1084 & ~n935 ) | ( n1084 & n1085 ) | ( ~n935 & n1085 ) ;
  assign n1088 = ( n927 & ~n1087 ) | ( n927 & n1086 ) | ( ~n1087 & n1086 ) ;
  assign n1062 = n1047 | n1061 ;
  assign n1068 = ( n181 & n1062 ) | ( n181 & n1067 ) | ( n1062 & n1067 ) ;
  assign n1069 = ~n145 & n1068 ;
  assign n1072 = n1067 &  n1071 ;
  assign n1076 = ( n145 & ~n1075 ) | ( n145 & 1'b0 ) | ( ~n1075 & 1'b0 ) ;
  assign n1077 = ~n1072 & n1076 ;
  assign n1078 = ( n920 & ~n933 ) | ( n920 & n929 ) | ( ~n933 & n929 ) ;
  assign n1079 = ( n976 & ~n929 ) | ( n976 & n1078 ) | ( ~n929 & n1078 ) ;
  assign n1080 = ( n933 & ~n976 ) | ( n933 & n1078 ) | ( ~n976 & n1078 ) ;
  assign n1081 = ( n1079 & ~n920 ) | ( n1079 & n1080 ) | ( ~n920 & n1080 ) ;
  assign n1082 = ~n1077 & n1081 ;
  assign n1083 = n1069 | n1082 ;
  assign n1089 = ( n150 & ~n1088 ) | ( n150 & n1083 ) | ( ~n1088 & n1083 ) ;
  assign n1090 = ( n942 & ~n961 ) | ( n942 & 1'b0 ) | ( ~n961 & 1'b0 ) ;
  assign n1091 = ( n958 & ~n976 ) | ( n958 & n1090 ) | ( ~n976 & n1090 ) ;
  assign n1092 = ~n958 & n1091 ;
  assign n1093 = n958 | n961 ;
  assign n1094 = ~n1093 & n976 ;
  assign n1095 = ( n1094 & ~n942 ) | ( n1094 & n1093 ) | ( ~n942 & n1093 ) ;
  assign n1096 = n1092 | n1095 ;
  assign n1097 = n943 | n950 ;
  assign n1098 = ~n1097 & n976 ;
  assign n1099 = ( n1098 & ~n964 ) | ( n1098 & n1097 ) | ( ~n964 & n1097 ) ;
  assign n1100 = n1096 &  n1099 ;
  assign n1101 = ~n1089 & n1100 ;
  assign n1102 = ( n133 & ~n1101 ) | ( n133 & n1100 ) | ( ~n1101 & n1100 ) ;
  assign n1105 = n1072 | n1075 ;
  assign n1106 = ( n1081 & ~n145 ) | ( n1081 & n1105 ) | ( ~n145 & n1105 ) ;
  assign n1107 = n150 &  n1106 ;
  assign n1108 = n1096 | n1107 ;
  assign n1103 = n150 | n1069 ;
  assign n1104 = n1082 | n1103 ;
  assign n1109 = n1088 | n1104 ;
  assign n1110 = ( n1108 & ~n1088 ) | ( n1108 & n1109 ) | ( ~n1088 & n1109 ) ;
  assign n1112 = ( n943 & ~n133 ) | ( n943 & n950 ) | ( ~n133 & n950 ) ;
  assign n1111 = ( n943 & ~n976 ) | ( n943 & n950 ) | ( ~n976 & n950 ) ;
  assign n1113 = ~n950 & n1111 ;
  assign n1114 = ( n950 & ~n1112 ) | ( n950 & n1113 ) | ( ~n1112 & n1113 ) ;
  assign n1115 = n946 | n973 ;
  assign n1116 = ( n949 & n968 ) | ( n949 & n1115 ) | ( n968 & n1115 ) ;
  assign n1117 = ( n949 & ~n1116 ) | ( n949 & 1'b0 ) | ( ~n1116 & 1'b0 ) ;
  assign n1118 = ( n956 & ~n964 ) | ( n956 & n1117 ) | ( ~n964 & n1117 ) ;
  assign n1119 = ~n956 & n1118 ;
  assign n1120 = n1114 | n1119 ;
  assign n1121 = ( n1110 & ~n1120 ) | ( n1110 & 1'b0 ) | ( ~n1120 & 1'b0 ) ;
  assign n1122 = n1102 &  n1121 ;
  assign n1231 = ~n1075 & n1122 ;
  assign n1233 = ( n1071 & ~n1232 ) | ( n1071 & n1231 ) | ( ~n1232 & n1231 ) ;
  assign n1234 = ( n1231 & ~n1075 ) | ( n1231 & n1232 ) | ( ~n1075 & n1232 ) ;
  assign n1235 = ( n1067 & ~n1233 ) | ( n1067 & n1234 ) | ( ~n1233 & n1234 ) ;
  assign n1224 = ~n1047 & n1122 ;
  assign n1225 = ( n1047 & n1052 ) | ( n1047 & n1060 ) | ( n1052 & n1060 ) ;
  assign n1227 = ( n1224 & ~n1047 ) | ( n1224 & n1225 ) | ( ~n1047 & n1225 ) ;
  assign n1226 = ( n1060 & ~n1225 ) | ( n1060 & n1224 ) | ( ~n1225 & n1224 ) ;
  assign n1228 = ( n1052 & ~n1227 ) | ( n1052 & n1226 ) | ( ~n1227 & n1226 ) ;
  assign n1210 = ( n1054 & ~n1045 ) | ( n1054 & n1058 ) | ( ~n1045 & n1058 ) ;
  assign n1209 = ~n1058 & n1122 ;
  assign n1211 = ( n1054 & ~n1210 ) | ( n1054 & n1209 ) | ( ~n1210 & n1209 ) ;
  assign n1212 = ( n1209 & ~n1058 ) | ( n1209 & n1210 ) | ( ~n1058 & n1210 ) ;
  assign n1213 = ( n1045 & ~n1211 ) | ( n1045 & n1212 ) | ( ~n1211 & n1212 ) ;
  assign n1202 = n1038 | n1122 ;
  assign n1203 = ( n1025 & ~n1122 ) | ( n1025 & n1202 ) | ( ~n1122 & n1202 ) ;
  assign n1204 = ( n1025 & ~n1203 ) | ( n1025 & n1030 ) | ( ~n1203 & n1030 ) ;
  assign n1205 = ( n1030 & ~n1025 ) | ( n1030 & n1203 ) | ( ~n1025 & n1203 ) ;
  assign n1206 = ( n1204 & ~n1030 ) | ( n1204 & n1205 ) | ( ~n1030 & n1205 ) ;
  assign n1187 = ~n1036 & n1122 ;
  assign n1188 = ( n1023 & n1032 ) | ( n1023 & n1036 ) | ( n1032 & n1036 ) ;
  assign n1190 = ( n1187 & ~n1036 ) | ( n1187 & n1188 ) | ( ~n1036 & n1188 ) ;
  assign n1189 = ( n1032 & ~n1188 ) | ( n1032 & n1187 ) | ( ~n1188 & n1187 ) ;
  assign n1191 = ( n1023 & ~n1190 ) | ( n1023 & n1189 ) | ( ~n1190 & n1189 ) ;
  assign n1181 = ( n999 & ~n1009 ) | ( n999 & n1016 ) | ( ~n1009 & n1016 ) ;
  assign n1180 = ~n999 & n1122 ;
  assign n1182 = ( n1016 & ~n1181 ) | ( n1016 & n1180 ) | ( ~n1181 & n1180 ) ;
  assign n1183 = ( n1180 & ~n999 ) | ( n1180 & n1181 ) | ( ~n999 & n1181 ) ;
  assign n1184 = ( n1009 & ~n1182 ) | ( n1009 & n1183 ) | ( ~n1182 & n1183 ) ;
  assign n1165 = n1011 &  n1014 ;
  assign n1166 = ( n1011 & n1122 ) | ( n1011 & n1165 ) | ( n1122 & n1165 ) ;
  assign n1167 = ( n997 & ~n1011 ) | ( n997 & n1166 ) | ( ~n1011 & n1166 ) ;
  assign n1168 = ( n997 & ~n1166 ) | ( n997 & n1011 ) | ( ~n1166 & n1011 ) ;
  assign n1169 = ( n1167 & ~n997 ) | ( n1167 & n1168 ) | ( ~n997 & n1168 ) ;
  assign n1153 = ( x104 & ~n983 ) | ( x104 & n976 ) | ( ~n983 & n976 ) ;
  assign n1154 = ( x104 & ~n1153 ) | ( x104 & 1'b0 ) | ( ~n1153 & 1'b0 ) ;
  assign n1155 = ( n978 & ~n1154 ) | ( n978 & n983 ) | ( ~n1154 & n983 ) ;
  assign n1156 = x104 | n976 ;
  assign n1157 = x105 &  n1156 ;
  assign n1158 = ( n988 & ~n1157 ) | ( n988 & 1'b0 ) | ( ~n1157 & 1'b0 ) ;
  assign n1159 = ( n1155 & ~n1122 ) | ( n1155 & n1158 ) | ( ~n1122 & n1158 ) ;
  assign n1160 = ~n1155 & n1159 ;
  assign n1161 = n1122 | n1159 ;
  assign n1162 = ( n1160 & ~n1158 ) | ( n1160 & n1161 ) | ( ~n1158 & n1161 ) ;
  assign n1125 = x100 | x101 ;
  assign n1130 = ~x102 & n1125 ;
  assign n1131 = ( x102 & ~n974 ) | ( x102 & n1130 ) | ( ~n974 & n1130 ) ;
  assign n1132 = ( n956 & ~n964 ) | ( n956 & n1131 ) | ( ~n964 & n1131 ) ;
  assign n1133 = ~n956 & n1132 ;
  assign n1134 = ( x103 & ~n1133 ) | ( x103 & n1122 ) | ( ~n1133 & n1122 ) ;
  assign n1129 = ( x102 & x103 ) | ( x102 & n1122 ) | ( x103 & n1122 ) ;
  assign n1135 = ( x102 & ~x103 ) | ( x102 & 1'b0 ) | ( ~x103 & 1'b0 ) ;
  assign n1136 = ( n1134 & ~n1129 ) | ( n1134 & n1135 ) | ( ~n1129 & n1135 ) ;
  assign n1127 = ( x102 & ~n1122 ) | ( x102 & 1'b0 ) | ( ~n1122 & 1'b0 ) ;
  assign n1126 = x102 | n1125 ;
  assign n1128 = ( n976 & ~n1127 ) | ( n976 & n1126 ) | ( ~n1127 & n1126 ) ;
  assign n1139 = ~n837 & n1128 ;
  assign n1140 = ~n1136 & n1139 ;
  assign n1141 = n838 | n1122 ;
  assign n1142 = n976 | n1119 ;
  assign n1143 = ( n1110 & n1114 ) | ( n1110 & n1142 ) | ( n1114 & n1142 ) ;
  assign n1144 = ( n1110 & ~n1143 ) | ( n1110 & 1'b0 ) | ( ~n1143 & 1'b0 ) ;
  assign n1145 = n1102 &  n1144 ;
  assign n1146 = n1141 | n1145 ;
  assign n1147 = ( x104 & ~n1146 ) | ( x104 & n1145 ) | ( ~n1146 & n1145 ) ;
  assign n1148 = x104 | n1145 ;
  assign n1149 = ( n1141 & ~n1148 ) | ( n1141 & 1'b0 ) | ( ~n1148 & 1'b0 ) ;
  assign n1150 = n1147 | n1149 ;
  assign n1151 = ~n1140 & n1150 ;
  assign n1137 = n1128 | n1136 ;
  assign n1138 = ( n837 & ~n1137 ) | ( n837 & n1136 ) | ( ~n1137 & n1136 ) ;
  assign n1170 = n713 | n1138 ;
  assign n1171 = n1151 | n1170 ;
  assign n1172 = ~n1162 & n1171 ;
  assign n1173 = ( n1128 & ~n1136 ) | ( n1128 & 1'b0 ) | ( ~n1136 & 1'b0 ) ;
  assign n1174 = ( n837 & ~n1173 ) | ( n837 & n1150 ) | ( ~n1173 & n1150 ) ;
  assign n1175 = n713 &  n1174 ;
  assign n1176 = n595 | n1175 ;
  assign n1177 = n1172 | n1176 ;
  assign n1178 = n1169 &  n1177 ;
  assign n1152 = n1138 | n1151 ;
  assign n1163 = ( n713 & ~n1162 ) | ( n713 & n1152 ) | ( ~n1162 & n1152 ) ;
  assign n1164 = n595 &  n1163 ;
  assign n1192 = n492 | n1164 ;
  assign n1193 = n1178 | n1192 ;
  assign n1194 = n1184 &  n1193 ;
  assign n1195 = n1172 | n1175 ;
  assign n1196 = ( n595 & n1169 ) | ( n595 & n1195 ) | ( n1169 & n1195 ) ;
  assign n1197 = n492 &  n1196 ;
  assign n1198 = n396 | n1197 ;
  assign n1199 = n1194 | n1198 ;
  assign n1200 = n1191 &  n1199 ;
  assign n1179 = n1164 | n1178 ;
  assign n1185 = ( n492 & n1179 ) | ( n492 & n1184 ) | ( n1179 & n1184 ) ;
  assign n1186 = n396 &  n1185 ;
  assign n1214 = n315 | n1186 ;
  assign n1215 = n1200 | n1214 ;
  assign n1216 = n1206 &  n1215 ;
  assign n1217 = n1194 | n1197 ;
  assign n1218 = ( n396 & n1191 ) | ( n396 & n1217 ) | ( n1191 & n1217 ) ;
  assign n1219 = n315 &  n1218 ;
  assign n1220 = n240 | n1219 ;
  assign n1221 = n1216 | n1220 ;
  assign n1222 = n1213 &  n1221 ;
  assign n1201 = n1186 | n1200 ;
  assign n1207 = ( n315 & n1201 ) | ( n315 & n1206 ) | ( n1201 & n1206 ) ;
  assign n1208 = n240 &  n1207 ;
  assign n1236 = n181 | n1208 ;
  assign n1237 = n1222 | n1236 ;
  assign n1238 = n1228 &  n1237 ;
  assign n1239 = n1216 | n1219 ;
  assign n1240 = ( n240 & n1213 ) | ( n240 & n1239 ) | ( n1213 & n1239 ) ;
  assign n1241 = n181 &  n1240 ;
  assign n1242 = ( n145 & ~n1241 ) | ( n145 & 1'b0 ) | ( ~n1241 & 1'b0 ) ;
  assign n1243 = ~n1238 & n1242 ;
  assign n1244 = ( n1235 & ~n1243 ) | ( n1235 & 1'b0 ) | ( ~n1243 & 1'b0 ) ;
  assign n1223 = n1208 | n1222 ;
  assign n1229 = ( n181 & n1223 ) | ( n181 & n1228 ) | ( n1223 & n1228 ) ;
  assign n1230 = ~n145 & n1229 ;
  assign n1264 = n150 | n1230 ;
  assign n1265 = n1244 | n1264 ;
  assign n1246 = ( n1077 & ~n1069 ) | ( n1077 & n1081 ) | ( ~n1069 & n1081 ) ;
  assign n1247 = ( n1122 & ~n1077 ) | ( n1122 & n1246 ) | ( ~n1077 & n1246 ) ;
  assign n1248 = ( n1069 & ~n1122 ) | ( n1069 & n1246 ) | ( ~n1122 & n1246 ) ;
  assign n1249 = ( n1247 & ~n1081 ) | ( n1247 & n1248 ) | ( ~n1081 & n1248 ) ;
  assign n1245 = n1230 | n1244 ;
  assign n1250 = ( n150 & ~n1249 ) | ( n150 & n1245 ) | ( ~n1249 & n1245 ) ;
  assign n1251 = n1088 &  n1104 ;
  assign n1252 = ( n1107 & ~n1122 ) | ( n1107 & n1251 ) | ( ~n1122 & n1251 ) ;
  assign n1253 = ~n1107 & n1252 ;
  assign n1254 = ( n1104 & ~n1107 ) | ( n1104 & 1'b0 ) | ( ~n1107 & 1'b0 ) ;
  assign n1255 = n1122 &  n1254 ;
  assign n1256 = ( n1088 & ~n1255 ) | ( n1088 & n1254 ) | ( ~n1255 & n1254 ) ;
  assign n1257 = ~n1253 & n1256 ;
  assign n1258 = n1089 &  n1096 ;
  assign n1259 = n1122 &  n1258 ;
  assign n1260 = ( n1110 & ~n1258 ) | ( n1110 & n1259 ) | ( ~n1258 & n1259 ) ;
  assign n1261 = ~n1257 & n1260 ;
  assign n1262 = ~n1250 & n1261 ;
  assign n1263 = ( n133 & ~n1262 ) | ( n133 & n1261 ) | ( ~n1262 & n1261 ) ;
  assign n1270 = n1265 | n1249 ;
  assign n1266 = n1238 | n1241 ;
  assign n1267 = ( n1235 & ~n145 ) | ( n1235 & n1266 ) | ( ~n145 & n1266 ) ;
  assign n1268 = n150 &  n1267 ;
  assign n1269 = ( n1257 & ~n1268 ) | ( n1257 & 1'b0 ) | ( ~n1268 & 1'b0 ) ;
  assign n1271 = ( n1249 & ~n1270 ) | ( n1249 & n1269 ) | ( ~n1270 & n1269 ) ;
  assign n1273 = ( n133 & n1089 ) | ( n133 & n1096 ) | ( n1089 & n1096 ) ;
  assign n1272 = ( n1089 & n1096 ) | ( n1089 & n1122 ) | ( n1096 & n1122 ) ;
  assign n1274 = ( n1096 & ~n1272 ) | ( n1096 & 1'b0 ) | ( ~n1272 & 1'b0 ) ;
  assign n1275 = ( n1273 & ~n1096 ) | ( n1273 & n1274 ) | ( ~n1096 & n1274 ) ;
  assign n1276 = n1092 | n1119 ;
  assign n1277 = ( n1114 & ~n1095 ) | ( n1114 & n1276 ) | ( ~n1095 & n1276 ) ;
  assign n1278 = n1095 | n1277 ;
  assign n1279 = ( n1102 & ~n1110 ) | ( n1102 & n1278 ) | ( ~n1110 & n1278 ) ;
  assign n1280 = ( n1102 & ~n1279 ) | ( n1102 & 1'b0 ) | ( ~n1279 & 1'b0 ) ;
  assign n1281 = n1275 | n1280 ;
  assign n1282 = n1271 | n1281 ;
  assign n1283 = ~n1263 |  n1282 ;
  assign n1420 = ( n1249 & ~n1268 ) | ( n1249 & 1'b0 ) | ( ~n1268 & 1'b0 ) ;
  assign n1421 = ( n1283 & ~n1265 ) | ( n1283 & n1420 ) | ( ~n1265 & n1420 ) ;
  assign n1422 = n1265 &  n1421 ;
  assign n1423 = ( n1265 & ~n1268 ) | ( n1265 & 1'b0 ) | ( ~n1268 & 1'b0 ) ;
  assign n1424 = ~n1283 & n1423 ;
  assign n1425 = ( n1249 & ~n1424 ) | ( n1249 & n1423 ) | ( ~n1424 & n1423 ) ;
  assign n1426 = ~n1422 & n1425 ;
  assign n1427 = ( n1250 & ~n1257 ) | ( n1250 & 1'b0 ) | ( ~n1257 & 1'b0 ) ;
  assign n1428 = ~n1283 & n1427 ;
  assign n1429 = ( n1271 & ~n1428 ) | ( n1271 & n1427 ) | ( ~n1428 & n1427 ) ;
  assign n1430 = n1426 | n1429 ;
  assign n1284 = x100 &  n1283 ;
  assign n1123 = x98 | x99 ;
  assign n1124 = x100 | n1123 ;
  assign n1285 = ( n1122 & ~n1284 ) | ( n1122 & n1124 ) | ( ~n1284 & n1124 ) ;
  assign n1286 = ( x100 & ~n1283 ) | ( x100 & x101 ) | ( ~n1283 & x101 ) ;
  assign n1292 = ( x100 & ~x101 ) | ( x100 & 1'b0 ) | ( ~x101 & 1'b0 ) ;
  assign n1287 = ~x100 & n1123 ;
  assign n1288 = ( x100 & ~n1120 ) | ( x100 & n1287 ) | ( ~n1120 & n1287 ) ;
  assign n1289 = ( n1110 & ~n1102 ) | ( n1110 & n1288 ) | ( ~n1102 & n1288 ) ;
  assign n1290 = n1102 &  n1289 ;
  assign n1291 = ( n1283 & ~x101 ) | ( n1283 & n1290 ) | ( ~x101 & n1290 ) ;
  assign n1293 = ( n1286 & ~n1292 ) | ( n1286 & n1291 ) | ( ~n1292 & n1291 ) ;
  assign n1294 = n1285 &  n1293 ;
  assign n1296 = n1122 | n1280 ;
  assign n1297 = ( n1275 & ~n1271 ) | ( n1275 & n1296 ) | ( ~n1271 & n1296 ) ;
  assign n1298 = n1271 | n1297 ;
  assign n1299 = ( n1263 & ~n1298 ) | ( n1263 & 1'b0 ) | ( ~n1298 & 1'b0 ) ;
  assign n1295 = ~n1125 & n1283 ;
  assign n1300 = ( n1295 & ~n1299 ) | ( n1295 & 1'b0 ) | ( ~n1299 & 1'b0 ) ;
  assign n1301 = ( x102 & n1299 ) | ( x102 & n1300 ) | ( n1299 & n1300 ) ;
  assign n1302 = x102 | n1299 ;
  assign n1303 = n1295 | n1302 ;
  assign n1304 = ~n1301 & n1303 ;
  assign n1305 = ( n976 & n1294 ) | ( n976 & n1304 ) | ( n1294 & n1304 ) ;
  assign n1306 = ( n837 & ~n1305 ) | ( n837 & 1'b0 ) | ( ~n1305 & 1'b0 ) ;
  assign n1310 = x102 | n1122 ;
  assign n1311 = x103 &  n1310 ;
  assign n1312 = ( n1141 & ~n1311 ) | ( n1141 & 1'b0 ) | ( ~n1311 & 1'b0 ) ;
  assign n1307 = ( x102 & ~n1133 ) | ( x102 & n1122 ) | ( ~n1133 & n1122 ) ;
  assign n1308 = ( x102 & ~n1307 ) | ( x102 & 1'b0 ) | ( ~n1307 & 1'b0 ) ;
  assign n1309 = ( n1128 & ~n1133 ) | ( n1128 & n1308 ) | ( ~n1133 & n1308 ) ;
  assign n1313 = ( n1283 & ~n1309 ) | ( n1283 & n1312 ) | ( ~n1309 & n1312 ) ;
  assign n1314 = n1309 &  n1313 ;
  assign n1315 = ( n1283 & ~n1313 ) | ( n1283 & 1'b0 ) | ( ~n1313 & 1'b0 ) ;
  assign n1316 = ( n1312 & ~n1314 ) | ( n1312 & n1315 ) | ( ~n1314 & n1315 ) ;
  assign n1317 = n976 &  n1285 ;
  assign n1318 = n1293 &  n1317 ;
  assign n1319 = n1304 | n1318 ;
  assign n1320 = ~n1285 & n1293 ;
  assign n1321 = ( n976 & ~n1320 ) | ( n976 & n1293 ) | ( ~n1320 & n1293 ) ;
  assign n1322 = ~n837 & n1321 ;
  assign n1323 = n1319 &  n1322 ;
  assign n1324 = ( n1316 & ~n1323 ) | ( n1316 & 1'b0 ) | ( ~n1323 & 1'b0 ) ;
  assign n1325 = n1306 | n1324 ;
  assign n1326 = ( n1138 & ~n1140 ) | ( n1138 & 1'b0 ) | ( ~n1140 & 1'b0 ) ;
  assign n1327 = ( n1150 & ~n1140 ) | ( n1150 & n1326 ) | ( ~n1140 & n1326 ) ;
  assign n1328 = ( n1140 & n1283 ) | ( n1140 & n1327 ) | ( n1283 & n1327 ) ;
  assign n1329 = ( n1283 & ~n1327 ) | ( n1283 & n1326 ) | ( ~n1327 & n1326 ) ;
  assign n1330 = ( n1150 & ~n1328 ) | ( n1150 & n1329 ) | ( ~n1328 & n1329 ) ;
  assign n1331 = ( n713 & n1325 ) | ( n713 & n1330 ) | ( n1325 & n1330 ) ;
  assign n1332 = n595 &  n1331 ;
  assign n1333 = n1175 | n1283 ;
  assign n1334 = ( n1162 & n1171 ) | ( n1162 & n1175 ) | ( n1171 & n1175 ) ;
  assign n1335 = ( n1333 & ~n1171 ) | ( n1333 & n1334 ) | ( ~n1171 & n1334 ) ;
  assign n1336 = ( n1175 & ~n1334 ) | ( n1175 & n1333 ) | ( ~n1334 & n1333 ) ;
  assign n1337 = ( n1162 & ~n1335 ) | ( n1162 & n1336 ) | ( ~n1335 & n1336 ) ;
  assign n1338 = n713 | n1306 ;
  assign n1339 = n1324 | n1338 ;
  assign n1340 = n1330 &  n1339 ;
  assign n1341 = n1319 &  n1321 ;
  assign n1342 = ( n837 & ~n1341 ) | ( n837 & n1316 ) | ( ~n1341 & n1316 ) ;
  assign n1343 = n713 &  n1342 ;
  assign n1344 = n595 | n1343 ;
  assign n1345 = n1340 | n1344 ;
  assign n1346 = ~n1337 & n1345 ;
  assign n1347 = n1332 | n1346 ;
  assign n1348 = n1164 | n1283 ;
  assign n1349 = ( n1164 & n1169 ) | ( n1164 & n1177 ) | ( n1169 & n1177 ) ;
  assign n1350 = ( n1348 & ~n1177 ) | ( n1348 & n1349 ) | ( ~n1177 & n1349 ) ;
  assign n1351 = ( n1164 & ~n1349 ) | ( n1164 & n1348 ) | ( ~n1349 & n1348 ) ;
  assign n1352 = ( n1169 & ~n1350 ) | ( n1169 & n1351 ) | ( ~n1350 & n1351 ) ;
  assign n1353 = ( n492 & n1347 ) | ( n492 & n1352 ) | ( n1347 & n1352 ) ;
  assign n1354 = n396 &  n1353 ;
  assign n1356 = ( n1193 & ~n1184 ) | ( n1193 & n1197 ) | ( ~n1184 & n1197 ) ;
  assign n1355 = n1197 | n1283 ;
  assign n1358 = ( n1197 & ~n1356 ) | ( n1197 & n1355 ) | ( ~n1356 & n1355 ) ;
  assign n1357 = ( n1355 & ~n1193 ) | ( n1355 & n1356 ) | ( ~n1193 & n1356 ) ;
  assign n1359 = ( n1184 & ~n1358 ) | ( n1184 & n1357 ) | ( ~n1358 & n1357 ) ;
  assign n1360 = n492 | n1332 ;
  assign n1361 = n1346 | n1360 ;
  assign n1362 = n1352 &  n1361 ;
  assign n1363 = n1340 | n1343 ;
  assign n1364 = ( n595 & ~n1337 ) | ( n595 & n1363 ) | ( ~n1337 & n1363 ) ;
  assign n1365 = n492 &  n1364 ;
  assign n1366 = n396 | n1365 ;
  assign n1367 = n1362 | n1366 ;
  assign n1368 = n1359 &  n1367 ;
  assign n1369 = n1354 | n1368 ;
  assign n1371 = ( n1186 & ~n1191 ) | ( n1186 & n1199 ) | ( ~n1191 & n1199 ) ;
  assign n1370 = n1186 | n1283 ;
  assign n1373 = ( n1186 & ~n1371 ) | ( n1186 & n1370 ) | ( ~n1371 & n1370 ) ;
  assign n1372 = ( n1370 & ~n1199 ) | ( n1370 & n1371 ) | ( ~n1199 & n1371 ) ;
  assign n1374 = ( n1191 & ~n1373 ) | ( n1191 & n1372 ) | ( ~n1373 & n1372 ) ;
  assign n1375 = ( n315 & n1369 ) | ( n315 & n1374 ) | ( n1369 & n1374 ) ;
  assign n1376 = n240 &  n1375 ;
  assign n1377 = n1219 | n1283 ;
  assign n1378 = ( n1206 & n1215 ) | ( n1206 & n1219 ) | ( n1215 & n1219 ) ;
  assign n1379 = ( n1377 & ~n1215 ) | ( n1377 & n1378 ) | ( ~n1215 & n1378 ) ;
  assign n1380 = ( n1219 & ~n1378 ) | ( n1219 & n1377 ) | ( ~n1378 & n1377 ) ;
  assign n1381 = ( n1206 & ~n1379 ) | ( n1206 & n1380 ) | ( ~n1379 & n1380 ) ;
  assign n1382 = n315 | n1354 ;
  assign n1383 = n1368 | n1382 ;
  assign n1384 = n1374 &  n1383 ;
  assign n1385 = n1362 | n1365 ;
  assign n1386 = ( n396 & n1359 ) | ( n396 & n1385 ) | ( n1359 & n1385 ) ;
  assign n1387 = n315 &  n1386 ;
  assign n1388 = n240 | n1387 ;
  assign n1389 = n1384 | n1388 ;
  assign n1390 = n1381 &  n1389 ;
  assign n1391 = n1376 | n1390 ;
  assign n1392 = ~n1221 & n1283 ;
  assign n1393 = ( n1208 & ~n1392 ) | ( n1208 & n1283 ) | ( ~n1392 & n1283 ) ;
  assign n1394 = ( n1208 & ~n1393 ) | ( n1208 & n1213 ) | ( ~n1393 & n1213 ) ;
  assign n1395 = ( n1213 & ~n1208 ) | ( n1213 & n1393 ) | ( ~n1208 & n1393 ) ;
  assign n1396 = ( n1394 & ~n1213 ) | ( n1394 & n1395 ) | ( ~n1213 & n1395 ) ;
  assign n1397 = ( n181 & n1391 ) | ( n181 & n1396 ) | ( n1391 & n1396 ) ;
  assign n1398 = ~n145 & n1397 ;
  assign n1400 = ( n1237 & ~n1228 ) | ( n1237 & n1241 ) | ( ~n1228 & n1241 ) ;
  assign n1399 = n1241 | n1283 ;
  assign n1402 = ( n1241 & ~n1400 ) | ( n1241 & n1399 ) | ( ~n1400 & n1399 ) ;
  assign n1401 = ( n1399 & ~n1237 ) | ( n1399 & n1400 ) | ( ~n1237 & n1400 ) ;
  assign n1403 = ( n1228 & ~n1402 ) | ( n1228 & n1401 ) | ( ~n1402 & n1401 ) ;
  assign n1404 = n181 | n1376 ;
  assign n1405 = n1390 | n1404 ;
  assign n1406 = n1396 &  n1405 ;
  assign n1407 = n1384 | n1387 ;
  assign n1408 = ( n240 & n1381 ) | ( n240 & n1407 ) | ( n1381 & n1407 ) ;
  assign n1409 = n181 &  n1408 ;
  assign n1410 = ( n145 & ~n1409 ) | ( n145 & 1'b0 ) | ( ~n1409 & 1'b0 ) ;
  assign n1411 = ~n1406 & n1410 ;
  assign n1412 = ( n1403 & ~n1411 ) | ( n1403 & 1'b0 ) | ( ~n1411 & 1'b0 ) ;
  assign n1413 = n1398 | n1412 ;
  assign n1414 = n1243 &  n1283 ;
  assign n1415 = ( n1230 & ~n1414 ) | ( n1230 & n1283 ) | ( ~n1414 & n1283 ) ;
  assign n1416 = ( n1230 & ~n1415 ) | ( n1230 & n1235 ) | ( ~n1415 & n1235 ) ;
  assign n1417 = ( n1235 & ~n1230 ) | ( n1235 & n1415 ) | ( ~n1230 & n1415 ) ;
  assign n1418 = ( n1416 & ~n1235 ) | ( n1416 & n1417 ) | ( ~n1235 & n1417 ) ;
  assign n1419 = ( n150 & n1413 ) | ( n150 & n1418 ) | ( n1413 & n1418 ) ;
  assign n1431 = n1419 | n1430 ;
  assign n1432 = ( n133 & ~n1430 ) | ( n133 & n1431 ) | ( ~n1430 & n1431 ) ;
  assign n1435 = n1406 | n1409 ;
  assign n1436 = ( n1403 & ~n145 ) | ( n1403 & n1435 ) | ( ~n145 & n1435 ) ;
  assign n1437 = n150 &  n1436 ;
  assign n1438 = ( n1426 & ~n1437 ) | ( n1426 & 1'b0 ) | ( ~n1437 & 1'b0 ) ;
  assign n1433 = n150 | n1398 ;
  assign n1434 = n1412 | n1433 ;
  assign n1439 = ( n1418 & ~n1434 ) | ( n1418 & 1'b0 ) | ( ~n1434 & 1'b0 ) ;
  assign n1440 = ( n1438 & ~n1418 ) | ( n1438 & n1439 ) | ( ~n1418 & n1439 ) ;
  assign n1442 = ( n133 & ~n1257 ) | ( n133 & n1250 ) | ( ~n1257 & n1250 ) ;
  assign n1441 = ( n1257 & ~n1250 ) | ( n1257 & n1283 ) | ( ~n1250 & n1283 ) ;
  assign n1443 = ~n1257 & n1441 ;
  assign n1444 = ( n1257 & n1442 ) | ( n1257 & n1443 ) | ( n1442 & n1443 ) ;
  assign n1445 = n1253 | n1280 ;
  assign n1446 = ( n1256 & n1275 ) | ( n1256 & n1445 ) | ( n1275 & n1445 ) ;
  assign n1447 = ( n1256 & ~n1446 ) | ( n1256 & 1'b0 ) | ( ~n1446 & 1'b0 ) ;
  assign n1448 = ( n1263 & ~n1447 ) | ( n1263 & n1271 ) | ( ~n1447 & n1271 ) ;
  assign n1449 = ( n1263 & ~n1448 ) | ( n1263 & 1'b0 ) | ( ~n1448 & 1'b0 ) ;
  assign n1450 = n1444 | n1449 ;
  assign n1451 = n1440 | n1450 ;
  assign n1452 = n1432 &  ~n1451 ;
  assign n1598 = ~n1398 & n1452 ;
  assign n1599 = ( n1403 & ~n1398 ) | ( n1403 & n1411 ) | ( ~n1398 & n1411 ) ;
  assign n1600 = ( n1598 & ~n1411 ) | ( n1598 & n1599 ) | ( ~n1411 & n1599 ) ;
  assign n1601 = ( n1398 & ~n1598 ) | ( n1398 & n1599 ) | ( ~n1598 & n1599 ) ;
  assign n1602 = ( n1600 & ~n1403 ) | ( n1600 & n1601 ) | ( ~n1403 & n1601 ) ;
  assign n1532 = n1345 | n1452 ;
  assign n1533 = ( n1332 & ~n1452 ) | ( n1332 & n1337 ) | ( ~n1452 & n1337 ) ;
  assign n1534 = ( n1452 & n1532 ) | ( n1452 & n1533 ) | ( n1532 & n1533 ) ;
  assign n1535 = ( n1332 & ~n1533 ) | ( n1332 & n1532 ) | ( ~n1533 & n1532 ) ;
  assign n1536 = ( n1337 & ~n1534 ) | ( n1337 & n1535 ) | ( ~n1534 & n1535 ) ;
  assign n1455 = x96 | x97 ;
  assign n1460 = ~x98 & n1455 ;
  assign n1461 = ( x98 & ~n1281 ) | ( x98 & n1460 ) | ( ~n1281 & n1460 ) ;
  assign n1462 = ( n1263 & ~n1461 ) | ( n1263 & n1271 ) | ( ~n1461 & n1271 ) ;
  assign n1463 = ( n1263 & ~n1462 ) | ( n1263 & 1'b0 ) | ( ~n1462 & 1'b0 ) ;
  assign n1464 = ( x99 & ~n1463 ) | ( x99 & n1452 ) | ( ~n1463 & n1452 ) ;
  assign n1459 = ( x98 & x99 ) | ( x98 & n1452 ) | ( x99 & n1452 ) ;
  assign n1465 = ( x98 & ~x99 ) | ( x98 & 1'b0 ) | ( ~x99 & 1'b0 ) ;
  assign n1466 = ( n1464 & ~n1459 ) | ( n1464 & n1465 ) | ( ~n1459 & n1465 ) ;
  assign n1456 = x98 | n1455 ;
  assign n1457 = ( x98 & ~n1452 ) | ( x98 & 1'b0 ) | ( ~n1452 & 1'b0 ) ;
  assign n1458 = ( n1283 & ~n1456 ) | ( n1283 & n1457 ) | ( ~n1456 & n1457 ) ;
  assign n1467 = ( n1458 & ~n1466 ) | ( n1458 & 1'b0 ) | ( ~n1466 & 1'b0 ) ;
  assign n1468 = ( n1466 & ~n1122 ) | ( n1466 & n1467 ) | ( ~n1122 & n1467 ) ;
  assign n1469 = ( n1122 & ~n1458 ) | ( n1122 & 1'b0 ) | ( ~n1458 & 1'b0 ) ;
  assign n1470 = ~n1466 & n1469 ;
  assign n1471 = n1123 | n1452 ;
  assign n1472 = ( n1283 & ~n1449 ) | ( n1283 & 1'b0 ) | ( ~n1449 & 1'b0 ) ;
  assign n1473 = ( n1440 & ~n1444 ) | ( n1440 & n1472 ) | ( ~n1444 & n1472 ) ;
  assign n1474 = ~n1440 & n1473 ;
  assign n1475 = n1432 &  n1474 ;
  assign n1476 = n1471 | n1475 ;
  assign n1477 = ( x100 & ~n1476 ) | ( x100 & n1475 ) | ( ~n1476 & n1475 ) ;
  assign n1478 = x100 | n1475 ;
  assign n1479 = ( n1471 & ~n1478 ) | ( n1471 & 1'b0 ) | ( ~n1478 & 1'b0 ) ;
  assign n1480 = n1477 | n1479 ;
  assign n1481 = ~n1470 & n1480 ;
  assign n1482 = n1468 | n1481 ;
  assign n1486 = ~x100 & n1283 ;
  assign n1487 = ( x101 & ~n1486 ) | ( x101 & 1'b0 ) | ( ~n1486 & 1'b0 ) ;
  assign n1488 = n1295 | n1487 ;
  assign n1483 = ( n1283 & ~x100 ) | ( n1283 & n1290 ) | ( ~x100 & n1290 ) ;
  assign n1484 = x100 &  n1483 ;
  assign n1485 = ( n1285 & ~n1290 ) | ( n1285 & n1484 ) | ( ~n1290 & n1484 ) ;
  assign n1489 = ( n1452 & n1485 ) | ( n1452 & n1488 ) | ( n1485 & n1488 ) ;
  assign n1491 = ~n1452 & n1489 ;
  assign n1490 = ( n1485 & ~n1489 ) | ( n1485 & 1'b0 ) | ( ~n1489 & 1'b0 ) ;
  assign n1492 = ( n1488 & ~n1491 ) | ( n1488 & n1490 ) | ( ~n1491 & n1490 ) ;
  assign n1493 = ( n976 & ~n1482 ) | ( n976 & n1492 ) | ( ~n1482 & n1492 ) ;
  assign n1494 = ( n837 & ~n1493 ) | ( n837 & 1'b0 ) | ( ~n1493 & 1'b0 ) ;
  assign n1495 = n1318 | n1321 ;
  assign n1496 = ( n1318 & n1304 ) | ( n1318 & n1495 ) | ( n1304 & n1495 ) ;
  assign n1498 = ( n1452 & ~n1318 ) | ( n1452 & n1496 ) | ( ~n1318 & n1496 ) ;
  assign n1497 = ( n1452 & ~n1496 ) | ( n1452 & n1495 ) | ( ~n1496 & n1495 ) ;
  assign n1499 = ( n1304 & ~n1498 ) | ( n1304 & n1497 ) | ( ~n1498 & n1497 ) ;
  assign n1500 = ( n976 & ~n1468 ) | ( n976 & 1'b0 ) | ( ~n1468 & 1'b0 ) ;
  assign n1501 = ~n1481 & n1500 ;
  assign n1502 = n1492 | n1501 ;
  assign n1503 = n1458 | n1466 ;
  assign n1504 = ( n1480 & ~n1122 ) | ( n1480 & n1503 ) | ( ~n1122 & n1503 ) ;
  assign n1505 = ~n976 & n1504 ;
  assign n1506 = n837 | n1505 ;
  assign n1507 = ( n1502 & ~n1506 ) | ( n1502 & 1'b0 ) | ( ~n1506 & 1'b0 ) ;
  assign n1508 = n1499 | n1507 ;
  assign n1509 = ~n1494 & n1508 ;
  assign n1510 = ~n1452 & n1323 ;
  assign n1511 = ( n1510 & ~n1306 ) | ( n1510 & n1452 ) | ( ~n1306 & n1452 ) ;
  assign n1512 = ( n1306 & n1316 ) | ( n1306 & n1511 ) | ( n1316 & n1511 ) ;
  assign n1513 = ( n1306 & ~n1316 ) | ( n1306 & n1511 ) | ( ~n1316 & n1511 ) ;
  assign n1514 = ( n1316 & ~n1512 ) | ( n1316 & n1513 ) | ( ~n1512 & n1513 ) ;
  assign n1515 = ( n1509 & ~n713 ) | ( n1509 & n1514 ) | ( ~n713 & n1514 ) ;
  assign n1516 = ( n595 & ~n1515 ) | ( n595 & 1'b0 ) | ( ~n1515 & 1'b0 ) ;
  assign n1517 = ~n1343 & n1452 ;
  assign n1518 = ( n1330 & n1339 ) | ( n1330 & n1343 ) | ( n1339 & n1343 ) ;
  assign n1520 = ( n1517 & ~n1343 ) | ( n1517 & n1518 ) | ( ~n1343 & n1518 ) ;
  assign n1519 = ( n1339 & ~n1518 ) | ( n1339 & n1517 ) | ( ~n1518 & n1517 ) ;
  assign n1521 = ( n1330 & ~n1520 ) | ( n1330 & n1519 ) | ( ~n1520 & n1519 ) ;
  assign n1522 = n713 | n1494 ;
  assign n1523 = ( n1508 & ~n1522 ) | ( n1508 & 1'b0 ) | ( ~n1522 & 1'b0 ) ;
  assign n1524 = n1514 | n1523 ;
  assign n1525 = ( n1502 & ~n1505 ) | ( n1502 & 1'b0 ) | ( ~n1505 & 1'b0 ) ;
  assign n1526 = ( n1499 & ~n837 ) | ( n1499 & n1525 ) | ( ~n837 & n1525 ) ;
  assign n1527 = ( n713 & ~n1526 ) | ( n713 & 1'b0 ) | ( ~n1526 & 1'b0 ) ;
  assign n1528 = n595 | n1527 ;
  assign n1529 = ( n1524 & ~n1528 ) | ( n1524 & 1'b0 ) | ( ~n1528 & 1'b0 ) ;
  assign n1530 = ( n1521 & ~n1529 ) | ( n1521 & 1'b0 ) | ( ~n1529 & 1'b0 ) ;
  assign n1531 = n1516 | n1530 ;
  assign n1537 = ( n492 & ~n1536 ) | ( n492 & n1531 ) | ( ~n1536 & n1531 ) ;
  assign n1538 = n396 &  n1537 ;
  assign n1540 = ( n1361 & ~n1352 ) | ( n1361 & n1365 ) | ( ~n1352 & n1365 ) ;
  assign n1539 = ~n1365 & n1452 ;
  assign n1541 = ( n1361 & ~n1540 ) | ( n1361 & n1539 ) | ( ~n1540 & n1539 ) ;
  assign n1542 = ( n1539 & ~n1365 ) | ( n1539 & n1540 ) | ( ~n1365 & n1540 ) ;
  assign n1543 = ( n1352 & ~n1541 ) | ( n1352 & n1542 ) | ( ~n1541 & n1542 ) ;
  assign n1544 = n492 | n1516 ;
  assign n1545 = n1530 | n1544 ;
  assign n1546 = ~n1536 & n1545 ;
  assign n1547 = ( n1524 & ~n1527 ) | ( n1524 & 1'b0 ) | ( ~n1527 & 1'b0 ) ;
  assign n1548 = ( n595 & ~n1547 ) | ( n595 & n1521 ) | ( ~n1547 & n1521 ) ;
  assign n1549 = n492 &  n1548 ;
  assign n1550 = n396 | n1549 ;
  assign n1551 = n1546 | n1550 ;
  assign n1552 = n1543 &  n1551 ;
  assign n1553 = n1538 | n1552 ;
  assign n1554 = ~n1354 & n1452 ;
  assign n1555 = ( n1354 & n1359 ) | ( n1354 & n1367 ) | ( n1359 & n1367 ) ;
  assign n1557 = ( n1554 & ~n1354 ) | ( n1554 & n1555 ) | ( ~n1354 & n1555 ) ;
  assign n1556 = ( n1367 & ~n1555 ) | ( n1367 & n1554 ) | ( ~n1555 & n1554 ) ;
  assign n1558 = ( n1359 & ~n1557 ) | ( n1359 & n1556 ) | ( ~n1557 & n1556 ) ;
  assign n1559 = ( n315 & n1553 ) | ( n315 & n1558 ) | ( n1553 & n1558 ) ;
  assign n1560 = n240 &  n1559 ;
  assign n1562 = ( n1383 & ~n1374 ) | ( n1383 & n1387 ) | ( ~n1374 & n1387 ) ;
  assign n1561 = ~n1387 & n1452 ;
  assign n1563 = ( n1383 & ~n1562 ) | ( n1383 & n1561 ) | ( ~n1562 & n1561 ) ;
  assign n1564 = ( n1561 & ~n1387 ) | ( n1561 & n1562 ) | ( ~n1387 & n1562 ) ;
  assign n1565 = ( n1374 & ~n1563 ) | ( n1374 & n1564 ) | ( ~n1563 & n1564 ) ;
  assign n1566 = n315 | n1538 ;
  assign n1567 = n1552 | n1566 ;
  assign n1568 = n1558 &  n1567 ;
  assign n1569 = n1546 | n1549 ;
  assign n1570 = ( n396 & n1543 ) | ( n396 & n1569 ) | ( n1543 & n1569 ) ;
  assign n1571 = n315 &  n1570 ;
  assign n1572 = n240 | n1571 ;
  assign n1573 = n1568 | n1572 ;
  assign n1574 = n1565 &  n1573 ;
  assign n1575 = n1560 | n1574 ;
  assign n1577 = ( n1376 & ~n1381 ) | ( n1376 & n1389 ) | ( ~n1381 & n1389 ) ;
  assign n1576 = ~n1376 & n1452 ;
  assign n1578 = ( n1389 & ~n1577 ) | ( n1389 & n1576 ) | ( ~n1577 & n1576 ) ;
  assign n1579 = ( n1576 & ~n1376 ) | ( n1576 & n1577 ) | ( ~n1376 & n1577 ) ;
  assign n1580 = ( n1381 & ~n1578 ) | ( n1381 & n1579 ) | ( ~n1578 & n1579 ) ;
  assign n1581 = ( n181 & n1575 ) | ( n181 & n1580 ) | ( n1575 & n1580 ) ;
  assign n1582 = ~n145 & n1581 ;
  assign n1583 = ~n1409 & n1452 ;
  assign n1584 = ( n1396 & n1405 ) | ( n1396 & n1409 ) | ( n1405 & n1409 ) ;
  assign n1586 = ( n1583 & ~n1409 ) | ( n1583 & n1584 ) | ( ~n1409 & n1584 ) ;
  assign n1585 = ( n1405 & ~n1584 ) | ( n1405 & n1583 ) | ( ~n1584 & n1583 ) ;
  assign n1587 = ( n1396 & ~n1586 ) | ( n1396 & n1585 ) | ( ~n1586 & n1585 ) ;
  assign n1588 = n181 | n1560 ;
  assign n1589 = n1574 | n1588 ;
  assign n1590 = n1580 &  n1589 ;
  assign n1591 = n1568 | n1571 ;
  assign n1592 = ( n240 & n1565 ) | ( n240 & n1591 ) | ( n1565 & n1591 ) ;
  assign n1593 = n181 &  n1592 ;
  assign n1594 = ( n145 & ~n1593 ) | ( n145 & 1'b0 ) | ( ~n1593 & 1'b0 ) ;
  assign n1595 = ~n1590 & n1594 ;
  assign n1596 = ( n1587 & ~n1595 ) | ( n1587 & 1'b0 ) | ( ~n1595 & 1'b0 ) ;
  assign n1597 = n1582 | n1596 ;
  assign n1603 = ( n150 & ~n1602 ) | ( n150 & n1597 ) | ( ~n1602 & n1597 ) ;
  assign n1604 = ~n1418 & n1434 ;
  assign n1605 = ( n1437 & ~n1452 ) | ( n1437 & n1604 ) | ( ~n1452 & n1604 ) ;
  assign n1606 = ~n1437 & n1605 ;
  assign n1607 = ( n1434 & ~n1437 ) | ( n1434 & 1'b0 ) | ( ~n1437 & 1'b0 ) ;
  assign n1608 = n1452 &  n1607 ;
  assign n1609 = ( n1418 & ~n1607 ) | ( n1418 & n1608 ) | ( ~n1607 & n1608 ) ;
  assign n1610 = n1606 | n1609 ;
  assign n1611 = ( n1419 & ~n1426 ) | ( n1419 & 1'b0 ) | ( ~n1426 & 1'b0 ) ;
  assign n1612 = n1452 &  n1611 ;
  assign n1613 = ( n1440 & ~n1612 ) | ( n1440 & n1611 ) | ( ~n1612 & n1611 ) ;
  assign n1614 = ( n1610 & ~n1613 ) | ( n1610 & 1'b0 ) | ( ~n1613 & 1'b0 ) ;
  assign n1615 = ~n1603 & n1614 ;
  assign n1616 = ( n133 & ~n1615 ) | ( n133 & n1614 ) | ( ~n1615 & n1614 ) ;
  assign n1617 = n150 | n1582 ;
  assign n1618 = n1596 | n1617 ;
  assign n1623 = n1618 | n1602 ;
  assign n1619 = n1590 | n1593 ;
  assign n1620 = ( n1587 & ~n145 ) | ( n1587 & n1619 ) | ( ~n145 & n1619 ) ;
  assign n1621 = n150 &  n1620 ;
  assign n1622 = n1610 | n1621 ;
  assign n1624 = ( n1623 & ~n1602 ) | ( n1623 & n1622 ) | ( ~n1602 & n1622 ) ;
  assign n1625 = ( n1419 & ~n1426 ) | ( n1419 & n1452 ) | ( ~n1426 & n1452 ) ;
  assign n1627 = n1426 | n1625 ;
  assign n1626 = ( n133 & ~n1426 ) | ( n133 & n1419 ) | ( ~n1426 & n1419 ) ;
  assign n1628 = ( n1426 & ~n1627 ) | ( n1426 & n1626 ) | ( ~n1627 & n1626 ) ;
  assign n1629 = n1422 | n1449 ;
  assign n1630 = ( n1425 & n1444 ) | ( n1425 & n1629 ) | ( n1444 & n1629 ) ;
  assign n1631 = ( n1425 & ~n1630 ) | ( n1425 & 1'b0 ) | ( ~n1630 & 1'b0 ) ;
  assign n1632 = ( n1432 & ~n1631 ) | ( n1432 & n1440 ) | ( ~n1631 & n1440 ) ;
  assign n1633 = ( n1432 & ~n1632 ) | ( n1432 & 1'b0 ) | ( ~n1632 & 1'b0 ) ;
  assign n1634 = n1628 | n1633 ;
  assign n1635 = ( n1624 & ~n1634 ) | ( n1624 & 1'b0 ) | ( ~n1634 & 1'b0 ) ;
  assign n1636 = n1616 &  n1635 ;
  assign n5673 = x62 | x63 ;
  assign n2707 = x82 | x83 ;
  assign n1723 = ( n1529 & ~n1636 ) | ( n1529 & 1'b0 ) | ( ~n1636 & 1'b0 ) ;
  assign n1724 = ( n1516 & ~n1636 ) | ( n1516 & n1521 ) | ( ~n1636 & n1521 ) ;
  assign n1725 = ( n1636 & ~n1723 ) | ( n1636 & n1724 ) | ( ~n1723 & n1724 ) ;
  assign n1726 = ( n1723 & ~n1516 ) | ( n1723 & n1724 ) | ( ~n1516 & n1724 ) ;
  assign n1727 = ( n1725 & ~n1521 ) | ( n1725 & n1726 ) | ( ~n1521 & n1726 ) ;
  assign n1708 = ~n1527 & n1636 ;
  assign n1709 = ( n1514 & ~n1527 ) | ( n1514 & n1523 ) | ( ~n1527 & n1523 ) ;
  assign n1710 = ( n1708 & ~n1523 ) | ( n1708 & n1709 ) | ( ~n1523 & n1709 ) ;
  assign n1711 = ( n1527 & ~n1708 ) | ( n1527 & n1709 ) | ( ~n1708 & n1709 ) ;
  assign n1712 = ( n1710 & ~n1514 ) | ( n1710 & n1711 ) | ( ~n1514 & n1711 ) ;
  assign n1701 = ~n1494 & n1636 ;
  assign n1702 = ( n1499 & ~n1494 ) | ( n1499 & n1507 ) | ( ~n1494 & n1507 ) ;
  assign n1703 = ( n1701 & ~n1507 ) | ( n1701 & n1702 ) | ( ~n1507 & n1702 ) ;
  assign n1704 = ( n1494 & ~n1701 ) | ( n1494 & n1702 ) | ( ~n1701 & n1702 ) ;
  assign n1705 = ( n1703 & ~n1499 ) | ( n1703 & n1704 ) | ( ~n1499 & n1704 ) ;
  assign n1686 = ~n1505 & n1636 ;
  assign n1687 = ( n1492 & ~n1501 ) | ( n1492 & n1505 ) | ( ~n1501 & n1505 ) ;
  assign n1688 = ( n1501 & ~n1686 ) | ( n1501 & n1687 ) | ( ~n1686 & n1687 ) ;
  assign n1689 = ( n1686 & ~n1505 ) | ( n1686 & n1687 ) | ( ~n1505 & n1687 ) ;
  assign n1690 = ( n1688 & ~n1492 ) | ( n1688 & n1689 ) | ( ~n1492 & n1689 ) ;
  assign n1679 = ( n1468 & ~n1470 ) | ( n1468 & 1'b0 ) | ( ~n1470 & 1'b0 ) ;
  assign n1680 = ( n1470 & ~n1679 ) | ( n1470 & n1480 ) | ( ~n1679 & n1480 ) ;
  assign n1681 = ( n1636 & ~n1470 ) | ( n1636 & n1680 ) | ( ~n1470 & n1680 ) ;
  assign n1682 = ( n1679 & ~n1636 ) | ( n1679 & n1680 ) | ( ~n1636 & n1680 ) ;
  assign n1683 = ( n1681 & ~n1480 ) | ( n1681 & n1682 ) | ( ~n1480 & n1682 ) ;
  assign n1660 = ( x98 & ~n1463 ) | ( x98 & n1452 ) | ( ~n1463 & n1452 ) ;
  assign n1661 = ( x98 & ~n1660 ) | ( x98 & 1'b0 ) | ( ~n1660 & 1'b0 ) ;
  assign n1662 = ( n1458 & ~n1661 ) | ( n1458 & n1463 ) | ( ~n1661 & n1463 ) ;
  assign n1663 = x98 | n1452 ;
  assign n1664 = x99 &  n1663 ;
  assign n1665 = ( n1471 & ~n1664 ) | ( n1471 & 1'b0 ) | ( ~n1664 & 1'b0 ) ;
  assign n1666 = ( n1662 & ~n1636 ) | ( n1662 & n1665 ) | ( ~n1636 & n1665 ) ;
  assign n1667 = ~n1662 & n1666 ;
  assign n1668 = n1636 | n1666 ;
  assign n1669 = ( n1667 & ~n1665 ) | ( n1667 & n1668 ) | ( ~n1665 & n1668 ) ;
  assign n1648 = n1455 | n1636 ;
  assign n1649 = n1452 | n1633 ;
  assign n1650 = ( n1624 & n1628 ) | ( n1624 & n1649 ) | ( n1628 & n1649 ) ;
  assign n1651 = ( n1624 & ~n1650 ) | ( n1624 & 1'b0 ) | ( ~n1650 & 1'b0 ) ;
  assign n1652 = n1616 &  n1651 ;
  assign n1653 = n1648 | n1652 ;
  assign n1654 = ( x98 & ~n1653 ) | ( x98 & n1652 ) | ( ~n1653 & n1652 ) ;
  assign n1655 = x98 | n1652 ;
  assign n1656 = ( n1648 & ~n1655 ) | ( n1648 & 1'b0 ) | ( ~n1655 & 1'b0 ) ;
  assign n1657 = n1654 | n1656 ;
  assign n1453 = x94 | x95 ;
  assign n1640 = ~x96 & n1453 ;
  assign n1641 = ( x96 & ~n1450 ) | ( x96 & n1640 ) | ( ~n1450 & n1640 ) ;
  assign n1642 = ( n1432 & ~n1641 ) | ( n1432 & n1440 ) | ( ~n1641 & n1440 ) ;
  assign n1643 = ( n1432 & ~n1642 ) | ( n1432 & 1'b0 ) | ( ~n1642 & 1'b0 ) ;
  assign n1644 = ( x97 & ~n1643 ) | ( x97 & n1636 ) | ( ~n1643 & n1636 ) ;
  assign n1639 = ( x96 & x97 ) | ( x96 & n1636 ) | ( x97 & n1636 ) ;
  assign n1645 = ( x96 & ~x97 ) | ( x96 & 1'b0 ) | ( ~x97 & 1'b0 ) ;
  assign n1646 = ( n1644 & ~n1639 ) | ( n1644 & n1645 ) | ( ~n1639 & n1645 ) ;
  assign n1637 = ( x96 & ~n1636 ) | ( x96 & 1'b0 ) | ( ~n1636 & 1'b0 ) ;
  assign n1454 = x96 | n1453 ;
  assign n1638 = ( n1452 & ~n1637 ) | ( n1452 & n1454 ) | ( ~n1637 & n1454 ) ;
  assign n1670 = ~n1283 & n1638 ;
  assign n1671 = ~n1646 & n1670 ;
  assign n1672 = ( n1657 & ~n1671 ) | ( n1657 & 1'b0 ) | ( ~n1671 & 1'b0 ) ;
  assign n1673 = n1638 | n1646 ;
  assign n1674 = ( n1283 & ~n1673 ) | ( n1283 & n1646 ) | ( ~n1673 & n1646 ) ;
  assign n1675 = ( n1122 & ~n1674 ) | ( n1122 & 1'b0 ) | ( ~n1674 & 1'b0 ) ;
  assign n1676 = ~n1672 & n1675 ;
  assign n1677 = n1669 | n1676 ;
  assign n1647 = ( n1638 & ~n1646 ) | ( n1638 & 1'b0 ) | ( ~n1646 & 1'b0 ) ;
  assign n1658 = ( n1283 & ~n1647 ) | ( n1283 & n1657 ) | ( ~n1647 & n1657 ) ;
  assign n1659 = ~n1122 & n1658 ;
  assign n1691 = ( n976 & ~n1659 ) | ( n976 & 1'b0 ) | ( ~n1659 & 1'b0 ) ;
  assign n1692 = n1677 &  n1691 ;
  assign n1693 = n1683 | n1692 ;
  assign n1694 = n1672 | n1674 ;
  assign n1695 = ( n1122 & ~n1694 ) | ( n1122 & n1669 ) | ( ~n1694 & n1669 ) ;
  assign n1696 = n976 | n1695 ;
  assign n1697 = ~n837 & n1696 ;
  assign n1698 = n1693 &  n1697 ;
  assign n1699 = ( n1690 & ~n1698 ) | ( n1690 & 1'b0 ) | ( ~n1698 & 1'b0 ) ;
  assign n1678 = ~n1659 & n1677 ;
  assign n1684 = ( n976 & n1678 ) | ( n976 & n1683 ) | ( n1678 & n1683 ) ;
  assign n1685 = ( n837 & ~n1684 ) | ( n837 & 1'b0 ) | ( ~n1684 & 1'b0 ) ;
  assign n1713 = n713 | n1685 ;
  assign n1714 = n1699 | n1713 ;
  assign n1715 = n1705 &  n1714 ;
  assign n1716 = n1693 &  n1696 ;
  assign n1717 = ( n837 & ~n1716 ) | ( n837 & n1690 ) | ( ~n1716 & n1690 ) ;
  assign n1718 = n713 &  n1717 ;
  assign n1738 = n1715 | n1718 ;
  assign n1739 = ( n595 & n1712 ) | ( n595 & n1738 ) | ( n1712 & n1738 ) ;
  assign n1740 = n492 &  n1739 ;
  assign n1719 = n595 | n1718 ;
  assign n1720 = n1715 | n1719 ;
  assign n1721 = n1712 &  n1720 ;
  assign n1700 = n1685 | n1699 ;
  assign n1706 = ( n713 & n1700 ) | ( n713 & n1705 ) | ( n1700 & n1705 ) ;
  assign n1707 = n595 &  n1706 ;
  assign n1735 = n492 | n1707 ;
  assign n1736 = n1721 | n1735 ;
  assign n1937 = ( n1736 & ~n1727 ) | ( n1736 & n1740 ) | ( ~n1727 & n1740 ) ;
  assign n1789 = ~n1582 & n1636 ;
  assign n1790 = ( n1587 & ~n1582 ) | ( n1587 & n1595 ) | ( ~n1582 & n1595 ) ;
  assign n1791 = ( n1789 & ~n1595 ) | ( n1789 & n1790 ) | ( ~n1595 & n1790 ) ;
  assign n1792 = ( n1582 & ~n1789 ) | ( n1582 & n1790 ) | ( ~n1789 & n1790 ) ;
  assign n1793 = ( n1791 & ~n1587 ) | ( n1791 & n1792 ) | ( ~n1587 & n1792 ) ;
  assign n1722 = n1707 | n1721 ;
  assign n1728 = ( n492 & ~n1727 ) | ( n492 & n1722 ) | ( ~n1727 & n1722 ) ;
  assign n1729 = n396 &  n1728 ;
  assign n1731 = ( n1545 & ~n1536 ) | ( n1545 & n1549 ) | ( ~n1536 & n1549 ) ;
  assign n1730 = ~n1549 & n1636 ;
  assign n1732 = ( n1545 & ~n1731 ) | ( n1545 & n1730 ) | ( ~n1731 & n1730 ) ;
  assign n1733 = ( n1730 & ~n1549 ) | ( n1730 & n1731 ) | ( ~n1549 & n1731 ) ;
  assign n1734 = ( n1536 & ~n1732 ) | ( n1536 & n1733 ) | ( ~n1732 & n1733 ) ;
  assign n1737 = ~n1727 & n1736 ;
  assign n1741 = n396 | n1740 ;
  assign n1742 = n1737 | n1741 ;
  assign n1743 = ~n1734 & n1742 ;
  assign n1744 = n1729 | n1743 ;
  assign n1745 = n1551 | n1636 ;
  assign n1746 = ( n1538 & ~n1636 ) | ( n1538 & n1543 ) | ( ~n1636 & n1543 ) ;
  assign n1747 = ( n1636 & n1745 ) | ( n1636 & n1746 ) | ( n1745 & n1746 ) ;
  assign n1748 = ( n1538 & ~n1746 ) | ( n1538 & n1745 ) | ( ~n1746 & n1745 ) ;
  assign n1749 = ( n1543 & ~n1747 ) | ( n1543 & n1748 ) | ( ~n1747 & n1748 ) ;
  assign n1750 = ( n315 & n1744 ) | ( n315 & n1749 ) | ( n1744 & n1749 ) ;
  assign n1751 = n240 &  n1750 ;
  assign n1753 = ( n1567 & ~n1558 ) | ( n1567 & n1571 ) | ( ~n1558 & n1571 ) ;
  assign n1752 = ~n1571 & n1636 ;
  assign n1754 = ( n1567 & ~n1753 ) | ( n1567 & n1752 ) | ( ~n1753 & n1752 ) ;
  assign n1755 = ( n1752 & ~n1571 ) | ( n1752 & n1753 ) | ( ~n1571 & n1753 ) ;
  assign n1756 = ( n1558 & ~n1754 ) | ( n1558 & n1755 ) | ( ~n1754 & n1755 ) ;
  assign n1757 = n315 | n1729 ;
  assign n1758 = n1743 | n1757 ;
  assign n1759 = n1749 &  n1758 ;
  assign n1760 = n1737 | n1740 ;
  assign n1761 = ( n396 & ~n1734 ) | ( n396 & n1760 ) | ( ~n1734 & n1760 ) ;
  assign n1762 = n315 &  n1761 ;
  assign n1763 = n240 | n1762 ;
  assign n1764 = n1759 | n1763 ;
  assign n1765 = n1756 &  n1764 ;
  assign n1766 = n1751 | n1765 ;
  assign n1767 = n1573 | n1636 ;
  assign n1768 = ( n1560 & ~n1636 ) | ( n1560 & n1565 ) | ( ~n1636 & n1565 ) ;
  assign n1769 = ( n1636 & n1767 ) | ( n1636 & n1768 ) | ( n1767 & n1768 ) ;
  assign n1770 = ( n1560 & ~n1768 ) | ( n1560 & n1767 ) | ( ~n1768 & n1767 ) ;
  assign n1771 = ( n1565 & ~n1769 ) | ( n1565 & n1770 ) | ( ~n1769 & n1770 ) ;
  assign n1772 = ( n181 & n1766 ) | ( n181 & n1771 ) | ( n1766 & n1771 ) ;
  assign n1773 = ~n145 & n1772 ;
  assign n1774 = ~n1593 & n1636 ;
  assign n1775 = ( n1580 & n1589 ) | ( n1580 & n1593 ) | ( n1589 & n1593 ) ;
  assign n1777 = ( n1774 & ~n1593 ) | ( n1774 & n1775 ) | ( ~n1593 & n1775 ) ;
  assign n1776 = ( n1589 & ~n1775 ) | ( n1589 & n1774 ) | ( ~n1775 & n1774 ) ;
  assign n1778 = ( n1580 & ~n1777 ) | ( n1580 & n1776 ) | ( ~n1777 & n1776 ) ;
  assign n1779 = n181 | n1751 ;
  assign n1780 = n1765 | n1779 ;
  assign n1781 = n1771 &  n1780 ;
  assign n1782 = n1759 | n1762 ;
  assign n1783 = ( n240 & n1756 ) | ( n240 & n1782 ) | ( n1756 & n1782 ) ;
  assign n1784 = n181 &  n1783 ;
  assign n1785 = ( n145 & ~n1784 ) | ( n145 & 1'b0 ) | ( ~n1784 & 1'b0 ) ;
  assign n1786 = ~n1781 & n1785 ;
  assign n1787 = ( n1778 & ~n1786 ) | ( n1778 & 1'b0 ) | ( ~n1786 & 1'b0 ) ;
  assign n1788 = n1773 | n1787 ;
  assign n1794 = ( n150 & ~n1793 ) | ( n150 & n1788 ) | ( ~n1793 & n1788 ) ;
  assign n1795 = ( n1602 & ~n1621 ) | ( n1602 & 1'b0 ) | ( ~n1621 & 1'b0 ) ;
  assign n1796 = ( n1618 & ~n1795 ) | ( n1618 & n1636 ) | ( ~n1795 & n1636 ) ;
  assign n1797 = ( n1618 & ~n1796 ) | ( n1618 & 1'b0 ) | ( ~n1796 & 1'b0 ) ;
  assign n1798 = ( n1618 & ~n1621 ) | ( n1618 & 1'b0 ) | ( ~n1621 & 1'b0 ) ;
  assign n1799 = n1636 &  n1798 ;
  assign n1800 = ( n1602 & ~n1799 ) | ( n1602 & n1798 ) | ( ~n1799 & n1798 ) ;
  assign n1801 = ~n1797 & n1800 ;
  assign n1802 = n1603 &  n1610 ;
  assign n1803 = n1636 &  n1802 ;
  assign n1804 = ( n1624 & ~n1802 ) | ( n1624 & n1803 ) | ( ~n1802 & n1803 ) ;
  assign n1805 = ~n1801 & n1804 ;
  assign n1806 = ~n1794 & n1805 ;
  assign n1807 = ( n133 & ~n1806 ) | ( n133 & n1805 ) | ( ~n1806 & n1805 ) ;
  assign n1808 = n150 | n1773 ;
  assign n1809 = n1787 | n1808 ;
  assign n1814 = n1793 | n1809 ;
  assign n1810 = n1781 | n1784 ;
  assign n1811 = ( n1778 & ~n145 ) | ( n1778 & n1810 ) | ( ~n145 & n1810 ) ;
  assign n1812 = n150 &  n1811 ;
  assign n1813 = ( n1801 & ~n1812 ) | ( n1801 & 1'b0 ) | ( ~n1812 & 1'b0 ) ;
  assign n1815 = ( n1793 & ~n1814 ) | ( n1793 & n1813 ) | ( ~n1814 & n1813 ) ;
  assign n1817 = ( n133 & n1603 ) | ( n133 & n1610 ) | ( n1603 & n1610 ) ;
  assign n1816 = ( n1603 & n1610 ) | ( n1603 & n1636 ) | ( n1610 & n1636 ) ;
  assign n1818 = ( n1610 & ~n1816 ) | ( n1610 & 1'b0 ) | ( ~n1816 & 1'b0 ) ;
  assign n1819 = ( n1817 & ~n1610 ) | ( n1817 & n1818 ) | ( ~n1610 & n1818 ) ;
  assign n1820 = n1606 | n1633 ;
  assign n1821 = ( n1628 & ~n1609 ) | ( n1628 & n1820 ) | ( ~n1609 & n1820 ) ;
  assign n1822 = n1609 | n1821 ;
  assign n1823 = ( n1616 & ~n1624 ) | ( n1616 & n1822 ) | ( ~n1624 & n1822 ) ;
  assign n1824 = ( n1616 & ~n1823 ) | ( n1616 & 1'b0 ) | ( ~n1823 & 1'b0 ) ;
  assign n1825 = n1819 | n1824 ;
  assign n1826 = n1815 | n1825 ;
  assign n1827 = ~n1807 |  n1826 ;
  assign n1936 = n1740 | n1827 ;
  assign n1939 = ( n1740 & ~n1937 ) | ( n1740 & n1936 ) | ( ~n1937 & n1936 ) ;
  assign n1938 = ( n1936 & ~n1736 ) | ( n1936 & n1937 ) | ( ~n1736 & n1937 ) ;
  assign n1940 = ( n1727 & ~n1939 ) | ( n1727 & n1938 ) | ( ~n1939 & n1938 ) ;
  assign n2001 = n1793 &  n1809 ;
  assign n2002 = ( n1812 & n1827 ) | ( n1812 & n2001 ) | ( n1827 & n2001 ) ;
  assign n2003 = ~n1812 & n2002 ;
  assign n2004 = ( n1809 & ~n1812 ) | ( n1809 & 1'b0 ) | ( ~n1812 & 1'b0 ) ;
  assign n2005 = ~n1827 & n2004 ;
  assign n2006 = ( n1793 & ~n2005 ) | ( n1793 & n2004 ) | ( ~n2005 & n2004 ) ;
  assign n2007 = ~n2003 & n2006 ;
  assign n2008 = ( n1794 & ~n1801 ) | ( n1794 & 1'b0 ) | ( ~n1801 & 1'b0 ) ;
  assign n2009 = ~n1827 & n2008 ;
  assign n2010 = ( n1815 & ~n2009 ) | ( n1815 & n2008 ) | ( ~n2009 & n2008 ) ;
  assign n2011 = n2007 | n2010 ;
  assign n1951 = ~n1742 & n1827 ;
  assign n1952 = ( n1729 & n1734 ) | ( n1729 & n1827 ) | ( n1734 & n1827 ) ;
  assign n1954 = ( n1951 & ~n1729 ) | ( n1951 & n1952 ) | ( ~n1729 & n1952 ) ;
  assign n1953 = ( n1827 & ~n1952 ) | ( n1827 & n1951 ) | ( ~n1952 & n1951 ) ;
  assign n1955 = ( n1734 & ~n1954 ) | ( n1734 & n1953 ) | ( ~n1954 & n1953 ) ;
  assign n1832 = x94 &  n1827 ;
  assign n1830 = x92 | x93 ;
  assign n1831 = x94 | n1830 ;
  assign n1833 = ( n1636 & ~n1832 ) | ( n1636 & n1831 ) | ( ~n1832 & n1831 ) ;
  assign n1834 = ( x94 & ~n1827 ) | ( x94 & x95 ) | ( ~n1827 & x95 ) ;
  assign n1840 = ( x94 & ~x95 ) | ( x94 & 1'b0 ) | ( ~x95 & 1'b0 ) ;
  assign n1835 = ~x94 & n1830 ;
  assign n1836 = ( x94 & ~n1634 ) | ( x94 & n1835 ) | ( ~n1634 & n1835 ) ;
  assign n1837 = ( n1624 & ~n1616 ) | ( n1624 & n1836 ) | ( ~n1616 & n1836 ) ;
  assign n1838 = n1616 &  n1837 ;
  assign n1839 = ( n1827 & ~x95 ) | ( n1827 & n1838 ) | ( ~x95 & n1838 ) ;
  assign n1841 = ( n1834 & ~n1840 ) | ( n1834 & n1839 ) | ( ~n1840 & n1839 ) ;
  assign n1842 = ~n1833 & n1841 ;
  assign n1843 = ( n1452 & ~n1842 ) | ( n1452 & n1841 ) | ( ~n1842 & n1841 ) ;
  assign n1844 = n1452 &  n1833 ;
  assign n1845 = n1841 &  n1844 ;
  assign n1847 = n1636 | n1824 ;
  assign n1848 = ( n1819 & ~n1815 ) | ( n1819 & n1847 ) | ( ~n1815 & n1847 ) ;
  assign n1849 = n1815 | n1848 ;
  assign n1850 = ( n1807 & ~n1849 ) | ( n1807 & 1'b0 ) | ( ~n1849 & 1'b0 ) ;
  assign n1846 = ~n1453 & n1827 ;
  assign n1851 = ~n1850 & n1846 ;
  assign n1852 = ( x96 & n1851 ) | ( x96 & n1850 ) | ( n1851 & n1850 ) ;
  assign n1853 = x96 | n1850 ;
  assign n1854 = n1846 | n1853 ;
  assign n1855 = ~n1852 & n1854 ;
  assign n1856 = n1845 | n1855 ;
  assign n1857 = n1843 &  n1856 ;
  assign n1858 = x96 | n1636 ;
  assign n1859 = x97 | n1858 ;
  assign n1860 = x97 &  n1858 ;
  assign n1861 = ( n1859 & ~n1860 ) | ( n1859 & 1'b0 ) | ( ~n1860 & 1'b0 ) ;
  assign n1863 = ( n1638 & ~n1827 ) | ( n1638 & 1'b0 ) | ( ~n1827 & 1'b0 ) ;
  assign n1862 = ~n1637 & n1643 ;
  assign n1864 = ( n1638 & n1861 ) | ( n1638 & n1862 ) | ( n1861 & n1862 ) ;
  assign n1865 = ( n1863 & ~n1862 ) | ( n1863 & n1864 ) | ( ~n1862 & n1864 ) ;
  assign n1866 = ( n1638 & ~n1864 ) | ( n1638 & n1863 ) | ( ~n1864 & n1863 ) ;
  assign n1867 = ( n1861 & ~n1865 ) | ( n1861 & n1866 ) | ( ~n1865 & n1866 ) ;
  assign n1868 = ( n1283 & ~n1857 ) | ( n1283 & n1867 ) | ( ~n1857 & n1867 ) ;
  assign n1869 = ~n1122 & n1868 ;
  assign n1870 = ~n1671 & n1674 ;
  assign n1871 = ( n1657 & ~n1671 ) | ( n1657 & n1870 ) | ( ~n1671 & n1870 ) ;
  assign n1873 = ( n1671 & n1827 ) | ( n1671 & n1871 ) | ( n1827 & n1871 ) ;
  assign n1872 = ( n1827 & ~n1871 ) | ( n1827 & n1870 ) | ( ~n1871 & n1870 ) ;
  assign n1874 = ( n1657 & ~n1873 ) | ( n1657 & n1872 ) | ( ~n1873 & n1872 ) ;
  assign n1875 = ~n1283 & n1843 ;
  assign n1876 = n1856 &  n1875 ;
  assign n1877 = ( n1867 & ~n1876 ) | ( n1867 & 1'b0 ) | ( ~n1876 & 1'b0 ) ;
  assign n1878 = n1833 &  n1841 ;
  assign n1879 = ( n1452 & n1855 ) | ( n1452 & n1878 ) | ( n1855 & n1878 ) ;
  assign n1880 = ( n1283 & ~n1879 ) | ( n1283 & 1'b0 ) | ( ~n1879 & 1'b0 ) ;
  assign n1881 = ( n1122 & ~n1880 ) | ( n1122 & 1'b0 ) | ( ~n1880 & 1'b0 ) ;
  assign n1882 = ~n1877 & n1881 ;
  assign n1883 = ( n1874 & ~n1882 ) | ( n1874 & 1'b0 ) | ( ~n1882 & 1'b0 ) ;
  assign n1884 = n1869 | n1883 ;
  assign n1885 = n1659 | n1827 ;
  assign n1886 = ( n1669 & ~n1659 ) | ( n1669 & n1676 ) | ( ~n1659 & n1676 ) ;
  assign n1888 = ( n1659 & n1885 ) | ( n1659 & n1886 ) | ( n1885 & n1886 ) ;
  assign n1887 = ( n1676 & ~n1886 ) | ( n1676 & n1885 ) | ( ~n1886 & n1885 ) ;
  assign n1889 = ( n1669 & ~n1888 ) | ( n1669 & n1887 ) | ( ~n1888 & n1887 ) ;
  assign n1890 = ( n976 & ~n1884 ) | ( n976 & n1889 ) | ( ~n1884 & n1889 ) ;
  assign n1891 = ( n837 & ~n1890 ) | ( n837 & 1'b0 ) | ( ~n1890 & 1'b0 ) ;
  assign n1892 = ( n1696 & ~n1827 ) | ( n1696 & 1'b0 ) | ( ~n1827 & 1'b0 ) ;
  assign n1893 = ( n1683 & n1692 ) | ( n1683 & n1696 ) | ( n1692 & n1696 ) ;
  assign n1894 = ( n1892 & ~n1692 ) | ( n1892 & n1893 ) | ( ~n1692 & n1893 ) ;
  assign n1895 = ( n1696 & ~n1893 ) | ( n1696 & n1892 ) | ( ~n1893 & n1892 ) ;
  assign n1896 = ( n1683 & ~n1894 ) | ( n1683 & n1895 ) | ( ~n1894 & n1895 ) ;
  assign n1897 = ( n976 & ~n1869 ) | ( n976 & 1'b0 ) | ( ~n1869 & 1'b0 ) ;
  assign n1898 = ~n1883 & n1897 ;
  assign n1899 = n1889 | n1898 ;
  assign n1900 = n1877 | n1880 ;
  assign n1901 = ( n1874 & ~n1122 ) | ( n1874 & n1900 ) | ( ~n1122 & n1900 ) ;
  assign n1902 = ~n976 & n1901 ;
  assign n1903 = n837 | n1902 ;
  assign n1904 = ( n1899 & ~n1903 ) | ( n1899 & 1'b0 ) | ( ~n1903 & 1'b0 ) ;
  assign n1905 = n1896 | n1904 ;
  assign n1906 = ~n1891 & n1905 ;
  assign n1907 = n1698 &  n1827 ;
  assign n1908 = ( n1685 & n1690 ) | ( n1685 & n1827 ) | ( n1690 & n1827 ) ;
  assign n1910 = ( n1907 & ~n1685 ) | ( n1907 & n1908 ) | ( ~n1685 & n1908 ) ;
  assign n1909 = ( n1827 & ~n1908 ) | ( n1827 & n1907 ) | ( ~n1908 & n1907 ) ;
  assign n1911 = ( n1690 & ~n1910 ) | ( n1690 & n1909 ) | ( ~n1910 & n1909 ) ;
  assign n1912 = ( n713 & ~n1906 ) | ( n713 & n1911 ) | ( ~n1906 & n1911 ) ;
  assign n1913 = n595 &  n1912 ;
  assign n1915 = ( n1714 & ~n1705 ) | ( n1714 & n1718 ) | ( ~n1705 & n1718 ) ;
  assign n1914 = n1718 | n1827 ;
  assign n1917 = ( n1718 & ~n1915 ) | ( n1718 & n1914 ) | ( ~n1915 & n1914 ) ;
  assign n1916 = ( n1914 & ~n1714 ) | ( n1914 & n1915 ) | ( ~n1714 & n1915 ) ;
  assign n1918 = ( n1705 & ~n1917 ) | ( n1705 & n1916 ) | ( ~n1917 & n1916 ) ;
  assign n1919 = n713 | n1891 ;
  assign n1920 = ( n1905 & ~n1919 ) | ( n1905 & 1'b0 ) | ( ~n1919 & 1'b0 ) ;
  assign n1921 = ( n1911 & ~n1920 ) | ( n1911 & 1'b0 ) | ( ~n1920 & 1'b0 ) ;
  assign n1922 = ( n1899 & ~n1902 ) | ( n1899 & 1'b0 ) | ( ~n1902 & 1'b0 ) ;
  assign n1923 = ( n1896 & ~n837 ) | ( n1896 & n1922 ) | ( ~n837 & n1922 ) ;
  assign n1924 = ( n713 & ~n1923 ) | ( n713 & 1'b0 ) | ( ~n1923 & 1'b0 ) ;
  assign n1925 = n595 | n1924 ;
  assign n1926 = n1921 | n1925 ;
  assign n1927 = n1918 &  n1926 ;
  assign n1928 = n1913 | n1927 ;
  assign n1929 = n1707 | n1827 ;
  assign n1930 = ( n1707 & n1712 ) | ( n1707 & n1720 ) | ( n1712 & n1720 ) ;
  assign n1931 = ( n1929 & ~n1720 ) | ( n1929 & n1930 ) | ( ~n1720 & n1930 ) ;
  assign n1932 = ( n1707 & ~n1930 ) | ( n1707 & n1929 ) | ( ~n1930 & n1929 ) ;
  assign n1933 = ( n1712 & ~n1931 ) | ( n1712 & n1932 ) | ( ~n1931 & n1932 ) ;
  assign n1934 = ( n492 & n1928 ) | ( n492 & n1933 ) | ( n1928 & n1933 ) ;
  assign n1935 = n396 &  n1934 ;
  assign n1941 = n492 | n1913 ;
  assign n1942 = n1927 | n1941 ;
  assign n1943 = n1933 &  n1942 ;
  assign n1944 = n1921 | n1924 ;
  assign n1945 = ( n595 & n1918 ) | ( n595 & n1944 ) | ( n1918 & n1944 ) ;
  assign n1946 = n492 &  n1945 ;
  assign n1947 = n396 | n1946 ;
  assign n1948 = n1943 | n1947 ;
  assign n1949 = ~n1940 & n1948 ;
  assign n1950 = n1935 | n1949 ;
  assign n1956 = ( n315 & ~n1955 ) | ( n315 & n1950 ) | ( ~n1955 & n1950 ) ;
  assign n1957 = n240 &  n1956 ;
  assign n1958 = n1762 | n1827 ;
  assign n1959 = ( n1749 & n1758 ) | ( n1749 & n1762 ) | ( n1758 & n1762 ) ;
  assign n1960 = ( n1958 & ~n1758 ) | ( n1958 & n1959 ) | ( ~n1758 & n1959 ) ;
  assign n1961 = ( n1762 & ~n1959 ) | ( n1762 & n1958 ) | ( ~n1959 & n1958 ) ;
  assign n1962 = ( n1749 & ~n1960 ) | ( n1749 & n1961 ) | ( ~n1960 & n1961 ) ;
  assign n1963 = n315 | n1935 ;
  assign n1964 = n1949 | n1963 ;
  assign n1965 = ~n1955 & n1964 ;
  assign n1966 = n1943 | n1946 ;
  assign n1967 = ( n396 & ~n1940 ) | ( n396 & n1966 ) | ( ~n1940 & n1966 ) ;
  assign n1968 = n315 &  n1967 ;
  assign n1969 = n240 | n1968 ;
  assign n1970 = n1965 | n1969 ;
  assign n1971 = n1962 &  n1970 ;
  assign n1972 = n1957 | n1971 ;
  assign n1973 = ~n1764 & n1827 ;
  assign n1974 = ( n1751 & ~n1973 ) | ( n1751 & n1827 ) | ( ~n1973 & n1827 ) ;
  assign n1975 = ( n1751 & ~n1974 ) | ( n1751 & n1756 ) | ( ~n1974 & n1756 ) ;
  assign n1976 = ( n1756 & ~n1751 ) | ( n1756 & n1974 ) | ( ~n1751 & n1974 ) ;
  assign n1977 = ( n1975 & ~n1756 ) | ( n1975 & n1976 ) | ( ~n1756 & n1976 ) ;
  assign n1978 = ( n181 & n1972 ) | ( n181 & n1977 ) | ( n1972 & n1977 ) ;
  assign n1979 = ~n145 & n1978 ;
  assign n1981 = ( n1780 & ~n1771 ) | ( n1780 & n1784 ) | ( ~n1771 & n1784 ) ;
  assign n1980 = n1784 | n1827 ;
  assign n1983 = ( n1784 & ~n1981 ) | ( n1784 & n1980 ) | ( ~n1981 & n1980 ) ;
  assign n1982 = ( n1980 & ~n1780 ) | ( n1980 & n1981 ) | ( ~n1780 & n1981 ) ;
  assign n1984 = ( n1771 & ~n1983 ) | ( n1771 & n1982 ) | ( ~n1983 & n1982 ) ;
  assign n1985 = n181 | n1957 ;
  assign n1986 = n1971 | n1985 ;
  assign n1987 = n1977 &  n1986 ;
  assign n1988 = n1965 | n1968 ;
  assign n1989 = ( n240 & n1962 ) | ( n240 & n1988 ) | ( n1962 & n1988 ) ;
  assign n1990 = n181 &  n1989 ;
  assign n1991 = ( n145 & ~n1990 ) | ( n145 & 1'b0 ) | ( ~n1990 & 1'b0 ) ;
  assign n1992 = ~n1987 & n1991 ;
  assign n1993 = ( n1984 & ~n1992 ) | ( n1984 & 1'b0 ) | ( ~n1992 & 1'b0 ) ;
  assign n1994 = n1979 | n1993 ;
  assign n1995 = n1773 | n1827 ;
  assign n1996 = ( n1778 & ~n1773 ) | ( n1778 & n1786 ) | ( ~n1773 & n1786 ) ;
  assign n1998 = ( n1773 & n1995 ) | ( n1773 & n1996 ) | ( n1995 & n1996 ) ;
  assign n1997 = ( n1786 & ~n1996 ) | ( n1786 & n1995 ) | ( ~n1996 & n1995 ) ;
  assign n1999 = ( n1778 & ~n1998 ) | ( n1778 & n1997 ) | ( ~n1998 & n1997 ) ;
  assign n2000 = ( n150 & n1994 ) | ( n150 & n1999 ) | ( n1994 & n1999 ) ;
  assign n2012 = n2000 | n2011 ;
  assign n2013 = ( n133 & ~n2011 ) | ( n133 & n2012 ) | ( ~n2011 & n2012 ) ;
  assign n2014 = n150 | n1979 ;
  assign n2015 = n1993 | n2014 ;
  assign n2020 = ~n2015 & n1999 ;
  assign n2016 = n1987 | n1990 ;
  assign n2017 = ( n1984 & ~n145 ) | ( n1984 & n2016 ) | ( ~n145 & n2016 ) ;
  assign n2018 = n150 &  n2017 ;
  assign n2019 = ( n2007 & ~n2018 ) | ( n2007 & 1'b0 ) | ( ~n2018 & 1'b0 ) ;
  assign n2021 = ( n2020 & ~n1999 ) | ( n2020 & n2019 ) | ( ~n1999 & n2019 ) ;
  assign n2023 = ( n133 & ~n1801 ) | ( n133 & n1794 ) | ( ~n1801 & n1794 ) ;
  assign n2022 = ( n1801 & ~n1794 ) | ( n1801 & n1827 ) | ( ~n1794 & n1827 ) ;
  assign n2024 = ~n1801 & n2022 ;
  assign n2025 = ( n1801 & n2023 ) | ( n1801 & n2024 ) | ( n2023 & n2024 ) ;
  assign n2026 = n1797 | n1824 ;
  assign n2027 = ( n1800 & n1819 ) | ( n1800 & n2026 ) | ( n1819 & n2026 ) ;
  assign n2028 = ( n1800 & ~n2027 ) | ( n1800 & 1'b0 ) | ( ~n2027 & 1'b0 ) ;
  assign n2029 = ( n1807 & ~n2028 ) | ( n1807 & n1815 ) | ( ~n2028 & n1815 ) ;
  assign n2030 = ( n1807 & ~n2029 ) | ( n1807 & 1'b0 ) | ( ~n2029 & 1'b0 ) ;
  assign n2031 = n2025 | n2030 ;
  assign n2032 = n2021 | n2031 ;
  assign n2033 = n2013 &  ~n2032 ;
  assign n2163 = n1948 | n2033 ;
  assign n2164 = ( n1935 & ~n2033 ) | ( n1935 & n1940 ) | ( ~n2033 & n1940 ) ;
  assign n2165 = ( n2033 & n2163 ) | ( n2033 & n2164 ) | ( n2163 & n2164 ) ;
  assign n2166 = ( n1935 & ~n2164 ) | ( n1935 & n2163 ) | ( ~n2164 & n2163 ) ;
  assign n2167 = ( n1940 & ~n2165 ) | ( n1940 & n2166 ) | ( ~n2165 & n2166 ) ;
  assign n2149 = ( n1942 & ~n1933 ) | ( n1942 & n1946 ) | ( ~n1933 & n1946 ) ;
  assign n2148 = ~n1946 & n2033 ;
  assign n2150 = ( n1942 & ~n2149 ) | ( n1942 & n2148 ) | ( ~n2149 & n2148 ) ;
  assign n2151 = ( n2148 & ~n1946 ) | ( n2148 & n2149 ) | ( ~n1946 & n2149 ) ;
  assign n2152 = ( n1933 & ~n2150 ) | ( n1933 & n2151 ) | ( ~n2150 & n2151 ) ;
  assign n2141 = n1926 | n2033 ;
  assign n2142 = ( n1918 & ~n1913 ) | ( n1918 & n2033 ) | ( ~n1913 & n2033 ) ;
  assign n2144 = ( n1913 & n2141 ) | ( n1913 & n2142 ) | ( n2141 & n2142 ) ;
  assign n2143 = ( n2033 & ~n2142 ) | ( n2033 & n2141 ) | ( ~n2142 & n2141 ) ;
  assign n2145 = ( n1918 & ~n2144 ) | ( n1918 & n2143 ) | ( ~n2144 & n2143 ) ;
  assign n2126 = ~n1924 & n2033 ;
  assign n2127 = ( n1911 & ~n1920 ) | ( n1911 & n1924 ) | ( ~n1920 & n1924 ) ;
  assign n2128 = ( n1920 & ~n2126 ) | ( n1920 & n2127 ) | ( ~n2126 & n2127 ) ;
  assign n2129 = ( n2126 & ~n1924 ) | ( n2126 & n2127 ) | ( ~n1924 & n2127 ) ;
  assign n2130 = ( n2128 & ~n1911 ) | ( n2128 & n2129 ) | ( ~n1911 & n2129 ) ;
  assign n2119 = ( n1904 & ~n2033 ) | ( n1904 & 1'b0 ) | ( ~n2033 & 1'b0 ) ;
  assign n2120 = ( n2033 & ~n1891 ) | ( n2033 & n2119 ) | ( ~n1891 & n2119 ) ;
  assign n2122 = ( n1891 & n1896 ) | ( n1891 & n2120 ) | ( n1896 & n2120 ) ;
  assign n2121 = ( n1891 & ~n1896 ) | ( n1891 & n2120 ) | ( ~n1896 & n2120 ) ;
  assign n2123 = ( n1896 & ~n2122 ) | ( n1896 & n2121 ) | ( ~n2122 & n2121 ) ;
  assign n2104 = ~n1902 & n2033 ;
  assign n2105 = ( n1889 & ~n1898 ) | ( n1889 & n1902 ) | ( ~n1898 & n1902 ) ;
  assign n2106 = ( n1898 & ~n2104 ) | ( n1898 & n2105 ) | ( ~n2104 & n2105 ) ;
  assign n2107 = ( n2104 & ~n1902 ) | ( n2104 & n2105 ) | ( ~n1902 & n2105 ) ;
  assign n2108 = ( n2106 & ~n1889 ) | ( n2106 & n2107 ) | ( ~n1889 & n2107 ) ;
  assign n2097 = ~n2033 & n1882 ;
  assign n2098 = ( n2097 & ~n1869 ) | ( n2097 & n2033 ) | ( ~n1869 & n2033 ) ;
  assign n2099 = ( n1869 & n1874 ) | ( n1869 & n2098 ) | ( n1874 & n2098 ) ;
  assign n2100 = ( n1869 & ~n1874 ) | ( n1869 & n2098 ) | ( ~n1874 & n2098 ) ;
  assign n2101 = ( n1874 & ~n2099 ) | ( n1874 & n2100 ) | ( ~n2099 & n2100 ) ;
  assign n2076 = n1843 | n1845 ;
  assign n2077 = ( n1845 & n1855 ) | ( n1845 & n2076 ) | ( n1855 & n2076 ) ;
  assign n2078 = ( n2033 & ~n1845 ) | ( n2033 & n2077 ) | ( ~n1845 & n2077 ) ;
  assign n2079 = ( n2033 & ~n2077 ) | ( n2033 & n2076 ) | ( ~n2077 & n2076 ) ;
  assign n2080 = ( n1855 & ~n2078 ) | ( n1855 & n2079 ) | ( ~n2078 & n2079 ) ;
  assign n2060 = ~x94 & n1827 ;
  assign n2061 = ( x95 & ~n2060 ) | ( x95 & 1'b0 ) | ( ~n2060 & 1'b0 ) ;
  assign n2062 = n1846 | n2061 ;
  assign n2057 = ( n1827 & ~x94 ) | ( n1827 & n1838 ) | ( ~x94 & n1838 ) ;
  assign n2058 = x94 &  n2057 ;
  assign n2059 = ( n1833 & ~n1838 ) | ( n1833 & n2058 ) | ( ~n1838 & n2058 ) ;
  assign n2063 = ( n2033 & n2059 ) | ( n2033 & n2062 ) | ( n2059 & n2062 ) ;
  assign n2065 = ~n2033 & n2063 ;
  assign n2064 = ( n2059 & ~n2063 ) | ( n2059 & 1'b0 ) | ( ~n2063 & 1'b0 ) ;
  assign n2066 = ( n2062 & ~n2065 ) | ( n2062 & n2064 ) | ( ~n2065 & n2064 ) ;
  assign n2045 = n1830 | n2033 ;
  assign n2046 = ( n1827 & ~n2030 ) | ( n1827 & 1'b0 ) | ( ~n2030 & 1'b0 ) ;
  assign n2047 = ( n2021 & ~n2025 ) | ( n2021 & n2046 ) | ( ~n2025 & n2046 ) ;
  assign n2048 = ~n2021 & n2047 ;
  assign n2049 = n2013 &  n2048 ;
  assign n2050 = n2045 | n2049 ;
  assign n2051 = ( x94 & ~n2050 ) | ( x94 & n2049 ) | ( ~n2050 & n2049 ) ;
  assign n2052 = x94 | n2049 ;
  assign n2053 = ( n2045 & ~n2052 ) | ( n2045 & 1'b0 ) | ( ~n2052 & 1'b0 ) ;
  assign n2054 = n2051 | n2053 ;
  assign n1828 = x90 | x91 ;
  assign n2037 = ~x92 & n1828 ;
  assign n2038 = ( x92 & ~n1825 ) | ( x92 & n2037 ) | ( ~n1825 & n2037 ) ;
  assign n2039 = ( n1807 & ~n2038 ) | ( n1807 & n1815 ) | ( ~n2038 & n1815 ) ;
  assign n2040 = ( n1807 & ~n2039 ) | ( n1807 & 1'b0 ) | ( ~n2039 & 1'b0 ) ;
  assign n2041 = ( x93 & ~n2040 ) | ( x93 & n2033 ) | ( ~n2040 & n2033 ) ;
  assign n2036 = ( x92 & x93 ) | ( x92 & n2033 ) | ( x93 & n2033 ) ;
  assign n2042 = ( x92 & ~x93 ) | ( x92 & 1'b0 ) | ( ~x93 & 1'b0 ) ;
  assign n2043 = ( n2041 & ~n2036 ) | ( n2041 & n2042 ) | ( ~n2036 & n2042 ) ;
  assign n1829 = x92 | n1828 ;
  assign n2034 = ( x92 & ~n2033 ) | ( x92 & 1'b0 ) | ( ~n2033 & 1'b0 ) ;
  assign n2035 = ( n1827 & ~n1829 ) | ( n1827 & n2034 ) | ( ~n1829 & n2034 ) ;
  assign n2067 = ( n1636 & ~n2035 ) | ( n1636 & 1'b0 ) | ( ~n2035 & 1'b0 ) ;
  assign n2068 = ~n2043 & n2067 ;
  assign n2069 = ( n2054 & ~n2068 ) | ( n2054 & 1'b0 ) | ( ~n2068 & 1'b0 ) ;
  assign n2070 = ~n2043 & n2035 ;
  assign n2071 = ( n2070 & ~n1636 ) | ( n2070 & n2043 ) | ( ~n1636 & n2043 ) ;
  assign n2072 = ( n1452 & ~n2071 ) | ( n1452 & 1'b0 ) | ( ~n2071 & 1'b0 ) ;
  assign n2073 = ~n2069 & n2072 ;
  assign n2074 = n2066 | n2073 ;
  assign n2044 = n2035 | n2043 ;
  assign n2055 = ( n2044 & ~n1636 ) | ( n2044 & n2054 ) | ( ~n1636 & n2054 ) ;
  assign n2056 = ~n1452 & n2055 ;
  assign n2083 = n1283 | n2056 ;
  assign n2084 = ( n2074 & ~n2083 ) | ( n2074 & 1'b0 ) | ( ~n2083 & 1'b0 ) ;
  assign n2085 = n2080 | n2084 ;
  assign n2086 = n2069 | n2071 ;
  assign n2087 = ( n1452 & ~n2086 ) | ( n1452 & n2066 ) | ( ~n2086 & n2066 ) ;
  assign n2088 = ( n1283 & ~n2087 ) | ( n1283 & 1'b0 ) | ( ~n2087 & 1'b0 ) ;
  assign n2089 = ( n1122 & ~n2088 ) | ( n1122 & 1'b0 ) | ( ~n2088 & 1'b0 ) ;
  assign n2090 = n2085 &  n2089 ;
  assign n2091 = ( n1867 & ~n1876 ) | ( n1867 & n1880 ) | ( ~n1876 & n1880 ) ;
  assign n2092 = ( n2033 & ~n1880 ) | ( n2033 & n2091 ) | ( ~n1880 & n2091 ) ;
  assign n2093 = ( n1876 & ~n2033 ) | ( n1876 & n2091 ) | ( ~n2033 & n2091 ) ;
  assign n2094 = ( n2092 & ~n1867 ) | ( n2092 & n2093 ) | ( ~n1867 & n2093 ) ;
  assign n2095 = n2090 | n2094 ;
  assign n2075 = ~n2056 & n2074 ;
  assign n2081 = ( n2075 & ~n1283 ) | ( n2075 & n2080 ) | ( ~n1283 & n2080 ) ;
  assign n2082 = n1122 | n2081 ;
  assign n2109 = n976 &  n2082 ;
  assign n2110 = n2095 &  n2109 ;
  assign n2111 = n2101 | n2110 ;
  assign n2112 = ( n2085 & ~n2088 ) | ( n2085 & 1'b0 ) | ( ~n2088 & 1'b0 ) ;
  assign n2113 = ( n1122 & n2094 ) | ( n1122 & n2112 ) | ( n2094 & n2112 ) ;
  assign n2114 = n976 | n2113 ;
  assign n2115 = ~n837 & n2114 ;
  assign n2116 = n2111 &  n2115 ;
  assign n2117 = ( n2108 & ~n2116 ) | ( n2108 & 1'b0 ) | ( ~n2116 & 1'b0 ) ;
  assign n2096 = n2082 &  n2095 ;
  assign n2102 = ( n976 & n2096 ) | ( n976 & n2101 ) | ( n2096 & n2101 ) ;
  assign n2103 = ( n837 & ~n2102 ) | ( n837 & 1'b0 ) | ( ~n2102 & 1'b0 ) ;
  assign n2131 = n713 | n2103 ;
  assign n2132 = n2117 | n2131 ;
  assign n2133 = n2123 &  n2132 ;
  assign n2134 = n2111 &  n2114 ;
  assign n2135 = ( n837 & ~n2134 ) | ( n837 & n2108 ) | ( ~n2134 & n2108 ) ;
  assign n2136 = n713 &  n2135 ;
  assign n2137 = n595 | n2136 ;
  assign n2138 = n2133 | n2137 ;
  assign n2139 = ~n2130 & n2138 ;
  assign n2118 = n2103 | n2117 ;
  assign n2124 = ( n713 & n2118 ) | ( n713 & n2123 ) | ( n2118 & n2123 ) ;
  assign n2125 = n595 &  n2124 ;
  assign n2153 = n492 | n2125 ;
  assign n2154 = n2139 | n2153 ;
  assign n2155 = n2145 &  n2154 ;
  assign n2156 = n2133 | n2136 ;
  assign n2157 = ( n595 & ~n2130 ) | ( n595 & n2156 ) | ( ~n2130 & n2156 ) ;
  assign n2158 = n492 &  n2157 ;
  assign n2178 = n2155 | n2158 ;
  assign n2179 = ( n396 & n2152 ) | ( n396 & n2178 ) | ( n2152 & n2178 ) ;
  assign n2180 = n315 &  n2179 ;
  assign n2159 = n396 | n2158 ;
  assign n2160 = n2155 | n2159 ;
  assign n2161 = n2152 &  n2160 ;
  assign n2140 = n2125 | n2139 ;
  assign n2146 = ( n492 & n2140 ) | ( n492 & n2145 ) | ( n2140 & n2145 ) ;
  assign n2147 = n396 &  n2146 ;
  assign n2175 = n315 | n2147 ;
  assign n2176 = n2161 | n2175 ;
  assign n2398 = ( n2176 & ~n2167 ) | ( n2176 & n2180 ) | ( ~n2167 & n2180 ) ;
  assign n2207 = ~n1979 & n2033 ;
  assign n2208 = ( n1984 & ~n1979 ) | ( n1984 & n1992 ) | ( ~n1979 & n1992 ) ;
  assign n2209 = ( n2207 & ~n1992 ) | ( n2207 & n2208 ) | ( ~n1992 & n2208 ) ;
  assign n2210 = ( n1979 & ~n2207 ) | ( n1979 & n2208 ) | ( ~n2207 & n2208 ) ;
  assign n2211 = ( n2209 & ~n1984 ) | ( n2209 & n2210 ) | ( ~n1984 & n2210 ) ;
  assign n2162 = n2147 | n2161 ;
  assign n2168 = ( n315 & ~n2167 ) | ( n315 & n2162 ) | ( ~n2167 & n2162 ) ;
  assign n2169 = n240 &  n2168 ;
  assign n2171 = ( n1964 & ~n1955 ) | ( n1964 & n1968 ) | ( ~n1955 & n1968 ) ;
  assign n2170 = ~n1968 & n2033 ;
  assign n2172 = ( n1964 & ~n2171 ) | ( n1964 & n2170 ) | ( ~n2171 & n2170 ) ;
  assign n2173 = ( n2170 & ~n1968 ) | ( n2170 & n2171 ) | ( ~n1968 & n2171 ) ;
  assign n2174 = ( n1955 & ~n2172 ) | ( n1955 & n2173 ) | ( ~n2172 & n2173 ) ;
  assign n2177 = ~n2167 & n2176 ;
  assign n2181 = n240 | n2180 ;
  assign n2182 = n2177 | n2181 ;
  assign n2183 = ~n2174 & n2182 ;
  assign n2184 = n2169 | n2183 ;
  assign n2185 = n1970 | n2033 ;
  assign n2186 = ( n1957 & ~n2033 ) | ( n1957 & n1962 ) | ( ~n2033 & n1962 ) ;
  assign n2187 = ( n2033 & n2185 ) | ( n2033 & n2186 ) | ( n2185 & n2186 ) ;
  assign n2188 = ( n1957 & ~n2186 ) | ( n1957 & n2185 ) | ( ~n2186 & n2185 ) ;
  assign n2189 = ( n1962 & ~n2187 ) | ( n1962 & n2188 ) | ( ~n2187 & n2188 ) ;
  assign n2190 = ( n181 & n2184 ) | ( n181 & n2189 ) | ( n2184 & n2189 ) ;
  assign n2191 = ~n145 & n2190 ;
  assign n2193 = ( n1986 & ~n1977 ) | ( n1986 & n1990 ) | ( ~n1977 & n1990 ) ;
  assign n2192 = ~n1990 & n2033 ;
  assign n2194 = ( n1986 & ~n2193 ) | ( n1986 & n2192 ) | ( ~n2193 & n2192 ) ;
  assign n2195 = ( n2192 & ~n1990 ) | ( n2192 & n2193 ) | ( ~n1990 & n2193 ) ;
  assign n2196 = ( n1977 & ~n2194 ) | ( n1977 & n2195 ) | ( ~n2194 & n2195 ) ;
  assign n2197 = n181 | n2169 ;
  assign n2198 = n2183 | n2197 ;
  assign n2199 = n2189 &  n2198 ;
  assign n2200 = n2177 | n2180 ;
  assign n2201 = ( n240 & ~n2174 ) | ( n240 & n2200 ) | ( ~n2174 & n2200 ) ;
  assign n2202 = n181 &  n2201 ;
  assign n2203 = ( n145 & ~n2202 ) | ( n145 & 1'b0 ) | ( ~n2202 & 1'b0 ) ;
  assign n2204 = ~n2199 & n2203 ;
  assign n2205 = ( n2196 & ~n2204 ) | ( n2196 & 1'b0 ) | ( ~n2204 & 1'b0 ) ;
  assign n2206 = n2191 | n2205 ;
  assign n2212 = ( n150 & ~n2211 ) | ( n150 & n2206 ) | ( ~n2211 & n2206 ) ;
  assign n2213 = n1999 | n2018 ;
  assign n2214 = ( n2015 & n2033 ) | ( n2015 & n2213 ) | ( n2033 & n2213 ) ;
  assign n2215 = ( n2015 & ~n2214 ) | ( n2015 & 1'b0 ) | ( ~n2214 & 1'b0 ) ;
  assign n2216 = ( n2015 & ~n2018 ) | ( n2015 & 1'b0 ) | ( ~n2018 & 1'b0 ) ;
  assign n2217 = n2033 &  n2216 ;
  assign n2218 = ( n1999 & ~n2216 ) | ( n1999 & n2217 ) | ( ~n2216 & n2217 ) ;
  assign n2219 = n2215 | n2218 ;
  assign n2220 = ( n2000 & ~n2007 ) | ( n2000 & 1'b0 ) | ( ~n2007 & 1'b0 ) ;
  assign n2221 = n2033 &  n2220 ;
  assign n2222 = ( n2021 & ~n2221 ) | ( n2021 & n2220 ) | ( ~n2221 & n2220 ) ;
  assign n2223 = ( n2219 & ~n2222 ) | ( n2219 & 1'b0 ) | ( ~n2222 & 1'b0 ) ;
  assign n2224 = ~n2212 & n2223 ;
  assign n2225 = ( n133 & ~n2224 ) | ( n133 & n2223 ) | ( ~n2224 & n2223 ) ;
  assign n2228 = n2199 | n2202 ;
  assign n2229 = ( n2196 & ~n145 ) | ( n2196 & n2228 ) | ( ~n145 & n2228 ) ;
  assign n2230 = n150 &  n2229 ;
  assign n2231 = n2219 | n2230 ;
  assign n2226 = n150 | n2191 ;
  assign n2227 = n2205 | n2226 ;
  assign n2232 = n2211 | n2227 ;
  assign n2233 = ( n2231 & ~n2211 ) | ( n2231 & n2232 ) | ( ~n2211 & n2232 ) ;
  assign n2234 = ( n2000 & ~n2007 ) | ( n2000 & n2033 ) | ( ~n2007 & n2033 ) ;
  assign n2236 = n2007 | n2234 ;
  assign n2235 = ( n133 & ~n2007 ) | ( n133 & n2000 ) | ( ~n2007 & n2000 ) ;
  assign n2237 = ( n2007 & ~n2236 ) | ( n2007 & n2235 ) | ( ~n2236 & n2235 ) ;
  assign n2238 = n2003 | n2030 ;
  assign n2239 = ( n2006 & n2025 ) | ( n2006 & n2238 ) | ( n2025 & n2238 ) ;
  assign n2240 = ( n2006 & ~n2239 ) | ( n2006 & 1'b0 ) | ( ~n2239 & 1'b0 ) ;
  assign n2241 = ( n2013 & ~n2240 ) | ( n2013 & n2021 ) | ( ~n2240 & n2021 ) ;
  assign n2242 = ( n2013 & ~n2241 ) | ( n2013 & 1'b0 ) | ( ~n2241 & 1'b0 ) ;
  assign n2243 = n2237 | n2242 ;
  assign n2244 = ( n2233 & ~n2243 ) | ( n2233 & 1'b0 ) | ( ~n2243 & 1'b0 ) ;
  assign n2245 = ~n2225 | ~n2244 ;
  assign n2397 = n2180 | n2245 ;
  assign n2400 = ( n2180 & ~n2398 ) | ( n2180 & n2397 ) | ( ~n2398 & n2397 ) ;
  assign n2399 = ( n2397 & ~n2176 ) | ( n2397 & n2398 ) | ( ~n2176 & n2398 ) ;
  assign n2401 = ( n2167 & ~n2400 ) | ( n2167 & n2399 ) | ( ~n2400 & n2399 ) ;
  assign n2412 = ~n2182 & n2245 ;
  assign n2413 = ( n2169 & n2174 ) | ( n2169 & n2245 ) | ( n2174 & n2245 ) ;
  assign n2415 = ( n2412 & ~n2169 ) | ( n2412 & n2413 ) | ( ~n2169 & n2413 ) ;
  assign n2414 = ( n2245 & ~n2413 ) | ( n2245 & n2412 ) | ( ~n2413 & n2412 ) ;
  assign n2416 = ( n2174 & ~n2415 ) | ( n2174 & n2414 ) | ( ~n2415 & n2414 ) ;
  assign n2368 = ~n2138 & n2245 ;
  assign n2369 = ( n2125 & n2130 ) | ( n2125 & n2245 ) | ( n2130 & n2245 ) ;
  assign n2371 = ( n2368 & ~n2125 ) | ( n2368 & n2369 ) | ( ~n2125 & n2369 ) ;
  assign n2370 = ( n2245 & ~n2369 ) | ( n2245 & n2368 ) | ( ~n2369 & n2368 ) ;
  assign n2372 = ( n2130 & ~n2371 ) | ( n2130 & n2370 ) | ( ~n2371 & n2370 ) ;
  assign n2279 = x92 | n2033 ;
  assign n2280 = x93 &  n2279 ;
  assign n2281 = ( n2045 & ~n2280 ) | ( n2045 & 1'b0 ) | ( ~n2280 & 1'b0 ) ;
  assign n2276 = ( x92 & ~n2040 ) | ( x92 & n2033 ) | ( ~n2040 & n2033 ) ;
  assign n2277 = ( x92 & ~n2276 ) | ( x92 & 1'b0 ) | ( ~n2276 & 1'b0 ) ;
  assign n2278 = ( n2035 & ~n2277 ) | ( n2035 & n2040 ) | ( ~n2277 & n2040 ) ;
  assign n2282 = ( n2245 & n2278 ) | ( n2245 & n2281 ) | ( n2278 & n2281 ) ;
  assign n2283 = ~n2278 & n2282 ;
  assign n2284 = ( n2245 & ~n2282 ) | ( n2245 & 1'b0 ) | ( ~n2282 & 1'b0 ) ;
  assign n2285 = ( n2281 & ~n2283 ) | ( n2281 & n2284 ) | ( ~n2283 & n2284 ) ;
  assign n2252 = ( x90 & ~n2245 ) | ( x90 & x91 ) | ( ~n2245 & x91 ) ;
  assign n2258 = ( x90 & ~x91 ) | ( x90 & 1'b0 ) | ( ~x91 & 1'b0 ) ;
  assign n2248 = x88 | x89 ;
  assign n2253 = ~x90 & n2248 ;
  assign n2254 = ( x90 & ~n2031 ) | ( x90 & n2253 ) | ( ~n2031 & n2253 ) ;
  assign n2255 = ( n2013 & ~n2254 ) | ( n2013 & n2021 ) | ( ~n2254 & n2021 ) ;
  assign n2256 = ( n2013 & ~n2255 ) | ( n2013 & 1'b0 ) | ( ~n2255 & 1'b0 ) ;
  assign n2257 = ( n2245 & ~x91 ) | ( n2245 & n2256 ) | ( ~x91 & n2256 ) ;
  assign n2259 = ( n2252 & ~n2258 ) | ( n2252 & n2257 ) | ( ~n2258 & n2257 ) ;
  assign n2250 = x90 &  n2245 ;
  assign n2249 = x90 | n2248 ;
  assign n2251 = ( n2033 & ~n2250 ) | ( n2033 & n2249 ) | ( ~n2250 & n2249 ) ;
  assign n2260 = ~n2251 & n2259 ;
  assign n2261 = ( n1827 & ~n2259 ) | ( n1827 & n2260 ) | ( ~n2259 & n2260 ) ;
  assign n2262 = ~n1827 & n2251 ;
  assign n2263 = n2259 &  n2262 ;
  assign n2265 = n2033 | n2242 ;
  assign n2266 = ( n2233 & n2237 ) | ( n2233 & n2265 ) | ( n2237 & n2265 ) ;
  assign n2267 = ( n2233 & ~n2266 ) | ( n2233 & 1'b0 ) | ( ~n2266 & 1'b0 ) ;
  assign n2268 = n2225 &  n2267 ;
  assign n2264 = ~n1828 & n2245 ;
  assign n2269 = ( n2264 & ~n2268 ) | ( n2264 & 1'b0 ) | ( ~n2268 & 1'b0 ) ;
  assign n2270 = ( x92 & n2268 ) | ( x92 & n2269 ) | ( n2268 & n2269 ) ;
  assign n2271 = x92 | n2268 ;
  assign n2272 = n2264 | n2271 ;
  assign n2273 = ~n2270 & n2272 ;
  assign n2274 = n2263 | n2273 ;
  assign n2275 = ~n2261 & n2274 ;
  assign n2286 = ( n1636 & ~n2285 ) | ( n1636 & n2275 ) | ( ~n2285 & n2275 ) ;
  assign n2287 = n1452 | n2286 ;
  assign n2288 = ~n2068 & n2071 ;
  assign n2289 = ( n2068 & ~n2288 ) | ( n2068 & n2245 ) | ( ~n2288 & n2245 ) ;
  assign n2290 = ( n2054 & ~n2289 ) | ( n2054 & n2068 ) | ( ~n2289 & n2068 ) ;
  assign n2291 = ( n2054 & ~n2068 ) | ( n2054 & n2289 ) | ( ~n2068 & n2289 ) ;
  assign n2292 = ( n2290 & ~n2054 ) | ( n2290 & n2291 ) | ( ~n2054 & n2291 ) ;
  assign n2293 = ( n1636 & ~n2261 ) | ( n1636 & 1'b0 ) | ( ~n2261 & 1'b0 ) ;
  assign n2294 = n2274 &  n2293 ;
  assign n2295 = ( n2285 & ~n2294 ) | ( n2285 & 1'b0 ) | ( ~n2294 & 1'b0 ) ;
  assign n2296 = n2251 &  n2259 ;
  assign n2297 = ( n2273 & ~n1827 ) | ( n2273 & n2296 ) | ( ~n1827 & n2296 ) ;
  assign n2298 = n1636 | n2297 ;
  assign n2299 = n1452 &  n2298 ;
  assign n2300 = ~n2295 & n2299 ;
  assign n2301 = ( n2292 & ~n2300 ) | ( n2292 & 1'b0 ) | ( ~n2300 & 1'b0 ) ;
  assign n2302 = ( n2287 & ~n2301 ) | ( n2287 & 1'b0 ) | ( ~n2301 & 1'b0 ) ;
  assign n2303 = n2056 | n2245 ;
  assign n2304 = ( n2056 & ~n2073 ) | ( n2056 & n2066 ) | ( ~n2073 & n2066 ) ;
  assign n2305 = ( n2073 & n2303 ) | ( n2073 & n2304 ) | ( n2303 & n2304 ) ;
  assign n2306 = ( n2056 & ~n2304 ) | ( n2056 & n2303 ) | ( ~n2304 & n2303 ) ;
  assign n2307 = ( n2066 & ~n2305 ) | ( n2066 & n2306 ) | ( ~n2305 & n2306 ) ;
  assign n2308 = ( n2302 & ~n1283 ) | ( n2302 & n2307 ) | ( ~n1283 & n2307 ) ;
  assign n2309 = n1122 | n2308 ;
  assign n2310 = n2088 | n2245 ;
  assign n2311 = ( n2080 & ~n2088 ) | ( n2080 & n2084 ) | ( ~n2088 & n2084 ) ;
  assign n2313 = ( n2088 & n2310 ) | ( n2088 & n2311 ) | ( n2310 & n2311 ) ;
  assign n2312 = ( n2084 & ~n2311 ) | ( n2084 & n2310 ) | ( ~n2311 & n2310 ) ;
  assign n2314 = ( n2080 & ~n2313 ) | ( n2080 & n2312 ) | ( ~n2313 & n2312 ) ;
  assign n2315 = ~n1283 & n2287 ;
  assign n2316 = ~n2301 & n2315 ;
  assign n2317 = n2307 | n2316 ;
  assign n2318 = ~n2295 & n2298 ;
  assign n2319 = ( n1452 & ~n2292 ) | ( n1452 & n2318 ) | ( ~n2292 & n2318 ) ;
  assign n2320 = ( n1283 & ~n2319 ) | ( n1283 & 1'b0 ) | ( ~n2319 & 1'b0 ) ;
  assign n2321 = ( n1122 & ~n2320 ) | ( n1122 & 1'b0 ) | ( ~n2320 & 1'b0 ) ;
  assign n2322 = n2317 &  n2321 ;
  assign n2323 = n2314 | n2322 ;
  assign n2324 = n2309 &  n2323 ;
  assign n2325 = ( n2082 & ~n2094 ) | ( n2082 & n2090 ) | ( ~n2094 & n2090 ) ;
  assign n2326 = ( n2090 & ~n2325 ) | ( n2090 & n2245 ) | ( ~n2325 & n2245 ) ;
  assign n2327 = ( n2245 & ~n2082 ) | ( n2245 & n2325 ) | ( ~n2082 & n2325 ) ;
  assign n2328 = ( n2094 & ~n2326 ) | ( n2094 & n2327 ) | ( ~n2326 & n2327 ) ;
  assign n2329 = ( n976 & n2324 ) | ( n976 & n2328 ) | ( n2324 & n2328 ) ;
  assign n2330 = ( n837 & ~n2329 ) | ( n837 & 1'b0 ) | ( ~n2329 & 1'b0 ) ;
  assign n2331 = ( n2114 & ~n2245 ) | ( n2114 & 1'b0 ) | ( ~n2245 & 1'b0 ) ;
  assign n2332 = ( n2101 & n2110 ) | ( n2101 & n2114 ) | ( n2110 & n2114 ) ;
  assign n2333 = ( n2331 & ~n2110 ) | ( n2331 & n2332 ) | ( ~n2110 & n2332 ) ;
  assign n2334 = ( n2114 & ~n2332 ) | ( n2114 & n2331 ) | ( ~n2332 & n2331 ) ;
  assign n2335 = ( n2101 & ~n2333 ) | ( n2101 & n2334 ) | ( ~n2333 & n2334 ) ;
  assign n2336 = n976 &  n2309 ;
  assign n2337 = n2323 &  n2336 ;
  assign n2338 = n2328 | n2337 ;
  assign n2339 = ( n2317 & ~n2320 ) | ( n2317 & 1'b0 ) | ( ~n2320 & 1'b0 ) ;
  assign n2340 = ( n1122 & n2314 ) | ( n1122 & n2339 ) | ( n2314 & n2339 ) ;
  assign n2341 = n976 | n2340 ;
  assign n2342 = ~n837 & n2341 ;
  assign n2343 = n2338 &  n2342 ;
  assign n2344 = n2335 | n2343 ;
  assign n2345 = ~n2330 & n2344 ;
  assign n2346 = n2116 &  n2245 ;
  assign n2347 = ( n2103 & n2108 ) | ( n2103 & n2245 ) | ( n2108 & n2245 ) ;
  assign n2349 = ( n2346 & ~n2103 ) | ( n2346 & n2347 ) | ( ~n2103 & n2347 ) ;
  assign n2348 = ( n2245 & ~n2347 ) | ( n2245 & n2346 ) | ( ~n2347 & n2346 ) ;
  assign n2350 = ( n2108 & ~n2349 ) | ( n2108 & n2348 ) | ( ~n2349 & n2348 ) ;
  assign n2351 = ( n713 & ~n2345 ) | ( n713 & n2350 ) | ( ~n2345 & n2350 ) ;
  assign n2352 = n595 &  n2351 ;
  assign n2353 = n2136 | n2245 ;
  assign n2354 = ( n2123 & n2132 ) | ( n2123 & n2136 ) | ( n2132 & n2136 ) ;
  assign n2355 = ( n2353 & ~n2132 ) | ( n2353 & n2354 ) | ( ~n2132 & n2354 ) ;
  assign n2356 = ( n2136 & ~n2354 ) | ( n2136 & n2353 ) | ( ~n2354 & n2353 ) ;
  assign n2357 = ( n2123 & ~n2355 ) | ( n2123 & n2356 ) | ( ~n2355 & n2356 ) ;
  assign n2358 = n713 | n2330 ;
  assign n2359 = ( n2344 & ~n2358 ) | ( n2344 & 1'b0 ) | ( ~n2358 & 1'b0 ) ;
  assign n2360 = ( n2350 & ~n2359 ) | ( n2350 & 1'b0 ) | ( ~n2359 & 1'b0 ) ;
  assign n2361 = n2338 &  n2341 ;
  assign n2362 = ( n2335 & ~n837 ) | ( n2335 & n2361 ) | ( ~n837 & n2361 ) ;
  assign n2363 = ( n713 & ~n2362 ) | ( n713 & 1'b0 ) | ( ~n2362 & 1'b0 ) ;
  assign n2364 = n595 | n2363 ;
  assign n2365 = n2360 | n2364 ;
  assign n2366 = n2357 &  n2365 ;
  assign n2367 = n2352 | n2366 ;
  assign n2373 = ( n492 & ~n2372 ) | ( n492 & n2367 ) | ( ~n2372 & n2367 ) ;
  assign n2374 = n396 &  n2373 ;
  assign n2375 = n2158 | n2245 ;
  assign n2376 = ( n2145 & n2154 ) | ( n2145 & n2158 ) | ( n2154 & n2158 ) ;
  assign n2377 = ( n2375 & ~n2154 ) | ( n2375 & n2376 ) | ( ~n2154 & n2376 ) ;
  assign n2378 = ( n2158 & ~n2376 ) | ( n2158 & n2375 ) | ( ~n2376 & n2375 ) ;
  assign n2379 = ( n2145 & ~n2377 ) | ( n2145 & n2378 ) | ( ~n2377 & n2378 ) ;
  assign n2380 = n492 | n2352 ;
  assign n2381 = n2366 | n2380 ;
  assign n2382 = ~n2372 & n2381 ;
  assign n2383 = n2360 | n2363 ;
  assign n2384 = ( n595 & n2357 ) | ( n595 & n2383 ) | ( n2357 & n2383 ) ;
  assign n2385 = n492 &  n2384 ;
  assign n2386 = n396 | n2385 ;
  assign n2387 = n2382 | n2386 ;
  assign n2388 = n2379 &  n2387 ;
  assign n2389 = n2374 | n2388 ;
  assign n2390 = ~n2160 & n2245 ;
  assign n2391 = ( n2147 & n2152 ) | ( n2147 & n2245 ) | ( n2152 & n2245 ) ;
  assign n2393 = ( n2390 & ~n2147 ) | ( n2390 & n2391 ) | ( ~n2147 & n2391 ) ;
  assign n2392 = ( n2245 & ~n2391 ) | ( n2245 & n2390 ) | ( ~n2391 & n2390 ) ;
  assign n2394 = ( n2152 & ~n2393 ) | ( n2152 & n2392 ) | ( ~n2393 & n2392 ) ;
  assign n2395 = ( n315 & n2389 ) | ( n315 & n2394 ) | ( n2389 & n2394 ) ;
  assign n2396 = n240 &  n2395 ;
  assign n2402 = n315 | n2374 ;
  assign n2403 = n2388 | n2402 ;
  assign n2404 = n2394 &  n2403 ;
  assign n2405 = n2382 | n2385 ;
  assign n2406 = ( n396 & n2379 ) | ( n396 & n2405 ) | ( n2379 & n2405 ) ;
  assign n2407 = n315 &  n2406 ;
  assign n2408 = n240 | n2407 ;
  assign n2409 = n2404 | n2408 ;
  assign n2410 = ~n2401 & n2409 ;
  assign n2411 = n2396 | n2410 ;
  assign n2417 = ( n181 & ~n2416 ) | ( n181 & n2411 ) | ( ~n2416 & n2411 ) ;
  assign n2418 = ~n145 & n2417 ;
  assign n2420 = ( n2198 & ~n2189 ) | ( n2198 & n2202 ) | ( ~n2189 & n2202 ) ;
  assign n2419 = n2202 | n2245 ;
  assign n2422 = ( n2202 & ~n2420 ) | ( n2202 & n2419 ) | ( ~n2420 & n2419 ) ;
  assign n2421 = ( n2419 & ~n2198 ) | ( n2419 & n2420 ) | ( ~n2198 & n2420 ) ;
  assign n2423 = ( n2189 & ~n2422 ) | ( n2189 & n2421 ) | ( ~n2422 & n2421 ) ;
  assign n2424 = n181 | n2396 ;
  assign n2425 = n2410 | n2424 ;
  assign n2426 = ~n2416 & n2425 ;
  assign n2427 = n2404 | n2407 ;
  assign n2428 = ( n240 & ~n2401 ) | ( n240 & n2427 ) | ( ~n2401 & n2427 ) ;
  assign n2429 = n181 &  n2428 ;
  assign n2430 = ( n145 & ~n2429 ) | ( n145 & 1'b0 ) | ( ~n2429 & 1'b0 ) ;
  assign n2431 = ~n2426 & n2430 ;
  assign n2432 = ( n2423 & ~n2431 ) | ( n2423 & 1'b0 ) | ( ~n2431 & 1'b0 ) ;
  assign n2433 = n2418 | n2432 ;
  assign n2434 = n2191 | n2245 ;
  assign n2435 = ( n2196 & ~n2191 ) | ( n2196 & n2204 ) | ( ~n2191 & n2204 ) ;
  assign n2437 = ( n2191 & n2434 ) | ( n2191 & n2435 ) | ( n2434 & n2435 ) ;
  assign n2436 = ( n2204 & ~n2435 ) | ( n2204 & n2434 ) | ( ~n2435 & n2434 ) ;
  assign n2438 = ( n2196 & ~n2437 ) | ( n2196 & n2436 ) | ( ~n2437 & n2436 ) ;
  assign n2439 = ( n150 & n2433 ) | ( n150 & n2438 ) | ( n2433 & n2438 ) ;
  assign n2440 = n2211 &  n2227 ;
  assign n2441 = ( n2230 & n2245 ) | ( n2230 & n2440 ) | ( n2245 & n2440 ) ;
  assign n2442 = ~n2230 & n2441 ;
  assign n2443 = ( n2227 & ~n2230 ) | ( n2227 & 1'b0 ) | ( ~n2230 & 1'b0 ) ;
  assign n2444 = ~n2245 & n2443 ;
  assign n2445 = ( n2211 & ~n2444 ) | ( n2211 & n2443 ) | ( ~n2444 & n2443 ) ;
  assign n2446 = ~n2442 & n2445 ;
  assign n2447 = n2212 &  n2219 ;
  assign n2448 = ~n2245 & n2447 ;
  assign n2449 = ( n2233 & ~n2447 ) | ( n2233 & n2448 ) | ( ~n2447 & n2448 ) ;
  assign n2450 = ~n2446 & n2449 ;
  assign n2451 = ~n2439 & n2450 ;
  assign n2452 = ( n133 & ~n2451 ) | ( n133 & n2450 ) | ( ~n2451 & n2450 ) ;
  assign n2455 = n2426 | n2429 ;
  assign n2456 = ( n2423 & ~n145 ) | ( n2423 & n2455 ) | ( ~n145 & n2455 ) ;
  assign n2457 = n150 &  n2456 ;
  assign n2458 = ( n2446 & ~n2457 ) | ( n2446 & 1'b0 ) | ( ~n2457 & 1'b0 ) ;
  assign n2453 = n150 | n2418 ;
  assign n2454 = n2432 | n2453 ;
  assign n2459 = ( n2438 & ~n2454 ) | ( n2438 & 1'b0 ) | ( ~n2454 & 1'b0 ) ;
  assign n2460 = ( n2458 & ~n2438 ) | ( n2458 & n2459 ) | ( ~n2438 & n2459 ) ;
  assign n2462 = ( n133 & n2212 ) | ( n133 & n2219 ) | ( n2212 & n2219 ) ;
  assign n2461 = ( n2212 & ~n2245 ) | ( n2212 & n2219 ) | ( ~n2245 & n2219 ) ;
  assign n2463 = ( n2219 & ~n2461 ) | ( n2219 & 1'b0 ) | ( ~n2461 & 1'b0 ) ;
  assign n2464 = ( n2462 & ~n2219 ) | ( n2462 & n2463 ) | ( ~n2219 & n2463 ) ;
  assign n2465 = n2215 | n2242 ;
  assign n2466 = ( n2237 & ~n2218 ) | ( n2237 & n2465 ) | ( ~n2218 & n2465 ) ;
  assign n2467 = n2218 | n2466 ;
  assign n2468 = ( n2225 & ~n2233 ) | ( n2225 & n2467 ) | ( ~n2233 & n2467 ) ;
  assign n2469 = ( n2225 & ~n2468 ) | ( n2225 & 1'b0 ) | ( ~n2468 & 1'b0 ) ;
  assign n2470 = n2464 | n2469 ;
  assign n2471 = n2460 | n2470 ;
  assign n2472 = ~n2452 |  n2471 ;
  assign n2647 = ( n2396 & ~n2401 ) | ( n2396 & n2472 ) | ( ~n2401 & n2472 ) ;
  assign n2646 = ~n2409 & n2472 ;
  assign n2648 = ( n2472 & ~n2647 ) | ( n2472 & n2646 ) | ( ~n2647 & n2646 ) ;
  assign n2649 = ( n2646 & ~n2396 ) | ( n2646 & n2647 ) | ( ~n2396 & n2647 ) ;
  assign n2650 = ( n2401 & ~n2648 ) | ( n2401 & n2649 ) | ( ~n2648 & n2649 ) ;
  assign n2631 = n2407 | n2472 ;
  assign n2632 = ( n2394 & n2403 ) | ( n2394 & n2407 ) | ( n2403 & n2407 ) ;
  assign n2633 = ( n2631 & ~n2403 ) | ( n2631 & n2632 ) | ( ~n2403 & n2632 ) ;
  assign n2634 = ( n2407 & ~n2632 ) | ( n2407 & n2631 ) | ( ~n2632 & n2631 ) ;
  assign n2635 = ( n2394 & ~n2633 ) | ( n2394 & n2634 ) | ( ~n2633 & n2634 ) ;
  assign n2624 = ~n2387 & n2472 ;
  assign n2625 = ( n2374 & ~n2624 ) | ( n2374 & n2472 ) | ( ~n2624 & n2472 ) ;
  assign n2626 = ( n2374 & ~n2625 ) | ( n2374 & n2379 ) | ( ~n2625 & n2379 ) ;
  assign n2627 = ( n2379 & ~n2374 ) | ( n2379 & n2625 ) | ( ~n2374 & n2625 ) ;
  assign n2628 = ( n2626 & ~n2379 ) | ( n2626 & n2627 ) | ( ~n2379 & n2627 ) ;
  assign n2610 = ( n2381 & ~n2372 ) | ( n2381 & n2385 ) | ( ~n2372 & n2385 ) ;
  assign n2609 = n2385 | n2472 ;
  assign n2612 = ( n2385 & ~n2610 ) | ( n2385 & n2609 ) | ( ~n2610 & n2609 ) ;
  assign n2611 = ( n2609 & ~n2381 ) | ( n2609 & n2610 ) | ( ~n2381 & n2610 ) ;
  assign n2613 = ( n2372 & ~n2612 ) | ( n2372 & n2611 ) | ( ~n2612 & n2611 ) ;
  assign n2602 = ~n2365 & n2472 ;
  assign n2603 = ( n2352 & n2357 ) | ( n2352 & n2472 ) | ( n2357 & n2472 ) ;
  assign n2605 = ( n2602 & ~n2352 ) | ( n2602 & n2603 ) | ( ~n2352 & n2603 ) ;
  assign n2604 = ( n2472 & ~n2603 ) | ( n2472 & n2602 ) | ( ~n2603 & n2602 ) ;
  assign n2606 = ( n2357 & ~n2605 ) | ( n2357 & n2604 ) | ( ~n2605 & n2604 ) ;
  assign n2587 = n2363 | n2472 ;
  assign n2588 = ( n2350 & ~n2359 ) | ( n2350 & n2363 ) | ( ~n2359 & n2363 ) ;
  assign n2589 = ( n2359 & n2587 ) | ( n2359 & n2588 ) | ( n2587 & n2588 ) ;
  assign n2590 = ( n2363 & ~n2588 ) | ( n2363 & n2587 ) | ( ~n2588 & n2587 ) ;
  assign n2591 = ( n2350 & ~n2589 ) | ( n2350 & n2590 ) | ( ~n2589 & n2590 ) ;
  assign n2580 = n2343 &  n2472 ;
  assign n2581 = ( n2330 & ~n2580 ) | ( n2330 & n2472 ) | ( ~n2580 & n2472 ) ;
  assign n2582 = ( n2335 & ~n2330 ) | ( n2335 & n2581 ) | ( ~n2330 & n2581 ) ;
  assign n2583 = ( n2330 & ~n2581 ) | ( n2330 & n2335 ) | ( ~n2581 & n2335 ) ;
  assign n2584 = ( n2582 & ~n2335 ) | ( n2582 & n2583 ) | ( ~n2335 & n2583 ) ;
  assign n2560 = ( n2309 & ~n2314 ) | ( n2309 & n2322 ) | ( ~n2314 & n2322 ) ;
  assign n2559 = ( n2309 & ~n2472 ) | ( n2309 & 1'b0 ) | ( ~n2472 & 1'b0 ) ;
  assign n2562 = ( n2309 & ~n2560 ) | ( n2309 & n2559 ) | ( ~n2560 & n2559 ) ;
  assign n2561 = ( n2559 & ~n2322 ) | ( n2559 & n2560 ) | ( ~n2322 & n2560 ) ;
  assign n2563 = ( n2314 & ~n2562 ) | ( n2314 & n2561 ) | ( ~n2562 & n2561 ) ;
  assign n2544 = n2320 | n2472 ;
  assign n2545 = ( n2307 & ~n2316 ) | ( n2307 & n2320 ) | ( ~n2316 & n2320 ) ;
  assign n2546 = ( n2316 & n2544 ) | ( n2316 & n2545 ) | ( n2544 & n2545 ) ;
  assign n2547 = ( n2320 & ~n2545 ) | ( n2320 & n2544 ) | ( ~n2545 & n2544 ) ;
  assign n2548 = ( n2307 & ~n2546 ) | ( n2307 & n2547 ) | ( ~n2546 & n2547 ) ;
  assign n2538 = ( n2287 & ~n2292 ) | ( n2287 & n2300 ) | ( ~n2292 & n2300 ) ;
  assign n2537 = ( n2287 & ~n2472 ) | ( n2287 & 1'b0 ) | ( ~n2472 & 1'b0 ) ;
  assign n2540 = ( n2287 & ~n2538 ) | ( n2287 & n2537 ) | ( ~n2538 & n2537 ) ;
  assign n2539 = ( n2537 & ~n2300 ) | ( n2537 & n2538 ) | ( ~n2300 & n2538 ) ;
  assign n2541 = ( n2292 & ~n2540 ) | ( n2292 & n2539 ) | ( ~n2540 & n2539 ) ;
  assign n2522 = ( n2298 & ~n2472 ) | ( n2298 & 1'b0 ) | ( ~n2472 & 1'b0 ) ;
  assign n2523 = ( n2285 & n2294 ) | ( n2285 & n2298 ) | ( n2294 & n2298 ) ;
  assign n2524 = ( n2522 & ~n2294 ) | ( n2522 & n2523 ) | ( ~n2294 & n2523 ) ;
  assign n2525 = ( n2298 & ~n2523 ) | ( n2298 & n2522 ) | ( ~n2523 & n2522 ) ;
  assign n2526 = ( n2285 & ~n2524 ) | ( n2285 & n2525 ) | ( ~n2524 & n2525 ) ;
  assign n2515 = ( n2261 & ~n2263 ) | ( n2261 & 1'b0 ) | ( ~n2263 & 1'b0 ) ;
  assign n2516 = ( n2263 & ~n2515 ) | ( n2263 & n2273 ) | ( ~n2515 & n2273 ) ;
  assign n2518 = ( n2472 & n2515 ) | ( n2472 & n2516 ) | ( n2515 & n2516 ) ;
  assign n2517 = ( n2263 & ~n2516 ) | ( n2263 & n2472 ) | ( ~n2516 & n2472 ) ;
  assign n2519 = ( n2273 & ~n2518 ) | ( n2273 & n2517 ) | ( ~n2518 & n2517 ) ;
  assign n2499 = ~x90 & n2245 ;
  assign n2500 = ( x91 & ~n2499 ) | ( x91 & 1'b0 ) | ( ~n2499 & 1'b0 ) ;
  assign n2501 = n2264 | n2500 ;
  assign n2496 = ( n2245 & ~x90 ) | ( n2245 & n2256 ) | ( ~x90 & n2256 ) ;
  assign n2497 = x90 &  n2496 ;
  assign n2498 = ( n2251 & ~n2256 ) | ( n2251 & n2497 ) | ( ~n2256 & n2497 ) ;
  assign n2502 = ( n2498 & ~n2472 ) | ( n2498 & n2501 ) | ( ~n2472 & n2501 ) ;
  assign n2504 = n2472 &  n2502 ;
  assign n2503 = ( n2498 & ~n2502 ) | ( n2498 & 1'b0 ) | ( ~n2502 & 1'b0 ) ;
  assign n2505 = ( n2501 & ~n2504 ) | ( n2501 & n2503 ) | ( ~n2504 & n2503 ) ;
  assign n2485 = ( n2245 & ~n2469 ) | ( n2245 & 1'b0 ) | ( ~n2469 & 1'b0 ) ;
  assign n2486 = ( n2460 & ~n2464 ) | ( n2460 & n2485 ) | ( ~n2464 & n2485 ) ;
  assign n2487 = ~n2460 & n2486 ;
  assign n2488 = n2452 &  n2487 ;
  assign n2484 = ~n2248 & n2472 ;
  assign n2489 = ( n2484 & ~n2488 ) | ( n2484 & 1'b0 ) | ( ~n2488 & 1'b0 ) ;
  assign n2490 = ( x90 & n2488 ) | ( x90 & n2489 ) | ( n2488 & n2489 ) ;
  assign n2491 = x90 | n2488 ;
  assign n2492 = n2484 | n2491 ;
  assign n2493 = ~n2490 & n2492 ;
  assign n2475 = ( x88 & ~n2472 ) | ( x88 & x89 ) | ( ~n2472 & x89 ) ;
  assign n2481 = ( x88 & ~x89 ) | ( x88 & 1'b0 ) | ( ~x89 & 1'b0 ) ;
  assign n2246 = x86 | x87 ;
  assign n2476 = ~x88 & n2246 ;
  assign n2477 = ( x88 & ~n2243 ) | ( x88 & n2476 ) | ( ~n2243 & n2476 ) ;
  assign n2478 = ( n2233 & ~n2225 ) | ( n2233 & n2477 ) | ( ~n2225 & n2477 ) ;
  assign n2479 = n2225 &  n2478 ;
  assign n2480 = ( n2472 & ~x89 ) | ( n2472 & n2479 ) | ( ~x89 & n2479 ) ;
  assign n2482 = ( n2475 & ~n2481 ) | ( n2475 & n2480 ) | ( ~n2481 & n2480 ) ;
  assign n2247 = x88 | n2246 ;
  assign n2473 = x88 &  n2472 ;
  assign n2474 = ( n2245 & ~n2247 ) | ( n2245 & n2473 ) | ( ~n2247 & n2473 ) ;
  assign n2506 = ( n2033 & ~n2474 ) | ( n2033 & 1'b0 ) | ( ~n2474 & 1'b0 ) ;
  assign n2507 = n2482 &  n2506 ;
  assign n2508 = n2493 | n2507 ;
  assign n2509 = n2474 &  n2482 ;
  assign n2510 = ( n2033 & ~n2509 ) | ( n2033 & n2482 ) | ( ~n2509 & n2482 ) ;
  assign n2511 = ~n1827 & n2510 ;
  assign n2512 = n2508 &  n2511 ;
  assign n2513 = n2505 | n2512 ;
  assign n2483 = ~n2474 & n2482 ;
  assign n2494 = ( n2033 & n2483 ) | ( n2033 & n2493 ) | ( n2483 & n2493 ) ;
  assign n2495 = ( n1827 & ~n2494 ) | ( n1827 & 1'b0 ) | ( ~n2494 & 1'b0 ) ;
  assign n2527 = ( n1636 & ~n2495 ) | ( n1636 & 1'b0 ) | ( ~n2495 & 1'b0 ) ;
  assign n2528 = n2513 &  n2527 ;
  assign n2529 = n2519 | n2528 ;
  assign n2530 = n2508 &  n2510 ;
  assign n2531 = ( n2505 & ~n1827 ) | ( n2505 & n2530 ) | ( ~n1827 & n2530 ) ;
  assign n2532 = n1636 | n2531 ;
  assign n2533 = n1452 &  n2532 ;
  assign n2534 = n2529 &  n2533 ;
  assign n2535 = ( n2526 & ~n2534 ) | ( n2526 & 1'b0 ) | ( ~n2534 & 1'b0 ) ;
  assign n2514 = ~n2495 & n2513 ;
  assign n2520 = ( n1636 & n2514 ) | ( n1636 & n2519 ) | ( n2514 & n2519 ) ;
  assign n2521 = n1452 | n2520 ;
  assign n2549 = ~n1283 & n2521 ;
  assign n2550 = ~n2535 & n2549 ;
  assign n2551 = ( n2541 & ~n2550 ) | ( n2541 & 1'b0 ) | ( ~n2550 & 1'b0 ) ;
  assign n2552 = n2529 &  n2532 ;
  assign n2553 = ( n1452 & ~n2526 ) | ( n1452 & n2552 ) | ( ~n2526 & n2552 ) ;
  assign n2554 = ( n1283 & ~n2553 ) | ( n1283 & 1'b0 ) | ( ~n2553 & 1'b0 ) ;
  assign n2555 = ( n1122 & ~n2554 ) | ( n1122 & 1'b0 ) | ( ~n2554 & 1'b0 ) ;
  assign n2556 = ~n2551 & n2555 ;
  assign n2557 = n2548 | n2556 ;
  assign n2536 = ( n2521 & ~n2535 ) | ( n2521 & 1'b0 ) | ( ~n2535 & 1'b0 ) ;
  assign n2542 = ( n1283 & ~n2536 ) | ( n1283 & n2541 ) | ( ~n2536 & n2541 ) ;
  assign n2543 = ~n1122 & n2542 ;
  assign n2566 = ( n976 & ~n2543 ) | ( n976 & 1'b0 ) | ( ~n2543 & 1'b0 ) ;
  assign n2567 = n2557 &  n2566 ;
  assign n2568 = n2563 | n2567 ;
  assign n2569 = n2551 | n2554 ;
  assign n2570 = ( n1122 & ~n2569 ) | ( n1122 & n2548 ) | ( ~n2569 & n2548 ) ;
  assign n2571 = n976 | n2570 ;
  assign n2572 = ~n837 & n2571 ;
  assign n2573 = n2568 &  n2572 ;
  assign n2574 = ( n2328 & n2337 ) | ( n2328 & n2341 ) | ( n2337 & n2341 ) ;
  assign n2575 = ( n2472 & ~n2341 ) | ( n2472 & n2574 ) | ( ~n2341 & n2574 ) ;
  assign n2576 = ( n2337 & ~n2574 ) | ( n2337 & n2472 ) | ( ~n2574 & n2472 ) ;
  assign n2577 = ( n2328 & ~n2575 ) | ( n2328 & n2576 ) | ( ~n2575 & n2576 ) ;
  assign n2578 = n2573 | n2577 ;
  assign n2558 = ~n2543 & n2557 ;
  assign n2564 = ( n976 & n2558 ) | ( n976 & n2563 ) | ( n2558 & n2563 ) ;
  assign n2565 = ( n837 & ~n2564 ) | ( n837 & 1'b0 ) | ( ~n2564 & 1'b0 ) ;
  assign n2592 = n713 | n2565 ;
  assign n2593 = ( n2578 & ~n2592 ) | ( n2578 & 1'b0 ) | ( ~n2592 & 1'b0 ) ;
  assign n2594 = n2584 | n2593 ;
  assign n2595 = n2568 &  n2571 ;
  assign n2596 = ( n2577 & ~n837 ) | ( n2577 & n2595 ) | ( ~n837 & n2595 ) ;
  assign n2597 = ( n713 & ~n2596 ) | ( n713 & 1'b0 ) | ( ~n2596 & 1'b0 ) ;
  assign n2598 = n595 | n2597 ;
  assign n2599 = ( n2594 & ~n2598 ) | ( n2594 & 1'b0 ) | ( ~n2598 & 1'b0 ) ;
  assign n2600 = ( n2591 & ~n2599 ) | ( n2591 & 1'b0 ) | ( ~n2599 & 1'b0 ) ;
  assign n2579 = ~n2565 & n2578 ;
  assign n2585 = ( n2579 & ~n713 ) | ( n2579 & n2584 ) | ( ~n713 & n2584 ) ;
  assign n2586 = ( n595 & ~n2585 ) | ( n595 & 1'b0 ) | ( ~n2585 & 1'b0 ) ;
  assign n2614 = n492 | n2586 ;
  assign n2615 = n2600 | n2614 ;
  assign n2616 = n2606 &  n2615 ;
  assign n2617 = ( n2594 & ~n2597 ) | ( n2594 & 1'b0 ) | ( ~n2597 & 1'b0 ) ;
  assign n2618 = ( n595 & ~n2617 ) | ( n595 & n2591 ) | ( ~n2617 & n2591 ) ;
  assign n2619 = n492 &  n2618 ;
  assign n2620 = n396 | n2619 ;
  assign n2621 = n2616 | n2620 ;
  assign n2622 = ~n2613 & n2621 ;
  assign n2601 = n2586 | n2600 ;
  assign n2607 = ( n492 & n2601 ) | ( n492 & n2606 ) | ( n2601 & n2606 ) ;
  assign n2608 = n396 &  n2607 ;
  assign n2636 = n315 | n2608 ;
  assign n2637 = n2622 | n2636 ;
  assign n2638 = n2628 &  n2637 ;
  assign n2639 = n2616 | n2619 ;
  assign n2640 = ( n396 & ~n2613 ) | ( n396 & n2639 ) | ( ~n2613 & n2639 ) ;
  assign n2641 = n315 &  n2640 ;
  assign n2661 = n2638 | n2641 ;
  assign n2662 = ( n240 & n2635 ) | ( n240 & n2661 ) | ( n2635 & n2661 ) ;
  assign n2663 = n181 &  n2662 ;
  assign n2623 = n2608 | n2622 ;
  assign n2629 = ( n315 & n2623 ) | ( n315 & n2628 ) | ( n2623 & n2628 ) ;
  assign n2630 = n240 &  n2629 ;
  assign n2642 = n240 | n2641 ;
  assign n2643 = n2638 | n2642 ;
  assign n2644 = n2635 &  n2643 ;
  assign n2645 = n2630 | n2644 ;
  assign n2651 = ( n181 & ~n2650 ) | ( n181 & n2645 ) | ( ~n2650 & n2645 ) ;
  assign n2652 = ~n145 & n2651 ;
  assign n2653 = n2429 | n2472 ;
  assign n2654 = ( n2416 & n2425 ) | ( n2416 & n2429 ) | ( n2425 & n2429 ) ;
  assign n2655 = ( n2653 & ~n2425 ) | ( n2653 & n2654 ) | ( ~n2425 & n2654 ) ;
  assign n2656 = ( n2429 & ~n2654 ) | ( n2429 & n2653 ) | ( ~n2654 & n2653 ) ;
  assign n2657 = ( n2416 & ~n2655 ) | ( n2416 & n2656 ) | ( ~n2655 & n2656 ) ;
  assign n2658 = n181 | n2630 ;
  assign n2659 = n2644 | n2658 ;
  assign n2660 = ~n2650 & n2659 ;
  assign n2664 = ( n145 & ~n2663 ) | ( n145 & 1'b0 ) | ( ~n2663 & 1'b0 ) ;
  assign n2665 = ~n2660 & n2664 ;
  assign n2666 = n2657 | n2665 ;
  assign n2667 = ~n2652 & n2666 ;
  assign n2668 = n2418 | n2472 ;
  assign n2669 = ( n2423 & ~n2418 ) | ( n2423 & n2431 ) | ( ~n2418 & n2431 ) ;
  assign n2671 = ( n2418 & n2668 ) | ( n2418 & n2669 ) | ( n2668 & n2669 ) ;
  assign n2670 = ( n2431 & ~n2669 ) | ( n2431 & n2668 ) | ( ~n2669 & n2668 ) ;
  assign n2672 = ( n2423 & ~n2671 ) | ( n2423 & n2670 ) | ( ~n2671 & n2670 ) ;
  assign n2673 = ( n150 & ~n2667 ) | ( n150 & n2672 ) | ( ~n2667 & n2672 ) ;
  assign n2674 = n2438 | n2457 ;
  assign n2675 = ( n2454 & ~n2472 ) | ( n2454 & n2674 ) | ( ~n2472 & n2674 ) ;
  assign n2676 = ( n2454 & ~n2675 ) | ( n2454 & 1'b0 ) | ( ~n2675 & 1'b0 ) ;
  assign n2677 = ( n2454 & ~n2457 ) | ( n2454 & 1'b0 ) | ( ~n2457 & 1'b0 ) ;
  assign n2678 = ~n2472 & n2677 ;
  assign n2679 = ( n2438 & ~n2677 ) | ( n2438 & n2678 ) | ( ~n2677 & n2678 ) ;
  assign n2680 = n2676 | n2679 ;
  assign n2681 = ( n2439 & ~n2446 ) | ( n2439 & 1'b0 ) | ( ~n2446 & 1'b0 ) ;
  assign n2682 = ~n2472 & n2681 ;
  assign n2683 = ( n2460 & ~n2682 ) | ( n2460 & n2681 ) | ( ~n2682 & n2681 ) ;
  assign n2684 = ( n2680 & ~n2683 ) | ( n2680 & 1'b0 ) | ( ~n2683 & 1'b0 ) ;
  assign n2685 = ~n2673 & n2684 ;
  assign n2686 = ( n133 & ~n2685 ) | ( n133 & n2684 ) | ( ~n2685 & n2684 ) ;
  assign n2687 = n150 | n2652 ;
  assign n2688 = ( n2666 & ~n2687 ) | ( n2666 & 1'b0 ) | ( ~n2687 & 1'b0 ) ;
  assign n2693 = n2688 &  n2672 ;
  assign n2689 = n2660 | n2663 ;
  assign n2690 = ( n145 & ~n2689 ) | ( n145 & n2657 ) | ( ~n2689 & n2657 ) ;
  assign n2691 = ( n150 & ~n2690 ) | ( n150 & 1'b0 ) | ( ~n2690 & 1'b0 ) ;
  assign n2692 = n2680 | n2691 ;
  assign n2694 = ( n2672 & ~n2693 ) | ( n2672 & n2692 ) | ( ~n2693 & n2692 ) ;
  assign n2696 = ( n133 & ~n2446 ) | ( n133 & n2439 ) | ( ~n2446 & n2439 ) ;
  assign n2695 = ( n2446 & ~n2439 ) | ( n2446 & n2472 ) | ( ~n2439 & n2472 ) ;
  assign n2697 = ~n2446 & n2695 ;
  assign n2698 = ( n2446 & n2696 ) | ( n2446 & n2697 ) | ( n2696 & n2697 ) ;
  assign n2699 = n2442 | n2469 ;
  assign n2700 = ( n2445 & n2464 ) | ( n2445 & n2699 ) | ( n2464 & n2699 ) ;
  assign n2701 = ( n2445 & ~n2700 ) | ( n2445 & 1'b0 ) | ( ~n2700 & 1'b0 ) ;
  assign n2702 = ( n2452 & ~n2701 ) | ( n2452 & n2460 ) | ( ~n2701 & n2460 ) ;
  assign n2703 = ( n2452 & ~n2702 ) | ( n2452 & 1'b0 ) | ( ~n2702 & 1'b0 ) ;
  assign n2704 = n2698 | n2703 ;
  assign n2705 = ( n2694 & ~n2704 ) | ( n2694 & 1'b0 ) | ( ~n2704 & 1'b0 ) ;
  assign n2706 = ~n2686 | ~n2705 ;
  assign n2902 = n2663 | n2706 ;
  assign n2903 = ( n2650 & n2659 ) | ( n2650 & n2663 ) | ( n2659 & n2663 ) ;
  assign n2904 = ( n2902 & ~n2659 ) | ( n2902 & n2903 ) | ( ~n2659 & n2903 ) ;
  assign n2905 = ( n2663 & ~n2903 ) | ( n2663 & n2902 ) | ( ~n2903 & n2902 ) ;
  assign n2906 = ( n2650 & ~n2904 ) | ( n2650 & n2905 ) | ( ~n2904 & n2905 ) ;
  assign n2895 = ~n2643 & n2706 ;
  assign n2896 = ( n2630 & ~n2895 ) | ( n2630 & n2706 ) | ( ~n2895 & n2706 ) ;
  assign n2897 = ( n2630 & ~n2896 ) | ( n2630 & n2635 ) | ( ~n2896 & n2635 ) ;
  assign n2898 = ( n2635 & ~n2630 ) | ( n2635 & n2896 ) | ( ~n2630 & n2896 ) ;
  assign n2899 = ( n2897 & ~n2635 ) | ( n2897 & n2898 ) | ( ~n2635 & n2898 ) ;
  assign n2880 = n2641 | n2706 ;
  assign n2881 = ( n2628 & n2637 ) | ( n2628 & n2641 ) | ( n2637 & n2641 ) ;
  assign n2882 = ( n2880 & ~n2637 ) | ( n2880 & n2881 ) | ( ~n2637 & n2881 ) ;
  assign n2883 = ( n2641 & ~n2881 ) | ( n2641 & n2880 ) | ( ~n2881 & n2880 ) ;
  assign n2884 = ( n2628 & ~n2882 ) | ( n2628 & n2883 ) | ( ~n2882 & n2883 ) ;
  assign n2873 = ~n2621 & n2706 ;
  assign n2874 = ( n2608 & ~n2873 ) | ( n2608 & n2706 ) | ( ~n2873 & n2706 ) ;
  assign n2875 = ( n2613 & ~n2608 ) | ( n2613 & n2874 ) | ( ~n2608 & n2874 ) ;
  assign n2876 = ( n2608 & ~n2874 ) | ( n2608 & n2613 ) | ( ~n2874 & n2613 ) ;
  assign n2877 = ( n2875 & ~n2613 ) | ( n2875 & n2876 ) | ( ~n2613 & n2876 ) ;
  assign n2858 = n2619 | n2706 ;
  assign n2859 = ( n2606 & n2615 ) | ( n2606 & n2619 ) | ( n2615 & n2619 ) ;
  assign n2860 = ( n2858 & ~n2615 ) | ( n2858 & n2859 ) | ( ~n2615 & n2859 ) ;
  assign n2861 = ( n2619 & ~n2859 ) | ( n2619 & n2858 ) | ( ~n2859 & n2858 ) ;
  assign n2862 = ( n2606 & ~n2860 ) | ( n2606 & n2861 ) | ( ~n2860 & n2861 ) ;
  assign n2851 = n2599 &  n2706 ;
  assign n2852 = ( n2586 & ~n2851 ) | ( n2586 & n2706 ) | ( ~n2851 & n2706 ) ;
  assign n2853 = ( n2586 & ~n2852 ) | ( n2586 & n2591 ) | ( ~n2852 & n2591 ) ;
  assign n2854 = ( n2591 & ~n2586 ) | ( n2591 & n2852 ) | ( ~n2586 & n2852 ) ;
  assign n2855 = ( n2853 & ~n2591 ) | ( n2853 & n2854 ) | ( ~n2591 & n2854 ) ;
  assign n2836 = n2597 | n2706 ;
  assign n2837 = ( n2584 & ~n2597 ) | ( n2584 & n2593 ) | ( ~n2597 & n2593 ) ;
  assign n2839 = ( n2597 & n2836 ) | ( n2597 & n2837 ) | ( n2836 & n2837 ) ;
  assign n2838 = ( n2593 & ~n2837 ) | ( n2593 & n2836 ) | ( ~n2837 & n2836 ) ;
  assign n2840 = ( n2584 & ~n2839 ) | ( n2584 & n2838 ) | ( ~n2839 & n2838 ) ;
  assign n2830 = ( n2565 & ~n2573 ) | ( n2565 & n2577 ) | ( ~n2573 & n2577 ) ;
  assign n2832 = ( n2573 & n2706 ) | ( n2573 & n2830 ) | ( n2706 & n2830 ) ;
  assign n2831 = ( n2565 & ~n2830 ) | ( n2565 & n2706 ) | ( ~n2830 & n2706 ) ;
  assign n2833 = ( n2577 & ~n2832 ) | ( n2577 & n2831 ) | ( ~n2832 & n2831 ) ;
  assign n2816 = ( n2567 & ~n2563 ) | ( n2567 & n2571 ) | ( ~n2563 & n2571 ) ;
  assign n2815 = ( n2571 & ~n2706 ) | ( n2571 & 1'b0 ) | ( ~n2706 & 1'b0 ) ;
  assign n2818 = ( n2571 & ~n2816 ) | ( n2571 & n2815 ) | ( ~n2816 & n2815 ) ;
  assign n2817 = ( n2815 & ~n2567 ) | ( n2815 & n2816 ) | ( ~n2567 & n2816 ) ;
  assign n2819 = ( n2563 & ~n2818 ) | ( n2563 & n2817 ) | ( ~n2818 & n2817 ) ;
  assign n2808 = n2543 | n2706 ;
  assign n2809 = ( n2548 & ~n2543 ) | ( n2548 & n2556 ) | ( ~n2543 & n2556 ) ;
  assign n2811 = ( n2543 & n2808 ) | ( n2543 & n2809 ) | ( n2808 & n2809 ) ;
  assign n2810 = ( n2556 & ~n2809 ) | ( n2556 & n2808 ) | ( ~n2809 & n2808 ) ;
  assign n2812 = ( n2548 & ~n2811 ) | ( n2548 & n2810 ) | ( ~n2811 & n2810 ) ;
  assign n2793 = n2554 | n2706 ;
  assign n2794 = ( n2541 & ~n2554 ) | ( n2541 & n2550 ) | ( ~n2554 & n2550 ) ;
  assign n2796 = ( n2554 & n2793 ) | ( n2554 & n2794 ) | ( n2793 & n2794 ) ;
  assign n2795 = ( n2550 & ~n2794 ) | ( n2550 & n2793 ) | ( ~n2794 & n2793 ) ;
  assign n2797 = ( n2541 & ~n2796 ) | ( n2541 & n2795 ) | ( ~n2796 & n2795 ) ;
  assign n2786 = n2534 &  n2706 ;
  assign n2787 = ( n2521 & ~n2706 ) | ( n2521 & n2786 ) | ( ~n2706 & n2786 ) ;
  assign n2788 = ( n2526 & ~n2521 ) | ( n2526 & n2787 ) | ( ~n2521 & n2787 ) ;
  assign n2789 = ( n2521 & ~n2787 ) | ( n2521 & n2526 ) | ( ~n2787 & n2526 ) ;
  assign n2790 = ( n2788 & ~n2526 ) | ( n2788 & n2789 ) | ( ~n2526 & n2789 ) ;
  assign n2771 = ( n2532 & ~n2706 ) | ( n2532 & 1'b0 ) | ( ~n2706 & 1'b0 ) ;
  assign n2772 = ( n2519 & n2528 ) | ( n2519 & n2532 ) | ( n2528 & n2532 ) ;
  assign n2773 = ( n2771 & ~n2528 ) | ( n2771 & n2772 ) | ( ~n2528 & n2772 ) ;
  assign n2774 = ( n2532 & ~n2772 ) | ( n2532 & n2771 ) | ( ~n2772 & n2771 ) ;
  assign n2775 = ( n2519 & ~n2773 ) | ( n2519 & n2774 ) | ( ~n2773 & n2774 ) ;
  assign n2764 = n2495 | n2706 ;
  assign n2765 = ( n2495 & ~n2512 ) | ( n2495 & n2505 ) | ( ~n2512 & n2505 ) ;
  assign n2766 = ( n2512 & n2764 ) | ( n2512 & n2765 ) | ( n2764 & n2765 ) ;
  assign n2767 = ( n2495 & ~n2765 ) | ( n2495 & n2764 ) | ( ~n2765 & n2764 ) ;
  assign n2768 = ( n2505 & ~n2766 ) | ( n2505 & n2767 ) | ( ~n2766 & n2767 ) ;
  assign n2749 = n2507 | n2510 ;
  assign n2750 = ( n2507 & n2706 ) | ( n2507 & n2749 ) | ( n2706 & n2749 ) ;
  assign n2751 = ( n2493 & ~n2507 ) | ( n2493 & n2750 ) | ( ~n2507 & n2750 ) ;
  assign n2752 = ( n2493 & ~n2750 ) | ( n2493 & n2507 ) | ( ~n2750 & n2507 ) ;
  assign n2753 = ( n2751 & ~n2493 ) | ( n2751 & n2752 ) | ( ~n2493 & n2752 ) ;
  assign n2740 = ~x88 & n2472 ;
  assign n2741 = ( x89 & ~n2740 ) | ( x89 & 1'b0 ) | ( ~n2740 & 1'b0 ) ;
  assign n2742 = n2484 | n2741 ;
  assign n2737 = ( n2472 & ~x88 ) | ( n2472 & n2479 ) | ( ~x88 & n2479 ) ;
  assign n2738 = x88 &  n2737 ;
  assign n2739 = ( n2474 & ~n2738 ) | ( n2474 & n2479 ) | ( ~n2738 & n2479 ) ;
  assign n2743 = ( n2706 & ~n2742 ) | ( n2706 & n2739 ) | ( ~n2742 & n2739 ) ;
  assign n2745 = ( n2706 & ~n2743 ) | ( n2706 & 1'b0 ) | ( ~n2743 & 1'b0 ) ;
  assign n2744 = ~n2739 & n2743 ;
  assign n2746 = ( n2742 & ~n2745 ) | ( n2742 & n2744 ) | ( ~n2745 & n2744 ) ;
  assign n2713 = ( x86 & ~n2706 ) | ( x86 & x87 ) | ( ~n2706 & x87 ) ;
  assign n2719 = ( x86 & ~x87 ) | ( x86 & 1'b0 ) | ( ~x87 & 1'b0 ) ;
  assign n2709 = x84 | x85 ;
  assign n2714 = ~x86 & n2709 ;
  assign n2715 = ( x86 & ~n2470 ) | ( x86 & n2714 ) | ( ~n2470 & n2714 ) ;
  assign n2716 = ( n2452 & ~n2715 ) | ( n2452 & n2460 ) | ( ~n2715 & n2460 ) ;
  assign n2717 = ( n2452 & ~n2716 ) | ( n2452 & 1'b0 ) | ( ~n2716 & 1'b0 ) ;
  assign n2718 = ( n2706 & ~x87 ) | ( n2706 & n2717 ) | ( ~x87 & n2717 ) ;
  assign n2720 = ( n2713 & ~n2719 ) | ( n2713 & n2718 ) | ( ~n2719 & n2718 ) ;
  assign n2710 = x86 | n2709 ;
  assign n2711 = x86 &  n2706 ;
  assign n2712 = ( n2472 & ~n2710 ) | ( n2472 & n2711 ) | ( ~n2710 & n2711 ) ;
  assign n2723 = n2245 | n2712 ;
  assign n2724 = ( n2720 & ~n2723 ) | ( n2720 & 1'b0 ) | ( ~n2723 & 1'b0 ) ;
  assign n2726 = ( n2472 & ~n2703 ) | ( n2472 & 1'b0 ) | ( ~n2703 & 1'b0 ) ;
  assign n2727 = ( n2694 & ~n2726 ) | ( n2694 & n2698 ) | ( ~n2726 & n2698 ) ;
  assign n2728 = ( n2694 & ~n2727 ) | ( n2694 & 1'b0 ) | ( ~n2727 & 1'b0 ) ;
  assign n2729 = n2686 &  n2728 ;
  assign n2725 = ~n2246 & n2706 ;
  assign n2730 = ( n2725 & ~n2729 ) | ( n2725 & 1'b0 ) | ( ~n2729 & 1'b0 ) ;
  assign n2731 = ( x88 & n2729 ) | ( x88 & n2730 ) | ( n2729 & n2730 ) ;
  assign n2732 = x88 | n2729 ;
  assign n2733 = n2725 | n2732 ;
  assign n2734 = ~n2731 & n2733 ;
  assign n2735 = n2724 | n2734 ;
  assign n2721 = n2712 &  n2720 ;
  assign n2722 = ( n2245 & ~n2720 ) | ( n2245 & n2721 ) | ( ~n2720 & n2721 ) ;
  assign n2754 = ( n2033 & ~n2722 ) | ( n2033 & 1'b0 ) | ( ~n2722 & 1'b0 ) ;
  assign n2755 = n2735 &  n2754 ;
  assign n2756 = n2746 | n2755 ;
  assign n2757 = ~n2712 & n2720 ;
  assign n2758 = ( n2734 & ~n2245 ) | ( n2734 & n2757 ) | ( ~n2245 & n2757 ) ;
  assign n2759 = n2033 | n2758 ;
  assign n2760 = ~n1827 & n2759 ;
  assign n2761 = n2756 &  n2760 ;
  assign n2762 = n2753 | n2761 ;
  assign n2736 = ~n2722 & n2735 ;
  assign n2747 = ( n2033 & n2736 ) | ( n2033 & n2746 ) | ( n2736 & n2746 ) ;
  assign n2748 = ( n1827 & ~n2747 ) | ( n1827 & 1'b0 ) | ( ~n2747 & 1'b0 ) ;
  assign n2776 = ( n1636 & ~n2748 ) | ( n1636 & 1'b0 ) | ( ~n2748 & 1'b0 ) ;
  assign n2777 = n2762 &  n2776 ;
  assign n2778 = n2768 | n2777 ;
  assign n2779 = n2756 &  n2759 ;
  assign n2780 = ( n2753 & ~n1827 ) | ( n2753 & n2779 ) | ( ~n1827 & n2779 ) ;
  assign n2781 = n1636 | n2780 ;
  assign n2782 = n1452 &  n2781 ;
  assign n2783 = n2778 &  n2782 ;
  assign n2784 = n2775 | n2783 ;
  assign n2763 = ~n2748 & n2762 ;
  assign n2769 = ( n1636 & n2763 ) | ( n1636 & n2768 ) | ( n2763 & n2768 ) ;
  assign n2770 = n1452 | n2769 ;
  assign n2798 = ~n1283 & n2770 ;
  assign n2799 = n2784 &  n2798 ;
  assign n2800 = ( n2790 & ~n2799 ) | ( n2790 & 1'b0 ) | ( ~n2799 & 1'b0 ) ;
  assign n2801 = n2778 &  n2781 ;
  assign n2802 = ( n1452 & n2775 ) | ( n1452 & n2801 ) | ( n2775 & n2801 ) ;
  assign n2803 = ( n1283 & ~n2802 ) | ( n1283 & 1'b0 ) | ( ~n2802 & 1'b0 ) ;
  assign n2804 = ( n1122 & ~n2803 ) | ( n1122 & 1'b0 ) | ( ~n2803 & 1'b0 ) ;
  assign n2805 = ~n2800 & n2804 ;
  assign n2806 = ( n2797 & ~n2805 ) | ( n2797 & 1'b0 ) | ( ~n2805 & 1'b0 ) ;
  assign n2785 = n2770 &  n2784 ;
  assign n2791 = ( n1283 & ~n2785 ) | ( n1283 & n2790 ) | ( ~n2785 & n2790 ) ;
  assign n2792 = ~n1122 & n2791 ;
  assign n2820 = ( n976 & ~n2792 ) | ( n976 & 1'b0 ) | ( ~n2792 & 1'b0 ) ;
  assign n2821 = ~n2806 & n2820 ;
  assign n2822 = n2812 | n2821 ;
  assign n2823 = n2800 | n2803 ;
  assign n2824 = ( n2797 & ~n1122 ) | ( n2797 & n2823 ) | ( ~n1122 & n2823 ) ;
  assign n2825 = ~n976 & n2824 ;
  assign n2826 = n837 | n2825 ;
  assign n2827 = ( n2822 & ~n2826 ) | ( n2822 & 1'b0 ) | ( ~n2826 & 1'b0 ) ;
  assign n2828 = n2819 | n2827 ;
  assign n2807 = n2792 | n2806 ;
  assign n2813 = ( n976 & ~n2807 ) | ( n976 & n2812 ) | ( ~n2807 & n2812 ) ;
  assign n2814 = ( n837 & ~n2813 ) | ( n837 & 1'b0 ) | ( ~n2813 & 1'b0 ) ;
  assign n2841 = n713 | n2814 ;
  assign n2842 = ( n2828 & ~n2841 ) | ( n2828 & 1'b0 ) | ( ~n2841 & 1'b0 ) ;
  assign n2843 = n2833 | n2842 ;
  assign n2844 = ( n2822 & ~n2825 ) | ( n2822 & 1'b0 ) | ( ~n2825 & 1'b0 ) ;
  assign n2845 = ( n2819 & ~n837 ) | ( n2819 & n2844 ) | ( ~n837 & n2844 ) ;
  assign n2846 = ( n713 & ~n2845 ) | ( n713 & 1'b0 ) | ( ~n2845 & 1'b0 ) ;
  assign n2847 = n595 | n2846 ;
  assign n2848 = ( n2843 & ~n2847 ) | ( n2843 & 1'b0 ) | ( ~n2847 & 1'b0 ) ;
  assign n2849 = n2840 | n2848 ;
  assign n2829 = ~n2814 & n2828 ;
  assign n2834 = ( n2829 & ~n713 ) | ( n2829 & n2833 ) | ( ~n713 & n2833 ) ;
  assign n2835 = ( n595 & ~n2834 ) | ( n595 & 1'b0 ) | ( ~n2834 & 1'b0 ) ;
  assign n2863 = n492 | n2835 ;
  assign n2864 = ( n2849 & ~n2863 ) | ( n2849 & 1'b0 ) | ( ~n2863 & 1'b0 ) ;
  assign n2865 = ( n2855 & ~n2864 ) | ( n2855 & 1'b0 ) | ( ~n2864 & 1'b0 ) ;
  assign n2866 = ( n2843 & ~n2846 ) | ( n2843 & 1'b0 ) | ( ~n2846 & 1'b0 ) ;
  assign n2867 = ( n2840 & ~n595 ) | ( n2840 & n2866 ) | ( ~n595 & n2866 ) ;
  assign n2868 = ( n492 & ~n2867 ) | ( n492 & 1'b0 ) | ( ~n2867 & 1'b0 ) ;
  assign n2869 = n396 | n2868 ;
  assign n2870 = n2865 | n2869 ;
  assign n2871 = n2862 &  n2870 ;
  assign n2850 = ~n2835 & n2849 ;
  assign n2856 = ( n492 & ~n2850 ) | ( n492 & n2855 ) | ( ~n2850 & n2855 ) ;
  assign n2857 = n396 &  n2856 ;
  assign n2885 = n315 | n2857 ;
  assign n2886 = n2871 | n2885 ;
  assign n2887 = ~n2877 & n2886 ;
  assign n2888 = n2865 | n2868 ;
  assign n2889 = ( n396 & n2862 ) | ( n396 & n2888 ) | ( n2862 & n2888 ) ;
  assign n2890 = n315 &  n2889 ;
  assign n2891 = n240 | n2890 ;
  assign n2892 = n2887 | n2891 ;
  assign n2893 = n2884 &  n2892 ;
  assign n2872 = n2857 | n2871 ;
  assign n2878 = ( n315 & ~n2877 ) | ( n315 & n2872 ) | ( ~n2877 & n2872 ) ;
  assign n2879 = n240 &  n2878 ;
  assign n2907 = n181 | n2879 ;
  assign n2908 = n2893 | n2907 ;
  assign n2909 = n2899 &  n2908 ;
  assign n2910 = n2887 | n2890 ;
  assign n2911 = ( n240 & n2884 ) | ( n240 & n2910 ) | ( n2884 & n2910 ) ;
  assign n2912 = n181 &  n2911 ;
  assign n2913 = ( n145 & ~n2912 ) | ( n145 & 1'b0 ) | ( ~n2912 & 1'b0 ) ;
  assign n2914 = ~n2909 & n2913 ;
  assign n2915 = n2906 | n2914 ;
  assign n2894 = n2879 | n2893 ;
  assign n2900 = ( n181 & n2894 ) | ( n181 & n2899 ) | ( n2894 & n2899 ) ;
  assign n2901 = ~n145 & n2900 ;
  assign n2936 = n150 | n2901 ;
  assign n2937 = ( n2915 & ~n2936 ) | ( n2915 & 1'b0 ) | ( ~n2936 & 1'b0 ) ;
  assign n2916 = ~n2901 & n2915 ;
  assign n2917 = n2652 | n2706 ;
  assign n2918 = ( n2652 & ~n2665 ) | ( n2652 & n2657 ) | ( ~n2665 & n2657 ) ;
  assign n2919 = ( n2665 & n2917 ) | ( n2665 & n2918 ) | ( n2917 & n2918 ) ;
  assign n2920 = ( n2652 & ~n2918 ) | ( n2652 & n2917 ) | ( ~n2918 & n2917 ) ;
  assign n2921 = ( n2657 & ~n2919 ) | ( n2657 & n2920 ) | ( ~n2919 & n2920 ) ;
  assign n2922 = ( n2916 & ~n150 ) | ( n2916 & n2921 ) | ( ~n150 & n2921 ) ;
  assign n2923 = n2672 | n2688 ;
  assign n2924 = ( n2691 & ~n2923 ) | ( n2691 & n2706 ) | ( ~n2923 & n2706 ) ;
  assign n2925 = ~n2691 & n2924 ;
  assign n2926 = n2688 | n2691 ;
  assign n2927 = n2706 | n2926 ;
  assign n2928 = ( n2672 & ~n2927 ) | ( n2672 & n2926 ) | ( ~n2927 & n2926 ) ;
  assign n2929 = n2925 | n2928 ;
  assign n2930 = n2673 &  n2680 ;
  assign n2931 = ~n2706 & n2930 ;
  assign n2932 = ( n2694 & ~n2930 ) | ( n2694 & n2931 ) | ( ~n2930 & n2931 ) ;
  assign n2933 = n2929 &  n2932 ;
  assign n2934 = n2922 &  n2933 ;
  assign n2935 = ( n133 & ~n2934 ) | ( n133 & n2933 ) | ( ~n2934 & n2933 ) ;
  assign n2938 = n2909 | n2912 ;
  assign n2939 = ( n145 & ~n2938 ) | ( n145 & n2906 ) | ( ~n2938 & n2906 ) ;
  assign n2940 = ( n150 & ~n2939 ) | ( n150 & 1'b0 ) | ( ~n2939 & 1'b0 ) ;
  assign n2941 = n2929 | n2940 ;
  assign n2942 = ~n2921 & n2937 ;
  assign n2943 = ( n2921 & ~n2941 ) | ( n2921 & n2942 ) | ( ~n2941 & n2942 ) ;
  assign n2945 = ( n133 & n2673 ) | ( n133 & n2680 ) | ( n2673 & n2680 ) ;
  assign n2944 = ( n2673 & ~n2706 ) | ( n2673 & n2680 ) | ( ~n2706 & n2680 ) ;
  assign n2946 = ( n2680 & ~n2944 ) | ( n2680 & 1'b0 ) | ( ~n2944 & 1'b0 ) ;
  assign n2947 = ( n2945 & ~n2680 ) | ( n2945 & n2946 ) | ( ~n2680 & n2946 ) ;
  assign n2948 = n2676 | n2703 ;
  assign n2949 = ( n2698 & ~n2679 ) | ( n2698 & n2948 ) | ( ~n2679 & n2948 ) ;
  assign n2950 = n2679 | n2949 ;
  assign n2951 = ( n2686 & ~n2694 ) | ( n2686 & n2950 ) | ( ~n2694 & n2950 ) ;
  assign n2952 = ( n2686 & ~n2951 ) | ( n2686 & 1'b0 ) | ( ~n2951 & 1'b0 ) ;
  assign n2953 = n2947 | n2952 ;
  assign n2954 = n2943 | n2953 ;
  assign n2955 = ~n2935 |  n2954 ;
  assign n3179 = ( n2921 & ~n2940 ) | ( n2921 & 1'b0 ) | ( ~n2940 & 1'b0 ) ;
  assign n3180 = ( n2937 & n2955 ) | ( n2937 & n3179 ) | ( n2955 & n3179 ) ;
  assign n3181 = ~n2937 & n3180 ;
  assign n3182 = n2937 | n2940 ;
  assign n3183 = n2955 | n3182 ;
  assign n3184 = ( n2921 & ~n3182 ) | ( n2921 & n3183 ) | ( ~n3182 & n3183 ) ;
  assign n3185 = ~n3181 & n3184 ;
  assign n3186 = ~n2922 & n2929 ;
  assign n3187 = ~n2955 & n3186 ;
  assign n3188 = ( n2943 & ~n3187 ) | ( n2943 & n3186 ) | ( ~n3187 & n3186 ) ;
  assign n3189 = n3185 | n3188 ;
  assign n3173 = n2901 | n2955 ;
  assign n3174 = ( n2901 & ~n2914 ) | ( n2901 & n2906 ) | ( ~n2914 & n2906 ) ;
  assign n3175 = ( n2914 & n3173 ) | ( n2914 & n3174 ) | ( n3173 & n3174 ) ;
  assign n3176 = ( n2901 & ~n3174 ) | ( n2901 & n3173 ) | ( ~n3174 & n3173 ) ;
  assign n3177 = ( n2906 & ~n3175 ) | ( n2906 & n3176 ) | ( ~n3175 & n3176 ) ;
  assign n3064 = n2805 &  n2955 ;
  assign n3065 = ( n2792 & ~n3064 ) | ( n2792 & n2955 ) | ( ~n3064 & n2955 ) ;
  assign n3066 = ( n2792 & ~n3065 ) | ( n2792 & n2797 ) | ( ~n3065 & n2797 ) ;
  assign n3067 = ( n2797 & ~n2792 ) | ( n2797 & n3065 ) | ( ~n2792 & n3065 ) ;
  assign n3068 = ( n3066 & ~n2797 ) | ( n3066 & n3067 ) | ( ~n2797 & n3067 ) ;
  assign n2708 = x84 | n2707 ;
  assign n2956 = x84 &  n2955 ;
  assign n2957 = ( n2706 & ~n2708 ) | ( n2706 & n2956 ) | ( ~n2708 & n2956 ) ;
  assign n2958 = ( x84 & ~n2955 ) | ( x84 & x85 ) | ( ~n2955 & x85 ) ;
  assign n2964 = ( x84 & ~x85 ) | ( x84 & 1'b0 ) | ( ~x85 & 1'b0 ) ;
  assign n2959 = ~x84 & n2707 ;
  assign n2960 = ( x84 & ~n2704 ) | ( x84 & n2959 ) | ( ~n2704 & n2959 ) ;
  assign n2961 = ( n2694 & ~n2686 ) | ( n2694 & n2960 ) | ( ~n2686 & n2960 ) ;
  assign n2962 = n2686 &  n2961 ;
  assign n2963 = ( n2955 & ~x85 ) | ( n2955 & n2962 ) | ( ~x85 & n2962 ) ;
  assign n2965 = ( n2958 & ~n2964 ) | ( n2958 & n2963 ) | ( ~n2964 & n2963 ) ;
  assign n2966 = ~n2957 & n2965 ;
  assign n2968 = ( n2706 & ~n2952 ) | ( n2706 & 1'b0 ) | ( ~n2952 & 1'b0 ) ;
  assign n2969 = ( n2943 & ~n2947 ) | ( n2943 & n2968 ) | ( ~n2947 & n2968 ) ;
  assign n2970 = ~n2943 & n2969 ;
  assign n2971 = n2935 &  n2970 ;
  assign n2967 = ~n2709 & n2955 ;
  assign n2972 = ( n2967 & ~n2971 ) | ( n2967 & 1'b0 ) | ( ~n2971 & 1'b0 ) ;
  assign n2973 = ( x86 & n2971 ) | ( x86 & n2972 ) | ( n2971 & n2972 ) ;
  assign n2974 = x86 | n2971 ;
  assign n2975 = n2967 | n2974 ;
  assign n2976 = ~n2973 & n2975 ;
  assign n2977 = ( n2966 & ~n2472 ) | ( n2966 & n2976 ) | ( ~n2472 & n2976 ) ;
  assign n2978 = ( n2245 & ~n2977 ) | ( n2245 & 1'b0 ) | ( ~n2977 & 1'b0 ) ;
  assign n2982 = ~x86 & n2706 ;
  assign n2983 = ( x87 & ~n2982 ) | ( x87 & 1'b0 ) | ( ~n2982 & 1'b0 ) ;
  assign n2984 = n2725 | n2983 ;
  assign n2979 = ( n2706 & ~x86 ) | ( n2706 & n2717 ) | ( ~x86 & n2717 ) ;
  assign n2980 = x86 &  n2979 ;
  assign n2981 = ( n2712 & ~n2980 ) | ( n2712 & n2717 ) | ( ~n2980 & n2717 ) ;
  assign n2985 = ( n2955 & ~n2984 ) | ( n2955 & n2981 ) | ( ~n2984 & n2981 ) ;
  assign n2987 = ( n2955 & ~n2985 ) | ( n2955 & 1'b0 ) | ( ~n2985 & 1'b0 ) ;
  assign n2986 = ~n2981 & n2985 ;
  assign n2988 = ( n2984 & ~n2987 ) | ( n2984 & n2986 ) | ( ~n2987 & n2986 ) ;
  assign n2989 = n2472 | n2957 ;
  assign n2990 = ( n2965 & ~n2989 ) | ( n2965 & 1'b0 ) | ( ~n2989 & 1'b0 ) ;
  assign n2991 = n2976 | n2990 ;
  assign n2992 = n2957 &  n2965 ;
  assign n2993 = ( n2472 & ~n2965 ) | ( n2472 & n2992 ) | ( ~n2965 & n2992 ) ;
  assign n2994 = n2245 | n2993 ;
  assign n2995 = ( n2991 & ~n2994 ) | ( n2991 & 1'b0 ) | ( ~n2994 & 1'b0 ) ;
  assign n2996 = n2988 | n2995 ;
  assign n2997 = ~n2978 & n2996 ;
  assign n2998 = ( n2722 & ~n2724 ) | ( n2722 & 1'b0 ) | ( ~n2724 & 1'b0 ) ;
  assign n2999 = ( n2724 & ~n2998 ) | ( n2724 & n2734 ) | ( ~n2998 & n2734 ) ;
  assign n3001 = ( n2955 & n2998 ) | ( n2955 & n2999 ) | ( n2998 & n2999 ) ;
  assign n3000 = ( n2724 & ~n2999 ) | ( n2724 & n2955 ) | ( ~n2999 & n2955 ) ;
  assign n3002 = ( n2734 & ~n3001 ) | ( n2734 & n3000 ) | ( ~n3001 & n3000 ) ;
  assign n3003 = ( n2033 & n2997 ) | ( n2033 & n3002 ) | ( n2997 & n3002 ) ;
  assign n3004 = ( n1827 & ~n3003 ) | ( n1827 & 1'b0 ) | ( ~n3003 & 1'b0 ) ;
  assign n3006 = ( n2755 & ~n2746 ) | ( n2755 & n2759 ) | ( ~n2746 & n2759 ) ;
  assign n3005 = ( n2759 & ~n2955 ) | ( n2759 & 1'b0 ) | ( ~n2955 & 1'b0 ) ;
  assign n3008 = ( n2759 & ~n3006 ) | ( n2759 & n3005 ) | ( ~n3006 & n3005 ) ;
  assign n3007 = ( n3005 & ~n2755 ) | ( n3005 & n3006 ) | ( ~n2755 & n3006 ) ;
  assign n3009 = ( n2746 & ~n3008 ) | ( n2746 & n3007 ) | ( ~n3008 & n3007 ) ;
  assign n3010 = ( n2033 & ~n2978 ) | ( n2033 & 1'b0 ) | ( ~n2978 & 1'b0 ) ;
  assign n3011 = n2996 &  n3010 ;
  assign n3012 = n3002 | n3011 ;
  assign n3013 = ( n2991 & ~n2993 ) | ( n2991 & 1'b0 ) | ( ~n2993 & 1'b0 ) ;
  assign n3014 = ( n2988 & ~n2245 ) | ( n2988 & n3013 ) | ( ~n2245 & n3013 ) ;
  assign n3015 = n2033 | n3014 ;
  assign n3016 = ~n1827 & n3015 ;
  assign n3017 = n3012 &  n3016 ;
  assign n3018 = n3009 | n3017 ;
  assign n3019 = ~n3004 & n3018 ;
  assign n3020 = n2748 | n2955 ;
  assign n3021 = ( n2753 & ~n2748 ) | ( n2753 & n2761 ) | ( ~n2748 & n2761 ) ;
  assign n3023 = ( n2748 & n3020 ) | ( n2748 & n3021 ) | ( n3020 & n3021 ) ;
  assign n3022 = ( n2761 & ~n3021 ) | ( n2761 & n3020 ) | ( ~n3021 & n3020 ) ;
  assign n3024 = ( n2753 & ~n3023 ) | ( n2753 & n3022 ) | ( ~n3023 & n3022 ) ;
  assign n3025 = ( n1636 & n3019 ) | ( n1636 & n3024 ) | ( n3019 & n3024 ) ;
  assign n3026 = n1452 | n3025 ;
  assign n3028 = ( n2777 & ~n2768 ) | ( n2777 & n2781 ) | ( ~n2768 & n2781 ) ;
  assign n3027 = ( n2781 & ~n2955 ) | ( n2781 & 1'b0 ) | ( ~n2955 & 1'b0 ) ;
  assign n3030 = ( n2781 & ~n3028 ) | ( n2781 & n3027 ) | ( ~n3028 & n3027 ) ;
  assign n3029 = ( n3027 & ~n2777 ) | ( n3027 & n3028 ) | ( ~n2777 & n3028 ) ;
  assign n3031 = ( n2768 & ~n3030 ) | ( n2768 & n3029 ) | ( ~n3030 & n3029 ) ;
  assign n3032 = ( n1636 & ~n3004 ) | ( n1636 & 1'b0 ) | ( ~n3004 & 1'b0 ) ;
  assign n3033 = n3018 &  n3032 ;
  assign n3034 = n3024 | n3033 ;
  assign n3035 = n3012 &  n3015 ;
  assign n3036 = ( n3009 & ~n1827 ) | ( n3009 & n3035 ) | ( ~n1827 & n3035 ) ;
  assign n3037 = n1636 | n3036 ;
  assign n3038 = n1452 &  n3037 ;
  assign n3039 = n3034 &  n3038 ;
  assign n3040 = n3031 | n3039 ;
  assign n3041 = n3026 &  n3040 ;
  assign n3043 = ( n2770 & ~n2775 ) | ( n2770 & n2783 ) | ( ~n2775 & n2783 ) ;
  assign n3042 = ( n2770 & ~n2955 ) | ( n2770 & 1'b0 ) | ( ~n2955 & 1'b0 ) ;
  assign n3045 = ( n2770 & ~n3043 ) | ( n2770 & n3042 ) | ( ~n3043 & n3042 ) ;
  assign n3044 = ( n3042 & ~n2783 ) | ( n3042 & n3043 ) | ( ~n2783 & n3043 ) ;
  assign n3046 = ( n2775 & ~n3045 ) | ( n2775 & n3044 ) | ( ~n3045 & n3044 ) ;
  assign n3047 = ( n3041 & ~n1283 ) | ( n3041 & n3046 ) | ( ~n1283 & n3046 ) ;
  assign n3048 = n1122 | n3047 ;
  assign n3049 = n2803 | n2955 ;
  assign n3050 = ( n2790 & ~n2799 ) | ( n2790 & n2803 ) | ( ~n2799 & n2803 ) ;
  assign n3051 = ( n2799 & n3049 ) | ( n2799 & n3050 ) | ( n3049 & n3050 ) ;
  assign n3052 = ( n2803 & ~n3050 ) | ( n2803 & n3049 ) | ( ~n3050 & n3049 ) ;
  assign n3053 = ( n2790 & ~n3051 ) | ( n2790 & n3052 ) | ( ~n3051 & n3052 ) ;
  assign n3054 = ~n1283 & n3026 ;
  assign n3055 = n3040 &  n3054 ;
  assign n3056 = n3046 | n3055 ;
  assign n3057 = n3034 &  n3037 ;
  assign n3058 = ( n1452 & n3031 ) | ( n1452 & n3057 ) | ( n3031 & n3057 ) ;
  assign n3059 = ( n1283 & ~n3058 ) | ( n1283 & 1'b0 ) | ( ~n3058 & 1'b0 ) ;
  assign n3060 = ( n1122 & ~n3059 ) | ( n1122 & 1'b0 ) | ( ~n3059 & 1'b0 ) ;
  assign n3061 = n3056 &  n3060 ;
  assign n3062 = ( n3053 & ~n3061 ) | ( n3053 & 1'b0 ) | ( ~n3061 & 1'b0 ) ;
  assign n3063 = ( n3048 & ~n3062 ) | ( n3048 & 1'b0 ) | ( ~n3062 & 1'b0 ) ;
  assign n3069 = ( n976 & ~n3068 ) | ( n976 & n3063 ) | ( ~n3068 & n3063 ) ;
  assign n3070 = ( n837 & ~n3069 ) | ( n837 & 1'b0 ) | ( ~n3069 & 1'b0 ) ;
  assign n3071 = n2825 | n2955 ;
  assign n3072 = ( n2812 & ~n2821 ) | ( n2812 & n2825 ) | ( ~n2821 & n2825 ) ;
  assign n3073 = ( n2821 & n3071 ) | ( n2821 & n3072 ) | ( n3071 & n3072 ) ;
  assign n3074 = ( n2825 & ~n3072 ) | ( n2825 & n3071 ) | ( ~n3072 & n3071 ) ;
  assign n3075 = ( n2812 & ~n3073 ) | ( n2812 & n3074 ) | ( ~n3073 & n3074 ) ;
  assign n3076 = n976 &  n3048 ;
  assign n3077 = ~n3062 & n3076 ;
  assign n3078 = ( n3068 & ~n3077 ) | ( n3068 & 1'b0 ) | ( ~n3077 & 1'b0 ) ;
  assign n3079 = ( n3056 & ~n3059 ) | ( n3056 & 1'b0 ) | ( ~n3059 & 1'b0 ) ;
  assign n3080 = ( n1122 & ~n3053 ) | ( n1122 & n3079 ) | ( ~n3053 & n3079 ) ;
  assign n3081 = n976 | n3080 ;
  assign n3082 = ~n837 & n3081 ;
  assign n3083 = ~n3078 & n3082 ;
  assign n3084 = n3075 | n3083 ;
  assign n3085 = ~n3070 & n3084 ;
  assign n3086 = n2814 | n2955 ;
  assign n3087 = ( n2819 & ~n2814 ) | ( n2819 & n2827 ) | ( ~n2814 & n2827 ) ;
  assign n3089 = ( n2814 & n3086 ) | ( n2814 & n3087 ) | ( n3086 & n3087 ) ;
  assign n3088 = ( n2827 & ~n3087 ) | ( n2827 & n3086 ) | ( ~n3087 & n3086 ) ;
  assign n3090 = ( n2819 & ~n3089 ) | ( n2819 & n3088 ) | ( ~n3089 & n3088 ) ;
  assign n3091 = ( n3085 & ~n713 ) | ( n3085 & n3090 ) | ( ~n713 & n3090 ) ;
  assign n3092 = ( n595 & ~n3091 ) | ( n595 & 1'b0 ) | ( ~n3091 & 1'b0 ) ;
  assign n3093 = n713 | n3070 ;
  assign n3094 = ( n3084 & ~n3093 ) | ( n3084 & 1'b0 ) | ( ~n3093 & 1'b0 ) ;
  assign n3095 = n3090 | n3094 ;
  assign n3096 = ~n3078 & n3081 ;
  assign n3097 = ( n3075 & ~n837 ) | ( n3075 & n3096 ) | ( ~n837 & n3096 ) ;
  assign n3098 = ( n713 & ~n3097 ) | ( n713 & 1'b0 ) | ( ~n3097 & 1'b0 ) ;
  assign n3099 = n595 | n3098 ;
  assign n3100 = ( n3095 & ~n3099 ) | ( n3095 & 1'b0 ) | ( ~n3099 & 1'b0 ) ;
  assign n3101 = ( n2833 & ~n2842 ) | ( n2833 & n2846 ) | ( ~n2842 & n2846 ) ;
  assign n3102 = ( n2842 & n2955 ) | ( n2842 & n3101 ) | ( n2955 & n3101 ) ;
  assign n3103 = ( n2846 & ~n3101 ) | ( n2846 & n2955 ) | ( ~n3101 & n2955 ) ;
  assign n3104 = ( n2833 & ~n3102 ) | ( n2833 & n3103 ) | ( ~n3102 & n3103 ) ;
  assign n3105 = n3100 | n3104 ;
  assign n3106 = ~n3092 & n3105 ;
  assign n3108 = ( n2835 & ~n2840 ) | ( n2835 & n2955 ) | ( ~n2840 & n2955 ) ;
  assign n3107 = n2848 &  n2955 ;
  assign n3109 = ( n2955 & ~n3108 ) | ( n2955 & n3107 ) | ( ~n3108 & n3107 ) ;
  assign n3110 = ( n3107 & ~n2835 ) | ( n3107 & n3108 ) | ( ~n2835 & n3108 ) ;
  assign n3111 = ( n2840 & ~n3109 ) | ( n2840 & n3110 ) | ( ~n3109 & n3110 ) ;
  assign n3112 = ( n3106 & ~n492 ) | ( n3106 & n3111 ) | ( ~n492 & n3111 ) ;
  assign n3113 = ( n396 & ~n3112 ) | ( n396 & 1'b0 ) | ( ~n3112 & 1'b0 ) ;
  assign n3114 = n2868 | n2955 ;
  assign n3115 = ( n2855 & ~n2864 ) | ( n2855 & n2868 ) | ( ~n2864 & n2868 ) ;
  assign n3116 = ( n2864 & n3114 ) | ( n2864 & n3115 ) | ( n3114 & n3115 ) ;
  assign n3117 = ( n2868 & ~n3115 ) | ( n2868 & n3114 ) | ( ~n3115 & n3114 ) ;
  assign n3118 = ( n2855 & ~n3116 ) | ( n2855 & n3117 ) | ( ~n3116 & n3117 ) ;
  assign n3119 = n492 | n3092 ;
  assign n3120 = ( n3105 & ~n3119 ) | ( n3105 & 1'b0 ) | ( ~n3119 & 1'b0 ) ;
  assign n3121 = n3111 | n3120 ;
  assign n3122 = ( n3095 & ~n3098 ) | ( n3095 & 1'b0 ) | ( ~n3098 & 1'b0 ) ;
  assign n3123 = ( n3104 & ~n595 ) | ( n3104 & n3122 ) | ( ~n595 & n3122 ) ;
  assign n3124 = ( n492 & ~n3123 ) | ( n492 & 1'b0 ) | ( ~n3123 & 1'b0 ) ;
  assign n3125 = n396 | n3124 ;
  assign n3126 = ( n3121 & ~n3125 ) | ( n3121 & 1'b0 ) | ( ~n3125 & 1'b0 ) ;
  assign n3127 = ( n3118 & ~n3126 ) | ( n3118 & 1'b0 ) | ( ~n3126 & 1'b0 ) ;
  assign n3128 = n3113 | n3127 ;
  assign n3129 = ~n2870 & n2955 ;
  assign n3130 = ( n2857 & ~n3129 ) | ( n2857 & n2955 ) | ( ~n3129 & n2955 ) ;
  assign n3131 = ( n2857 & ~n3130 ) | ( n2857 & n2862 ) | ( ~n3130 & n2862 ) ;
  assign n3132 = ( n2862 & ~n2857 ) | ( n2862 & n3130 ) | ( ~n2857 & n3130 ) ;
  assign n3133 = ( n3131 & ~n2862 ) | ( n3131 & n3132 ) | ( ~n2862 & n3132 ) ;
  assign n3134 = ( n315 & n3128 ) | ( n315 & n3133 ) | ( n3128 & n3133 ) ;
  assign n3135 = n240 &  n3134 ;
  assign n3137 = ( n2886 & ~n2877 ) | ( n2886 & n2890 ) | ( ~n2877 & n2890 ) ;
  assign n3136 = n2890 | n2955 ;
  assign n3139 = ( n2890 & ~n3137 ) | ( n2890 & n3136 ) | ( ~n3137 & n3136 ) ;
  assign n3138 = ( n3136 & ~n2886 ) | ( n3136 & n3137 ) | ( ~n2886 & n3137 ) ;
  assign n3140 = ( n2877 & ~n3139 ) | ( n2877 & n3138 ) | ( ~n3139 & n3138 ) ;
  assign n3141 = n315 | n3113 ;
  assign n3142 = n3127 | n3141 ;
  assign n3143 = n3133 &  n3142 ;
  assign n3144 = ( n3121 & ~n3124 ) | ( n3121 & 1'b0 ) | ( ~n3124 & 1'b0 ) ;
  assign n3145 = ( n396 & ~n3144 ) | ( n396 & n3118 ) | ( ~n3144 & n3118 ) ;
  assign n3146 = n315 &  n3145 ;
  assign n3147 = n240 | n3146 ;
  assign n3148 = n3143 | n3147 ;
  assign n3149 = ~n3140 & n3148 ;
  assign n3150 = n3135 | n3149 ;
  assign n3151 = ~n2892 & n2955 ;
  assign n3152 = ( n2879 & n2884 ) | ( n2879 & n2955 ) | ( n2884 & n2955 ) ;
  assign n3154 = ( n3151 & ~n2879 ) | ( n3151 & n3152 ) | ( ~n2879 & n3152 ) ;
  assign n3153 = ( n2955 & ~n3152 ) | ( n2955 & n3151 ) | ( ~n3152 & n3151 ) ;
  assign n3155 = ( n2884 & ~n3154 ) | ( n2884 & n3153 ) | ( ~n3154 & n3153 ) ;
  assign n3156 = ( n181 & n3150 ) | ( n181 & n3155 ) | ( n3150 & n3155 ) ;
  assign n3157 = ~n145 & n3156 ;
  assign n3159 = ( n2908 & ~n2899 ) | ( n2908 & n2912 ) | ( ~n2899 & n2912 ) ;
  assign n3158 = n2912 | n2955 ;
  assign n3161 = ( n2912 & ~n3159 ) | ( n2912 & n3158 ) | ( ~n3159 & n3158 ) ;
  assign n3160 = ( n3158 & ~n2908 ) | ( n3158 & n3159 ) | ( ~n2908 & n3159 ) ;
  assign n3162 = ( n2899 & ~n3161 ) | ( n2899 & n3160 ) | ( ~n3161 & n3160 ) ;
  assign n3163 = n181 | n3135 ;
  assign n3164 = n3149 | n3163 ;
  assign n3165 = n3155 &  n3164 ;
  assign n3166 = n3143 | n3146 ;
  assign n3167 = ( n240 & ~n3140 ) | ( n240 & n3166 ) | ( ~n3140 & n3166 ) ;
  assign n3168 = n181 &  n3167 ;
  assign n3169 = ( n145 & ~n3168 ) | ( n145 & 1'b0 ) | ( ~n3168 & 1'b0 ) ;
  assign n3170 = ~n3165 & n3169 ;
  assign n3171 = ( n3162 & ~n3170 ) | ( n3162 & 1'b0 ) | ( ~n3170 & 1'b0 ) ;
  assign n3172 = n3157 | n3171 ;
  assign n3178 = ( n150 & ~n3177 ) | ( n150 & n3172 ) | ( ~n3177 & n3172 ) ;
  assign n3190 = n3178 | n3189 ;
  assign n3191 = ( n133 & ~n3189 ) | ( n133 & n3190 ) | ( ~n3189 & n3190 ) ;
  assign n3192 = n150 | n3157 ;
  assign n3193 = n3171 | n3192 ;
  assign n3198 = n3193 | n3177 ;
  assign n3194 = n3165 | n3168 ;
  assign n3195 = ( n3162 & ~n145 ) | ( n3162 & n3194 ) | ( ~n145 & n3194 ) ;
  assign n3196 = n150 &  n3195 ;
  assign n3197 = ( n3185 & ~n3196 ) | ( n3185 & 1'b0 ) | ( ~n3196 & 1'b0 ) ;
  assign n3199 = ( n3177 & ~n3198 ) | ( n3177 & n3197 ) | ( ~n3198 & n3197 ) ;
  assign n3201 = ( n133 & ~n2922 ) | ( n133 & n2929 ) | ( ~n2922 & n2929 ) ;
  assign n3200 = ( n2922 & ~n2929 ) | ( n2922 & n2955 ) | ( ~n2929 & n2955 ) ;
  assign n3202 = n2929 &  n3200 ;
  assign n3203 = ( n3201 & ~n2929 ) | ( n3201 & n3202 ) | ( ~n2929 & n3202 ) ;
  assign n3204 = n2925 | n2952 ;
  assign n3205 = ( n2947 & ~n2928 ) | ( n2947 & n3204 ) | ( ~n2928 & n3204 ) ;
  assign n3206 = n2928 | n3205 ;
  assign n3207 = ( n2935 & n2943 ) | ( n2935 & n3206 ) | ( n2943 & n3206 ) ;
  assign n3208 = ( n2935 & ~n3207 ) | ( n2935 & 1'b0 ) | ( ~n3207 & 1'b0 ) ;
  assign n3209 = n3203 | n3208 ;
  assign n3210 = n3199 | n3209 ;
  assign n3211 = ~n3191 |  n3210 ;
  assign n3230 = ~n2707 & n3211 ;
  assign n3509 = ~x82 & n3211 ;
  assign n3510 = ( x83 & ~n3509 ) | ( x83 & 1'b0 ) | ( ~n3509 & 1'b0 ) ;
  assign n3511 = n3230 | n3510 ;
  assign n3450 = n3177 &  n3193 ;
  assign n3451 = ( n3196 & n3211 ) | ( n3196 & n3450 ) | ( n3211 & n3450 ) ;
  assign n3452 = ~n3196 & n3451 ;
  assign n3453 = ( n3193 & ~n3196 ) | ( n3193 & 1'b0 ) | ( ~n3196 & 1'b0 ) ;
  assign n3454 = ~n3211 & n3453 ;
  assign n3455 = ( n3177 & ~n3454 ) | ( n3177 & n3453 ) | ( ~n3454 & n3453 ) ;
  assign n3456 = ~n3452 & n3455 ;
  assign n3457 = ( n3178 & ~n3185 ) | ( n3178 & 1'b0 ) | ( ~n3185 & 1'b0 ) ;
  assign n3458 = ~n3211 & n3457 ;
  assign n3459 = ( n3199 & ~n3458 ) | ( n3199 & n3457 ) | ( ~n3458 & n3457 ) ;
  assign n3460 = n3456 | n3459 ;
  assign n3422 = ~n3148 & n3211 ;
  assign n3423 = ( n3135 & ~n3422 ) | ( n3135 & n3211 ) | ( ~n3422 & n3211 ) ;
  assign n3424 = ( n3140 & ~n3135 ) | ( n3140 & n3423 ) | ( ~n3135 & n3423 ) ;
  assign n3425 = ( n3135 & ~n3423 ) | ( n3135 & n3140 ) | ( ~n3423 & n3140 ) ;
  assign n3426 = ( n3424 & ~n3140 ) | ( n3424 & n3425 ) | ( ~n3140 & n3425 ) ;
  assign n3379 = ( n3100 & ~n3092 ) | ( n3100 & n3104 ) | ( ~n3092 & n3104 ) ;
  assign n3380 = ( n3092 & n3211 ) | ( n3092 & n3379 ) | ( n3211 & n3379 ) ;
  assign n3381 = ( n3100 & ~n3379 ) | ( n3100 & n3211 ) | ( ~n3379 & n3211 ) ;
  assign n3382 = ( n3104 & ~n3380 ) | ( n3104 & n3381 ) | ( ~n3380 & n3381 ) ;
  assign n3358 = ( n3070 & ~n3075 ) | ( n3070 & n3211 ) | ( ~n3075 & n3211 ) ;
  assign n3357 = n3083 &  n3211 ;
  assign n3359 = ( n3211 & ~n3358 ) | ( n3211 & n3357 ) | ( ~n3358 & n3357 ) ;
  assign n3360 = ( n3357 & ~n3070 ) | ( n3357 & n3358 ) | ( ~n3070 & n3358 ) ;
  assign n3361 = ( n3075 & ~n3359 ) | ( n3075 & n3360 ) | ( ~n3359 & n3360 ) ;
  assign n3335 = ( n3048 & ~n3211 ) | ( n3048 & 1'b0 ) | ( ~n3211 & 1'b0 ) ;
  assign n3336 = ( n3048 & n3053 ) | ( n3048 & n3061 ) | ( n3053 & n3061 ) ;
  assign n3337 = ( n3335 & ~n3061 ) | ( n3335 & n3336 ) | ( ~n3061 & n3336 ) ;
  assign n3338 = ( n3048 & ~n3336 ) | ( n3048 & n3335 ) | ( ~n3336 & n3335 ) ;
  assign n3339 = ( n3053 & ~n3337 ) | ( n3053 & n3338 ) | ( ~n3337 & n3338 ) ;
  assign n3218 = ( x82 & ~n3211 ) | ( x82 & x83 ) | ( ~n3211 & x83 ) ;
  assign n3224 = ( x82 & ~x83 ) | ( x82 & 1'b0 ) | ( ~x83 & 1'b0 ) ;
  assign n3214 = x80 | x81 ;
  assign n3219 = ~x82 & n3214 ;
  assign n3220 = ( x82 & ~n2953 ) | ( x82 & n3219 ) | ( ~n2953 & n3219 ) ;
  assign n3221 = ( n2935 & ~n3220 ) | ( n2935 & n2943 ) | ( ~n3220 & n2943 ) ;
  assign n3222 = ( n2935 & ~n3221 ) | ( n2935 & 1'b0 ) | ( ~n3221 & 1'b0 ) ;
  assign n3223 = ( n3211 & ~x83 ) | ( n3211 & n3222 ) | ( ~x83 & n3222 ) ;
  assign n3225 = ( n3218 & ~n3224 ) | ( n3218 & n3223 ) | ( ~n3224 & n3223 ) ;
  assign n3215 = x82 | n3214 ;
  assign n3216 = x82 &  n3211 ;
  assign n3217 = ( n2955 & ~n3215 ) | ( n2955 & n3216 ) | ( ~n3215 & n3216 ) ;
  assign n3226 = n3217 &  n3225 ;
  assign n3227 = ( n2706 & ~n3225 ) | ( n2706 & n3226 ) | ( ~n3225 & n3226 ) ;
  assign n3228 = n2706 | n3217 ;
  assign n3229 = ( n3225 & ~n3228 ) | ( n3225 & 1'b0 ) | ( ~n3228 & 1'b0 ) ;
  assign n3231 = ( n2955 & ~n3208 ) | ( n2955 & 1'b0 ) | ( ~n3208 & 1'b0 ) ;
  assign n3232 = ( n3199 & ~n3203 ) | ( n3199 & n3231 ) | ( ~n3203 & n3231 ) ;
  assign n3233 = ~n3199 & n3232 ;
  assign n3234 = n3191 &  n3233 ;
  assign n3235 = ( n3230 & ~n3234 ) | ( n3230 & 1'b0 ) | ( ~n3234 & 1'b0 ) ;
  assign n3236 = ( x84 & n3234 ) | ( x84 & n3235 ) | ( n3234 & n3235 ) ;
  assign n3237 = x84 | n3234 ;
  assign n3238 = n3230 | n3237 ;
  assign n3239 = ~n3236 & n3238 ;
  assign n3240 = n3229 | n3239 ;
  assign n3241 = ~n3227 & n3240 ;
  assign n3245 = ~x84 & n2955 ;
  assign n3246 = ( x85 & ~n3245 ) | ( x85 & 1'b0 ) | ( ~n3245 & 1'b0 ) ;
  assign n3247 = n2967 | n3246 ;
  assign n3242 = ( n2955 & ~x84 ) | ( n2955 & n2962 ) | ( ~x84 & n2962 ) ;
  assign n3243 = x84 &  n3242 ;
  assign n3244 = ( n2957 & ~n3243 ) | ( n2957 & n2962 ) | ( ~n3243 & n2962 ) ;
  assign n3248 = ( n3211 & ~n3247 ) | ( n3211 & n3244 ) | ( ~n3247 & n3244 ) ;
  assign n3250 = ( n3211 & ~n3248 ) | ( n3211 & 1'b0 ) | ( ~n3248 & 1'b0 ) ;
  assign n3249 = ~n3244 & n3248 ;
  assign n3251 = ( n3247 & ~n3250 ) | ( n3247 & n3249 ) | ( ~n3250 & n3249 ) ;
  assign n3252 = ( n3241 & ~n2472 ) | ( n3241 & n3251 ) | ( ~n2472 & n3251 ) ;
  assign n3253 = ( n2245 & ~n3252 ) | ( n2245 & 1'b0 ) | ( ~n3252 & 1'b0 ) ;
  assign n3254 = ~n2990 & n2993 ;
  assign n3255 = ( n2976 & ~n3254 ) | ( n2976 & n2990 ) | ( ~n3254 & n2990 ) ;
  assign n3256 = ( n3211 & n3254 ) | ( n3211 & n3255 ) | ( n3254 & n3255 ) ;
  assign n3257 = ( n2990 & ~n3255 ) | ( n2990 & n3211 ) | ( ~n3255 & n3211 ) ;
  assign n3258 = ( n2976 & ~n3256 ) | ( n2976 & n3257 ) | ( ~n3256 & n3257 ) ;
  assign n3259 = n2472 | n3227 ;
  assign n3260 = ( n3240 & ~n3259 ) | ( n3240 & 1'b0 ) | ( ~n3259 & 1'b0 ) ;
  assign n3261 = n3251 | n3260 ;
  assign n3262 = ~n3217 & n3225 ;
  assign n3263 = ( n3239 & ~n2706 ) | ( n3239 & n3262 ) | ( ~n2706 & n3262 ) ;
  assign n3264 = ( n2472 & ~n3263 ) | ( n2472 & 1'b0 ) | ( ~n3263 & 1'b0 ) ;
  assign n3265 = n2245 | n3264 ;
  assign n3266 = ( n3261 & ~n3265 ) | ( n3261 & 1'b0 ) | ( ~n3265 & 1'b0 ) ;
  assign n3267 = n3258 | n3266 ;
  assign n3268 = ~n3253 & n3267 ;
  assign n3269 = n2978 | n3211 ;
  assign n3270 = ( n2978 & ~n2995 ) | ( n2978 & n2988 ) | ( ~n2995 & n2988 ) ;
  assign n3271 = ( n2995 & n3269 ) | ( n2995 & n3270 ) | ( n3269 & n3270 ) ;
  assign n3272 = ( n2978 & ~n3270 ) | ( n2978 & n3269 ) | ( ~n3270 & n3269 ) ;
  assign n3273 = ( n2988 & ~n3271 ) | ( n2988 & n3272 ) | ( ~n3271 & n3272 ) ;
  assign n3274 = ( n2033 & n3268 ) | ( n2033 & n3273 ) | ( n3268 & n3273 ) ;
  assign n3275 = ( n1827 & ~n3274 ) | ( n1827 & 1'b0 ) | ( ~n3274 & 1'b0 ) ;
  assign n3276 = ( n3015 & ~n3211 ) | ( n3015 & 1'b0 ) | ( ~n3211 & 1'b0 ) ;
  assign n3277 = ( n3002 & n3011 ) | ( n3002 & n3015 ) | ( n3011 & n3015 ) ;
  assign n3278 = ( n3276 & ~n3011 ) | ( n3276 & n3277 ) | ( ~n3011 & n3277 ) ;
  assign n3279 = ( n3015 & ~n3277 ) | ( n3015 & n3276 ) | ( ~n3277 & n3276 ) ;
  assign n3280 = ( n3002 & ~n3278 ) | ( n3002 & n3279 ) | ( ~n3278 & n3279 ) ;
  assign n3281 = ( n2033 & ~n3253 ) | ( n2033 & 1'b0 ) | ( ~n3253 & 1'b0 ) ;
  assign n3282 = n3267 &  n3281 ;
  assign n3283 = n3273 | n3282 ;
  assign n3284 = ( n3261 & ~n3264 ) | ( n3261 & 1'b0 ) | ( ~n3264 & 1'b0 ) ;
  assign n3285 = ( n3258 & ~n2245 ) | ( n3258 & n3284 ) | ( ~n2245 & n3284 ) ;
  assign n3286 = n2033 | n3285 ;
  assign n3287 = ~n1827 & n3286 ;
  assign n3288 = n3283 &  n3287 ;
  assign n3289 = n3280 | n3288 ;
  assign n3290 = ~n3275 & n3289 ;
  assign n3291 = n3017 &  n3211 ;
  assign n3292 = ( n3004 & ~n3291 ) | ( n3004 & n3211 ) | ( ~n3291 & n3211 ) ;
  assign n3293 = ( n3009 & ~n3004 ) | ( n3009 & n3292 ) | ( ~n3004 & n3292 ) ;
  assign n3294 = ( n3004 & ~n3292 ) | ( n3004 & n3009 ) | ( ~n3292 & n3009 ) ;
  assign n3295 = ( n3293 & ~n3009 ) | ( n3293 & n3294 ) | ( ~n3009 & n3294 ) ;
  assign n3296 = ( n1636 & n3290 ) | ( n1636 & n3295 ) | ( n3290 & n3295 ) ;
  assign n3297 = n1452 | n3296 ;
  assign n3299 = ( n3033 & ~n3024 ) | ( n3033 & n3037 ) | ( ~n3024 & n3037 ) ;
  assign n3298 = ( n3037 & ~n3211 ) | ( n3037 & 1'b0 ) | ( ~n3211 & 1'b0 ) ;
  assign n3301 = ( n3037 & ~n3299 ) | ( n3037 & n3298 ) | ( ~n3299 & n3298 ) ;
  assign n3300 = ( n3298 & ~n3033 ) | ( n3298 & n3299 ) | ( ~n3033 & n3299 ) ;
  assign n3302 = ( n3024 & ~n3301 ) | ( n3024 & n3300 ) | ( ~n3301 & n3300 ) ;
  assign n3303 = ( n1636 & ~n3275 ) | ( n1636 & 1'b0 ) | ( ~n3275 & 1'b0 ) ;
  assign n3304 = n3289 &  n3303 ;
  assign n3305 = n3295 | n3304 ;
  assign n3306 = n3283 &  n3286 ;
  assign n3307 = ( n3280 & ~n1827 ) | ( n3280 & n3306 ) | ( ~n1827 & n3306 ) ;
  assign n3308 = n1636 | n3307 ;
  assign n3309 = n1452 &  n3308 ;
  assign n3310 = n3305 &  n3309 ;
  assign n3311 = n3302 | n3310 ;
  assign n3312 = n3297 &  n3311 ;
  assign n3313 = ( n3026 & ~n3211 ) | ( n3026 & 1'b0 ) | ( ~n3211 & 1'b0 ) ;
  assign n3314 = ( n3026 & n3031 ) | ( n3026 & n3039 ) | ( n3031 & n3039 ) ;
  assign n3315 = ( n3313 & ~n3039 ) | ( n3313 & n3314 ) | ( ~n3039 & n3314 ) ;
  assign n3316 = ( n3026 & ~n3314 ) | ( n3026 & n3313 ) | ( ~n3314 & n3313 ) ;
  assign n3317 = ( n3031 & ~n3315 ) | ( n3031 & n3316 ) | ( ~n3315 & n3316 ) ;
  assign n3318 = ( n3312 & ~n1283 ) | ( n3312 & n3317 ) | ( ~n1283 & n3317 ) ;
  assign n3319 = n1122 | n3318 ;
  assign n3320 = n3059 | n3211 ;
  assign n3321 = ( n3046 & ~n3055 ) | ( n3046 & n3059 ) | ( ~n3055 & n3059 ) ;
  assign n3322 = ( n3055 & n3320 ) | ( n3055 & n3321 ) | ( n3320 & n3321 ) ;
  assign n3323 = ( n3059 & ~n3321 ) | ( n3059 & n3320 ) | ( ~n3321 & n3320 ) ;
  assign n3324 = ( n3046 & ~n3322 ) | ( n3046 & n3323 ) | ( ~n3322 & n3323 ) ;
  assign n3325 = ~n1283 & n3297 ;
  assign n3326 = n3311 &  n3325 ;
  assign n3327 = n3317 | n3326 ;
  assign n3328 = n3305 &  n3308 ;
  assign n3329 = ( n1452 & n3302 ) | ( n1452 & n3328 ) | ( n3302 & n3328 ) ;
  assign n3330 = ( n1283 & ~n3329 ) | ( n1283 & 1'b0 ) | ( ~n3329 & 1'b0 ) ;
  assign n3331 = ( n1122 & ~n3330 ) | ( n1122 & 1'b0 ) | ( ~n3330 & 1'b0 ) ;
  assign n3332 = n3327 &  n3331 ;
  assign n3333 = n3324 | n3332 ;
  assign n3334 = n3319 &  n3333 ;
  assign n3340 = ( n976 & ~n3339 ) | ( n976 & n3334 ) | ( ~n3339 & n3334 ) ;
  assign n3341 = ( n837 & ~n3340 ) | ( n837 & 1'b0 ) | ( ~n3340 & 1'b0 ) ;
  assign n3343 = ( n3077 & ~n3068 ) | ( n3077 & n3081 ) | ( ~n3068 & n3081 ) ;
  assign n3342 = ( n3081 & ~n3211 ) | ( n3081 & 1'b0 ) | ( ~n3211 & 1'b0 ) ;
  assign n3345 = ( n3081 & ~n3343 ) | ( n3081 & n3342 ) | ( ~n3343 & n3342 ) ;
  assign n3344 = ( n3342 & ~n3077 ) | ( n3342 & n3343 ) | ( ~n3077 & n3343 ) ;
  assign n3346 = ( n3068 & ~n3345 ) | ( n3068 & n3344 ) | ( ~n3345 & n3344 ) ;
  assign n3347 = n976 &  n3319 ;
  assign n3348 = n3333 &  n3347 ;
  assign n3349 = ( n3339 & ~n3348 ) | ( n3339 & 1'b0 ) | ( ~n3348 & 1'b0 ) ;
  assign n3350 = ( n3327 & ~n3330 ) | ( n3327 & 1'b0 ) | ( ~n3330 & 1'b0 ) ;
  assign n3351 = ( n1122 & n3324 ) | ( n1122 & n3350 ) | ( n3324 & n3350 ) ;
  assign n3352 = n976 | n3351 ;
  assign n3353 = ~n837 & n3352 ;
  assign n3354 = ~n3349 & n3353 ;
  assign n3355 = ( n3346 & ~n3354 ) | ( n3346 & 1'b0 ) | ( ~n3354 & 1'b0 ) ;
  assign n3356 = n3341 | n3355 ;
  assign n3362 = ( n713 & ~n3361 ) | ( n713 & n3356 ) | ( ~n3361 & n3356 ) ;
  assign n3363 = n595 &  n3362 ;
  assign n3364 = n3098 | n3211 ;
  assign n3365 = ( n3090 & ~n3094 ) | ( n3090 & n3098 ) | ( ~n3094 & n3098 ) ;
  assign n3366 = ( n3094 & n3364 ) | ( n3094 & n3365 ) | ( n3364 & n3365 ) ;
  assign n3367 = ( n3098 & ~n3365 ) | ( n3098 & n3364 ) | ( ~n3365 & n3364 ) ;
  assign n3368 = ( n3090 & ~n3366 ) | ( n3090 & n3367 ) | ( ~n3366 & n3367 ) ;
  assign n3369 = n713 | n3341 ;
  assign n3370 = n3355 | n3369 ;
  assign n3371 = ~n3361 & n3370 ;
  assign n3372 = ~n3349 & n3352 ;
  assign n3373 = ( n837 & ~n3372 ) | ( n837 & n3346 ) | ( ~n3372 & n3346 ) ;
  assign n3374 = n713 &  n3373 ;
  assign n3375 = n595 | n3374 ;
  assign n3376 = n3371 | n3375 ;
  assign n3377 = ~n3368 & n3376 ;
  assign n3378 = n3363 | n3377 ;
  assign n3383 = ( n492 & ~n3382 ) | ( n492 & n3378 ) | ( ~n3382 & n3378 ) ;
  assign n3384 = n396 &  n3383 ;
  assign n3385 = n3124 | n3211 ;
  assign n3386 = ( n3111 & ~n3124 ) | ( n3111 & n3120 ) | ( ~n3124 & n3120 ) ;
  assign n3388 = ( n3124 & n3385 ) | ( n3124 & n3386 ) | ( n3385 & n3386 ) ;
  assign n3387 = ( n3120 & ~n3386 ) | ( n3120 & n3385 ) | ( ~n3386 & n3385 ) ;
  assign n3389 = ( n3111 & ~n3388 ) | ( n3111 & n3387 ) | ( ~n3388 & n3387 ) ;
  assign n3390 = n492 | n3363 ;
  assign n3391 = n3377 | n3390 ;
  assign n3392 = ~n3382 & n3391 ;
  assign n3393 = n3371 | n3374 ;
  assign n3394 = ( n595 & ~n3368 ) | ( n595 & n3393 ) | ( ~n3368 & n3393 ) ;
  assign n3395 = n492 &  n3394 ;
  assign n3396 = n396 | n3395 ;
  assign n3397 = n3392 | n3396 ;
  assign n3398 = ~n3389 & n3397 ;
  assign n3399 = n3384 | n3398 ;
  assign n3401 = ( n3113 & ~n3118 ) | ( n3113 & n3211 ) | ( ~n3118 & n3211 ) ;
  assign n3400 = n3126 &  n3211 ;
  assign n3402 = ( n3211 & ~n3401 ) | ( n3211 & n3400 ) | ( ~n3401 & n3400 ) ;
  assign n3403 = ( n3400 & ~n3113 ) | ( n3400 & n3401 ) | ( ~n3113 & n3401 ) ;
  assign n3404 = ( n3118 & ~n3402 ) | ( n3118 & n3403 ) | ( ~n3402 & n3403 ) ;
  assign n3405 = ( n315 & n3399 ) | ( n315 & n3404 ) | ( n3399 & n3404 ) ;
  assign n3406 = n240 &  n3405 ;
  assign n3407 = n3146 | n3211 ;
  assign n3408 = ( n3133 & n3142 ) | ( n3133 & n3146 ) | ( n3142 & n3146 ) ;
  assign n3409 = ( n3407 & ~n3142 ) | ( n3407 & n3408 ) | ( ~n3142 & n3408 ) ;
  assign n3410 = ( n3146 & ~n3408 ) | ( n3146 & n3407 ) | ( ~n3408 & n3407 ) ;
  assign n3411 = ( n3133 & ~n3409 ) | ( n3133 & n3410 ) | ( ~n3409 & n3410 ) ;
  assign n3412 = n315 | n3384 ;
  assign n3413 = n3398 | n3412 ;
  assign n3414 = n3404 &  n3413 ;
  assign n3415 = n3392 | n3395 ;
  assign n3416 = ( n396 & ~n3389 ) | ( n396 & n3415 ) | ( ~n3389 & n3415 ) ;
  assign n3417 = n315 &  n3416 ;
  assign n3418 = n240 | n3417 ;
  assign n3419 = n3414 | n3418 ;
  assign n3420 = n3411 &  n3419 ;
  assign n3421 = n3406 | n3420 ;
  assign n3427 = ( n181 & ~n3426 ) | ( n181 & n3421 ) | ( ~n3426 & n3421 ) ;
  assign n3428 = ~n145 & n3427 ;
  assign n3430 = ( n3164 & ~n3155 ) | ( n3164 & n3168 ) | ( ~n3155 & n3168 ) ;
  assign n3429 = n3168 | n3211 ;
  assign n3432 = ( n3168 & ~n3430 ) | ( n3168 & n3429 ) | ( ~n3430 & n3429 ) ;
  assign n3431 = ( n3429 & ~n3164 ) | ( n3429 & n3430 ) | ( ~n3164 & n3430 ) ;
  assign n3433 = ( n3155 & ~n3432 ) | ( n3155 & n3431 ) | ( ~n3432 & n3431 ) ;
  assign n3434 = n181 | n3406 ;
  assign n3435 = n3420 | n3434 ;
  assign n3436 = ~n3426 & n3435 ;
  assign n3437 = n3414 | n3417 ;
  assign n3438 = ( n240 & n3411 ) | ( n240 & n3437 ) | ( n3411 & n3437 ) ;
  assign n3439 = n181 &  n3438 ;
  assign n3440 = ( n145 & ~n3439 ) | ( n145 & 1'b0 ) | ( ~n3439 & 1'b0 ) ;
  assign n3441 = ~n3436 & n3440 ;
  assign n3442 = ( n3433 & ~n3441 ) | ( n3433 & 1'b0 ) | ( ~n3441 & 1'b0 ) ;
  assign n3443 = n3428 | n3442 ;
  assign n3444 = n3157 | n3211 ;
  assign n3445 = ( n3162 & ~n3157 ) | ( n3162 & n3170 ) | ( ~n3157 & n3170 ) ;
  assign n3447 = ( n3157 & n3444 ) | ( n3157 & n3445 ) | ( n3444 & n3445 ) ;
  assign n3446 = ( n3170 & ~n3445 ) | ( n3170 & n3444 ) | ( ~n3445 & n3444 ) ;
  assign n3448 = ( n3162 & ~n3447 ) | ( n3162 & n3446 ) | ( ~n3447 & n3446 ) ;
  assign n3449 = ( n150 & n3443 ) | ( n150 & n3448 ) | ( n3443 & n3448 ) ;
  assign n3461 = n3449 | n3460 ;
  assign n3462 = ( n133 & ~n3460 ) | ( n133 & n3461 ) | ( ~n3460 & n3461 ) ;
  assign n3465 = n3436 | n3439 ;
  assign n3466 = ( n3433 & ~n145 ) | ( n3433 & n3465 ) | ( ~n145 & n3465 ) ;
  assign n3467 = n150 &  n3466 ;
  assign n3468 = ( n3456 & ~n3467 ) | ( n3456 & 1'b0 ) | ( ~n3467 & 1'b0 ) ;
  assign n3463 = n150 | n3428 ;
  assign n3464 = n3442 | n3463 ;
  assign n3469 = ( n3448 & ~n3464 ) | ( n3448 & 1'b0 ) | ( ~n3464 & 1'b0 ) ;
  assign n3470 = ( n3468 & ~n3448 ) | ( n3468 & n3469 ) | ( ~n3448 & n3469 ) ;
  assign n3472 = ( n133 & ~n3185 ) | ( n133 & n3178 ) | ( ~n3185 & n3178 ) ;
  assign n3471 = ( n3185 & ~n3178 ) | ( n3185 & n3211 ) | ( ~n3178 & n3211 ) ;
  assign n3473 = ~n3185 & n3471 ;
  assign n3474 = ( n3185 & n3472 ) | ( n3185 & n3473 ) | ( n3472 & n3473 ) ;
  assign n3475 = n3181 | n3208 ;
  assign n3476 = ( n3184 & n3203 ) | ( n3184 & n3475 ) | ( n3203 & n3475 ) ;
  assign n3477 = ( n3184 & ~n3476 ) | ( n3184 & 1'b0 ) | ( ~n3476 & 1'b0 ) ;
  assign n3478 = ( n3191 & ~n3477 ) | ( n3191 & n3199 ) | ( ~n3477 & n3199 ) ;
  assign n3479 = ( n3191 & ~n3478 ) | ( n3191 & 1'b0 ) | ( ~n3478 & 1'b0 ) ;
  assign n3480 = n3474 | n3479 ;
  assign n3481 = n3470 | n3480 ;
  assign n3482 = ~n3462 |  n3481 ;
  assign n3506 = ( n3211 & ~x82 ) | ( n3211 & n3222 ) | ( ~x82 & n3222 ) ;
  assign n3507 = x82 &  n3506 ;
  assign n3508 = ( n3217 & ~n3507 ) | ( n3217 & n3222 ) | ( ~n3507 & n3222 ) ;
  assign n3512 = ( n3482 & ~n3511 ) | ( n3482 & n3508 ) | ( ~n3511 & n3508 ) ;
  assign n3514 = ( n3482 & ~n3512 ) | ( n3482 & 1'b0 ) | ( ~n3512 & 1'b0 ) ;
  assign n3513 = ~n3508 & n3512 ;
  assign n3515 = ( n3511 & ~n3514 ) | ( n3511 & n3513 ) | ( ~n3514 & n3513 ) ;
  assign n3495 = ( n3211 & ~n3479 ) | ( n3211 & 1'b0 ) | ( ~n3479 & 1'b0 ) ;
  assign n3496 = ( n3470 & ~n3474 ) | ( n3470 & n3495 ) | ( ~n3474 & n3495 ) ;
  assign n3497 = ~n3470 & n3496 ;
  assign n3498 = n3462 &  n3497 ;
  assign n3494 = ~n3214 & n3482 ;
  assign n3499 = ( n3494 & ~n3498 ) | ( n3494 & 1'b0 ) | ( ~n3498 & 1'b0 ) ;
  assign n3500 = ( x82 & n3498 ) | ( x82 & n3499 ) | ( n3498 & n3499 ) ;
  assign n3501 = x82 | n3498 ;
  assign n3502 = n3494 | n3501 ;
  assign n3503 = ~n3500 & n3502 ;
  assign n3485 = ( x80 & ~n3482 ) | ( x80 & x81 ) | ( ~n3482 & x81 ) ;
  assign n3491 = ( x80 & ~x81 ) | ( x80 & 1'b0 ) | ( ~x81 & 1'b0 ) ;
  assign n3212 = x78 | x79 ;
  assign n3486 = ~x80 & n3212 ;
  assign n3487 = ( x80 & ~n3209 ) | ( x80 & n3486 ) | ( ~n3209 & n3486 ) ;
  assign n3488 = ( n3191 & ~n3487 ) | ( n3191 & n3199 ) | ( ~n3487 & n3199 ) ;
  assign n3489 = ( n3191 & ~n3488 ) | ( n3191 & 1'b0 ) | ( ~n3488 & 1'b0 ) ;
  assign n3490 = ( n3482 & ~x81 ) | ( n3482 & n3489 ) | ( ~x81 & n3489 ) ;
  assign n3492 = ( n3485 & ~n3491 ) | ( n3485 & n3490 ) | ( ~n3491 & n3490 ) ;
  assign n3213 = x80 | n3212 ;
  assign n3483 = x80 &  n3482 ;
  assign n3484 = ( n3211 & ~n3213 ) | ( n3211 & n3483 ) | ( ~n3213 & n3483 ) ;
  assign n3516 = n2955 | n3484 ;
  assign n3517 = ( n3492 & ~n3516 ) | ( n3492 & 1'b0 ) | ( ~n3516 & 1'b0 ) ;
  assign n3518 = n3503 | n3517 ;
  assign n3519 = n3484 &  n3492 ;
  assign n3520 = ( n2955 & ~n3492 ) | ( n2955 & n3519 ) | ( ~n3492 & n3519 ) ;
  assign n3521 = n2706 | n3520 ;
  assign n3522 = ( n3518 & ~n3521 ) | ( n3518 & 1'b0 ) | ( ~n3521 & 1'b0 ) ;
  assign n3493 = ~n3484 & n3492 ;
  assign n3504 = ( n3493 & ~n2955 ) | ( n3493 & n3503 ) | ( ~n2955 & n3503 ) ;
  assign n3505 = ( n2706 & ~n3504 ) | ( n2706 & 1'b0 ) | ( ~n3504 & 1'b0 ) ;
  assign n3678 = ~n3397 & n3482 ;
  assign n3679 = ( n3384 & ~n3678 ) | ( n3384 & n3482 ) | ( ~n3678 & n3482 ) ;
  assign n3680 = ( n3389 & ~n3384 ) | ( n3389 & n3679 ) | ( ~n3384 & n3679 ) ;
  assign n3681 = ( n3384 & ~n3679 ) | ( n3384 & n3389 ) | ( ~n3679 & n3389 ) ;
  assign n3682 = ( n3680 & ~n3389 ) | ( n3680 & n3681 ) | ( ~n3389 & n3681 ) ;
  assign n3657 = ~n3376 & n3482 ;
  assign n3658 = ( n3363 & ~n3657 ) | ( n3363 & n3482 ) | ( ~n3657 & n3482 ) ;
  assign n3659 = ( n3368 & ~n3363 ) | ( n3368 & n3658 ) | ( ~n3363 & n3658 ) ;
  assign n3660 = ( n3363 & ~n3658 ) | ( n3363 & n3368 ) | ( ~n3658 & n3368 ) ;
  assign n3661 = ( n3659 & ~n3368 ) | ( n3659 & n3660 ) | ( ~n3368 & n3660 ) ;
  assign n3523 = n3515 | n3522 ;
  assign n3524 = ~n3505 & n3523 ;
  assign n3525 = ( n3227 & ~n3229 ) | ( n3227 & 1'b0 ) | ( ~n3229 & 1'b0 ) ;
  assign n3526 = ( n3229 & ~n3525 ) | ( n3229 & n3239 ) | ( ~n3525 & n3239 ) ;
  assign n3528 = ( n3482 & n3525 ) | ( n3482 & n3526 ) | ( n3525 & n3526 ) ;
  assign n3527 = ( n3229 & ~n3526 ) | ( n3229 & n3482 ) | ( ~n3526 & n3482 ) ;
  assign n3529 = ( n3239 & ~n3528 ) | ( n3239 & n3527 ) | ( ~n3528 & n3527 ) ;
  assign n3530 = ( n3524 & ~n2472 ) | ( n3524 & n3529 ) | ( ~n2472 & n3529 ) ;
  assign n3531 = ( n2245 & ~n3530 ) | ( n2245 & 1'b0 ) | ( ~n3530 & 1'b0 ) ;
  assign n3532 = n3264 | n3482 ;
  assign n3533 = ( n3251 & ~n3260 ) | ( n3251 & n3264 ) | ( ~n3260 & n3264 ) ;
  assign n3534 = ( n3260 & n3532 ) | ( n3260 & n3533 ) | ( n3532 & n3533 ) ;
  assign n3535 = ( n3264 & ~n3533 ) | ( n3264 & n3532 ) | ( ~n3533 & n3532 ) ;
  assign n3536 = ( n3251 & ~n3534 ) | ( n3251 & n3535 ) | ( ~n3534 & n3535 ) ;
  assign n3537 = n2472 | n3505 ;
  assign n3538 = ( n3523 & ~n3537 ) | ( n3523 & 1'b0 ) | ( ~n3537 & 1'b0 ) ;
  assign n3539 = n3529 | n3538 ;
  assign n3540 = ( n3518 & ~n3520 ) | ( n3518 & 1'b0 ) | ( ~n3520 & 1'b0 ) ;
  assign n3541 = ( n3515 & ~n2706 ) | ( n3515 & n3540 ) | ( ~n2706 & n3540 ) ;
  assign n3542 = ( n2472 & ~n3541 ) | ( n2472 & 1'b0 ) | ( ~n3541 & 1'b0 ) ;
  assign n3543 = n2245 | n3542 ;
  assign n3544 = ( n3539 & ~n3543 ) | ( n3539 & 1'b0 ) | ( ~n3543 & 1'b0 ) ;
  assign n3545 = n3536 | n3544 ;
  assign n3546 = ~n3531 & n3545 ;
  assign n3547 = n3253 | n3482 ;
  assign n3548 = ( n3258 & ~n3253 ) | ( n3258 & n3266 ) | ( ~n3253 & n3266 ) ;
  assign n3550 = ( n3253 & n3547 ) | ( n3253 & n3548 ) | ( n3547 & n3548 ) ;
  assign n3549 = ( n3266 & ~n3548 ) | ( n3266 & n3547 ) | ( ~n3548 & n3547 ) ;
  assign n3551 = ( n3258 & ~n3550 ) | ( n3258 & n3549 ) | ( ~n3550 & n3549 ) ;
  assign n3552 = ( n2033 & n3546 ) | ( n2033 & n3551 ) | ( n3546 & n3551 ) ;
  assign n3553 = ( n1827 & ~n3552 ) | ( n1827 & 1'b0 ) | ( ~n3552 & 1'b0 ) ;
  assign n3555 = ( n3282 & ~n3273 ) | ( n3282 & n3286 ) | ( ~n3273 & n3286 ) ;
  assign n3554 = ( n3286 & ~n3482 ) | ( n3286 & 1'b0 ) | ( ~n3482 & 1'b0 ) ;
  assign n3557 = ( n3286 & ~n3555 ) | ( n3286 & n3554 ) | ( ~n3555 & n3554 ) ;
  assign n3556 = ( n3554 & ~n3282 ) | ( n3554 & n3555 ) | ( ~n3282 & n3555 ) ;
  assign n3558 = ( n3273 & ~n3557 ) | ( n3273 & n3556 ) | ( ~n3557 & n3556 ) ;
  assign n3559 = ( n2033 & ~n3531 ) | ( n2033 & 1'b0 ) | ( ~n3531 & 1'b0 ) ;
  assign n3560 = n3545 &  n3559 ;
  assign n3561 = n3551 | n3560 ;
  assign n3562 = ( n3539 & ~n3542 ) | ( n3539 & 1'b0 ) | ( ~n3542 & 1'b0 ) ;
  assign n3563 = ( n3536 & ~n2245 ) | ( n3536 & n3562 ) | ( ~n2245 & n3562 ) ;
  assign n3564 = n2033 | n3563 ;
  assign n3565 = ~n1827 & n3564 ;
  assign n3566 = n3561 &  n3565 ;
  assign n3567 = n3558 | n3566 ;
  assign n3568 = ~n3553 & n3567 ;
  assign n3569 = n3275 | n3482 ;
  assign n3570 = ( n3275 & ~n3288 ) | ( n3275 & n3280 ) | ( ~n3288 & n3280 ) ;
  assign n3571 = ( n3288 & n3569 ) | ( n3288 & n3570 ) | ( n3569 & n3570 ) ;
  assign n3572 = ( n3275 & ~n3570 ) | ( n3275 & n3569 ) | ( ~n3570 & n3569 ) ;
  assign n3573 = ( n3280 & ~n3571 ) | ( n3280 & n3572 ) | ( ~n3571 & n3572 ) ;
  assign n3574 = ( n1636 & n3568 ) | ( n1636 & n3573 ) | ( n3568 & n3573 ) ;
  assign n3575 = n1452 | n3574 ;
  assign n3576 = ( n3308 & ~n3482 ) | ( n3308 & 1'b0 ) | ( ~n3482 & 1'b0 ) ;
  assign n3577 = ( n3295 & n3304 ) | ( n3295 & n3308 ) | ( n3304 & n3308 ) ;
  assign n3578 = ( n3576 & ~n3304 ) | ( n3576 & n3577 ) | ( ~n3304 & n3577 ) ;
  assign n3579 = ( n3308 & ~n3577 ) | ( n3308 & n3576 ) | ( ~n3577 & n3576 ) ;
  assign n3580 = ( n3295 & ~n3578 ) | ( n3295 & n3579 ) | ( ~n3578 & n3579 ) ;
  assign n3581 = ( n1636 & ~n3553 ) | ( n1636 & 1'b0 ) | ( ~n3553 & 1'b0 ) ;
  assign n3582 = n3567 &  n3581 ;
  assign n3583 = n3573 | n3582 ;
  assign n3584 = n3561 &  n3564 ;
  assign n3585 = ( n3558 & ~n1827 ) | ( n3558 & n3584 ) | ( ~n1827 & n3584 ) ;
  assign n3586 = n1636 | n3585 ;
  assign n3587 = n1452 &  n3586 ;
  assign n3588 = n3583 &  n3587 ;
  assign n3589 = n3580 | n3588 ;
  assign n3590 = n3575 &  n3589 ;
  assign n3591 = n3310 &  n3482 ;
  assign n3592 = ( n3297 & ~n3482 ) | ( n3297 & n3591 ) | ( ~n3482 & n3591 ) ;
  assign n3593 = ( n3297 & ~n3592 ) | ( n3297 & n3302 ) | ( ~n3592 & n3302 ) ;
  assign n3594 = ( n3302 & ~n3297 ) | ( n3302 & n3592 ) | ( ~n3297 & n3592 ) ;
  assign n3595 = ( n3593 & ~n3302 ) | ( n3593 & n3594 ) | ( ~n3302 & n3594 ) ;
  assign n3596 = ( n3590 & ~n1283 ) | ( n3590 & n3595 ) | ( ~n1283 & n3595 ) ;
  assign n3597 = n1122 | n3596 ;
  assign n3598 = n3330 | n3482 ;
  assign n3599 = ( n3317 & ~n3326 ) | ( n3317 & n3330 ) | ( ~n3326 & n3330 ) ;
  assign n3600 = ( n3326 & n3598 ) | ( n3326 & n3599 ) | ( n3598 & n3599 ) ;
  assign n3601 = ( n3330 & ~n3599 ) | ( n3330 & n3598 ) | ( ~n3599 & n3598 ) ;
  assign n3602 = ( n3317 & ~n3600 ) | ( n3317 & n3601 ) | ( ~n3600 & n3601 ) ;
  assign n3603 = ~n1283 & n3575 ;
  assign n3604 = n3589 &  n3603 ;
  assign n3605 = n3595 | n3604 ;
  assign n3606 = n3583 &  n3586 ;
  assign n3607 = ( n1452 & n3580 ) | ( n1452 & n3606 ) | ( n3580 & n3606 ) ;
  assign n3608 = ( n1283 & ~n3607 ) | ( n1283 & 1'b0 ) | ( ~n3607 & 1'b0 ) ;
  assign n3609 = ( n1122 & ~n3608 ) | ( n1122 & 1'b0 ) | ( ~n3608 & 1'b0 ) ;
  assign n3610 = n3605 &  n3609 ;
  assign n3611 = n3602 | n3610 ;
  assign n3612 = n3597 &  n3611 ;
  assign n3613 = ( n3319 & ~n3482 ) | ( n3319 & 1'b0 ) | ( ~n3482 & 1'b0 ) ;
  assign n3614 = ( n3319 & n3324 ) | ( n3319 & n3332 ) | ( n3324 & n3332 ) ;
  assign n3615 = ( n3613 & ~n3332 ) | ( n3613 & n3614 ) | ( ~n3332 & n3614 ) ;
  assign n3616 = ( n3319 & ~n3614 ) | ( n3319 & n3613 ) | ( ~n3614 & n3613 ) ;
  assign n3617 = ( n3324 & ~n3615 ) | ( n3324 & n3616 ) | ( ~n3615 & n3616 ) ;
  assign n3618 = ( n976 & n3612 ) | ( n976 & n3617 ) | ( n3612 & n3617 ) ;
  assign n3619 = ( n837 & ~n3618 ) | ( n837 & 1'b0 ) | ( ~n3618 & 1'b0 ) ;
  assign n3620 = ( n3352 & ~n3482 ) | ( n3352 & 1'b0 ) | ( ~n3482 & 1'b0 ) ;
  assign n3621 = ( n3339 & n3348 ) | ( n3339 & n3352 ) | ( n3348 & n3352 ) ;
  assign n3622 = ( n3620 & ~n3348 ) | ( n3620 & n3621 ) | ( ~n3348 & n3621 ) ;
  assign n3623 = ( n3352 & ~n3621 ) | ( n3352 & n3620 ) | ( ~n3621 & n3620 ) ;
  assign n3624 = ( n3339 & ~n3622 ) | ( n3339 & n3623 ) | ( ~n3622 & n3623 ) ;
  assign n3625 = n976 &  n3597 ;
  assign n3626 = n3611 &  n3625 ;
  assign n3627 = n3617 | n3626 ;
  assign n3628 = ( n3605 & ~n3608 ) | ( n3605 & 1'b0 ) | ( ~n3608 & 1'b0 ) ;
  assign n3629 = ( n1122 & n3602 ) | ( n1122 & n3628 ) | ( n3602 & n3628 ) ;
  assign n3630 = n976 | n3629 ;
  assign n3631 = ~n837 & n3630 ;
  assign n3632 = n3627 &  n3631 ;
  assign n3633 = ( n3624 & ~n3632 ) | ( n3624 & 1'b0 ) | ( ~n3632 & 1'b0 ) ;
  assign n3634 = n3619 | n3633 ;
  assign n3635 = n3341 | n3482 ;
  assign n3636 = ( n3346 & ~n3341 ) | ( n3346 & n3354 ) | ( ~n3341 & n3354 ) ;
  assign n3638 = ( n3341 & n3635 ) | ( n3341 & n3636 ) | ( n3635 & n3636 ) ;
  assign n3637 = ( n3354 & ~n3636 ) | ( n3354 & n3635 ) | ( ~n3636 & n3635 ) ;
  assign n3639 = ( n3346 & ~n3638 ) | ( n3346 & n3637 ) | ( ~n3638 & n3637 ) ;
  assign n3640 = ( n713 & n3634 ) | ( n713 & n3639 ) | ( n3634 & n3639 ) ;
  assign n3641 = n595 &  n3640 ;
  assign n3643 = ( n3370 & ~n3361 ) | ( n3370 & n3374 ) | ( ~n3361 & n3374 ) ;
  assign n3642 = n3374 | n3482 ;
  assign n3645 = ( n3374 & ~n3643 ) | ( n3374 & n3642 ) | ( ~n3643 & n3642 ) ;
  assign n3644 = ( n3642 & ~n3370 ) | ( n3642 & n3643 ) | ( ~n3370 & n3643 ) ;
  assign n3646 = ( n3361 & ~n3645 ) | ( n3361 & n3644 ) | ( ~n3645 & n3644 ) ;
  assign n3647 = n713 | n3619 ;
  assign n3648 = n3633 | n3647 ;
  assign n3649 = n3639 &  n3648 ;
  assign n3650 = n3627 &  n3630 ;
  assign n3651 = ( n837 & ~n3650 ) | ( n837 & n3624 ) | ( ~n3650 & n3624 ) ;
  assign n3652 = n713 &  n3651 ;
  assign n3653 = n595 | n3652 ;
  assign n3654 = n3649 | n3653 ;
  assign n3655 = ~n3646 & n3654 ;
  assign n3656 = n3641 | n3655 ;
  assign n3662 = ( n492 & ~n3661 ) | ( n492 & n3656 ) | ( ~n3661 & n3656 ) ;
  assign n3663 = n396 &  n3662 ;
  assign n3664 = n492 | n3641 ;
  assign n3665 = n3655 | n3664 ;
  assign n3666 = ~n3661 & n3665 ;
  assign n3667 = n3649 | n3652 ;
  assign n3668 = ( n595 & ~n3646 ) | ( n595 & n3667 ) | ( ~n3646 & n3667 ) ;
  assign n3669 = n492 &  n3668 ;
  assign n3670 = n396 | n3669 ;
  assign n3671 = n3666 | n3670 ;
  assign n3672 = ( n3391 & ~n3382 ) | ( n3391 & n3395 ) | ( ~n3382 & n3395 ) ;
  assign n3673 = ( n3395 & ~n3672 ) | ( n3395 & n3482 ) | ( ~n3672 & n3482 ) ;
  assign n3674 = ( n3482 & ~n3391 ) | ( n3482 & n3672 ) | ( ~n3391 & n3672 ) ;
  assign n3675 = ( n3382 & ~n3673 ) | ( n3382 & n3674 ) | ( ~n3673 & n3674 ) ;
  assign n3676 = ( n3671 & ~n3675 ) | ( n3671 & 1'b0 ) | ( ~n3675 & 1'b0 ) ;
  assign n3677 = n3663 | n3676 ;
  assign n3683 = ( n315 & ~n3682 ) | ( n315 & n3677 ) | ( ~n3682 & n3677 ) ;
  assign n3684 = n240 &  n3683 ;
  assign n3685 = n3417 | n3482 ;
  assign n3686 = ( n3404 & n3413 ) | ( n3404 & n3417 ) | ( n3413 & n3417 ) ;
  assign n3687 = ( n3685 & ~n3413 ) | ( n3685 & n3686 ) | ( ~n3413 & n3686 ) ;
  assign n3688 = ( n3417 & ~n3686 ) | ( n3417 & n3685 ) | ( ~n3686 & n3685 ) ;
  assign n3689 = ( n3404 & ~n3687 ) | ( n3404 & n3688 ) | ( ~n3687 & n3688 ) ;
  assign n3690 = n315 | n3663 ;
  assign n3691 = n3676 | n3690 ;
  assign n3692 = ~n3682 & n3691 ;
  assign n3693 = n3666 | n3669 ;
  assign n3694 = ( n396 & ~n3675 ) | ( n396 & n3693 ) | ( ~n3675 & n3693 ) ;
  assign n3695 = n315 &  n3694 ;
  assign n3696 = n240 | n3695 ;
  assign n3697 = n3692 | n3696 ;
  assign n3698 = n3689 &  n3697 ;
  assign n3699 = n3684 | n3698 ;
  assign n3700 = ~n3419 & n3482 ;
  assign n3701 = ( n3406 & ~n3700 ) | ( n3406 & n3482 ) | ( ~n3700 & n3482 ) ;
  assign n3702 = ( n3406 & ~n3701 ) | ( n3406 & n3411 ) | ( ~n3701 & n3411 ) ;
  assign n3703 = ( n3411 & ~n3406 ) | ( n3411 & n3701 ) | ( ~n3406 & n3701 ) ;
  assign n3704 = ( n3702 & ~n3411 ) | ( n3702 & n3703 ) | ( ~n3411 & n3703 ) ;
  assign n3705 = ( n181 & n3699 ) | ( n181 & n3704 ) | ( n3699 & n3704 ) ;
  assign n3706 = ~n145 & n3705 ;
  assign n3707 = n3439 | n3482 ;
  assign n3708 = ( n3426 & n3435 ) | ( n3426 & n3439 ) | ( n3435 & n3439 ) ;
  assign n3709 = ( n3707 & ~n3435 ) | ( n3707 & n3708 ) | ( ~n3435 & n3708 ) ;
  assign n3710 = ( n3439 & ~n3708 ) | ( n3439 & n3707 ) | ( ~n3708 & n3707 ) ;
  assign n3711 = ( n3426 & ~n3709 ) | ( n3426 & n3710 ) | ( ~n3709 & n3710 ) ;
  assign n3712 = n181 | n3684 ;
  assign n3713 = n3698 | n3712 ;
  assign n3714 = n3704 &  n3713 ;
  assign n3715 = n3692 | n3695 ;
  assign n3716 = ( n240 & n3689 ) | ( n240 & n3715 ) | ( n3689 & n3715 ) ;
  assign n3717 = n181 &  n3716 ;
  assign n3718 = ( n145 & ~n3717 ) | ( n145 & 1'b0 ) | ( ~n3717 & 1'b0 ) ;
  assign n3719 = ~n3714 & n3718 ;
  assign n3720 = n3711 | n3719 ;
  assign n3721 = ~n3706 & n3720 ;
  assign n3722 = n3428 | n3482 ;
  assign n3723 = ( n3433 & ~n3428 ) | ( n3433 & n3441 ) | ( ~n3428 & n3441 ) ;
  assign n3725 = ( n3428 & n3722 ) | ( n3428 & n3723 ) | ( n3722 & n3723 ) ;
  assign n3724 = ( n3441 & ~n3723 ) | ( n3441 & n3722 ) | ( ~n3723 & n3722 ) ;
  assign n3726 = ( n3433 & ~n3725 ) | ( n3433 & n3724 ) | ( ~n3725 & n3724 ) ;
  assign n3727 = ( n150 & ~n3721 ) | ( n150 & n3726 ) | ( ~n3721 & n3726 ) ;
  assign n3728 = n3448 | n3467 ;
  assign n3729 = ( n3464 & ~n3482 ) | ( n3464 & n3728 ) | ( ~n3482 & n3728 ) ;
  assign n3730 = ( n3464 & ~n3729 ) | ( n3464 & 1'b0 ) | ( ~n3729 & 1'b0 ) ;
  assign n3731 = ( n3464 & ~n3467 ) | ( n3464 & 1'b0 ) | ( ~n3467 & 1'b0 ) ;
  assign n3732 = ~n3482 & n3731 ;
  assign n3733 = ( n3448 & ~n3731 ) | ( n3448 & n3732 ) | ( ~n3731 & n3732 ) ;
  assign n3734 = n3730 | n3733 ;
  assign n3735 = ( n3449 & ~n3456 ) | ( n3449 & 1'b0 ) | ( ~n3456 & 1'b0 ) ;
  assign n3736 = ~n3482 & n3735 ;
  assign n3737 = ( n3470 & ~n3736 ) | ( n3470 & n3735 ) | ( ~n3736 & n3735 ) ;
  assign n3738 = ( n3734 & ~n3737 ) | ( n3734 & 1'b0 ) | ( ~n3737 & 1'b0 ) ;
  assign n3739 = ~n3727 & n3738 ;
  assign n3740 = ( n133 & ~n3739 ) | ( n133 & n3738 ) | ( ~n3739 & n3738 ) ;
  assign n3741 = n150 | n3706 ;
  assign n3742 = ( n3720 & ~n3741 ) | ( n3720 & 1'b0 ) | ( ~n3741 & 1'b0 ) ;
  assign n3747 = n3726 &  n3742 ;
  assign n3743 = n3714 | n3717 ;
  assign n3744 = ( n145 & ~n3743 ) | ( n145 & n3711 ) | ( ~n3743 & n3711 ) ;
  assign n3745 = ( n150 & ~n3744 ) | ( n150 & 1'b0 ) | ( ~n3744 & 1'b0 ) ;
  assign n3746 = n3734 | n3745 ;
  assign n3748 = ( n3726 & ~n3747 ) | ( n3726 & n3746 ) | ( ~n3747 & n3746 ) ;
  assign n3750 = ( n133 & ~n3456 ) | ( n133 & n3449 ) | ( ~n3456 & n3449 ) ;
  assign n3749 = ( n3456 & ~n3449 ) | ( n3456 & n3482 ) | ( ~n3449 & n3482 ) ;
  assign n3751 = ~n3456 & n3749 ;
  assign n3752 = ( n3456 & n3750 ) | ( n3456 & n3751 ) | ( n3750 & n3751 ) ;
  assign n3753 = n3452 | n3479 ;
  assign n3754 = ( n3455 & n3474 ) | ( n3455 & n3753 ) | ( n3474 & n3753 ) ;
  assign n3755 = ( n3455 & ~n3754 ) | ( n3455 & 1'b0 ) | ( ~n3754 & 1'b0 ) ;
  assign n3756 = ( n3462 & ~n3755 ) | ( n3462 & n3470 ) | ( ~n3755 & n3470 ) ;
  assign n3757 = ( n3462 & ~n3756 ) | ( n3462 & 1'b0 ) | ( ~n3756 & 1'b0 ) ;
  assign n3758 = n3752 | n3757 ;
  assign n3759 = ( n3748 & ~n3758 ) | ( n3748 & 1'b0 ) | ( ~n3758 & 1'b0 ) ;
  assign n3760 = ~n3740 | ~n3759 ;
  assign n3818 = n3505 | n3760 ;
  assign n3819 = ( n3505 & ~n3522 ) | ( n3505 & n3515 ) | ( ~n3522 & n3515 ) ;
  assign n3820 = ( n3522 & n3818 ) | ( n3522 & n3819 ) | ( n3818 & n3819 ) ;
  assign n3821 = ( n3505 & ~n3819 ) | ( n3505 & n3818 ) | ( ~n3819 & n3818 ) ;
  assign n3822 = ( n3515 & ~n3820 ) | ( n3515 & n3821 ) | ( ~n3820 & n3821 ) ;
  assign n3803 = ~n3517 & n3520 ;
  assign n3804 = ( n3517 & ~n3803 ) | ( n3517 & n3760 ) | ( ~n3803 & n3760 ) ;
  assign n3805 = ( n3503 & ~n3517 ) | ( n3503 & n3804 ) | ( ~n3517 & n3804 ) ;
  assign n3806 = ( n3503 & ~n3804 ) | ( n3503 & n3517 ) | ( ~n3804 & n3517 ) ;
  assign n3807 = ( n3805 & ~n3503 ) | ( n3805 & n3806 ) | ( ~n3503 & n3806 ) ;
  assign n3794 = ~x80 & n3482 ;
  assign n3795 = ( x81 & ~n3794 ) | ( x81 & 1'b0 ) | ( ~n3794 & 1'b0 ) ;
  assign n3796 = n3494 | n3795 ;
  assign n3791 = ( n3482 & ~x80 ) | ( n3482 & n3489 ) | ( ~x80 & n3489 ) ;
  assign n3792 = x80 &  n3791 ;
  assign n3793 = ( n3484 & ~n3792 ) | ( n3484 & n3489 ) | ( ~n3792 & n3489 ) ;
  assign n3797 = ( n3760 & ~n3796 ) | ( n3760 & n3793 ) | ( ~n3796 & n3793 ) ;
  assign n3799 = ( n3760 & ~n3797 ) | ( n3760 & 1'b0 ) | ( ~n3797 & 1'b0 ) ;
  assign n3798 = ~n3793 & n3797 ;
  assign n3800 = ( n3796 & ~n3799 ) | ( n3796 & n3798 ) | ( ~n3799 & n3798 ) ;
  assign n3767 = ( x78 & ~n3760 ) | ( x78 & x79 ) | ( ~n3760 & x79 ) ;
  assign n3773 = ( x78 & ~x79 ) | ( x78 & 1'b0 ) | ( ~x79 & 1'b0 ) ;
  assign n3763 = x76 | x77 ;
  assign n3768 = ~x78 & n3763 ;
  assign n3769 = ( x78 & ~n3480 ) | ( x78 & n3768 ) | ( ~n3480 & n3768 ) ;
  assign n3770 = ( n3462 & ~n3769 ) | ( n3462 & n3470 ) | ( ~n3769 & n3470 ) ;
  assign n3771 = ( n3462 & ~n3770 ) | ( n3462 & 1'b0 ) | ( ~n3770 & 1'b0 ) ;
  assign n3772 = ( n3760 & ~x79 ) | ( n3760 & n3771 ) | ( ~x79 & n3771 ) ;
  assign n3774 = ( n3767 & ~n3773 ) | ( n3767 & n3772 ) | ( ~n3773 & n3772 ) ;
  assign n3764 = x78 | n3763 ;
  assign n3765 = x78 &  n3760 ;
  assign n3766 = ( n3482 & ~n3764 ) | ( n3482 & n3765 ) | ( ~n3764 & n3765 ) ;
  assign n3777 = n3211 | n3766 ;
  assign n3778 = ( n3774 & ~n3777 ) | ( n3774 & 1'b0 ) | ( ~n3777 & 1'b0 ) ;
  assign n3780 = ( n3482 & ~n3757 ) | ( n3482 & 1'b0 ) | ( ~n3757 & 1'b0 ) ;
  assign n3781 = ( n3748 & ~n3780 ) | ( n3748 & n3752 ) | ( ~n3780 & n3752 ) ;
  assign n3782 = ( n3748 & ~n3781 ) | ( n3748 & 1'b0 ) | ( ~n3781 & 1'b0 ) ;
  assign n3783 = n3740 &  n3782 ;
  assign n3779 = ~n3212 & n3760 ;
  assign n3784 = ( n3779 & ~n3783 ) | ( n3779 & 1'b0 ) | ( ~n3783 & 1'b0 ) ;
  assign n3785 = ( x80 & n3783 ) | ( x80 & n3784 ) | ( n3783 & n3784 ) ;
  assign n3786 = x80 | n3783 ;
  assign n3787 = n3779 | n3786 ;
  assign n3788 = ~n3785 & n3787 ;
  assign n3789 = n3778 | n3788 ;
  assign n3775 = n3766 &  n3774 ;
  assign n3776 = ( n3211 & ~n3774 ) | ( n3211 & n3775 ) | ( ~n3774 & n3775 ) ;
  assign n3808 = n2955 | n3776 ;
  assign n3809 = ( n3789 & ~n3808 ) | ( n3789 & 1'b0 ) | ( ~n3808 & 1'b0 ) ;
  assign n3810 = n3800 | n3809 ;
  assign n3811 = ~n3766 & n3774 ;
  assign n3812 = ( n3788 & ~n3211 ) | ( n3788 & n3811 ) | ( ~n3211 & n3811 ) ;
  assign n3813 = ( n2955 & ~n3812 ) | ( n2955 & 1'b0 ) | ( ~n3812 & 1'b0 ) ;
  assign n3814 = n2706 | n3813 ;
  assign n3815 = ( n3810 & ~n3814 ) | ( n3810 & 1'b0 ) | ( ~n3814 & 1'b0 ) ;
  assign n3816 = n3807 | n3815 ;
  assign n3790 = ~n3776 & n3789 ;
  assign n3801 = ( n3790 & ~n2955 ) | ( n3790 & n3800 ) | ( ~n2955 & n3800 ) ;
  assign n3802 = ( n2706 & ~n3801 ) | ( n2706 & 1'b0 ) | ( ~n3801 & 1'b0 ) ;
  assign n3830 = n2472 | n3802 ;
  assign n3831 = ( n3816 & ~n3830 ) | ( n3816 & 1'b0 ) | ( ~n3830 & 1'b0 ) ;
  assign n3833 = ( n3810 & ~n3813 ) | ( n3810 & 1'b0 ) | ( ~n3813 & 1'b0 ) ;
  assign n3834 = ( n3807 & ~n2706 ) | ( n3807 & n3833 ) | ( ~n2706 & n3833 ) ;
  assign n3835 = ( n2472 & ~n3834 ) | ( n2472 & 1'b0 ) | ( ~n3834 & 1'b0 ) ;
  assign n4015 = n3706 | n3760 ;
  assign n4016 = ( n3706 & ~n3719 ) | ( n3706 & n3711 ) | ( ~n3719 & n3711 ) ;
  assign n4017 = ( n3719 & n4015 ) | ( n3719 & n4016 ) | ( n4015 & n4016 ) ;
  assign n4018 = ( n3706 & ~n4016 ) | ( n3706 & n4015 ) | ( ~n4016 & n4015 ) ;
  assign n4019 = ( n3711 & ~n4017 ) | ( n3711 & n4018 ) | ( ~n4017 & n4018 ) ;
  assign n3972 = ( n3663 & n3671 ) | ( n3663 & n3675 ) | ( n3671 & n3675 ) ;
  assign n3973 = ( n3760 & ~n3671 ) | ( n3760 & n3972 ) | ( ~n3671 & n3972 ) ;
  assign n3974 = ( n3663 & ~n3972 ) | ( n3663 & n3760 ) | ( ~n3972 & n3760 ) ;
  assign n3975 = ( n3675 & ~n3973 ) | ( n3675 & n3974 ) | ( ~n3973 & n3974 ) ;
  assign n3950 = n3641 | n3760 ;
  assign n3951 = ( n3641 & n3646 ) | ( n3641 & n3654 ) | ( n3646 & n3654 ) ;
  assign n3952 = ( n3950 & ~n3654 ) | ( n3950 & n3951 ) | ( ~n3654 & n3951 ) ;
  assign n3953 = ( n3641 & ~n3951 ) | ( n3641 & n3950 ) | ( ~n3951 & n3950 ) ;
  assign n3954 = ( n3646 & ~n3952 ) | ( n3646 & n3953 ) | ( ~n3952 & n3953 ) ;
  assign n3817 = ~n3802 & n3816 ;
  assign n3823 = ( n3817 & ~n2472 ) | ( n3817 & n3822 ) | ( ~n2472 & n3822 ) ;
  assign n3824 = ( n2245 & ~n3823 ) | ( n2245 & 1'b0 ) | ( ~n3823 & 1'b0 ) ;
  assign n3825 = n3542 | n3760 ;
  assign n3826 = ( n3529 & ~n3542 ) | ( n3529 & n3538 ) | ( ~n3542 & n3538 ) ;
  assign n3828 = ( n3542 & n3825 ) | ( n3542 & n3826 ) | ( n3825 & n3826 ) ;
  assign n3827 = ( n3538 & ~n3826 ) | ( n3538 & n3825 ) | ( ~n3826 & n3825 ) ;
  assign n3829 = ( n3529 & ~n3828 ) | ( n3529 & n3827 ) | ( ~n3828 & n3827 ) ;
  assign n3832 = n3822 | n3831 ;
  assign n3836 = n2245 | n3835 ;
  assign n3837 = ( n3832 & ~n3836 ) | ( n3832 & 1'b0 ) | ( ~n3836 & 1'b0 ) ;
  assign n3838 = n3829 | n3837 ;
  assign n3839 = ~n3824 & n3838 ;
  assign n3840 = n3544 &  n3760 ;
  assign n3841 = ( n3531 & n3536 ) | ( n3531 & n3760 ) | ( n3536 & n3760 ) ;
  assign n3843 = ( n3840 & ~n3531 ) | ( n3840 & n3841 ) | ( ~n3531 & n3841 ) ;
  assign n3842 = ( n3760 & ~n3841 ) | ( n3760 & n3840 ) | ( ~n3841 & n3840 ) ;
  assign n3844 = ( n3536 & ~n3843 ) | ( n3536 & n3842 ) | ( ~n3843 & n3842 ) ;
  assign n3845 = ( n2033 & n3839 ) | ( n2033 & n3844 ) | ( n3839 & n3844 ) ;
  assign n3846 = ( n1827 & ~n3845 ) | ( n1827 & 1'b0 ) | ( ~n3845 & 1'b0 ) ;
  assign n3848 = ( n3560 & ~n3551 ) | ( n3560 & n3564 ) | ( ~n3551 & n3564 ) ;
  assign n3847 = ( n3564 & ~n3760 ) | ( n3564 & 1'b0 ) | ( ~n3760 & 1'b0 ) ;
  assign n3850 = ( n3564 & ~n3848 ) | ( n3564 & n3847 ) | ( ~n3848 & n3847 ) ;
  assign n3849 = ( n3847 & ~n3560 ) | ( n3847 & n3848 ) | ( ~n3560 & n3848 ) ;
  assign n3851 = ( n3551 & ~n3850 ) | ( n3551 & n3849 ) | ( ~n3850 & n3849 ) ;
  assign n3852 = ( n2033 & ~n3824 ) | ( n2033 & 1'b0 ) | ( ~n3824 & 1'b0 ) ;
  assign n3853 = n3838 &  n3852 ;
  assign n3854 = n3844 | n3853 ;
  assign n3855 = ( n3832 & ~n3835 ) | ( n3832 & 1'b0 ) | ( ~n3835 & 1'b0 ) ;
  assign n3856 = ( n3829 & ~n2245 ) | ( n3829 & n3855 ) | ( ~n2245 & n3855 ) ;
  assign n3857 = n2033 | n3856 ;
  assign n3858 = ~n1827 & n3857 ;
  assign n3859 = n3854 &  n3858 ;
  assign n3860 = n3851 | n3859 ;
  assign n3861 = ~n3846 & n3860 ;
  assign n3862 = n3553 | n3760 ;
  assign n3863 = ( n3558 & ~n3553 ) | ( n3558 & n3566 ) | ( ~n3553 & n3566 ) ;
  assign n3865 = ( n3553 & n3862 ) | ( n3553 & n3863 ) | ( n3862 & n3863 ) ;
  assign n3864 = ( n3566 & ~n3863 ) | ( n3566 & n3862 ) | ( ~n3863 & n3862 ) ;
  assign n3866 = ( n3558 & ~n3865 ) | ( n3558 & n3864 ) | ( ~n3865 & n3864 ) ;
  assign n3867 = ( n1636 & n3861 ) | ( n1636 & n3866 ) | ( n3861 & n3866 ) ;
  assign n3868 = n1452 | n3867 ;
  assign n3870 = ( n3582 & ~n3573 ) | ( n3582 & n3586 ) | ( ~n3573 & n3586 ) ;
  assign n3869 = ( n3586 & ~n3760 ) | ( n3586 & 1'b0 ) | ( ~n3760 & 1'b0 ) ;
  assign n3872 = ( n3586 & ~n3870 ) | ( n3586 & n3869 ) | ( ~n3870 & n3869 ) ;
  assign n3871 = ( n3869 & ~n3582 ) | ( n3869 & n3870 ) | ( ~n3582 & n3870 ) ;
  assign n3873 = ( n3573 & ~n3872 ) | ( n3573 & n3871 ) | ( ~n3872 & n3871 ) ;
  assign n3874 = ( n1636 & ~n3846 ) | ( n1636 & 1'b0 ) | ( ~n3846 & 1'b0 ) ;
  assign n3875 = n3860 &  n3874 ;
  assign n3876 = n3866 | n3875 ;
  assign n3877 = n3854 &  n3857 ;
  assign n3878 = ( n3851 & ~n1827 ) | ( n3851 & n3877 ) | ( ~n1827 & n3877 ) ;
  assign n3879 = n1636 | n3878 ;
  assign n3880 = n1452 &  n3879 ;
  assign n3881 = n3876 &  n3880 ;
  assign n3882 = n3873 | n3881 ;
  assign n3883 = n3868 &  n3882 ;
  assign n3885 = ( n3575 & ~n3580 ) | ( n3575 & n3588 ) | ( ~n3580 & n3588 ) ;
  assign n3884 = ( n3575 & ~n3760 ) | ( n3575 & 1'b0 ) | ( ~n3760 & 1'b0 ) ;
  assign n3887 = ( n3575 & ~n3885 ) | ( n3575 & n3884 ) | ( ~n3885 & n3884 ) ;
  assign n3886 = ( n3884 & ~n3588 ) | ( n3884 & n3885 ) | ( ~n3588 & n3885 ) ;
  assign n3888 = ( n3580 & ~n3887 ) | ( n3580 & n3886 ) | ( ~n3887 & n3886 ) ;
  assign n3889 = ( n3883 & ~n1283 ) | ( n3883 & n3888 ) | ( ~n1283 & n3888 ) ;
  assign n3890 = n1122 | n3889 ;
  assign n3891 = n3608 | n3760 ;
  assign n3892 = ( n3595 & ~n3608 ) | ( n3595 & n3604 ) | ( ~n3608 & n3604 ) ;
  assign n3894 = ( n3608 & n3891 ) | ( n3608 & n3892 ) | ( n3891 & n3892 ) ;
  assign n3893 = ( n3604 & ~n3892 ) | ( n3604 & n3891 ) | ( ~n3892 & n3891 ) ;
  assign n3895 = ( n3595 & ~n3894 ) | ( n3595 & n3893 ) | ( ~n3894 & n3893 ) ;
  assign n3896 = ~n1283 & n3868 ;
  assign n3897 = n3882 &  n3896 ;
  assign n3898 = n3888 | n3897 ;
  assign n3899 = n3876 &  n3879 ;
  assign n3900 = ( n1452 & n3873 ) | ( n1452 & n3899 ) | ( n3873 & n3899 ) ;
  assign n3901 = ( n1283 & ~n3900 ) | ( n1283 & 1'b0 ) | ( ~n3900 & 1'b0 ) ;
  assign n3902 = ( n1122 & ~n3901 ) | ( n1122 & 1'b0 ) | ( ~n3901 & 1'b0 ) ;
  assign n3903 = n3898 &  n3902 ;
  assign n3904 = n3895 | n3903 ;
  assign n3905 = n3890 &  n3904 ;
  assign n3906 = n3610 &  n3760 ;
  assign n3907 = ( n3602 & ~n3597 ) | ( n3602 & n3760 ) | ( ~n3597 & n3760 ) ;
  assign n3909 = ( n3597 & n3906 ) | ( n3597 & n3907 ) | ( n3906 & n3907 ) ;
  assign n3908 = ( n3760 & ~n3907 ) | ( n3760 & n3906 ) | ( ~n3907 & n3906 ) ;
  assign n3910 = ( n3602 & ~n3909 ) | ( n3602 & n3908 ) | ( ~n3909 & n3908 ) ;
  assign n3911 = ( n976 & n3905 ) | ( n976 & n3910 ) | ( n3905 & n3910 ) ;
  assign n3912 = ( n837 & ~n3911 ) | ( n837 & 1'b0 ) | ( ~n3911 & 1'b0 ) ;
  assign n3914 = ( n3626 & ~n3617 ) | ( n3626 & n3630 ) | ( ~n3617 & n3630 ) ;
  assign n3913 = ( n3630 & ~n3760 ) | ( n3630 & 1'b0 ) | ( ~n3760 & 1'b0 ) ;
  assign n3916 = ( n3630 & ~n3914 ) | ( n3630 & n3913 ) | ( ~n3914 & n3913 ) ;
  assign n3915 = ( n3913 & ~n3626 ) | ( n3913 & n3914 ) | ( ~n3626 & n3914 ) ;
  assign n3917 = ( n3617 & ~n3916 ) | ( n3617 & n3915 ) | ( ~n3916 & n3915 ) ;
  assign n3918 = n976 &  n3890 ;
  assign n3919 = n3904 &  n3918 ;
  assign n3920 = n3910 | n3919 ;
  assign n3921 = ( n3898 & ~n3901 ) | ( n3898 & 1'b0 ) | ( ~n3901 & 1'b0 ) ;
  assign n3922 = ( n1122 & n3895 ) | ( n1122 & n3921 ) | ( n3895 & n3921 ) ;
  assign n3923 = n976 | n3922 ;
  assign n3924 = ~n837 & n3923 ;
  assign n3925 = n3920 &  n3924 ;
  assign n3926 = n3917 | n3925 ;
  assign n3927 = ~n3912 & n3926 ;
  assign n3928 = n3619 | n3760 ;
  assign n3929 = ( n3619 & ~n3632 ) | ( n3619 & n3624 ) | ( ~n3632 & n3624 ) ;
  assign n3930 = ( n3632 & n3928 ) | ( n3632 & n3929 ) | ( n3928 & n3929 ) ;
  assign n3931 = ( n3619 & ~n3929 ) | ( n3619 & n3928 ) | ( ~n3929 & n3928 ) ;
  assign n3932 = ( n3624 & ~n3930 ) | ( n3624 & n3931 ) | ( ~n3930 & n3931 ) ;
  assign n3933 = ( n713 & ~n3927 ) | ( n713 & n3932 ) | ( ~n3927 & n3932 ) ;
  assign n3934 = n595 &  n3933 ;
  assign n3936 = ( n3648 & ~n3639 ) | ( n3648 & n3652 ) | ( ~n3639 & n3652 ) ;
  assign n3935 = n3652 | n3760 ;
  assign n3938 = ( n3652 & ~n3936 ) | ( n3652 & n3935 ) | ( ~n3936 & n3935 ) ;
  assign n3937 = ( n3935 & ~n3648 ) | ( n3935 & n3936 ) | ( ~n3648 & n3936 ) ;
  assign n3939 = ( n3639 & ~n3938 ) | ( n3639 & n3937 ) | ( ~n3938 & n3937 ) ;
  assign n3940 = n713 | n3912 ;
  assign n3941 = ( n3926 & ~n3940 ) | ( n3926 & 1'b0 ) | ( ~n3940 & 1'b0 ) ;
  assign n3942 = ( n3932 & ~n3941 ) | ( n3932 & 1'b0 ) | ( ~n3941 & 1'b0 ) ;
  assign n3943 = n3920 &  n3923 ;
  assign n3944 = ( n3917 & ~n837 ) | ( n3917 & n3943 ) | ( ~n837 & n3943 ) ;
  assign n3945 = ( n713 & ~n3944 ) | ( n713 & 1'b0 ) | ( ~n3944 & 1'b0 ) ;
  assign n3946 = n595 | n3945 ;
  assign n3947 = n3942 | n3946 ;
  assign n3948 = n3939 &  n3947 ;
  assign n3949 = n3934 | n3948 ;
  assign n3955 = ( n492 & ~n3954 ) | ( n492 & n3949 ) | ( ~n3954 & n3949 ) ;
  assign n3956 = n396 &  n3955 ;
  assign n3958 = ( n3665 & ~n3661 ) | ( n3665 & n3669 ) | ( ~n3661 & n3669 ) ;
  assign n3957 = n3669 | n3760 ;
  assign n3960 = ( n3669 & ~n3958 ) | ( n3669 & n3957 ) | ( ~n3958 & n3957 ) ;
  assign n3959 = ( n3957 & ~n3665 ) | ( n3957 & n3958 ) | ( ~n3665 & n3958 ) ;
  assign n3961 = ( n3661 & ~n3960 ) | ( n3661 & n3959 ) | ( ~n3960 & n3959 ) ;
  assign n3962 = n492 | n3934 ;
  assign n3963 = n3948 | n3962 ;
  assign n3964 = ~n3954 & n3963 ;
  assign n3965 = n3942 | n3945 ;
  assign n3966 = ( n595 & n3939 ) | ( n595 & n3965 ) | ( n3939 & n3965 ) ;
  assign n3967 = n492 &  n3966 ;
  assign n3968 = n396 | n3967 ;
  assign n3969 = n3964 | n3968 ;
  assign n3970 = ~n3961 & n3969 ;
  assign n3971 = n3956 | n3970 ;
  assign n3976 = ( n315 & ~n3975 ) | ( n315 & n3971 ) | ( ~n3975 & n3971 ) ;
  assign n3977 = n240 &  n3976 ;
  assign n3979 = ( n3691 & ~n3682 ) | ( n3691 & n3695 ) | ( ~n3682 & n3695 ) ;
  assign n3978 = n3695 | n3760 ;
  assign n3981 = ( n3695 & ~n3979 ) | ( n3695 & n3978 ) | ( ~n3979 & n3978 ) ;
  assign n3980 = ( n3978 & ~n3691 ) | ( n3978 & n3979 ) | ( ~n3691 & n3979 ) ;
  assign n3982 = ( n3682 & ~n3981 ) | ( n3682 & n3980 ) | ( ~n3981 & n3980 ) ;
  assign n3983 = n315 | n3956 ;
  assign n3984 = n3970 | n3983 ;
  assign n3985 = ~n3975 & n3984 ;
  assign n3986 = n3964 | n3967 ;
  assign n3987 = ( n396 & ~n3961 ) | ( n396 & n3986 ) | ( ~n3961 & n3986 ) ;
  assign n3988 = n315 &  n3987 ;
  assign n3989 = n240 | n3988 ;
  assign n3990 = n3985 | n3989 ;
  assign n3991 = ~n3982 & n3990 ;
  assign n3992 = n3977 | n3991 ;
  assign n3993 = ~n3697 & n3760 ;
  assign n3994 = ( n3684 & n3689 ) | ( n3684 & n3760 ) | ( n3689 & n3760 ) ;
  assign n3996 = ( n3993 & ~n3684 ) | ( n3993 & n3994 ) | ( ~n3684 & n3994 ) ;
  assign n3995 = ( n3760 & ~n3994 ) | ( n3760 & n3993 ) | ( ~n3994 & n3993 ) ;
  assign n3997 = ( n3689 & ~n3996 ) | ( n3689 & n3995 ) | ( ~n3996 & n3995 ) ;
  assign n3998 = ( n181 & n3992 ) | ( n181 & n3997 ) | ( n3992 & n3997 ) ;
  assign n3999 = ~n145 & n3998 ;
  assign n4001 = ( n3713 & ~n3704 ) | ( n3713 & n3717 ) | ( ~n3704 & n3717 ) ;
  assign n4000 = n3717 | n3760 ;
  assign n4003 = ( n3717 & ~n4001 ) | ( n3717 & n4000 ) | ( ~n4001 & n4000 ) ;
  assign n4002 = ( n4000 & ~n3713 ) | ( n4000 & n4001 ) | ( ~n3713 & n4001 ) ;
  assign n4004 = ( n3704 & ~n4003 ) | ( n3704 & n4002 ) | ( ~n4003 & n4002 ) ;
  assign n4005 = n181 | n3977 ;
  assign n4006 = n3991 | n4005 ;
  assign n4007 = n3997 &  n4006 ;
  assign n4008 = n3985 | n3988 ;
  assign n4009 = ( n240 & ~n3982 ) | ( n240 & n4008 ) | ( ~n3982 & n4008 ) ;
  assign n4010 = n181 &  n4009 ;
  assign n4011 = ( n145 & ~n4010 ) | ( n145 & 1'b0 ) | ( ~n4010 & 1'b0 ) ;
  assign n4012 = ~n4007 & n4011 ;
  assign n4013 = ( n4004 & ~n4012 ) | ( n4004 & 1'b0 ) | ( ~n4012 & 1'b0 ) ;
  assign n4014 = n3999 | n4013 ;
  assign n4020 = ( n150 & ~n4019 ) | ( n150 & n4014 ) | ( ~n4019 & n4014 ) ;
  assign n4021 = n3726 | n3742 ;
  assign n4022 = ( n3745 & ~n4021 ) | ( n3745 & n3760 ) | ( ~n4021 & n3760 ) ;
  assign n4023 = ~n3745 & n4022 ;
  assign n4024 = n3742 | n3745 ;
  assign n4025 = n3760 | n4024 ;
  assign n4026 = ( n3726 & ~n4025 ) | ( n3726 & n4024 ) | ( ~n4025 & n4024 ) ;
  assign n4027 = n4023 | n4026 ;
  assign n4028 = n3727 &  n3734 ;
  assign n4029 = ~n3760 & n4028 ;
  assign n4030 = ( n3748 & ~n4028 ) | ( n3748 & n4029 ) | ( ~n4028 & n4029 ) ;
  assign n4031 = n4027 &  n4030 ;
  assign n4032 = ~n4020 & n4031 ;
  assign n4033 = ( n133 & ~n4032 ) | ( n133 & n4031 ) | ( ~n4032 & n4031 ) ;
  assign n4036 = n4007 | n4010 ;
  assign n4037 = ( n4004 & ~n145 ) | ( n4004 & n4036 ) | ( ~n145 & n4036 ) ;
  assign n4038 = n150 &  n4037 ;
  assign n4039 = n4027 | n4038 ;
  assign n4034 = n150 | n3999 ;
  assign n4035 = n4013 | n4034 ;
  assign n4040 = n4019 | n4035 ;
  assign n4041 = ( n4039 & ~n4019 ) | ( n4039 & n4040 ) | ( ~n4019 & n4040 ) ;
  assign n4043 = ( n133 & n3727 ) | ( n133 & n3734 ) | ( n3727 & n3734 ) ;
  assign n4042 = ( n3727 & ~n3760 ) | ( n3727 & n3734 ) | ( ~n3760 & n3734 ) ;
  assign n4044 = ( n3734 & ~n4042 ) | ( n3734 & 1'b0 ) | ( ~n4042 & 1'b0 ) ;
  assign n4045 = ( n4043 & ~n3734 ) | ( n4043 & n4044 ) | ( ~n3734 & n4044 ) ;
  assign n4046 = n3730 | n3757 ;
  assign n4047 = ( n3752 & ~n3733 ) | ( n3752 & n4046 ) | ( ~n3733 & n4046 ) ;
  assign n4048 = n3733 | n4047 ;
  assign n4049 = ( n3740 & ~n3748 ) | ( n3740 & n4048 ) | ( ~n3748 & n4048 ) ;
  assign n4050 = ( n3740 & ~n4049 ) | ( n3740 & 1'b0 ) | ( ~n4049 & 1'b0 ) ;
  assign n4051 = n4045 | n4050 ;
  assign n4052 = ( n4041 & ~n4051 ) | ( n4041 & 1'b0 ) | ( ~n4051 & 1'b0 ) ;
  assign n4053 = ~n4033 | ~n4052 ;
  assign n4125 = n3835 | n4053 ;
  assign n4126 = ( n3822 & ~n3831 ) | ( n3822 & n3835 ) | ( ~n3831 & n3835 ) ;
  assign n4127 = ( n3831 & n4125 ) | ( n3831 & n4126 ) | ( n4125 & n4126 ) ;
  assign n4128 = ( n3835 & ~n4126 ) | ( n3835 & n4125 ) | ( ~n4126 & n4125 ) ;
  assign n4129 = ( n3822 & ~n4127 ) | ( n3822 & n4128 ) | ( ~n4127 & n4128 ) ;
  assign n3761 = x74 | x75 ;
  assign n3762 = x76 | n3761 ;
  assign n4054 = x76 &  n4053 ;
  assign n4055 = ( n3760 & ~n3762 ) | ( n3760 & n4054 ) | ( ~n3762 & n4054 ) ;
  assign n4056 = ( x76 & ~n4053 ) | ( x76 & x77 ) | ( ~n4053 & x77 ) ;
  assign n4062 = ( x76 & ~x77 ) | ( x76 & 1'b0 ) | ( ~x77 & 1'b0 ) ;
  assign n4057 = ~x76 & n3761 ;
  assign n4058 = ( x76 & ~n3758 ) | ( x76 & n4057 ) | ( ~n3758 & n4057 ) ;
  assign n4059 = ( n3748 & ~n3740 ) | ( n3748 & n4058 ) | ( ~n3740 & n4058 ) ;
  assign n4060 = n3740 &  n4059 ;
  assign n4061 = ( n4053 & ~x77 ) | ( n4053 & n4060 ) | ( ~x77 & n4060 ) ;
  assign n4063 = ( n4056 & ~n4062 ) | ( n4056 & n4061 ) | ( ~n4062 & n4061 ) ;
  assign n4064 = ~n4055 & n4063 ;
  assign n4066 = ( n3760 & ~n4050 ) | ( n3760 & 1'b0 ) | ( ~n4050 & 1'b0 ) ;
  assign n4067 = ( n4041 & ~n4066 ) | ( n4041 & n4045 ) | ( ~n4066 & n4045 ) ;
  assign n4068 = ( n4041 & ~n4067 ) | ( n4041 & 1'b0 ) | ( ~n4067 & 1'b0 ) ;
  assign n4069 = n4033 &  n4068 ;
  assign n4065 = ~n3763 & n4053 ;
  assign n4070 = ( n4065 & ~n4069 ) | ( n4065 & 1'b0 ) | ( ~n4069 & 1'b0 ) ;
  assign n4071 = ( x78 & n4069 ) | ( x78 & n4070 ) | ( n4069 & n4070 ) ;
  assign n4072 = x78 | n4069 ;
  assign n4073 = n4065 | n4072 ;
  assign n4074 = ~n4071 & n4073 ;
  assign n4075 = ( n4064 & ~n3482 ) | ( n4064 & n4074 ) | ( ~n3482 & n4074 ) ;
  assign n4076 = ( n3211 & ~n4075 ) | ( n3211 & 1'b0 ) | ( ~n4075 & 1'b0 ) ;
  assign n4080 = ~x78 & n3760 ;
  assign n4081 = ( x79 & ~n4080 ) | ( x79 & 1'b0 ) | ( ~n4080 & 1'b0 ) ;
  assign n4082 = n3779 | n4081 ;
  assign n4077 = ( n3760 & ~x78 ) | ( n3760 & n3771 ) | ( ~x78 & n3771 ) ;
  assign n4078 = x78 &  n4077 ;
  assign n4079 = ( n3766 & ~n4078 ) | ( n3766 & n3771 ) | ( ~n4078 & n3771 ) ;
  assign n4083 = ( n4053 & ~n4082 ) | ( n4053 & n4079 ) | ( ~n4082 & n4079 ) ;
  assign n4085 = ( n4053 & ~n4083 ) | ( n4053 & 1'b0 ) | ( ~n4083 & 1'b0 ) ;
  assign n4084 = ~n4079 & n4083 ;
  assign n4086 = ( n4082 & ~n4085 ) | ( n4082 & n4084 ) | ( ~n4085 & n4084 ) ;
  assign n4087 = n3482 | n4055 ;
  assign n4088 = ( n4063 & ~n4087 ) | ( n4063 & 1'b0 ) | ( ~n4087 & 1'b0 ) ;
  assign n4089 = n4074 | n4088 ;
  assign n4090 = n4055 &  n4063 ;
  assign n4091 = ( n3482 & ~n4063 ) | ( n3482 & n4090 ) | ( ~n4063 & n4090 ) ;
  assign n4092 = n3211 | n4091 ;
  assign n4093 = ( n4089 & ~n4092 ) | ( n4089 & 1'b0 ) | ( ~n4092 & 1'b0 ) ;
  assign n4094 = n4086 | n4093 ;
  assign n4095 = ~n4076 & n4094 ;
  assign n4096 = ( n3776 & ~n3778 ) | ( n3776 & 1'b0 ) | ( ~n3778 & 1'b0 ) ;
  assign n4097 = ( n3778 & ~n4096 ) | ( n3778 & n3788 ) | ( ~n4096 & n3788 ) ;
  assign n4099 = ( n4053 & n4096 ) | ( n4053 & n4097 ) | ( n4096 & n4097 ) ;
  assign n4098 = ( n3778 & ~n4097 ) | ( n3778 & n4053 ) | ( ~n4097 & n4053 ) ;
  assign n4100 = ( n3788 & ~n4099 ) | ( n3788 & n4098 ) | ( ~n4099 & n4098 ) ;
  assign n4101 = ( n4095 & ~n2955 ) | ( n4095 & n4100 ) | ( ~n2955 & n4100 ) ;
  assign n4102 = ( n2706 & ~n4101 ) | ( n2706 & 1'b0 ) | ( ~n4101 & 1'b0 ) ;
  assign n4103 = n3813 | n4053 ;
  assign n4104 = ( n3800 & ~n3809 ) | ( n3800 & n3813 ) | ( ~n3809 & n3813 ) ;
  assign n4105 = ( n3809 & n4103 ) | ( n3809 & n4104 ) | ( n4103 & n4104 ) ;
  assign n4106 = ( n3813 & ~n4104 ) | ( n3813 & n4103 ) | ( ~n4104 & n4103 ) ;
  assign n4107 = ( n3800 & ~n4105 ) | ( n3800 & n4106 ) | ( ~n4105 & n4106 ) ;
  assign n4108 = n2955 | n4076 ;
  assign n4109 = ( n4094 & ~n4108 ) | ( n4094 & 1'b0 ) | ( ~n4108 & 1'b0 ) ;
  assign n4110 = n4100 | n4109 ;
  assign n4111 = ( n4089 & ~n4091 ) | ( n4089 & 1'b0 ) | ( ~n4091 & 1'b0 ) ;
  assign n4112 = ( n4086 & ~n3211 ) | ( n4086 & n4111 ) | ( ~n3211 & n4111 ) ;
  assign n4113 = ( n2955 & ~n4112 ) | ( n2955 & 1'b0 ) | ( ~n4112 & 1'b0 ) ;
  assign n4114 = n2706 | n4113 ;
  assign n4115 = ( n4110 & ~n4114 ) | ( n4110 & 1'b0 ) | ( ~n4114 & 1'b0 ) ;
  assign n4116 = n4107 | n4115 ;
  assign n4117 = ~n4102 & n4116 ;
  assign n4118 = n3802 | n4053 ;
  assign n4119 = ( n3807 & ~n3802 ) | ( n3807 & n3815 ) | ( ~n3802 & n3815 ) ;
  assign n4121 = ( n3802 & n4118 ) | ( n3802 & n4119 ) | ( n4118 & n4119 ) ;
  assign n4120 = ( n3815 & ~n4119 ) | ( n3815 & n4118 ) | ( ~n4119 & n4118 ) ;
  assign n4122 = ( n3807 & ~n4121 ) | ( n3807 & n4120 ) | ( ~n4121 & n4120 ) ;
  assign n4123 = ( n4117 & ~n2472 ) | ( n4117 & n4122 ) | ( ~n2472 & n4122 ) ;
  assign n4124 = ( n2245 & ~n4123 ) | ( n2245 & 1'b0 ) | ( ~n4123 & 1'b0 ) ;
  assign n4294 = ( n3977 & ~n3982 ) | ( n3977 & n4053 ) | ( ~n3982 & n4053 ) ;
  assign n4293 = ~n3990 & n4053 ;
  assign n4295 = ( n4053 & ~n4294 ) | ( n4053 & n4293 ) | ( ~n4294 & n4293 ) ;
  assign n4296 = ( n4293 & ~n3977 ) | ( n4293 & n4294 ) | ( ~n3977 & n4294 ) ;
  assign n4297 = ( n3982 & ~n4295 ) | ( n3982 & n4296 ) | ( ~n4295 & n4296 ) ;
  assign n4272 = n3956 | n4053 ;
  assign n4273 = ( n3956 & n3961 ) | ( n3956 & n3969 ) | ( n3961 & n3969 ) ;
  assign n4274 = ( n4272 & ~n3969 ) | ( n4272 & n4273 ) | ( ~n3969 & n4273 ) ;
  assign n4275 = ( n3956 & ~n4273 ) | ( n3956 & n4272 ) | ( ~n4273 & n4272 ) ;
  assign n4276 = ( n3961 & ~n4274 ) | ( n3961 & n4275 ) | ( ~n4274 & n4275 ) ;
  assign n4130 = n2472 | n4102 ;
  assign n4131 = ( n4116 & ~n4130 ) | ( n4116 & 1'b0 ) | ( ~n4130 & 1'b0 ) ;
  assign n4132 = n4122 | n4131 ;
  assign n4133 = ( n4110 & ~n4113 ) | ( n4110 & 1'b0 ) | ( ~n4113 & 1'b0 ) ;
  assign n4134 = ( n4107 & ~n2706 ) | ( n4107 & n4133 ) | ( ~n2706 & n4133 ) ;
  assign n4135 = ( n2472 & ~n4134 ) | ( n2472 & 1'b0 ) | ( ~n4134 & 1'b0 ) ;
  assign n4136 = n2245 | n4135 ;
  assign n4137 = ( n4132 & ~n4136 ) | ( n4132 & 1'b0 ) | ( ~n4136 & 1'b0 ) ;
  assign n4138 = n4129 | n4137 ;
  assign n4139 = ~n4124 & n4138 ;
  assign n4140 = n3824 | n4053 ;
  assign n4141 = ( n3824 & ~n3837 ) | ( n3824 & n3829 ) | ( ~n3837 & n3829 ) ;
  assign n4142 = ( n3837 & n4140 ) | ( n3837 & n4141 ) | ( n4140 & n4141 ) ;
  assign n4143 = ( n3824 & ~n4141 ) | ( n3824 & n4140 ) | ( ~n4141 & n4140 ) ;
  assign n4144 = ( n3829 & ~n4142 ) | ( n3829 & n4143 ) | ( ~n4142 & n4143 ) ;
  assign n4145 = ( n2033 & n4139 ) | ( n2033 & n4144 ) | ( n4139 & n4144 ) ;
  assign n4146 = ( n1827 & ~n4145 ) | ( n1827 & 1'b0 ) | ( ~n4145 & 1'b0 ) ;
  assign n4147 = ( n3857 & ~n4053 ) | ( n3857 & 1'b0 ) | ( ~n4053 & 1'b0 ) ;
  assign n4148 = ( n3844 & n3853 ) | ( n3844 & n3857 ) | ( n3853 & n3857 ) ;
  assign n4149 = ( n4147 & ~n3853 ) | ( n4147 & n4148 ) | ( ~n3853 & n4148 ) ;
  assign n4150 = ( n3857 & ~n4148 ) | ( n3857 & n4147 ) | ( ~n4148 & n4147 ) ;
  assign n4151 = ( n3844 & ~n4149 ) | ( n3844 & n4150 ) | ( ~n4149 & n4150 ) ;
  assign n4152 = ( n2033 & ~n4124 ) | ( n2033 & 1'b0 ) | ( ~n4124 & 1'b0 ) ;
  assign n4153 = n4138 &  n4152 ;
  assign n4154 = n4144 | n4153 ;
  assign n4155 = ( n4132 & ~n4135 ) | ( n4132 & 1'b0 ) | ( ~n4135 & 1'b0 ) ;
  assign n4156 = ( n4129 & ~n2245 ) | ( n4129 & n4155 ) | ( ~n2245 & n4155 ) ;
  assign n4157 = n2033 | n4156 ;
  assign n4158 = ~n1827 & n4157 ;
  assign n4159 = n4154 &  n4158 ;
  assign n4160 = n4151 | n4159 ;
  assign n4161 = ~n4146 & n4160 ;
  assign n4162 = n3859 &  n4053 ;
  assign n4163 = ( n3846 & ~n4162 ) | ( n3846 & n4053 ) | ( ~n4162 & n4053 ) ;
  assign n4164 = ( n3851 & ~n3846 ) | ( n3851 & n4163 ) | ( ~n3846 & n4163 ) ;
  assign n4165 = ( n3846 & ~n4163 ) | ( n3846 & n3851 ) | ( ~n4163 & n3851 ) ;
  assign n4166 = ( n4164 & ~n3851 ) | ( n4164 & n4165 ) | ( ~n3851 & n4165 ) ;
  assign n4167 = ( n1636 & n4161 ) | ( n1636 & n4166 ) | ( n4161 & n4166 ) ;
  assign n4168 = n1452 | n4167 ;
  assign n4170 = ( n3875 & ~n3866 ) | ( n3875 & n3879 ) | ( ~n3866 & n3879 ) ;
  assign n4169 = ( n3879 & ~n4053 ) | ( n3879 & 1'b0 ) | ( ~n4053 & 1'b0 ) ;
  assign n4172 = ( n3879 & ~n4170 ) | ( n3879 & n4169 ) | ( ~n4170 & n4169 ) ;
  assign n4171 = ( n4169 & ~n3875 ) | ( n4169 & n4170 ) | ( ~n3875 & n4170 ) ;
  assign n4173 = ( n3866 & ~n4172 ) | ( n3866 & n4171 ) | ( ~n4172 & n4171 ) ;
  assign n4174 = ( n1636 & ~n4146 ) | ( n1636 & 1'b0 ) | ( ~n4146 & 1'b0 ) ;
  assign n4175 = n4160 &  n4174 ;
  assign n4176 = n4166 | n4175 ;
  assign n4177 = n4154 &  n4157 ;
  assign n4178 = ( n4151 & ~n1827 ) | ( n4151 & n4177 ) | ( ~n1827 & n4177 ) ;
  assign n4179 = n1636 | n4178 ;
  assign n4180 = n1452 &  n4179 ;
  assign n4181 = n4176 &  n4180 ;
  assign n4182 = n4173 | n4181 ;
  assign n4183 = n4168 &  n4182 ;
  assign n4184 = ( n3868 & ~n4053 ) | ( n3868 & 1'b0 ) | ( ~n4053 & 1'b0 ) ;
  assign n4185 = ( n3868 & n3873 ) | ( n3868 & n3881 ) | ( n3873 & n3881 ) ;
  assign n4186 = ( n4184 & ~n3881 ) | ( n4184 & n4185 ) | ( ~n3881 & n4185 ) ;
  assign n4187 = ( n3868 & ~n4185 ) | ( n3868 & n4184 ) | ( ~n4185 & n4184 ) ;
  assign n4188 = ( n3873 & ~n4186 ) | ( n3873 & n4187 ) | ( ~n4186 & n4187 ) ;
  assign n4189 = ( n4183 & ~n1283 ) | ( n4183 & n4188 ) | ( ~n1283 & n4188 ) ;
  assign n4190 = n1122 | n4189 ;
  assign n4191 = n3901 | n4053 ;
  assign n4192 = ( n3888 & ~n3897 ) | ( n3888 & n3901 ) | ( ~n3897 & n3901 ) ;
  assign n4193 = ( n3897 & n4191 ) | ( n3897 & n4192 ) | ( n4191 & n4192 ) ;
  assign n4194 = ( n3901 & ~n4192 ) | ( n3901 & n4191 ) | ( ~n4192 & n4191 ) ;
  assign n4195 = ( n3888 & ~n4193 ) | ( n3888 & n4194 ) | ( ~n4193 & n4194 ) ;
  assign n4196 = ~n1283 & n4168 ;
  assign n4197 = n4182 &  n4196 ;
  assign n4198 = n4188 | n4197 ;
  assign n4199 = n4176 &  n4179 ;
  assign n4200 = ( n1452 & n4173 ) | ( n1452 & n4199 ) | ( n4173 & n4199 ) ;
  assign n4201 = ( n1283 & ~n4200 ) | ( n1283 & 1'b0 ) | ( ~n4200 & 1'b0 ) ;
  assign n4202 = ( n1122 & ~n4201 ) | ( n1122 & 1'b0 ) | ( ~n4201 & 1'b0 ) ;
  assign n4203 = n4198 &  n4202 ;
  assign n4204 = n4195 | n4203 ;
  assign n4205 = n4190 &  n4204 ;
  assign n4207 = ( n3890 & ~n3895 ) | ( n3890 & n3903 ) | ( ~n3895 & n3903 ) ;
  assign n4206 = ( n3890 & ~n4053 ) | ( n3890 & 1'b0 ) | ( ~n4053 & 1'b0 ) ;
  assign n4209 = ( n3890 & ~n4207 ) | ( n3890 & n4206 ) | ( ~n4207 & n4206 ) ;
  assign n4208 = ( n4206 & ~n3903 ) | ( n4206 & n4207 ) | ( ~n3903 & n4207 ) ;
  assign n4210 = ( n3895 & ~n4209 ) | ( n3895 & n4208 ) | ( ~n4209 & n4208 ) ;
  assign n4211 = ( n976 & n4205 ) | ( n976 & n4210 ) | ( n4205 & n4210 ) ;
  assign n4212 = ( n837 & ~n4211 ) | ( n837 & 1'b0 ) | ( ~n4211 & 1'b0 ) ;
  assign n4213 = ( n3923 & ~n4053 ) | ( n3923 & 1'b0 ) | ( ~n4053 & 1'b0 ) ;
  assign n4214 = ( n3910 & n3919 ) | ( n3910 & n3923 ) | ( n3919 & n3923 ) ;
  assign n4215 = ( n4213 & ~n3919 ) | ( n4213 & n4214 ) | ( ~n3919 & n4214 ) ;
  assign n4216 = ( n3923 & ~n4214 ) | ( n3923 & n4213 ) | ( ~n4214 & n4213 ) ;
  assign n4217 = ( n3910 & ~n4215 ) | ( n3910 & n4216 ) | ( ~n4215 & n4216 ) ;
  assign n4218 = n976 &  n4190 ;
  assign n4219 = n4204 &  n4218 ;
  assign n4220 = n4210 | n4219 ;
  assign n4221 = ( n4198 & ~n4201 ) | ( n4198 & 1'b0 ) | ( ~n4201 & 1'b0 ) ;
  assign n4222 = ( n1122 & n4195 ) | ( n1122 & n4221 ) | ( n4195 & n4221 ) ;
  assign n4223 = n976 | n4222 ;
  assign n4224 = ~n837 & n4223 ;
  assign n4225 = n4220 &  n4224 ;
  assign n4226 = n4217 | n4225 ;
  assign n4227 = ~n4212 & n4226 ;
  assign n4229 = ( n3912 & ~n3917 ) | ( n3912 & n4053 ) | ( ~n3917 & n4053 ) ;
  assign n4228 = n3925 &  n4053 ;
  assign n4230 = ( n4053 & ~n4229 ) | ( n4053 & n4228 ) | ( ~n4229 & n4228 ) ;
  assign n4231 = ( n4228 & ~n3912 ) | ( n4228 & n4229 ) | ( ~n3912 & n4229 ) ;
  assign n4232 = ( n3917 & ~n4230 ) | ( n3917 & n4231 ) | ( ~n4230 & n4231 ) ;
  assign n4233 = ( n4227 & ~n713 ) | ( n4227 & n4232 ) | ( ~n713 & n4232 ) ;
  assign n4234 = ( n595 & ~n4233 ) | ( n595 & 1'b0 ) | ( ~n4233 & 1'b0 ) ;
  assign n4235 = n3945 | n4053 ;
  assign n4236 = ( n3932 & ~n3945 ) | ( n3932 & n3941 ) | ( ~n3945 & n3941 ) ;
  assign n4238 = ( n3945 & n4235 ) | ( n3945 & n4236 ) | ( n4235 & n4236 ) ;
  assign n4237 = ( n3941 & ~n4236 ) | ( n3941 & n4235 ) | ( ~n4236 & n4235 ) ;
  assign n4239 = ( n3932 & ~n4238 ) | ( n3932 & n4237 ) | ( ~n4238 & n4237 ) ;
  assign n4240 = n713 | n4212 ;
  assign n4241 = ( n4226 & ~n4240 ) | ( n4226 & 1'b0 ) | ( ~n4240 & 1'b0 ) ;
  assign n4242 = n4232 | n4241 ;
  assign n4243 = n4220 &  n4223 ;
  assign n4244 = ( n4217 & ~n837 ) | ( n4217 & n4243 ) | ( ~n837 & n4243 ) ;
  assign n4245 = ( n713 & ~n4244 ) | ( n713 & 1'b0 ) | ( ~n4244 & 1'b0 ) ;
  assign n4246 = n595 | n4245 ;
  assign n4247 = ( n4242 & ~n4246 ) | ( n4242 & 1'b0 ) | ( ~n4246 & 1'b0 ) ;
  assign n4248 = ( n4239 & ~n4247 ) | ( n4239 & 1'b0 ) | ( ~n4247 & 1'b0 ) ;
  assign n4249 = n4234 | n4248 ;
  assign n4250 = n3934 | n4053 ;
  assign n4251 = ( n3934 & n3939 ) | ( n3934 & n3947 ) | ( n3939 & n3947 ) ;
  assign n4252 = ( n4250 & ~n3947 ) | ( n4250 & n4251 ) | ( ~n3947 & n4251 ) ;
  assign n4253 = ( n3934 & ~n4251 ) | ( n3934 & n4250 ) | ( ~n4251 & n4250 ) ;
  assign n4254 = ( n3939 & ~n4252 ) | ( n3939 & n4253 ) | ( ~n4252 & n4253 ) ;
  assign n4255 = ( n492 & n4249 ) | ( n492 & n4254 ) | ( n4249 & n4254 ) ;
  assign n4256 = n396 &  n4255 ;
  assign n4257 = n3967 | n4053 ;
  assign n4258 = ( n3954 & n3963 ) | ( n3954 & n3967 ) | ( n3963 & n3967 ) ;
  assign n4259 = ( n4257 & ~n3963 ) | ( n4257 & n4258 ) | ( ~n3963 & n4258 ) ;
  assign n4260 = ( n3967 & ~n4258 ) | ( n3967 & n4257 ) | ( ~n4258 & n4257 ) ;
  assign n4261 = ( n3954 & ~n4259 ) | ( n3954 & n4260 ) | ( ~n4259 & n4260 ) ;
  assign n4262 = n492 | n4234 ;
  assign n4263 = n4248 | n4262 ;
  assign n4264 = n4254 &  n4263 ;
  assign n4265 = ( n4242 & ~n4245 ) | ( n4242 & 1'b0 ) | ( ~n4245 & 1'b0 ) ;
  assign n4266 = ( n595 & ~n4265 ) | ( n595 & n4239 ) | ( ~n4265 & n4239 ) ;
  assign n4267 = n492 &  n4266 ;
  assign n4268 = n396 | n4267 ;
  assign n4269 = n4264 | n4268 ;
  assign n4270 = ~n4261 & n4269 ;
  assign n4271 = n4256 | n4270 ;
  assign n4277 = ( n315 & ~n4276 ) | ( n315 & n4271 ) | ( ~n4276 & n4271 ) ;
  assign n4278 = n240 &  n4277 ;
  assign n4279 = n315 | n4256 ;
  assign n4280 = n4270 | n4279 ;
  assign n4281 = ~n4276 & n4280 ;
  assign n4282 = n4264 | n4267 ;
  assign n4283 = ( n396 & ~n4261 ) | ( n396 & n4282 ) | ( ~n4261 & n4282 ) ;
  assign n4284 = n315 &  n4283 ;
  assign n4285 = n240 | n4284 ;
  assign n4286 = n4281 | n4285 ;
  assign n4287 = ( n3984 & ~n3975 ) | ( n3984 & n3988 ) | ( ~n3975 & n3988 ) ;
  assign n4288 = ( n3988 & ~n4287 ) | ( n3988 & n4053 ) | ( ~n4287 & n4053 ) ;
  assign n4289 = ( n4053 & ~n3984 ) | ( n4053 & n4287 ) | ( ~n3984 & n4287 ) ;
  assign n4290 = ( n3975 & ~n4288 ) | ( n3975 & n4289 ) | ( ~n4288 & n4289 ) ;
  assign n4291 = ( n4286 & ~n4290 ) | ( n4286 & 1'b0 ) | ( ~n4290 & 1'b0 ) ;
  assign n4292 = n4278 | n4291 ;
  assign n4298 = ( n181 & ~n4297 ) | ( n181 & n4292 ) | ( ~n4297 & n4292 ) ;
  assign n4299 = ~n145 & n4298 ;
  assign n4301 = ( n4006 & ~n3997 ) | ( n4006 & n4010 ) | ( ~n3997 & n4010 ) ;
  assign n4300 = n4010 | n4053 ;
  assign n4303 = ( n4010 & ~n4301 ) | ( n4010 & n4300 ) | ( ~n4301 & n4300 ) ;
  assign n4302 = ( n4300 & ~n4006 ) | ( n4300 & n4301 ) | ( ~n4006 & n4301 ) ;
  assign n4304 = ( n3997 & ~n4303 ) | ( n3997 & n4302 ) | ( ~n4303 & n4302 ) ;
  assign n4305 = n181 | n4278 ;
  assign n4306 = n4291 | n4305 ;
  assign n4307 = ~n4297 & n4306 ;
  assign n4308 = n4281 | n4284 ;
  assign n4309 = ( n240 & ~n4290 ) | ( n240 & n4308 ) | ( ~n4290 & n4308 ) ;
  assign n4310 = n181 &  n4309 ;
  assign n4311 = ( n145 & ~n4310 ) | ( n145 & 1'b0 ) | ( ~n4310 & 1'b0 ) ;
  assign n4312 = ~n4307 & n4311 ;
  assign n4313 = ( n4304 & ~n4312 ) | ( n4304 & 1'b0 ) | ( ~n4312 & 1'b0 ) ;
  assign n4314 = n4299 | n4313 ;
  assign n4315 = n3999 | n4053 ;
  assign n4316 = ( n4004 & ~n3999 ) | ( n4004 & n4012 ) | ( ~n3999 & n4012 ) ;
  assign n4318 = ( n3999 & n4315 ) | ( n3999 & n4316 ) | ( n4315 & n4316 ) ;
  assign n4317 = ( n4012 & ~n4316 ) | ( n4012 & n4315 ) | ( ~n4316 & n4315 ) ;
  assign n4319 = ( n4004 & ~n4318 ) | ( n4004 & n4317 ) | ( ~n4318 & n4317 ) ;
  assign n4320 = ( n150 & n4314 ) | ( n150 & n4319 ) | ( n4314 & n4319 ) ;
  assign n4321 = ( n4019 & ~n4038 ) | ( n4019 & 1'b0 ) | ( ~n4038 & 1'b0 ) ;
  assign n4322 = ( n4053 & ~n4035 ) | ( n4053 & n4321 ) | ( ~n4035 & n4321 ) ;
  assign n4323 = n4035 &  n4322 ;
  assign n4324 = ( n4035 & ~n4038 ) | ( n4035 & 1'b0 ) | ( ~n4038 & 1'b0 ) ;
  assign n4325 = ~n4053 & n4324 ;
  assign n4326 = ( n4019 & ~n4325 ) | ( n4019 & n4324 ) | ( ~n4325 & n4324 ) ;
  assign n4327 = ~n4323 & n4326 ;
  assign n4328 = n4020 &  n4027 ;
  assign n4329 = ~n4053 & n4328 ;
  assign n4330 = ( n4041 & ~n4328 ) | ( n4041 & n4329 ) | ( ~n4328 & n4329 ) ;
  assign n4331 = ~n4327 & n4330 ;
  assign n4332 = ~n4320 & n4331 ;
  assign n4333 = ( n133 & ~n4332 ) | ( n133 & n4331 ) | ( ~n4332 & n4331 ) ;
  assign n4336 = n4307 | n4310 ;
  assign n4337 = ( n4304 & ~n145 ) | ( n4304 & n4336 ) | ( ~n145 & n4336 ) ;
  assign n4338 = n150 &  n4337 ;
  assign n4339 = ( n4327 & ~n4338 ) | ( n4327 & 1'b0 ) | ( ~n4338 & 1'b0 ) ;
  assign n4334 = n150 | n4299 ;
  assign n4335 = n4313 | n4334 ;
  assign n4340 = ( n4319 & ~n4335 ) | ( n4319 & 1'b0 ) | ( ~n4335 & 1'b0 ) ;
  assign n4341 = ( n4339 & ~n4319 ) | ( n4339 & n4340 ) | ( ~n4319 & n4340 ) ;
  assign n4343 = ( n133 & n4020 ) | ( n133 & n4027 ) | ( n4020 & n4027 ) ;
  assign n4342 = ( n4020 & ~n4053 ) | ( n4020 & n4027 ) | ( ~n4053 & n4027 ) ;
  assign n4344 = ( n4027 & ~n4342 ) | ( n4027 & 1'b0 ) | ( ~n4342 & 1'b0 ) ;
  assign n4345 = ( n4343 & ~n4027 ) | ( n4343 & n4344 ) | ( ~n4027 & n4344 ) ;
  assign n4346 = n4023 | n4050 ;
  assign n4347 = ( n4045 & ~n4026 ) | ( n4045 & n4346 ) | ( ~n4026 & n4346 ) ;
  assign n4348 = n4026 | n4347 ;
  assign n4349 = ( n4033 & ~n4041 ) | ( n4033 & n4348 ) | ( ~n4041 & n4348 ) ;
  assign n4350 = ( n4033 & ~n4349 ) | ( n4033 & 1'b0 ) | ( ~n4349 & 1'b0 ) ;
  assign n4351 = n4345 | n4350 ;
  assign n4352 = n4341 | n4351 ;
  assign n4353 = ~n4333 |  n4352 ;
  assign n4455 = n4124 | n4353 ;
  assign n4456 = ( n4129 & ~n4124 ) | ( n4129 & n4137 ) | ( ~n4124 & n4137 ) ;
  assign n4458 = ( n4124 & n4455 ) | ( n4124 & n4456 ) | ( n4455 & n4456 ) ;
  assign n4457 = ( n4137 & ~n4456 ) | ( n4137 & n4455 ) | ( ~n4456 & n4455 ) ;
  assign n4459 = ( n4129 & ~n4458 ) | ( n4129 & n4457 ) | ( ~n4458 & n4457 ) ;
  assign n4440 = n4135 | n4353 ;
  assign n4441 = ( n4122 & ~n4131 ) | ( n4122 & n4135 ) | ( ~n4131 & n4135 ) ;
  assign n4442 = ( n4131 & n4440 ) | ( n4131 & n4441 ) | ( n4440 & n4441 ) ;
  assign n4443 = ( n4135 & ~n4441 ) | ( n4135 & n4440 ) | ( ~n4441 & n4440 ) ;
  assign n4444 = ( n4122 & ~n4442 ) | ( n4122 & n4443 ) | ( ~n4442 & n4443 ) ;
  assign n4433 = n4115 &  n4353 ;
  assign n4434 = ( n4102 & n4107 ) | ( n4102 & n4353 ) | ( n4107 & n4353 ) ;
  assign n4436 = ( n4433 & ~n4102 ) | ( n4433 & n4434 ) | ( ~n4102 & n4434 ) ;
  assign n4435 = ( n4353 & ~n4434 ) | ( n4353 & n4433 ) | ( ~n4434 & n4433 ) ;
  assign n4437 = ( n4107 & ~n4436 ) | ( n4107 & n4435 ) | ( ~n4436 & n4435 ) ;
  assign n4418 = n4113 | n4353 ;
  assign n4419 = ( n4100 & ~n4113 ) | ( n4100 & n4109 ) | ( ~n4113 & n4109 ) ;
  assign n4421 = ( n4113 & n4418 ) | ( n4113 & n4419 ) | ( n4418 & n4419 ) ;
  assign n4420 = ( n4109 & ~n4419 ) | ( n4109 & n4418 ) | ( ~n4419 & n4418 ) ;
  assign n4422 = ( n4100 & ~n4421 ) | ( n4100 & n4420 ) | ( ~n4421 & n4420 ) ;
  assign n4411 = n4076 | n4353 ;
  assign n4412 = ( n4076 & ~n4093 ) | ( n4076 & n4086 ) | ( ~n4093 & n4086 ) ;
  assign n4413 = ( n4093 & n4411 ) | ( n4093 & n4412 ) | ( n4411 & n4412 ) ;
  assign n4414 = ( n4076 & ~n4412 ) | ( n4076 & n4411 ) | ( ~n4412 & n4411 ) ;
  assign n4415 = ( n4086 & ~n4413 ) | ( n4086 & n4414 ) | ( ~n4413 & n4414 ) ;
  assign n4396 = ~n4088 & n4091 ;
  assign n4397 = ( n4074 & ~n4088 ) | ( n4074 & n4396 ) | ( ~n4088 & n4396 ) ;
  assign n4399 = ( n4353 & n4088 ) | ( n4353 & n4397 ) | ( n4088 & n4397 ) ;
  assign n4398 = ( n4353 & ~n4397 ) | ( n4353 & n4396 ) | ( ~n4397 & n4396 ) ;
  assign n4400 = ( n4074 & ~n4399 ) | ( n4074 & n4398 ) | ( ~n4399 & n4398 ) ;
  assign n4387 = ~x76 & n4053 ;
  assign n4388 = ( x77 & ~n4387 ) | ( x77 & 1'b0 ) | ( ~n4387 & 1'b0 ) ;
  assign n4389 = n4065 | n4388 ;
  assign n4384 = ( n4053 & ~x76 ) | ( n4053 & n4060 ) | ( ~x76 & n4060 ) ;
  assign n4385 = x76 &  n4384 ;
  assign n4386 = ( n4055 & ~n4385 ) | ( n4055 & n4060 ) | ( ~n4385 & n4060 ) ;
  assign n4390 = ( n4353 & ~n4389 ) | ( n4353 & n4386 ) | ( ~n4389 & n4386 ) ;
  assign n4392 = ( n4353 & ~n4390 ) | ( n4353 & 1'b0 ) | ( ~n4390 & 1'b0 ) ;
  assign n4391 = ~n4386 & n4390 ;
  assign n4393 = ( n4389 & ~n4392 ) | ( n4389 & n4391 ) | ( ~n4392 & n4391 ) ;
  assign n4360 = ( x74 & ~n4353 ) | ( x74 & x75 ) | ( ~n4353 & x75 ) ;
  assign n4366 = ( x74 & ~x75 ) | ( x74 & 1'b0 ) | ( ~x75 & 1'b0 ) ;
  assign n4356 = x72 | x73 ;
  assign n4361 = ~x74 & n4356 ;
  assign n4362 = ( x74 & ~n4051 ) | ( x74 & n4361 ) | ( ~n4051 & n4361 ) ;
  assign n4363 = ( n4041 & ~n4033 ) | ( n4041 & n4362 ) | ( ~n4033 & n4362 ) ;
  assign n4364 = n4033 &  n4363 ;
  assign n4365 = ( n4353 & ~x75 ) | ( n4353 & n4364 ) | ( ~x75 & n4364 ) ;
  assign n4367 = ( n4360 & ~n4366 ) | ( n4360 & n4365 ) | ( ~n4366 & n4365 ) ;
  assign n4357 = x74 | n4356 ;
  assign n4358 = x74 &  n4353 ;
  assign n4359 = ( n4053 & ~n4357 ) | ( n4053 & n4358 ) | ( ~n4357 & n4358 ) ;
  assign n4370 = n3760 | n4359 ;
  assign n4371 = ( n4367 & ~n4370 ) | ( n4367 & 1'b0 ) | ( ~n4370 & 1'b0 ) ;
  assign n4373 = ( n4053 & ~n4350 ) | ( n4053 & 1'b0 ) | ( ~n4350 & 1'b0 ) ;
  assign n4374 = ( n4341 & ~n4345 ) | ( n4341 & n4373 ) | ( ~n4345 & n4373 ) ;
  assign n4375 = ~n4341 & n4374 ;
  assign n4376 = n4333 &  n4375 ;
  assign n4372 = ~n3761 & n4353 ;
  assign n4377 = ( n4372 & ~n4376 ) | ( n4372 & 1'b0 ) | ( ~n4376 & 1'b0 ) ;
  assign n4378 = ( x76 & n4376 ) | ( x76 & n4377 ) | ( n4376 & n4377 ) ;
  assign n4379 = x76 | n4376 ;
  assign n4380 = n4372 | n4379 ;
  assign n4381 = ~n4378 & n4380 ;
  assign n4382 = n4371 | n4381 ;
  assign n4368 = n4359 &  n4367 ;
  assign n4369 = ( n3760 & ~n4367 ) | ( n3760 & n4368 ) | ( ~n4367 & n4368 ) ;
  assign n4401 = n3482 | n4369 ;
  assign n4402 = ( n4382 & ~n4401 ) | ( n4382 & 1'b0 ) | ( ~n4401 & 1'b0 ) ;
  assign n4403 = n4393 | n4402 ;
  assign n4404 = ~n4359 & n4367 ;
  assign n4405 = ( n4381 & ~n3760 ) | ( n4381 & n4404 ) | ( ~n3760 & n4404 ) ;
  assign n4406 = ( n3482 & ~n4405 ) | ( n3482 & 1'b0 ) | ( ~n4405 & 1'b0 ) ;
  assign n4407 = n3211 | n4406 ;
  assign n4408 = ( n4403 & ~n4407 ) | ( n4403 & 1'b0 ) | ( ~n4407 & 1'b0 ) ;
  assign n4409 = n4400 | n4408 ;
  assign n4383 = ~n4369 & n4382 ;
  assign n4394 = ( n4383 & ~n3482 ) | ( n4383 & n4393 ) | ( ~n3482 & n4393 ) ;
  assign n4395 = ( n3211 & ~n4394 ) | ( n3211 & 1'b0 ) | ( ~n4394 & 1'b0 ) ;
  assign n4423 = n2955 | n4395 ;
  assign n4424 = ( n4409 & ~n4423 ) | ( n4409 & 1'b0 ) | ( ~n4423 & 1'b0 ) ;
  assign n4425 = n4415 | n4424 ;
  assign n4426 = ( n4403 & ~n4406 ) | ( n4403 & 1'b0 ) | ( ~n4406 & 1'b0 ) ;
  assign n4427 = ( n4400 & ~n3211 ) | ( n4400 & n4426 ) | ( ~n3211 & n4426 ) ;
  assign n4428 = ( n2955 & ~n4427 ) | ( n2955 & 1'b0 ) | ( ~n4427 & 1'b0 ) ;
  assign n4429 = n2706 | n4428 ;
  assign n4430 = ( n4425 & ~n4429 ) | ( n4425 & 1'b0 ) | ( ~n4429 & 1'b0 ) ;
  assign n4431 = n4422 | n4430 ;
  assign n4410 = ~n4395 & n4409 ;
  assign n4416 = ( n4410 & ~n2955 ) | ( n4410 & n4415 ) | ( ~n2955 & n4415 ) ;
  assign n4417 = ( n2706 & ~n4416 ) | ( n2706 & 1'b0 ) | ( ~n4416 & 1'b0 ) ;
  assign n4445 = n2472 | n4417 ;
  assign n4446 = ( n4431 & ~n4445 ) | ( n4431 & 1'b0 ) | ( ~n4445 & 1'b0 ) ;
  assign n4447 = n4437 | n4446 ;
  assign n4448 = ( n4425 & ~n4428 ) | ( n4425 & 1'b0 ) | ( ~n4428 & 1'b0 ) ;
  assign n4449 = ( n4422 & ~n2706 ) | ( n4422 & n4448 ) | ( ~n2706 & n4448 ) ;
  assign n4450 = ( n2472 & ~n4449 ) | ( n2472 & 1'b0 ) | ( ~n4449 & 1'b0 ) ;
  assign n4470 = ( n4447 & ~n4450 ) | ( n4447 & 1'b0 ) | ( ~n4450 & 1'b0 ) ;
  assign n4471 = ( n4444 & ~n2245 ) | ( n4444 & n4470 ) | ( ~n2245 & n4470 ) ;
  assign n4472 = n2033 | n4471 ;
  assign n4451 = n2245 | n4450 ;
  assign n4452 = ( n4447 & ~n4451 ) | ( n4447 & 1'b0 ) | ( ~n4451 & 1'b0 ) ;
  assign n4453 = n4444 | n4452 ;
  assign n4432 = ~n4417 & n4431 ;
  assign n4438 = ( n4432 & ~n2472 ) | ( n4432 & n4437 ) | ( ~n2472 & n4437 ) ;
  assign n4439 = ( n2245 & ~n4438 ) | ( n2245 & 1'b0 ) | ( ~n4438 & 1'b0 ) ;
  assign n4467 = ( n2033 & ~n4439 ) | ( n2033 & 1'b0 ) | ( ~n4439 & 1'b0 ) ;
  assign n4468 = n4453 &  n4467 ;
  assign n4785 = ( n4468 & ~n4459 ) | ( n4468 & n4472 ) | ( ~n4459 & n4472 ) ;
  assign n4609 = ( n4278 & n4286 ) | ( n4278 & n4290 ) | ( n4286 & n4290 ) ;
  assign n4611 = ( n4353 & ~n4286 ) | ( n4353 & n4609 ) | ( ~n4286 & n4609 ) ;
  assign n4610 = ( n4278 & ~n4609 ) | ( n4278 & n4353 ) | ( ~n4609 & n4353 ) ;
  assign n4612 = ( n4290 & ~n4611 ) | ( n4290 & n4610 ) | ( ~n4611 & n4610 ) ;
  assign n4588 = ( n4256 & ~n4261 ) | ( n4256 & n4269 ) | ( ~n4261 & n4269 ) ;
  assign n4587 = n4256 | n4353 ;
  assign n4590 = ( n4256 & ~n4588 ) | ( n4256 & n4587 ) | ( ~n4588 & n4587 ) ;
  assign n4589 = ( n4587 & ~n4269 ) | ( n4587 & n4588 ) | ( ~n4269 & n4588 ) ;
  assign n4591 = ( n4261 & ~n4590 ) | ( n4261 & n4589 ) | ( ~n4590 & n4589 ) ;
  assign n4454 = ~n4439 & n4453 ;
  assign n4460 = ( n2033 & n4454 ) | ( n2033 & n4459 ) | ( n4454 & n4459 ) ;
  assign n4461 = ( n1827 & ~n4460 ) | ( n1827 & 1'b0 ) | ( ~n4460 & 1'b0 ) ;
  assign n4463 = ( n4153 & ~n4144 ) | ( n4153 & n4157 ) | ( ~n4144 & n4157 ) ;
  assign n4462 = ( n4157 & ~n4353 ) | ( n4157 & 1'b0 ) | ( ~n4353 & 1'b0 ) ;
  assign n4465 = ( n4157 & ~n4463 ) | ( n4157 & n4462 ) | ( ~n4463 & n4462 ) ;
  assign n4464 = ( n4462 & ~n4153 ) | ( n4462 & n4463 ) | ( ~n4153 & n4463 ) ;
  assign n4466 = ( n4144 & ~n4465 ) | ( n4144 & n4464 ) | ( ~n4465 & n4464 ) ;
  assign n4469 = n4459 | n4468 ;
  assign n4473 = ~n1827 & n4472 ;
  assign n4474 = n4469 &  n4473 ;
  assign n4475 = n4466 | n4474 ;
  assign n4476 = ~n4461 & n4475 ;
  assign n4477 = n4146 | n4353 ;
  assign n4478 = ( n4146 & ~n4159 ) | ( n4146 & n4151 ) | ( ~n4159 & n4151 ) ;
  assign n4479 = ( n4159 & n4477 ) | ( n4159 & n4478 ) | ( n4477 & n4478 ) ;
  assign n4480 = ( n4146 & ~n4478 ) | ( n4146 & n4477 ) | ( ~n4478 & n4477 ) ;
  assign n4481 = ( n4151 & ~n4479 ) | ( n4151 & n4480 ) | ( ~n4479 & n4480 ) ;
  assign n4482 = ( n1636 & n4476 ) | ( n1636 & n4481 ) | ( n4476 & n4481 ) ;
  assign n4483 = n1452 | n4482 ;
  assign n4484 = ( n4179 & ~n4353 ) | ( n4179 & 1'b0 ) | ( ~n4353 & 1'b0 ) ;
  assign n4485 = ( n4166 & n4175 ) | ( n4166 & n4179 ) | ( n4175 & n4179 ) ;
  assign n4486 = ( n4484 & ~n4175 ) | ( n4484 & n4485 ) | ( ~n4175 & n4485 ) ;
  assign n4487 = ( n4179 & ~n4485 ) | ( n4179 & n4484 ) | ( ~n4485 & n4484 ) ;
  assign n4488 = ( n4166 & ~n4486 ) | ( n4166 & n4487 ) | ( ~n4486 & n4487 ) ;
  assign n4489 = ( n1636 & ~n4461 ) | ( n1636 & 1'b0 ) | ( ~n4461 & 1'b0 ) ;
  assign n4490 = n4475 &  n4489 ;
  assign n4491 = n4481 | n4490 ;
  assign n4492 = n4469 &  n4472 ;
  assign n4493 = ( n4466 & ~n1827 ) | ( n4466 & n4492 ) | ( ~n1827 & n4492 ) ;
  assign n4494 = n1636 | n4493 ;
  assign n4495 = n1452 &  n4494 ;
  assign n4496 = n4491 &  n4495 ;
  assign n4497 = n4488 | n4496 ;
  assign n4498 = n4483 &  n4497 ;
  assign n4499 = n4181 &  n4353 ;
  assign n4500 = ( n4173 & ~n4168 ) | ( n4173 & n4353 ) | ( ~n4168 & n4353 ) ;
  assign n4502 = ( n4499 & n4168 ) | ( n4499 & n4500 ) | ( n4168 & n4500 ) ;
  assign n4501 = ( n4353 & ~n4500 ) | ( n4353 & n4499 ) | ( ~n4500 & n4499 ) ;
  assign n4503 = ( n4173 & ~n4502 ) | ( n4173 & n4501 ) | ( ~n4502 & n4501 ) ;
  assign n4504 = ( n4498 & ~n1283 ) | ( n4498 & n4503 ) | ( ~n1283 & n4503 ) ;
  assign n4505 = n1122 | n4504 ;
  assign n4506 = n4201 | n4353 ;
  assign n4507 = ( n4188 & ~n4197 ) | ( n4188 & n4201 ) | ( ~n4197 & n4201 ) ;
  assign n4508 = ( n4197 & n4506 ) | ( n4197 & n4507 ) | ( n4506 & n4507 ) ;
  assign n4509 = ( n4201 & ~n4507 ) | ( n4201 & n4506 ) | ( ~n4507 & n4506 ) ;
  assign n4510 = ( n4188 & ~n4508 ) | ( n4188 & n4509 ) | ( ~n4508 & n4509 ) ;
  assign n4511 = ~n1283 & n4483 ;
  assign n4512 = n4497 &  n4511 ;
  assign n4513 = n4503 | n4512 ;
  assign n4514 = n4491 &  n4494 ;
  assign n4515 = ( n1452 & n4488 ) | ( n1452 & n4514 ) | ( n4488 & n4514 ) ;
  assign n4516 = ( n1283 & ~n4515 ) | ( n1283 & 1'b0 ) | ( ~n4515 & 1'b0 ) ;
  assign n4517 = ( n1122 & ~n4516 ) | ( n1122 & 1'b0 ) | ( ~n4516 & 1'b0 ) ;
  assign n4518 = n4513 &  n4517 ;
  assign n4519 = n4510 | n4518 ;
  assign n4520 = n4505 &  n4519 ;
  assign n4521 = ( n4190 & ~n4353 ) | ( n4190 & 1'b0 ) | ( ~n4353 & 1'b0 ) ;
  assign n4522 = ( n4190 & n4195 ) | ( n4190 & n4203 ) | ( n4195 & n4203 ) ;
  assign n4523 = ( n4521 & ~n4203 ) | ( n4521 & n4522 ) | ( ~n4203 & n4522 ) ;
  assign n4524 = ( n4190 & ~n4522 ) | ( n4190 & n4521 ) | ( ~n4522 & n4521 ) ;
  assign n4525 = ( n4195 & ~n4523 ) | ( n4195 & n4524 ) | ( ~n4523 & n4524 ) ;
  assign n4526 = ( n976 & n4520 ) | ( n976 & n4525 ) | ( n4520 & n4525 ) ;
  assign n4527 = ( n837 & ~n4526 ) | ( n837 & 1'b0 ) | ( ~n4526 & 1'b0 ) ;
  assign n4529 = ( n4219 & ~n4210 ) | ( n4219 & n4223 ) | ( ~n4210 & n4223 ) ;
  assign n4528 = ( n4223 & ~n4353 ) | ( n4223 & 1'b0 ) | ( ~n4353 & 1'b0 ) ;
  assign n4531 = ( n4223 & ~n4529 ) | ( n4223 & n4528 ) | ( ~n4529 & n4528 ) ;
  assign n4530 = ( n4528 & ~n4219 ) | ( n4528 & n4529 ) | ( ~n4219 & n4529 ) ;
  assign n4532 = ( n4210 & ~n4531 ) | ( n4210 & n4530 ) | ( ~n4531 & n4530 ) ;
  assign n4533 = n976 &  n4505 ;
  assign n4534 = n4519 &  n4533 ;
  assign n4535 = n4525 | n4534 ;
  assign n4536 = ( n4513 & ~n4516 ) | ( n4513 & 1'b0 ) | ( ~n4516 & 1'b0 ) ;
  assign n4537 = ( n1122 & n4510 ) | ( n1122 & n4536 ) | ( n4510 & n4536 ) ;
  assign n4538 = n976 | n4537 ;
  assign n4539 = ~n837 & n4538 ;
  assign n4540 = n4535 &  n4539 ;
  assign n4541 = n4532 | n4540 ;
  assign n4542 = ~n4527 & n4541 ;
  assign n4543 = n4212 | n4353 ;
  assign n4544 = ( n4212 & ~n4225 ) | ( n4212 & n4217 ) | ( ~n4225 & n4217 ) ;
  assign n4545 = ( n4225 & n4543 ) | ( n4225 & n4544 ) | ( n4543 & n4544 ) ;
  assign n4546 = ( n4212 & ~n4544 ) | ( n4212 & n4543 ) | ( ~n4544 & n4543 ) ;
  assign n4547 = ( n4217 & ~n4545 ) | ( n4217 & n4546 ) | ( ~n4545 & n4546 ) ;
  assign n4548 = ( n4542 & ~n713 ) | ( n4542 & n4547 ) | ( ~n713 & n4547 ) ;
  assign n4549 = ( n595 & ~n4548 ) | ( n595 & 1'b0 ) | ( ~n4548 & 1'b0 ) ;
  assign n4550 = n4245 | n4353 ;
  assign n4551 = ( n4232 & ~n4245 ) | ( n4232 & n4241 ) | ( ~n4245 & n4241 ) ;
  assign n4553 = ( n4245 & n4550 ) | ( n4245 & n4551 ) | ( n4550 & n4551 ) ;
  assign n4552 = ( n4241 & ~n4551 ) | ( n4241 & n4550 ) | ( ~n4551 & n4550 ) ;
  assign n4554 = ( n4232 & ~n4553 ) | ( n4232 & n4552 ) | ( ~n4553 & n4552 ) ;
  assign n4555 = n713 | n4527 ;
  assign n4556 = ( n4541 & ~n4555 ) | ( n4541 & 1'b0 ) | ( ~n4555 & 1'b0 ) ;
  assign n4557 = n4547 | n4556 ;
  assign n4558 = n4535 &  n4538 ;
  assign n4559 = ( n4532 & ~n837 ) | ( n4532 & n4558 ) | ( ~n837 & n4558 ) ;
  assign n4560 = ( n713 & ~n4559 ) | ( n713 & 1'b0 ) | ( ~n4559 & 1'b0 ) ;
  assign n4561 = n595 | n4560 ;
  assign n4562 = ( n4557 & ~n4561 ) | ( n4557 & 1'b0 ) | ( ~n4561 & 1'b0 ) ;
  assign n4563 = n4554 | n4562 ;
  assign n4564 = ~n4549 & n4563 ;
  assign n4565 = n4247 &  n4353 ;
  assign n4566 = ( n4234 & n4239 ) | ( n4234 & n4353 ) | ( n4239 & n4353 ) ;
  assign n4568 = ( n4565 & ~n4234 ) | ( n4565 & n4566 ) | ( ~n4234 & n4566 ) ;
  assign n4567 = ( n4353 & ~n4566 ) | ( n4353 & n4565 ) | ( ~n4566 & n4565 ) ;
  assign n4569 = ( n4239 & ~n4568 ) | ( n4239 & n4567 ) | ( ~n4568 & n4567 ) ;
  assign n4570 = ( n492 & ~n4564 ) | ( n492 & n4569 ) | ( ~n4564 & n4569 ) ;
  assign n4571 = n396 &  n4570 ;
  assign n4573 = ( n4263 & ~n4254 ) | ( n4263 & n4267 ) | ( ~n4254 & n4267 ) ;
  assign n4572 = n4267 | n4353 ;
  assign n4575 = ( n4267 & ~n4573 ) | ( n4267 & n4572 ) | ( ~n4573 & n4572 ) ;
  assign n4574 = ( n4572 & ~n4263 ) | ( n4572 & n4573 ) | ( ~n4263 & n4573 ) ;
  assign n4576 = ( n4254 & ~n4575 ) | ( n4254 & n4574 ) | ( ~n4575 & n4574 ) ;
  assign n4577 = n492 | n4549 ;
  assign n4578 = ( n4563 & ~n4577 ) | ( n4563 & 1'b0 ) | ( ~n4577 & 1'b0 ) ;
  assign n4579 = ( n4569 & ~n4578 ) | ( n4569 & 1'b0 ) | ( ~n4578 & 1'b0 ) ;
  assign n4580 = ( n4557 & ~n4560 ) | ( n4557 & 1'b0 ) | ( ~n4560 & 1'b0 ) ;
  assign n4581 = ( n4554 & ~n595 ) | ( n4554 & n4580 ) | ( ~n595 & n4580 ) ;
  assign n4582 = ( n492 & ~n4581 ) | ( n492 & 1'b0 ) | ( ~n4581 & 1'b0 ) ;
  assign n4583 = n396 | n4582 ;
  assign n4584 = n4579 | n4583 ;
  assign n4585 = n4576 &  n4584 ;
  assign n4586 = n4571 | n4585 ;
  assign n4592 = ( n315 & ~n4591 ) | ( n315 & n4586 ) | ( ~n4591 & n4586 ) ;
  assign n4593 = n240 &  n4592 ;
  assign n4594 = n4284 | n4353 ;
  assign n4595 = ( n4276 & n4280 ) | ( n4276 & n4284 ) | ( n4280 & n4284 ) ;
  assign n4596 = ( n4594 & ~n4280 ) | ( n4594 & n4595 ) | ( ~n4280 & n4595 ) ;
  assign n4597 = ( n4284 & ~n4595 ) | ( n4284 & n4594 ) | ( ~n4595 & n4594 ) ;
  assign n4598 = ( n4276 & ~n4596 ) | ( n4276 & n4597 ) | ( ~n4596 & n4597 ) ;
  assign n4599 = n315 | n4571 ;
  assign n4600 = n4585 | n4599 ;
  assign n4601 = ~n4591 & n4600 ;
  assign n4602 = n4579 | n4582 ;
  assign n4603 = ( n396 & n4576 ) | ( n396 & n4602 ) | ( n4576 & n4602 ) ;
  assign n4604 = n315 &  n4603 ;
  assign n4605 = n240 | n4604 ;
  assign n4606 = n4601 | n4605 ;
  assign n4607 = ~n4598 & n4606 ;
  assign n4608 = n4593 | n4607 ;
  assign n4613 = ( n181 & ~n4612 ) | ( n181 & n4608 ) | ( ~n4612 & n4608 ) ;
  assign n4614 = ~n145 & n4613 ;
  assign n4616 = ( n4306 & ~n4297 ) | ( n4306 & n4310 ) | ( ~n4297 & n4310 ) ;
  assign n4615 = n4310 | n4353 ;
  assign n4618 = ( n4310 & ~n4616 ) | ( n4310 & n4615 ) | ( ~n4616 & n4615 ) ;
  assign n4617 = ( n4615 & ~n4306 ) | ( n4615 & n4616 ) | ( ~n4306 & n4616 ) ;
  assign n4619 = ( n4297 & ~n4618 ) | ( n4297 & n4617 ) | ( ~n4618 & n4617 ) ;
  assign n4620 = n181 | n4593 ;
  assign n4621 = n4607 | n4620 ;
  assign n4622 = ~n4612 & n4621 ;
  assign n4623 = n4601 | n4604 ;
  assign n4624 = ( n240 & ~n4598 ) | ( n240 & n4623 ) | ( ~n4598 & n4623 ) ;
  assign n4625 = n181 &  n4624 ;
  assign n4626 = ( n145 & ~n4625 ) | ( n145 & 1'b0 ) | ( ~n4625 & 1'b0 ) ;
  assign n4627 = ~n4622 & n4626 ;
  assign n4628 = n4619 | n4627 ;
  assign n4629 = ~n4614 & n4628 ;
  assign n4630 = n4299 | n4353 ;
  assign n4631 = ( n4304 & ~n4299 ) | ( n4304 & n4312 ) | ( ~n4299 & n4312 ) ;
  assign n4633 = ( n4299 & n4630 ) | ( n4299 & n4631 ) | ( n4630 & n4631 ) ;
  assign n4632 = ( n4312 & ~n4631 ) | ( n4312 & n4630 ) | ( ~n4631 & n4630 ) ;
  assign n4634 = ( n4304 & ~n4633 ) | ( n4304 & n4632 ) | ( ~n4633 & n4632 ) ;
  assign n4635 = ( n150 & ~n4629 ) | ( n150 & n4634 ) | ( ~n4629 & n4634 ) ;
  assign n4636 = ~n4319 & n4335 ;
  assign n4637 = ( n4338 & n4353 ) | ( n4338 & n4636 ) | ( n4353 & n4636 ) ;
  assign n4638 = ~n4338 & n4637 ;
  assign n4639 = ( n4335 & ~n4338 ) | ( n4335 & 1'b0 ) | ( ~n4338 & 1'b0 ) ;
  assign n4640 = ~n4353 & n4639 ;
  assign n4641 = ( n4319 & ~n4639 ) | ( n4319 & n4640 ) | ( ~n4639 & n4640 ) ;
  assign n4642 = n4638 | n4641 ;
  assign n4643 = ( n4320 & ~n4327 ) | ( n4320 & 1'b0 ) | ( ~n4327 & 1'b0 ) ;
  assign n4644 = ~n4353 & n4643 ;
  assign n4645 = ( n4341 & ~n4644 ) | ( n4341 & n4643 ) | ( ~n4644 & n4643 ) ;
  assign n4646 = ( n4642 & ~n4645 ) | ( n4642 & 1'b0 ) | ( ~n4645 & 1'b0 ) ;
  assign n4647 = ~n4635 & n4646 ;
  assign n4648 = ( n133 & ~n4647 ) | ( n133 & n4646 ) | ( ~n4647 & n4646 ) ;
  assign n4649 = n150 | n4614 ;
  assign n4650 = ( n4628 & ~n4649 ) | ( n4628 & 1'b0 ) | ( ~n4649 & 1'b0 ) ;
  assign n4655 = n4634 &  n4650 ;
  assign n4651 = n4622 | n4625 ;
  assign n4652 = ( n145 & ~n4651 ) | ( n145 & n4619 ) | ( ~n4651 & n4619 ) ;
  assign n4653 = ( n150 & ~n4652 ) | ( n150 & 1'b0 ) | ( ~n4652 & 1'b0 ) ;
  assign n4654 = n4642 | n4653 ;
  assign n4656 = ( n4634 & ~n4655 ) | ( n4634 & n4654 ) | ( ~n4655 & n4654 ) ;
  assign n4658 = ( n133 & ~n4327 ) | ( n133 & n4320 ) | ( ~n4327 & n4320 ) ;
  assign n4657 = ( n4327 & ~n4320 ) | ( n4327 & n4353 ) | ( ~n4320 & n4353 ) ;
  assign n4659 = ~n4327 & n4657 ;
  assign n4660 = ( n4327 & n4658 ) | ( n4327 & n4659 ) | ( n4658 & n4659 ) ;
  assign n4661 = n4323 | n4350 ;
  assign n4662 = ( n4326 & n4345 ) | ( n4326 & n4661 ) | ( n4345 & n4661 ) ;
  assign n4663 = ( n4326 & ~n4662 ) | ( n4326 & 1'b0 ) | ( ~n4662 & 1'b0 ) ;
  assign n4664 = ( n4333 & ~n4663 ) | ( n4333 & n4341 ) | ( ~n4663 & n4341 ) ;
  assign n4665 = ( n4333 & ~n4664 ) | ( n4333 & 1'b0 ) | ( ~n4664 & 1'b0 ) ;
  assign n4666 = n4660 | n4665 ;
  assign n4667 = ( n4656 & ~n4666 ) | ( n4656 & 1'b0 ) | ( ~n4666 & 1'b0 ) ;
  assign n4668 = ~n4648 | ~n4667 ;
  assign n4784 = ( n4472 & ~n4668 ) | ( n4472 & 1'b0 ) | ( ~n4668 & 1'b0 ) ;
  assign n4787 = ( n4472 & ~n4785 ) | ( n4472 & n4784 ) | ( ~n4785 & n4784 ) ;
  assign n4786 = ( n4784 & ~n4468 ) | ( n4784 & n4785 ) | ( ~n4468 & n4785 ) ;
  assign n4788 = ( n4459 & ~n4787 ) | ( n4459 & n4786 ) | ( ~n4787 & n4786 ) ;
  assign n4354 = x70 | x71 ;
  assign n4355 = x72 | n4354 ;
  assign n4669 = x72 &  n4668 ;
  assign n4670 = ( n4353 & ~n4355 ) | ( n4353 & n4669 ) | ( ~n4355 & n4669 ) ;
  assign n4671 = ( x72 & ~n4668 ) | ( x72 & x73 ) | ( ~n4668 & x73 ) ;
  assign n4677 = ( x72 & ~x73 ) | ( x72 & 1'b0 ) | ( ~x73 & 1'b0 ) ;
  assign n4672 = ~x72 & n4354 ;
  assign n4673 = ( x72 & ~n4351 ) | ( x72 & n4672 ) | ( ~n4351 & n4672 ) ;
  assign n4674 = ( n4333 & ~n4673 ) | ( n4333 & n4341 ) | ( ~n4673 & n4341 ) ;
  assign n4675 = ( n4333 & ~n4674 ) | ( n4333 & 1'b0 ) | ( ~n4674 & 1'b0 ) ;
  assign n4676 = ( n4668 & ~x73 ) | ( n4668 & n4675 ) | ( ~x73 & n4675 ) ;
  assign n4678 = ( n4671 & ~n4677 ) | ( n4671 & n4676 ) | ( ~n4677 & n4676 ) ;
  assign n4679 = ~n4670 & n4678 ;
  assign n4681 = ( n4353 & ~n4665 ) | ( n4353 & 1'b0 ) | ( ~n4665 & 1'b0 ) ;
  assign n4682 = ( n4656 & ~n4681 ) | ( n4656 & n4660 ) | ( ~n4681 & n4660 ) ;
  assign n4683 = ( n4656 & ~n4682 ) | ( n4656 & 1'b0 ) | ( ~n4682 & 1'b0 ) ;
  assign n4684 = n4648 &  n4683 ;
  assign n4680 = ~n4356 & n4668 ;
  assign n4685 = ( n4680 & ~n4684 ) | ( n4680 & 1'b0 ) | ( ~n4684 & 1'b0 ) ;
  assign n4686 = ( x74 & n4684 ) | ( x74 & n4685 ) | ( n4684 & n4685 ) ;
  assign n4687 = x74 | n4684 ;
  assign n4688 = n4680 | n4687 ;
  assign n4689 = ~n4686 & n4688 ;
  assign n4690 = ( n4679 & ~n4053 ) | ( n4679 & n4689 ) | ( ~n4053 & n4689 ) ;
  assign n4691 = ( n3760 & ~n4690 ) | ( n3760 & 1'b0 ) | ( ~n4690 & 1'b0 ) ;
  assign n4695 = ~x74 & n4353 ;
  assign n4696 = ( x75 & ~n4695 ) | ( x75 & 1'b0 ) | ( ~n4695 & 1'b0 ) ;
  assign n4697 = n4372 | n4696 ;
  assign n4692 = ( n4353 & ~x74 ) | ( n4353 & n4364 ) | ( ~x74 & n4364 ) ;
  assign n4693 = x74 &  n4692 ;
  assign n4694 = ( n4359 & ~n4693 ) | ( n4359 & n4364 ) | ( ~n4693 & n4364 ) ;
  assign n4698 = ( n4668 & ~n4697 ) | ( n4668 & n4694 ) | ( ~n4697 & n4694 ) ;
  assign n4700 = ( n4668 & ~n4698 ) | ( n4668 & 1'b0 ) | ( ~n4698 & 1'b0 ) ;
  assign n4699 = ~n4694 & n4698 ;
  assign n4701 = ( n4697 & ~n4700 ) | ( n4697 & n4699 ) | ( ~n4700 & n4699 ) ;
  assign n4702 = n4053 | n4670 ;
  assign n4703 = ( n4678 & ~n4702 ) | ( n4678 & 1'b0 ) | ( ~n4702 & 1'b0 ) ;
  assign n4704 = n4689 | n4703 ;
  assign n4705 = n4670 &  n4678 ;
  assign n4706 = ( n4053 & ~n4678 ) | ( n4053 & n4705 ) | ( ~n4678 & n4705 ) ;
  assign n4707 = n3760 | n4706 ;
  assign n4708 = ( n4704 & ~n4707 ) | ( n4704 & 1'b0 ) | ( ~n4707 & 1'b0 ) ;
  assign n4709 = n4701 | n4708 ;
  assign n4710 = ~n4691 & n4709 ;
  assign n4711 = ( n4369 & ~n4371 ) | ( n4369 & 1'b0 ) | ( ~n4371 & 1'b0 ) ;
  assign n4712 = ( n4371 & ~n4711 ) | ( n4371 & n4381 ) | ( ~n4711 & n4381 ) ;
  assign n4714 = ( n4668 & n4711 ) | ( n4668 & n4712 ) | ( n4711 & n4712 ) ;
  assign n4713 = ( n4371 & ~n4712 ) | ( n4371 & n4668 ) | ( ~n4712 & n4668 ) ;
  assign n4715 = ( n4381 & ~n4714 ) | ( n4381 & n4713 ) | ( ~n4714 & n4713 ) ;
  assign n4716 = ( n4710 & ~n3482 ) | ( n4710 & n4715 ) | ( ~n3482 & n4715 ) ;
  assign n4717 = ( n3211 & ~n4716 ) | ( n3211 & 1'b0 ) | ( ~n4716 & 1'b0 ) ;
  assign n4718 = n4406 | n4668 ;
  assign n4719 = ( n4393 & ~n4402 ) | ( n4393 & n4406 ) | ( ~n4402 & n4406 ) ;
  assign n4720 = ( n4402 & n4718 ) | ( n4402 & n4719 ) | ( n4718 & n4719 ) ;
  assign n4721 = ( n4406 & ~n4719 ) | ( n4406 & n4718 ) | ( ~n4719 & n4718 ) ;
  assign n4722 = ( n4393 & ~n4720 ) | ( n4393 & n4721 ) | ( ~n4720 & n4721 ) ;
  assign n4723 = n3482 | n4691 ;
  assign n4724 = ( n4709 & ~n4723 ) | ( n4709 & 1'b0 ) | ( ~n4723 & 1'b0 ) ;
  assign n4725 = n4715 | n4724 ;
  assign n4726 = ( n4704 & ~n4706 ) | ( n4704 & 1'b0 ) | ( ~n4706 & 1'b0 ) ;
  assign n4727 = ( n4701 & ~n3760 ) | ( n4701 & n4726 ) | ( ~n3760 & n4726 ) ;
  assign n4728 = ( n3482 & ~n4727 ) | ( n3482 & 1'b0 ) | ( ~n4727 & 1'b0 ) ;
  assign n4729 = n3211 | n4728 ;
  assign n4730 = ( n4725 & ~n4729 ) | ( n4725 & 1'b0 ) | ( ~n4729 & 1'b0 ) ;
  assign n4731 = n4722 | n4730 ;
  assign n4732 = ~n4717 & n4731 ;
  assign n4733 = n4395 | n4668 ;
  assign n4734 = ( n4400 & ~n4395 ) | ( n4400 & n4408 ) | ( ~n4395 & n4408 ) ;
  assign n4736 = ( n4395 & n4733 ) | ( n4395 & n4734 ) | ( n4733 & n4734 ) ;
  assign n4735 = ( n4408 & ~n4734 ) | ( n4408 & n4733 ) | ( ~n4734 & n4733 ) ;
  assign n4737 = ( n4400 & ~n4736 ) | ( n4400 & n4735 ) | ( ~n4736 & n4735 ) ;
  assign n4738 = ( n4732 & ~n2955 ) | ( n4732 & n4737 ) | ( ~n2955 & n4737 ) ;
  assign n4739 = ( n2706 & ~n4738 ) | ( n2706 & 1'b0 ) | ( ~n4738 & 1'b0 ) ;
  assign n4740 = n4428 | n4668 ;
  assign n4741 = ( n4415 & ~n4424 ) | ( n4415 & n4428 ) | ( ~n4424 & n4428 ) ;
  assign n4742 = ( n4424 & n4740 ) | ( n4424 & n4741 ) | ( n4740 & n4741 ) ;
  assign n4743 = ( n4428 & ~n4741 ) | ( n4428 & n4740 ) | ( ~n4741 & n4740 ) ;
  assign n4744 = ( n4415 & ~n4742 ) | ( n4415 & n4743 ) | ( ~n4742 & n4743 ) ;
  assign n4745 = n2955 | n4717 ;
  assign n4746 = ( n4731 & ~n4745 ) | ( n4731 & 1'b0 ) | ( ~n4745 & 1'b0 ) ;
  assign n4747 = n4737 | n4746 ;
  assign n4748 = ( n4725 & ~n4728 ) | ( n4725 & 1'b0 ) | ( ~n4728 & 1'b0 ) ;
  assign n4749 = ( n4722 & ~n3211 ) | ( n4722 & n4748 ) | ( ~n3211 & n4748 ) ;
  assign n4750 = ( n2955 & ~n4749 ) | ( n2955 & 1'b0 ) | ( ~n4749 & 1'b0 ) ;
  assign n4751 = n2706 | n4750 ;
  assign n4752 = ( n4747 & ~n4751 ) | ( n4747 & 1'b0 ) | ( ~n4751 & 1'b0 ) ;
  assign n4753 = n4744 | n4752 ;
  assign n4754 = ~n4739 & n4753 ;
  assign n4755 = n4417 | n4668 ;
  assign n4756 = ( n4417 & ~n4430 ) | ( n4417 & n4422 ) | ( ~n4430 & n4422 ) ;
  assign n4757 = ( n4430 & n4755 ) | ( n4430 & n4756 ) | ( n4755 & n4756 ) ;
  assign n4758 = ( n4417 & ~n4756 ) | ( n4417 & n4755 ) | ( ~n4756 & n4755 ) ;
  assign n4759 = ( n4422 & ~n4757 ) | ( n4422 & n4758 ) | ( ~n4757 & n4758 ) ;
  assign n4760 = ( n4754 & ~n2472 ) | ( n4754 & n4759 ) | ( ~n2472 & n4759 ) ;
  assign n4761 = ( n2245 & ~n4760 ) | ( n2245 & 1'b0 ) | ( ~n4760 & 1'b0 ) ;
  assign n4762 = n4450 | n4668 ;
  assign n4763 = ( n4437 & ~n4450 ) | ( n4437 & n4446 ) | ( ~n4450 & n4446 ) ;
  assign n4765 = ( n4450 & n4762 ) | ( n4450 & n4763 ) | ( n4762 & n4763 ) ;
  assign n4764 = ( n4446 & ~n4763 ) | ( n4446 & n4762 ) | ( ~n4763 & n4762 ) ;
  assign n4766 = ( n4437 & ~n4765 ) | ( n4437 & n4764 ) | ( ~n4765 & n4764 ) ;
  assign n4767 = n2472 | n4739 ;
  assign n4768 = ( n4753 & ~n4767 ) | ( n4753 & 1'b0 ) | ( ~n4767 & 1'b0 ) ;
  assign n4769 = n4759 | n4768 ;
  assign n4770 = ( n4747 & ~n4750 ) | ( n4747 & 1'b0 ) | ( ~n4750 & 1'b0 ) ;
  assign n4771 = ( n4744 & ~n2706 ) | ( n4744 & n4770 ) | ( ~n2706 & n4770 ) ;
  assign n4772 = ( n2472 & ~n4771 ) | ( n2472 & 1'b0 ) | ( ~n4771 & 1'b0 ) ;
  assign n4773 = n2245 | n4772 ;
  assign n4774 = ( n4769 & ~n4773 ) | ( n4769 & 1'b0 ) | ( ~n4773 & 1'b0 ) ;
  assign n4775 = n4766 | n4774 ;
  assign n4776 = ~n4761 & n4775 ;
  assign n4777 = n4452 &  n4668 ;
  assign n4778 = ( n4439 & n4444 ) | ( n4439 & n4668 ) | ( n4444 & n4668 ) ;
  assign n4780 = ( n4777 & ~n4439 ) | ( n4777 & n4778 ) | ( ~n4439 & n4778 ) ;
  assign n4779 = ( n4668 & ~n4778 ) | ( n4668 & n4777 ) | ( ~n4778 & n4777 ) ;
  assign n4781 = ( n4444 & ~n4780 ) | ( n4444 & n4779 ) | ( ~n4780 & n4779 ) ;
  assign n4782 = ( n2033 & n4776 ) | ( n2033 & n4781 ) | ( n4776 & n4781 ) ;
  assign n4783 = ( n1827 & ~n4782 ) | ( n1827 & 1'b0 ) | ( ~n4782 & 1'b0 ) ;
  assign n4789 = ( n2033 & ~n4761 ) | ( n2033 & 1'b0 ) | ( ~n4761 & 1'b0 ) ;
  assign n4790 = n4775 &  n4789 ;
  assign n4791 = n4781 | n4790 ;
  assign n4792 = ( n4769 & ~n4772 ) | ( n4769 & 1'b0 ) | ( ~n4772 & 1'b0 ) ;
  assign n4793 = ( n4766 & ~n2245 ) | ( n4766 & n4792 ) | ( ~n2245 & n4792 ) ;
  assign n4794 = n2033 | n4793 ;
  assign n4795 = ~n1827 & n4794 ;
  assign n4796 = n4791 &  n4795 ;
  assign n4932 = ( n4593 & ~n4598 ) | ( n4593 & n4606 ) | ( ~n4598 & n4606 ) ;
  assign n4931 = n4593 | n4668 ;
  assign n4934 = ( n4593 & ~n4932 ) | ( n4593 & n4931 ) | ( ~n4932 & n4931 ) ;
  assign n4933 = ( n4931 & ~n4606 ) | ( n4931 & n4932 ) | ( ~n4606 & n4932 ) ;
  assign n4935 = ( n4598 & ~n4934 ) | ( n4598 & n4933 ) | ( ~n4934 & n4933 ) ;
  assign n4797 = n4788 | n4796 ;
  assign n4798 = ~n4783 & n4797 ;
  assign n4799 = n4461 | n4668 ;
  assign n4800 = ( n4466 & ~n4461 ) | ( n4466 & n4474 ) | ( ~n4461 & n4474 ) ;
  assign n4802 = ( n4461 & n4799 ) | ( n4461 & n4800 ) | ( n4799 & n4800 ) ;
  assign n4801 = ( n4474 & ~n4800 ) | ( n4474 & n4799 ) | ( ~n4800 & n4799 ) ;
  assign n4803 = ( n4466 & ~n4802 ) | ( n4466 & n4801 ) | ( ~n4802 & n4801 ) ;
  assign n4804 = ( n1636 & n4798 ) | ( n1636 & n4803 ) | ( n4798 & n4803 ) ;
  assign n4805 = n1452 | n4804 ;
  assign n4807 = ( n4490 & ~n4481 ) | ( n4490 & n4494 ) | ( ~n4481 & n4494 ) ;
  assign n4806 = ( n4494 & ~n4668 ) | ( n4494 & 1'b0 ) | ( ~n4668 & 1'b0 ) ;
  assign n4809 = ( n4494 & ~n4807 ) | ( n4494 & n4806 ) | ( ~n4807 & n4806 ) ;
  assign n4808 = ( n4806 & ~n4490 ) | ( n4806 & n4807 ) | ( ~n4490 & n4807 ) ;
  assign n4810 = ( n4481 & ~n4809 ) | ( n4481 & n4808 ) | ( ~n4809 & n4808 ) ;
  assign n4811 = ( n1636 & ~n4783 ) | ( n1636 & 1'b0 ) | ( ~n4783 & 1'b0 ) ;
  assign n4812 = n4797 &  n4811 ;
  assign n4813 = n4803 | n4812 ;
  assign n4814 = n4791 &  n4794 ;
  assign n4815 = ( n4788 & ~n1827 ) | ( n4788 & n4814 ) | ( ~n1827 & n4814 ) ;
  assign n4816 = n1636 | n4815 ;
  assign n4817 = n1452 &  n4816 ;
  assign n4818 = n4813 &  n4817 ;
  assign n4819 = n4810 | n4818 ;
  assign n4820 = n4805 &  n4819 ;
  assign n4822 = ( n4483 & ~n4488 ) | ( n4483 & n4496 ) | ( ~n4488 & n4496 ) ;
  assign n4821 = ( n4483 & ~n4668 ) | ( n4483 & 1'b0 ) | ( ~n4668 & 1'b0 ) ;
  assign n4824 = ( n4483 & ~n4822 ) | ( n4483 & n4821 ) | ( ~n4822 & n4821 ) ;
  assign n4823 = ( n4821 & ~n4496 ) | ( n4821 & n4822 ) | ( ~n4496 & n4822 ) ;
  assign n4825 = ( n4488 & ~n4824 ) | ( n4488 & n4823 ) | ( ~n4824 & n4823 ) ;
  assign n4826 = ( n4820 & ~n1283 ) | ( n4820 & n4825 ) | ( ~n1283 & n4825 ) ;
  assign n4827 = n1122 | n4826 ;
  assign n4828 = n4516 | n4668 ;
  assign n4829 = ( n4503 & ~n4516 ) | ( n4503 & n4512 ) | ( ~n4516 & n4512 ) ;
  assign n4831 = ( n4516 & n4828 ) | ( n4516 & n4829 ) | ( n4828 & n4829 ) ;
  assign n4830 = ( n4512 & ~n4829 ) | ( n4512 & n4828 ) | ( ~n4829 & n4828 ) ;
  assign n4832 = ( n4503 & ~n4831 ) | ( n4503 & n4830 ) | ( ~n4831 & n4830 ) ;
  assign n4833 = ~n1283 & n4805 ;
  assign n4834 = n4819 &  n4833 ;
  assign n4835 = n4825 | n4834 ;
  assign n4836 = n4813 &  n4816 ;
  assign n4837 = ( n1452 & n4810 ) | ( n1452 & n4836 ) | ( n4810 & n4836 ) ;
  assign n4838 = ( n1283 & ~n4837 ) | ( n1283 & 1'b0 ) | ( ~n4837 & 1'b0 ) ;
  assign n4839 = ( n1122 & ~n4838 ) | ( n1122 & 1'b0 ) | ( ~n4838 & 1'b0 ) ;
  assign n4840 = n4835 &  n4839 ;
  assign n4841 = n4832 | n4840 ;
  assign n4842 = n4827 &  n4841 ;
  assign n4843 = n4518 &  n4668 ;
  assign n4844 = ( n4505 & ~n4668 ) | ( n4505 & n4510 ) | ( ~n4668 & n4510 ) ;
  assign n4845 = ( n4668 & n4843 ) | ( n4668 & n4844 ) | ( n4843 & n4844 ) ;
  assign n4846 = ( n4505 & ~n4844 ) | ( n4505 & n4843 ) | ( ~n4844 & n4843 ) ;
  assign n4847 = ( n4510 & ~n4845 ) | ( n4510 & n4846 ) | ( ~n4845 & n4846 ) ;
  assign n4848 = ( n976 & n4842 ) | ( n976 & n4847 ) | ( n4842 & n4847 ) ;
  assign n4849 = ( n837 & ~n4848 ) | ( n837 & 1'b0 ) | ( ~n4848 & 1'b0 ) ;
  assign n4851 = ( n4534 & ~n4525 ) | ( n4534 & n4538 ) | ( ~n4525 & n4538 ) ;
  assign n4850 = ( n4538 & ~n4668 ) | ( n4538 & 1'b0 ) | ( ~n4668 & 1'b0 ) ;
  assign n4853 = ( n4538 & ~n4851 ) | ( n4538 & n4850 ) | ( ~n4851 & n4850 ) ;
  assign n4852 = ( n4850 & ~n4534 ) | ( n4850 & n4851 ) | ( ~n4534 & n4851 ) ;
  assign n4854 = ( n4525 & ~n4853 ) | ( n4525 & n4852 ) | ( ~n4853 & n4852 ) ;
  assign n4855 = n976 &  n4827 ;
  assign n4856 = n4841 &  n4855 ;
  assign n4857 = n4847 | n4856 ;
  assign n4858 = ( n4835 & ~n4838 ) | ( n4835 & 1'b0 ) | ( ~n4838 & 1'b0 ) ;
  assign n4859 = ( n1122 & n4832 ) | ( n1122 & n4858 ) | ( n4832 & n4858 ) ;
  assign n4860 = n976 | n4859 ;
  assign n4861 = ~n837 & n4860 ;
  assign n4862 = n4857 &  n4861 ;
  assign n4863 = n4854 | n4862 ;
  assign n4864 = ~n4849 & n4863 ;
  assign n4865 = n4527 | n4668 ;
  assign n4866 = ( n4532 & ~n4527 ) | ( n4532 & n4540 ) | ( ~n4527 & n4540 ) ;
  assign n4868 = ( n4527 & n4865 ) | ( n4527 & n4866 ) | ( n4865 & n4866 ) ;
  assign n4867 = ( n4540 & ~n4866 ) | ( n4540 & n4865 ) | ( ~n4866 & n4865 ) ;
  assign n4869 = ( n4532 & ~n4868 ) | ( n4532 & n4867 ) | ( ~n4868 & n4867 ) ;
  assign n4870 = ( n4864 & ~n713 ) | ( n4864 & n4869 ) | ( ~n713 & n4869 ) ;
  assign n4871 = ( n595 & ~n4870 ) | ( n595 & 1'b0 ) | ( ~n4870 & 1'b0 ) ;
  assign n4872 = n4560 | n4668 ;
  assign n4873 = ( n4547 & ~n4556 ) | ( n4547 & n4560 ) | ( ~n4556 & n4560 ) ;
  assign n4874 = ( n4556 & n4872 ) | ( n4556 & n4873 ) | ( n4872 & n4873 ) ;
  assign n4875 = ( n4560 & ~n4873 ) | ( n4560 & n4872 ) | ( ~n4873 & n4872 ) ;
  assign n4876 = ( n4547 & ~n4874 ) | ( n4547 & n4875 ) | ( ~n4874 & n4875 ) ;
  assign n4877 = n713 | n4849 ;
  assign n4878 = ( n4863 & ~n4877 ) | ( n4863 & 1'b0 ) | ( ~n4877 & 1'b0 ) ;
  assign n4879 = n4869 | n4878 ;
  assign n4880 = n4857 &  n4860 ;
  assign n4881 = ( n4854 & ~n837 ) | ( n4854 & n4880 ) | ( ~n837 & n4880 ) ;
  assign n4882 = ( n713 & ~n4881 ) | ( n713 & 1'b0 ) | ( ~n4881 & 1'b0 ) ;
  assign n4883 = n595 | n4882 ;
  assign n4884 = ( n4879 & ~n4883 ) | ( n4879 & 1'b0 ) | ( ~n4883 & 1'b0 ) ;
  assign n4885 = n4876 | n4884 ;
  assign n4886 = ~n4871 & n4885 ;
  assign n4887 = n4549 | n4668 ;
  assign n4888 = ( n4549 & ~n4562 ) | ( n4549 & n4554 ) | ( ~n4562 & n4554 ) ;
  assign n4889 = ( n4562 & n4887 ) | ( n4562 & n4888 ) | ( n4887 & n4888 ) ;
  assign n4890 = ( n4549 & ~n4888 ) | ( n4549 & n4887 ) | ( ~n4888 & n4887 ) ;
  assign n4891 = ( n4554 & ~n4889 ) | ( n4554 & n4890 ) | ( ~n4889 & n4890 ) ;
  assign n4892 = ( n4886 & ~n492 ) | ( n4886 & n4891 ) | ( ~n492 & n4891 ) ;
  assign n4893 = ( n396 & ~n4892 ) | ( n396 & 1'b0 ) | ( ~n4892 & 1'b0 ) ;
  assign n4894 = n4582 | n4668 ;
  assign n4895 = ( n4569 & ~n4578 ) | ( n4569 & n4582 ) | ( ~n4578 & n4582 ) ;
  assign n4896 = ( n4578 & n4894 ) | ( n4578 & n4895 ) | ( n4894 & n4895 ) ;
  assign n4897 = ( n4582 & ~n4895 ) | ( n4582 & n4894 ) | ( ~n4895 & n4894 ) ;
  assign n4898 = ( n4569 & ~n4896 ) | ( n4569 & n4897 ) | ( ~n4896 & n4897 ) ;
  assign n4899 = n492 | n4871 ;
  assign n4900 = ( n4885 & ~n4899 ) | ( n4885 & 1'b0 ) | ( ~n4899 & 1'b0 ) ;
  assign n4901 = n4891 | n4900 ;
  assign n4902 = ( n4879 & ~n4882 ) | ( n4879 & 1'b0 ) | ( ~n4882 & 1'b0 ) ;
  assign n4903 = ( n4876 & ~n595 ) | ( n4876 & n4902 ) | ( ~n595 & n4902 ) ;
  assign n4904 = ( n492 & ~n4903 ) | ( n492 & 1'b0 ) | ( ~n4903 & 1'b0 ) ;
  assign n4905 = n396 | n4904 ;
  assign n4906 = ( n4901 & ~n4905 ) | ( n4901 & 1'b0 ) | ( ~n4905 & 1'b0 ) ;
  assign n4907 = ( n4898 & ~n4906 ) | ( n4898 & 1'b0 ) | ( ~n4906 & 1'b0 ) ;
  assign n4908 = n4893 | n4907 ;
  assign n4909 = ~n4584 & n4668 ;
  assign n4910 = ( n4571 & n4576 ) | ( n4571 & n4668 ) | ( n4576 & n4668 ) ;
  assign n4912 = ( n4909 & ~n4571 ) | ( n4909 & n4910 ) | ( ~n4571 & n4910 ) ;
  assign n4911 = ( n4668 & ~n4910 ) | ( n4668 & n4909 ) | ( ~n4910 & n4909 ) ;
  assign n4913 = ( n4576 & ~n4912 ) | ( n4576 & n4911 ) | ( ~n4912 & n4911 ) ;
  assign n4914 = ( n315 & n4908 ) | ( n315 & n4913 ) | ( n4908 & n4913 ) ;
  assign n4915 = n240 &  n4914 ;
  assign n4916 = n4604 | n4668 ;
  assign n4917 = ( n4591 & n4600 ) | ( n4591 & n4604 ) | ( n4600 & n4604 ) ;
  assign n4918 = ( n4916 & ~n4600 ) | ( n4916 & n4917 ) | ( ~n4600 & n4917 ) ;
  assign n4919 = ( n4604 & ~n4917 ) | ( n4604 & n4916 ) | ( ~n4917 & n4916 ) ;
  assign n4920 = ( n4591 & ~n4918 ) | ( n4591 & n4919 ) | ( ~n4918 & n4919 ) ;
  assign n4921 = n315 | n4893 ;
  assign n4922 = n4907 | n4921 ;
  assign n4923 = n4913 &  n4922 ;
  assign n4924 = ( n4901 & ~n4904 ) | ( n4901 & 1'b0 ) | ( ~n4904 & 1'b0 ) ;
  assign n4925 = ( n396 & ~n4924 ) | ( n396 & n4898 ) | ( ~n4924 & n4898 ) ;
  assign n4926 = n315 &  n4925 ;
  assign n4927 = n240 | n4926 ;
  assign n4928 = n4923 | n4927 ;
  assign n4929 = ~n4920 & n4928 ;
  assign n4930 = n4915 | n4929 ;
  assign n4936 = ( n181 & ~n4935 ) | ( n181 & n4930 ) | ( ~n4935 & n4930 ) ;
  assign n4937 = ~n145 & n4936 ;
  assign n4938 = n181 | n4915 ;
  assign n4939 = n4929 | n4938 ;
  assign n4940 = ~n4935 & n4939 ;
  assign n4941 = n4923 | n4926 ;
  assign n4942 = ( n240 & ~n4920 ) | ( n240 & n4941 ) | ( ~n4920 & n4941 ) ;
  assign n4943 = n181 &  n4942 ;
  assign n4944 = ( n145 & ~n4943 ) | ( n145 & 1'b0 ) | ( ~n4943 & 1'b0 ) ;
  assign n4945 = ~n4940 & n4944 ;
  assign n4946 = ( n4621 & ~n4612 ) | ( n4621 & n4625 ) | ( ~n4612 & n4625 ) ;
  assign n4948 = ( n4668 & ~n4946 ) | ( n4668 & n4625 ) | ( ~n4946 & n4625 ) ;
  assign n4947 = ( n4946 & ~n4621 ) | ( n4946 & n4668 ) | ( ~n4621 & n4668 ) ;
  assign n4949 = ( n4612 & ~n4948 ) | ( n4612 & n4947 ) | ( ~n4948 & n4947 ) ;
  assign n4950 = n4945 | n4949 ;
  assign n4951 = ~n4937 & n4950 ;
  assign n4952 = n4614 | n4668 ;
  assign n4953 = ( n4614 & ~n4627 ) | ( n4614 & n4619 ) | ( ~n4627 & n4619 ) ;
  assign n4954 = ( n4627 & n4952 ) | ( n4627 & n4953 ) | ( n4952 & n4953 ) ;
  assign n4955 = ( n4614 & ~n4953 ) | ( n4614 & n4952 ) | ( ~n4953 & n4952 ) ;
  assign n4956 = ( n4619 & ~n4954 ) | ( n4619 & n4955 ) | ( ~n4954 & n4955 ) ;
  assign n4957 = ( n4951 & ~n150 ) | ( n4951 & n4956 ) | ( ~n150 & n4956 ) ;
  assign n4958 = n4634 | n4653 ;
  assign n4959 = ( n4650 & ~n4958 ) | ( n4650 & n4668 ) | ( ~n4958 & n4668 ) ;
  assign n4960 = ~n4650 & n4959 ;
  assign n4961 = n4650 | n4653 ;
  assign n4962 = n4668 | n4961 ;
  assign n4963 = ( n4634 & ~n4962 ) | ( n4634 & n4961 ) | ( ~n4962 & n4961 ) ;
  assign n4964 = n4960 | n4963 ;
  assign n4965 = n4635 &  n4642 ;
  assign n4966 = ~n4668 & n4965 ;
  assign n4967 = ( n4656 & ~n4965 ) | ( n4656 & n4966 ) | ( ~n4965 & n4966 ) ;
  assign n4968 = n4964 &  n4967 ;
  assign n4969 = n4957 &  n4968 ;
  assign n4970 = ( n133 & ~n4969 ) | ( n133 & n4968 ) | ( ~n4969 & n4968 ) ;
  assign n4973 = n4940 | n4943 ;
  assign n4974 = ( n145 & ~n4973 ) | ( n145 & n4949 ) | ( ~n4973 & n4949 ) ;
  assign n4975 = ( n150 & ~n4974 ) | ( n150 & 1'b0 ) | ( ~n4974 & 1'b0 ) ;
  assign n4976 = n4964 | n4975 ;
  assign n4971 = n150 | n4937 ;
  assign n4972 = ( n4950 & ~n4971 ) | ( n4950 & 1'b0 ) | ( ~n4971 & 1'b0 ) ;
  assign n4977 = ~n4956 & n4972 ;
  assign n4978 = ( n4956 & ~n4976 ) | ( n4956 & n4977 ) | ( ~n4976 & n4977 ) ;
  assign n4980 = ( n133 & n4635 ) | ( n133 & n4642 ) | ( n4635 & n4642 ) ;
  assign n4979 = ( n4635 & ~n4668 ) | ( n4635 & n4642 ) | ( ~n4668 & n4642 ) ;
  assign n4981 = ( n4642 & ~n4979 ) | ( n4642 & 1'b0 ) | ( ~n4979 & 1'b0 ) ;
  assign n4982 = ( n4980 & ~n4642 ) | ( n4980 & n4981 ) | ( ~n4642 & n4981 ) ;
  assign n4983 = n4638 | n4665 ;
  assign n4984 = ( n4660 & ~n4641 ) | ( n4660 & n4983 ) | ( ~n4641 & n4983 ) ;
  assign n4985 = n4641 | n4984 ;
  assign n4986 = ( n4648 & ~n4656 ) | ( n4648 & n4985 ) | ( ~n4656 & n4985 ) ;
  assign n4987 = ( n4648 & ~n4986 ) | ( n4648 & 1'b0 ) | ( ~n4986 & 1'b0 ) ;
  assign n4988 = n4982 | n4987 ;
  assign n4989 = n4978 | n4988 ;
  assign n4990 = ~n4970 |  n4989 ;
  assign n5136 = n4796 &  n4990 ;
  assign n5137 = ( n4783 & ~n5136 ) | ( n4783 & n4990 ) | ( ~n5136 & n4990 ) ;
  assign n5138 = ( n4788 & ~n4783 ) | ( n4788 & n5137 ) | ( ~n4783 & n5137 ) ;
  assign n5139 = ( n4783 & ~n5137 ) | ( n4783 & n4788 ) | ( ~n5137 & n4788 ) ;
  assign n5140 = ( n5138 & ~n4788 ) | ( n5138 & n5139 ) | ( ~n4788 & n5139 ) ;
  assign n5121 = ( n4794 & ~n4990 ) | ( n4794 & 1'b0 ) | ( ~n4990 & 1'b0 ) ;
  assign n5122 = ( n4781 & n4790 ) | ( n4781 & n4794 ) | ( n4790 & n4794 ) ;
  assign n5123 = ( n5121 & ~n4790 ) | ( n5121 & n5122 ) | ( ~n4790 & n5122 ) ;
  assign n5124 = ( n4794 & ~n5122 ) | ( n4794 & n5121 ) | ( ~n5122 & n5121 ) ;
  assign n5125 = ( n4781 & ~n5123 ) | ( n4781 & n5124 ) | ( ~n5123 & n5124 ) ;
  assign n5114 = n4761 | n4990 ;
  assign n5115 = ( n4761 & ~n4774 ) | ( n4761 & n4766 ) | ( ~n4774 & n4766 ) ;
  assign n5116 = ( n4774 & n5114 ) | ( n4774 & n5115 ) | ( n5114 & n5115 ) ;
  assign n5117 = ( n4761 & ~n5115 ) | ( n4761 & n5114 ) | ( ~n5115 & n5114 ) ;
  assign n5118 = ( n4766 & ~n5116 ) | ( n4766 & n5117 ) | ( ~n5116 & n5117 ) ;
  assign n5099 = n4772 | n4990 ;
  assign n5100 = ( n4759 & ~n4768 ) | ( n4759 & n4772 ) | ( ~n4768 & n4772 ) ;
  assign n5101 = ( n4768 & n5099 ) | ( n4768 & n5100 ) | ( n5099 & n5100 ) ;
  assign n5102 = ( n4772 & ~n5100 ) | ( n4772 & n5099 ) | ( ~n5100 & n5099 ) ;
  assign n5103 = ( n4759 & ~n5101 ) | ( n4759 & n5102 ) | ( ~n5101 & n5102 ) ;
  assign n5092 = n4739 | n4990 ;
  assign n5093 = ( n4744 & ~n4739 ) | ( n4744 & n4752 ) | ( ~n4739 & n4752 ) ;
  assign n5095 = ( n4739 & n5092 ) | ( n4739 & n5093 ) | ( n5092 & n5093 ) ;
  assign n5094 = ( n4752 & ~n5093 ) | ( n4752 & n5092 ) | ( ~n5093 & n5092 ) ;
  assign n5096 = ( n4744 & ~n5095 ) | ( n4744 & n5094 ) | ( ~n5095 & n5094 ) ;
  assign n5077 = n4750 | n4990 ;
  assign n5078 = ( n4737 & ~n4746 ) | ( n4737 & n4750 ) | ( ~n4746 & n4750 ) ;
  assign n5079 = ( n4746 & n5077 ) | ( n4746 & n5078 ) | ( n5077 & n5078 ) ;
  assign n5080 = ( n4750 & ~n5078 ) | ( n4750 & n5077 ) | ( ~n5078 & n5077 ) ;
  assign n5081 = ( n4737 & ~n5079 ) | ( n4737 & n5080 ) | ( ~n5079 & n5080 ) ;
  assign n5070 = n4730 &  n4990 ;
  assign n5071 = ( n4717 & n4722 ) | ( n4717 & n4990 ) | ( n4722 & n4990 ) ;
  assign n5073 = ( n5070 & ~n4717 ) | ( n5070 & n5071 ) | ( ~n4717 & n5071 ) ;
  assign n5072 = ( n4990 & ~n5071 ) | ( n4990 & n5070 ) | ( ~n5071 & n5070 ) ;
  assign n5074 = ( n4722 & ~n5073 ) | ( n4722 & n5072 ) | ( ~n5073 & n5072 ) ;
  assign n5055 = n4728 | n4990 ;
  assign n5056 = ( n4715 & ~n4728 ) | ( n4715 & n4724 ) | ( ~n4728 & n4724 ) ;
  assign n5058 = ( n4728 & n5055 ) | ( n4728 & n5056 ) | ( n5055 & n5056 ) ;
  assign n5057 = ( n4724 & ~n5056 ) | ( n4724 & n5055 ) | ( ~n5056 & n5055 ) ;
  assign n5059 = ( n4715 & ~n5058 ) | ( n4715 & n5057 ) | ( ~n5058 & n5057 ) ;
  assign n5048 = n4691 | n4990 ;
  assign n5049 = ( n4691 & ~n4708 ) | ( n4691 & n4701 ) | ( ~n4708 & n4701 ) ;
  assign n5050 = ( n4708 & n5048 ) | ( n4708 & n5049 ) | ( n5048 & n5049 ) ;
  assign n5051 = ( n4691 & ~n5049 ) | ( n4691 & n5048 ) | ( ~n5049 & n5048 ) ;
  assign n5052 = ( n4701 & ~n5050 ) | ( n4701 & n5051 ) | ( ~n5050 & n5051 ) ;
  assign n5033 = ~n4703 & n4706 ;
  assign n5034 = ( n4689 & ~n4703 ) | ( n4689 & n5033 ) | ( ~n4703 & n5033 ) ;
  assign n5036 = ( n4703 & n4990 ) | ( n4703 & n5034 ) | ( n4990 & n5034 ) ;
  assign n5035 = ( n4990 & ~n5034 ) | ( n4990 & n5033 ) | ( ~n5034 & n5033 ) ;
  assign n5037 = ( n4689 & ~n5036 ) | ( n4689 & n5035 ) | ( ~n5036 & n5035 ) ;
  assign n5024 = ~x72 & n4668 ;
  assign n5025 = ( x73 & ~n5024 ) | ( x73 & 1'b0 ) | ( ~n5024 & 1'b0 ) ;
  assign n5026 = n4680 | n5025 ;
  assign n5021 = ( n4668 & ~x72 ) | ( n4668 & n4675 ) | ( ~x72 & n4675 ) ;
  assign n5022 = x72 &  n5021 ;
  assign n5023 = ( n4670 & ~n5022 ) | ( n4670 & n4675 ) | ( ~n5022 & n4675 ) ;
  assign n5027 = ( n4990 & ~n5026 ) | ( n4990 & n5023 ) | ( ~n5026 & n5023 ) ;
  assign n5029 = ( n4990 & ~n5027 ) | ( n4990 & 1'b0 ) | ( ~n5027 & 1'b0 ) ;
  assign n5028 = ~n5023 & n5027 ;
  assign n5030 = ( n5026 & ~n5029 ) | ( n5026 & n5028 ) | ( ~n5029 & n5028 ) ;
  assign n4997 = ( x70 & ~n4990 ) | ( x70 & x71 ) | ( ~n4990 & x71 ) ;
  assign n5003 = ( x70 & ~x71 ) | ( x70 & 1'b0 ) | ( ~x71 & 1'b0 ) ;
  assign n4993 = x68 | x69 ;
  assign n4998 = ~x70 & n4993 ;
  assign n4999 = ( x70 & ~n4666 ) | ( x70 & n4998 ) | ( ~n4666 & n4998 ) ;
  assign n5000 = ( n4656 & ~n4648 ) | ( n4656 & n4999 ) | ( ~n4648 & n4999 ) ;
  assign n5001 = n4648 &  n5000 ;
  assign n5002 = ( n4990 & ~x71 ) | ( n4990 & n5001 ) | ( ~x71 & n5001 ) ;
  assign n5004 = ( n4997 & ~n5003 ) | ( n4997 & n5002 ) | ( ~n5003 & n5002 ) ;
  assign n4994 = x70 | n4993 ;
  assign n4995 = x70 &  n4990 ;
  assign n4996 = ( n4668 & ~n4994 ) | ( n4668 & n4995 ) | ( ~n4994 & n4995 ) ;
  assign n5007 = n4353 | n4996 ;
  assign n5008 = ( n5004 & ~n5007 ) | ( n5004 & 1'b0 ) | ( ~n5007 & 1'b0 ) ;
  assign n5010 = ( n4668 & ~n4987 ) | ( n4668 & 1'b0 ) | ( ~n4987 & 1'b0 ) ;
  assign n5011 = ( n4978 & ~n4982 ) | ( n4978 & n5010 ) | ( ~n4982 & n5010 ) ;
  assign n5012 = ~n4978 & n5011 ;
  assign n5013 = n4970 &  n5012 ;
  assign n5009 = ~n4354 & n4990 ;
  assign n5014 = ( n5009 & ~n5013 ) | ( n5009 & 1'b0 ) | ( ~n5013 & 1'b0 ) ;
  assign n5015 = ( x72 & n5013 ) | ( x72 & n5014 ) | ( n5013 & n5014 ) ;
  assign n5016 = x72 | n5013 ;
  assign n5017 = n5009 | n5016 ;
  assign n5018 = ~n5015 & n5017 ;
  assign n5019 = n5008 | n5018 ;
  assign n5005 = n4996 &  n5004 ;
  assign n5006 = ( n4353 & ~n5004 ) | ( n4353 & n5005 ) | ( ~n5004 & n5005 ) ;
  assign n5038 = n4053 | n5006 ;
  assign n5039 = ( n5019 & ~n5038 ) | ( n5019 & 1'b0 ) | ( ~n5038 & 1'b0 ) ;
  assign n5040 = n5030 | n5039 ;
  assign n5041 = ~n4996 & n5004 ;
  assign n5042 = ( n5018 & ~n4353 ) | ( n5018 & n5041 ) | ( ~n4353 & n5041 ) ;
  assign n5043 = ( n4053 & ~n5042 ) | ( n4053 & 1'b0 ) | ( ~n5042 & 1'b0 ) ;
  assign n5044 = n3760 | n5043 ;
  assign n5045 = ( n5040 & ~n5044 ) | ( n5040 & 1'b0 ) | ( ~n5044 & 1'b0 ) ;
  assign n5046 = n5037 | n5045 ;
  assign n5020 = ~n5006 & n5019 ;
  assign n5031 = ( n5020 & ~n4053 ) | ( n5020 & n5030 ) | ( ~n4053 & n5030 ) ;
  assign n5032 = ( n3760 & ~n5031 ) | ( n3760 & 1'b0 ) | ( ~n5031 & 1'b0 ) ;
  assign n5060 = n3482 | n5032 ;
  assign n5061 = ( n5046 & ~n5060 ) | ( n5046 & 1'b0 ) | ( ~n5060 & 1'b0 ) ;
  assign n5062 = n5052 | n5061 ;
  assign n5063 = ( n5040 & ~n5043 ) | ( n5040 & 1'b0 ) | ( ~n5043 & 1'b0 ) ;
  assign n5064 = ( n5037 & ~n3760 ) | ( n5037 & n5063 ) | ( ~n3760 & n5063 ) ;
  assign n5065 = ( n3482 & ~n5064 ) | ( n3482 & 1'b0 ) | ( ~n5064 & 1'b0 ) ;
  assign n5066 = n3211 | n5065 ;
  assign n5067 = ( n5062 & ~n5066 ) | ( n5062 & 1'b0 ) | ( ~n5066 & 1'b0 ) ;
  assign n5068 = n5059 | n5067 ;
  assign n5047 = ~n5032 & n5046 ;
  assign n5053 = ( n5047 & ~n3482 ) | ( n5047 & n5052 ) | ( ~n3482 & n5052 ) ;
  assign n5054 = ( n3211 & ~n5053 ) | ( n3211 & 1'b0 ) | ( ~n5053 & 1'b0 ) ;
  assign n5082 = n2955 | n5054 ;
  assign n5083 = ( n5068 & ~n5082 ) | ( n5068 & 1'b0 ) | ( ~n5082 & 1'b0 ) ;
  assign n5084 = n5074 | n5083 ;
  assign n5085 = ( n5062 & ~n5065 ) | ( n5062 & 1'b0 ) | ( ~n5065 & 1'b0 ) ;
  assign n5086 = ( n5059 & ~n3211 ) | ( n5059 & n5085 ) | ( ~n3211 & n5085 ) ;
  assign n5087 = ( n2955 & ~n5086 ) | ( n2955 & 1'b0 ) | ( ~n5086 & 1'b0 ) ;
  assign n5088 = n2706 | n5087 ;
  assign n5089 = ( n5084 & ~n5088 ) | ( n5084 & 1'b0 ) | ( ~n5088 & 1'b0 ) ;
  assign n5090 = n5081 | n5089 ;
  assign n5069 = ~n5054 & n5068 ;
  assign n5075 = ( n5069 & ~n2955 ) | ( n5069 & n5074 ) | ( ~n2955 & n5074 ) ;
  assign n5076 = ( n2706 & ~n5075 ) | ( n2706 & 1'b0 ) | ( ~n5075 & 1'b0 ) ;
  assign n5104 = n2472 | n5076 ;
  assign n5105 = ( n5090 & ~n5104 ) | ( n5090 & 1'b0 ) | ( ~n5104 & 1'b0 ) ;
  assign n5106 = n5096 | n5105 ;
  assign n5107 = ( n5084 & ~n5087 ) | ( n5084 & 1'b0 ) | ( ~n5087 & 1'b0 ) ;
  assign n5108 = ( n5081 & ~n2706 ) | ( n5081 & n5107 ) | ( ~n2706 & n5107 ) ;
  assign n5109 = ( n2472 & ~n5108 ) | ( n2472 & 1'b0 ) | ( ~n5108 & 1'b0 ) ;
  assign n5110 = n2245 | n5109 ;
  assign n5111 = ( n5106 & ~n5110 ) | ( n5106 & 1'b0 ) | ( ~n5110 & 1'b0 ) ;
  assign n5112 = n5103 | n5111 ;
  assign n5091 = ~n5076 & n5090 ;
  assign n5097 = ( n5091 & ~n2472 ) | ( n5091 & n5096 ) | ( ~n2472 & n5096 ) ;
  assign n5098 = ( n2245 & ~n5097 ) | ( n2245 & 1'b0 ) | ( ~n5097 & 1'b0 ) ;
  assign n5126 = ( n2033 & ~n5098 ) | ( n2033 & 1'b0 ) | ( ~n5098 & 1'b0 ) ;
  assign n5127 = n5112 &  n5126 ;
  assign n5128 = n5118 | n5127 ;
  assign n5129 = ( n5106 & ~n5109 ) | ( n5106 & 1'b0 ) | ( ~n5109 & 1'b0 ) ;
  assign n5130 = ( n5103 & ~n2245 ) | ( n5103 & n5129 ) | ( ~n2245 & n5129 ) ;
  assign n5131 = n2033 | n5130 ;
  assign n5151 = n5128 &  n5131 ;
  assign n5152 = ( n5125 & ~n1827 ) | ( n5125 & n5151 ) | ( ~n1827 & n5151 ) ;
  assign n5153 = n1636 | n5152 ;
  assign n5295 = ( n4956 & ~n4972 ) | ( n4956 & 1'b0 ) | ( ~n4972 & 1'b0 ) ;
  assign n5296 = ( n4975 & n4990 ) | ( n4975 & n5295 ) | ( n4990 & n5295 ) ;
  assign n5297 = ~n4975 & n5296 ;
  assign n5298 = n4972 | n4975 ;
  assign n5299 = n4990 | n5298 ;
  assign n5300 = ( n4956 & ~n5298 ) | ( n4956 & n5299 ) | ( ~n5298 & n5299 ) ;
  assign n5301 = ~n5297 & n5300 ;
  assign n5302 = ~n4957 & n4964 ;
  assign n5303 = ~n4990 & n5302 ;
  assign n5304 = ( n4978 & ~n5303 ) | ( n4978 & n5302 ) | ( ~n5303 & n5302 ) ;
  assign n5305 = n5301 | n5304 ;
  assign n5268 = ~n4928 & n4990 ;
  assign n5269 = ( n4915 & n4920 ) | ( n4915 & n4990 ) | ( n4920 & n4990 ) ;
  assign n5271 = ( n5268 & ~n4915 ) | ( n5268 & n5269 ) | ( ~n4915 & n5269 ) ;
  assign n5270 = ( n4990 & ~n5269 ) | ( n4990 & n5268 ) | ( ~n5269 & n5268 ) ;
  assign n5272 = ( n4920 & ~n5271 ) | ( n4920 & n5270 ) | ( ~n5271 & n5270 ) ;
  assign n5113 = ~n5098 & n5112 ;
  assign n5119 = ( n2033 & n5113 ) | ( n2033 & n5118 ) | ( n5113 & n5118 ) ;
  assign n5120 = ( n1827 & ~n5119 ) | ( n1827 & 1'b0 ) | ( ~n5119 & 1'b0 ) ;
  assign n5132 = ~n1827 & n5131 ;
  assign n5133 = n5128 &  n5132 ;
  assign n5134 = n5125 | n5133 ;
  assign n5135 = ~n5120 & n5134 ;
  assign n5141 = ( n1636 & n5135 ) | ( n1636 & n5140 ) | ( n5135 & n5140 ) ;
  assign n5142 = n1452 | n5141 ;
  assign n5144 = ( n4812 & ~n4803 ) | ( n4812 & n4816 ) | ( ~n4803 & n4816 ) ;
  assign n5143 = ( n4816 & ~n4990 ) | ( n4816 & 1'b0 ) | ( ~n4990 & 1'b0 ) ;
  assign n5146 = ( n4816 & ~n5144 ) | ( n4816 & n5143 ) | ( ~n5144 & n5143 ) ;
  assign n5145 = ( n5143 & ~n4812 ) | ( n5143 & n5144 ) | ( ~n4812 & n5144 ) ;
  assign n5147 = ( n4803 & ~n5146 ) | ( n4803 & n5145 ) | ( ~n5146 & n5145 ) ;
  assign n5148 = ( n1636 & ~n5120 ) | ( n1636 & 1'b0 ) | ( ~n5120 & 1'b0 ) ;
  assign n5149 = n5134 &  n5148 ;
  assign n5150 = n5140 | n5149 ;
  assign n5154 = n1452 &  n5153 ;
  assign n5155 = n5150 &  n5154 ;
  assign n5156 = n5147 | n5155 ;
  assign n5157 = n5142 &  n5156 ;
  assign n5158 = ( n4805 & ~n4990 ) | ( n4805 & 1'b0 ) | ( ~n4990 & 1'b0 ) ;
  assign n5159 = ( n4805 & n4810 ) | ( n4805 & n4818 ) | ( n4810 & n4818 ) ;
  assign n5160 = ( n5158 & ~n4818 ) | ( n5158 & n5159 ) | ( ~n4818 & n5159 ) ;
  assign n5161 = ( n4805 & ~n5159 ) | ( n4805 & n5158 ) | ( ~n5159 & n5158 ) ;
  assign n5162 = ( n4810 & ~n5160 ) | ( n4810 & n5161 ) | ( ~n5160 & n5161 ) ;
  assign n5163 = ( n5157 & ~n1283 ) | ( n5157 & n5162 ) | ( ~n1283 & n5162 ) ;
  assign n5164 = n1122 | n5163 ;
  assign n5165 = n4838 | n4990 ;
  assign n5166 = ( n4825 & ~n4834 ) | ( n4825 & n4838 ) | ( ~n4834 & n4838 ) ;
  assign n5167 = ( n4834 & n5165 ) | ( n4834 & n5166 ) | ( n5165 & n5166 ) ;
  assign n5168 = ( n4838 & ~n5166 ) | ( n4838 & n5165 ) | ( ~n5166 & n5165 ) ;
  assign n5169 = ( n4825 & ~n5167 ) | ( n4825 & n5168 ) | ( ~n5167 & n5168 ) ;
  assign n5170 = ~n1283 & n5142 ;
  assign n5171 = n5156 &  n5170 ;
  assign n5172 = n5162 | n5171 ;
  assign n5173 = n5150 &  n5153 ;
  assign n5174 = ( n1452 & n5147 ) | ( n1452 & n5173 ) | ( n5147 & n5173 ) ;
  assign n5175 = ( n1283 & ~n5174 ) | ( n1283 & 1'b0 ) | ( ~n5174 & 1'b0 ) ;
  assign n5176 = ( n1122 & ~n5175 ) | ( n1122 & 1'b0 ) | ( ~n5175 & 1'b0 ) ;
  assign n5177 = n5172 &  n5176 ;
  assign n5178 = n5169 | n5177 ;
  assign n5179 = n5164 &  n5178 ;
  assign n5181 = ( n4827 & ~n4832 ) | ( n4827 & n4840 ) | ( ~n4832 & n4840 ) ;
  assign n5180 = ( n4827 & ~n4990 ) | ( n4827 & 1'b0 ) | ( ~n4990 & 1'b0 ) ;
  assign n5183 = ( n4827 & ~n5181 ) | ( n4827 & n5180 ) | ( ~n5181 & n5180 ) ;
  assign n5182 = ( n5180 & ~n4840 ) | ( n5180 & n5181 ) | ( ~n4840 & n5181 ) ;
  assign n5184 = ( n4832 & ~n5183 ) | ( n4832 & n5182 ) | ( ~n5183 & n5182 ) ;
  assign n5185 = ( n976 & n5179 ) | ( n976 & n5184 ) | ( n5179 & n5184 ) ;
  assign n5186 = ( n837 & ~n5185 ) | ( n837 & 1'b0 ) | ( ~n5185 & 1'b0 ) ;
  assign n5187 = ( n4860 & ~n4990 ) | ( n4860 & 1'b0 ) | ( ~n4990 & 1'b0 ) ;
  assign n5188 = ( n4847 & n4856 ) | ( n4847 & n4860 ) | ( n4856 & n4860 ) ;
  assign n5189 = ( n5187 & ~n4856 ) | ( n5187 & n5188 ) | ( ~n4856 & n5188 ) ;
  assign n5190 = ( n4860 & ~n5188 ) | ( n4860 & n5187 ) | ( ~n5188 & n5187 ) ;
  assign n5191 = ( n4847 & ~n5189 ) | ( n4847 & n5190 ) | ( ~n5189 & n5190 ) ;
  assign n5192 = n976 &  n5164 ;
  assign n5193 = n5178 &  n5192 ;
  assign n5194 = n5184 | n5193 ;
  assign n5195 = ( n5172 & ~n5175 ) | ( n5172 & 1'b0 ) | ( ~n5175 & 1'b0 ) ;
  assign n5196 = ( n1122 & n5169 ) | ( n1122 & n5195 ) | ( n5169 & n5195 ) ;
  assign n5197 = n976 | n5196 ;
  assign n5198 = ~n837 & n5197 ;
  assign n5199 = n5194 &  n5198 ;
  assign n5200 = n5191 | n5199 ;
  assign n5201 = ~n5186 & n5200 ;
  assign n5203 = ( n4849 & ~n4854 ) | ( n4849 & n4990 ) | ( ~n4854 & n4990 ) ;
  assign n5202 = n4862 &  n4990 ;
  assign n5204 = ( n4990 & ~n5203 ) | ( n4990 & n5202 ) | ( ~n5203 & n5202 ) ;
  assign n5205 = ( n5202 & ~n4849 ) | ( n5202 & n5203 ) | ( ~n4849 & n5203 ) ;
  assign n5206 = ( n4854 & ~n5204 ) | ( n4854 & n5205 ) | ( ~n5204 & n5205 ) ;
  assign n5207 = ( n5201 & ~n713 ) | ( n5201 & n5206 ) | ( ~n713 & n5206 ) ;
  assign n5208 = ( n595 & ~n5207 ) | ( n595 & 1'b0 ) | ( ~n5207 & 1'b0 ) ;
  assign n5209 = n4882 | n4990 ;
  assign n5210 = ( n4869 & ~n4878 ) | ( n4869 & n4882 ) | ( ~n4878 & n4882 ) ;
  assign n5211 = ( n4878 & n5209 ) | ( n4878 & n5210 ) | ( n5209 & n5210 ) ;
  assign n5212 = ( n4882 & ~n5210 ) | ( n4882 & n5209 ) | ( ~n5210 & n5209 ) ;
  assign n5213 = ( n4869 & ~n5211 ) | ( n4869 & n5212 ) | ( ~n5211 & n5212 ) ;
  assign n5214 = n713 | n5186 ;
  assign n5215 = ( n5200 & ~n5214 ) | ( n5200 & 1'b0 ) | ( ~n5214 & 1'b0 ) ;
  assign n5216 = n5206 | n5215 ;
  assign n5217 = n5194 &  n5197 ;
  assign n5218 = ( n5191 & ~n837 ) | ( n5191 & n5217 ) | ( ~n837 & n5217 ) ;
  assign n5219 = ( n713 & ~n5218 ) | ( n713 & 1'b0 ) | ( ~n5218 & 1'b0 ) ;
  assign n5220 = n595 | n5219 ;
  assign n5221 = ( n5216 & ~n5220 ) | ( n5216 & 1'b0 ) | ( ~n5220 & 1'b0 ) ;
  assign n5222 = n5213 | n5221 ;
  assign n5223 = ~n5208 & n5222 ;
  assign n5224 = n4871 | n4990 ;
  assign n5225 = ( n4876 & ~n4871 ) | ( n4876 & n4884 ) | ( ~n4871 & n4884 ) ;
  assign n5227 = ( n4871 & n5224 ) | ( n4871 & n5225 ) | ( n5224 & n5225 ) ;
  assign n5226 = ( n4884 & ~n5225 ) | ( n4884 & n5224 ) | ( ~n5225 & n5224 ) ;
  assign n5228 = ( n4876 & ~n5227 ) | ( n4876 & n5226 ) | ( ~n5227 & n5226 ) ;
  assign n5229 = ( n5223 & ~n492 ) | ( n5223 & n5228 ) | ( ~n492 & n5228 ) ;
  assign n5230 = ( n396 & ~n5229 ) | ( n396 & 1'b0 ) | ( ~n5229 & 1'b0 ) ;
  assign n5231 = n4904 | n4990 ;
  assign n5232 = ( n4891 & ~n4900 ) | ( n4891 & n4904 ) | ( ~n4900 & n4904 ) ;
  assign n5233 = ( n4900 & n5231 ) | ( n4900 & n5232 ) | ( n5231 & n5232 ) ;
  assign n5234 = ( n4904 & ~n5232 ) | ( n4904 & n5231 ) | ( ~n5232 & n5231 ) ;
  assign n5235 = ( n4891 & ~n5233 ) | ( n4891 & n5234 ) | ( ~n5233 & n5234 ) ;
  assign n5236 = n492 | n5208 ;
  assign n5237 = ( n5222 & ~n5236 ) | ( n5222 & 1'b0 ) | ( ~n5236 & 1'b0 ) ;
  assign n5238 = n5228 | n5237 ;
  assign n5239 = ( n5216 & ~n5219 ) | ( n5216 & 1'b0 ) | ( ~n5219 & 1'b0 ) ;
  assign n5240 = ( n5213 & ~n595 ) | ( n5213 & n5239 ) | ( ~n595 & n5239 ) ;
  assign n5241 = ( n492 & ~n5240 ) | ( n492 & 1'b0 ) | ( ~n5240 & 1'b0 ) ;
  assign n5242 = n396 | n5241 ;
  assign n5243 = ( n5238 & ~n5242 ) | ( n5238 & 1'b0 ) | ( ~n5242 & 1'b0 ) ;
  assign n5244 = n5235 | n5243 ;
  assign n5245 = ~n5230 & n5244 ;
  assign n5246 = n4893 | n4990 ;
  assign n5247 = ( n4898 & ~n4893 ) | ( n4898 & n4906 ) | ( ~n4893 & n4906 ) ;
  assign n5249 = ( n4893 & n5246 ) | ( n4893 & n5247 ) | ( n5246 & n5247 ) ;
  assign n5248 = ( n4906 & ~n5247 ) | ( n4906 & n5246 ) | ( ~n5247 & n5246 ) ;
  assign n5250 = ( n4898 & ~n5249 ) | ( n4898 & n5248 ) | ( ~n5249 & n5248 ) ;
  assign n5251 = ( n315 & ~n5245 ) | ( n315 & n5250 ) | ( ~n5245 & n5250 ) ;
  assign n5252 = n240 &  n5251 ;
  assign n5253 = n4926 | n4990 ;
  assign n5254 = ( n4913 & n4922 ) | ( n4913 & n4926 ) | ( n4922 & n4926 ) ;
  assign n5255 = ( n5253 & ~n4922 ) | ( n5253 & n5254 ) | ( ~n4922 & n5254 ) ;
  assign n5256 = ( n4926 & ~n5254 ) | ( n4926 & n5253 ) | ( ~n5254 & n5253 ) ;
  assign n5257 = ( n4913 & ~n5255 ) | ( n4913 & n5256 ) | ( ~n5255 & n5256 ) ;
  assign n5258 = n315 | n5230 ;
  assign n5259 = ( n5244 & ~n5258 ) | ( n5244 & 1'b0 ) | ( ~n5258 & 1'b0 ) ;
  assign n5260 = ( n5250 & ~n5259 ) | ( n5250 & 1'b0 ) | ( ~n5259 & 1'b0 ) ;
  assign n5261 = ( n5238 & ~n5241 ) | ( n5238 & 1'b0 ) | ( ~n5241 & 1'b0 ) ;
  assign n5262 = ( n5235 & ~n396 ) | ( n5235 & n5261 ) | ( ~n396 & n5261 ) ;
  assign n5263 = ( n315 & ~n5262 ) | ( n315 & 1'b0 ) | ( ~n5262 & 1'b0 ) ;
  assign n5264 = n240 | n5263 ;
  assign n5265 = n5260 | n5264 ;
  assign n5266 = n5257 &  n5265 ;
  assign n5267 = n5252 | n5266 ;
  assign n5273 = ( n181 & ~n5272 ) | ( n181 & n5267 ) | ( ~n5272 & n5267 ) ;
  assign n5274 = ~n145 & n5273 ;
  assign n5275 = n4943 | n4990 ;
  assign n5276 = ( n4935 & n4939 ) | ( n4935 & n4943 ) | ( n4939 & n4943 ) ;
  assign n5277 = ( n5275 & ~n4939 ) | ( n5275 & n5276 ) | ( ~n4939 & n5276 ) ;
  assign n5278 = ( n4943 & ~n5276 ) | ( n4943 & n5275 ) | ( ~n5276 & n5275 ) ;
  assign n5279 = ( n4935 & ~n5277 ) | ( n4935 & n5278 ) | ( ~n5277 & n5278 ) ;
  assign n5280 = n181 | n5252 ;
  assign n5281 = n5266 | n5280 ;
  assign n5282 = ~n5272 & n5281 ;
  assign n5283 = n5260 | n5263 ;
  assign n5284 = ( n240 & n5257 ) | ( n240 & n5283 ) | ( n5257 & n5283 ) ;
  assign n5285 = n181 &  n5284 ;
  assign n5286 = ( n145 & ~n5285 ) | ( n145 & 1'b0 ) | ( ~n5285 & 1'b0 ) ;
  assign n5287 = ~n5282 & n5286 ;
  assign n5288 = n5279 | n5287 ;
  assign n5289 = ~n5274 & n5288 ;
  assign n5290 = ( n4937 & ~n4945 ) | ( n4937 & n4949 ) | ( ~n4945 & n4949 ) ;
  assign n5291 = ( n4945 & n4990 ) | ( n4945 & n5290 ) | ( n4990 & n5290 ) ;
  assign n5292 = ( n4937 & ~n5290 ) | ( n4937 & n4990 ) | ( ~n5290 & n4990 ) ;
  assign n5293 = ( n4949 & ~n5291 ) | ( n4949 & n5292 ) | ( ~n5291 & n5292 ) ;
  assign n5294 = ( n5289 & ~n150 ) | ( n5289 & n5293 ) | ( ~n150 & n5293 ) ;
  assign n5306 = ~n5305 & n5294 ;
  assign n5307 = ( n5306 & ~n133 ) | ( n5306 & n5305 ) | ( ~n133 & n5305 ) ;
  assign n5308 = n150 | n5274 ;
  assign n5309 = ( n5288 & ~n5308 ) | ( n5288 & 1'b0 ) | ( ~n5308 & 1'b0 ) ;
  assign n5314 = ~n5293 & n5309 ;
  assign n5310 = n5282 | n5285 ;
  assign n5311 = ( n145 & ~n5310 ) | ( n145 & n5279 ) | ( ~n5310 & n5279 ) ;
  assign n5312 = ( n150 & ~n5311 ) | ( n150 & 1'b0 ) | ( ~n5311 & 1'b0 ) ;
  assign n5313 = ( n5301 & ~n5312 ) | ( n5301 & 1'b0 ) | ( ~n5312 & 1'b0 ) ;
  assign n5315 = ( n5293 & n5314 ) | ( n5293 & n5313 ) | ( n5314 & n5313 ) ;
  assign n5317 = ( n133 & ~n4957 ) | ( n133 & n4964 ) | ( ~n4957 & n4964 ) ;
  assign n5316 = ( n4957 & ~n4964 ) | ( n4957 & n4990 ) | ( ~n4964 & n4990 ) ;
  assign n5318 = n4964 &  n5316 ;
  assign n5319 = ( n5317 & ~n4964 ) | ( n5317 & n5318 ) | ( ~n4964 & n5318 ) ;
  assign n5320 = n4960 | n4987 ;
  assign n5321 = ( n4982 & ~n4963 ) | ( n4982 & n5320 ) | ( ~n4963 & n5320 ) ;
  assign n5322 = n4963 | n5321 ;
  assign n5323 = ( n4970 & n4978 ) | ( n4970 & n5322 ) | ( n4978 & n5322 ) ;
  assign n5324 = ( n4970 & ~n5323 ) | ( n4970 & 1'b0 ) | ( ~n5323 & 1'b0 ) ;
  assign n5325 = n5319 | n5324 ;
  assign n5326 = n5315 | n5325 ;
  assign n5327 = n5307 | n5326 ;
  assign n5487 = ( n5153 & ~n5327 ) | ( n5153 & 1'b0 ) | ( ~n5327 & 1'b0 ) ;
  assign n5488 = ( n5140 & n5149 ) | ( n5140 & n5153 ) | ( n5149 & n5153 ) ;
  assign n5489 = ( n5487 & ~n5149 ) | ( n5487 & n5488 ) | ( ~n5149 & n5488 ) ;
  assign n5490 = ( n5153 & ~n5488 ) | ( n5153 & n5487 ) | ( ~n5488 & n5487 ) ;
  assign n5491 = ( n5140 & ~n5489 ) | ( n5140 & n5490 ) | ( ~n5489 & n5490 ) ;
  assign n5480 = n5120 | n5327 ;
  assign n5481 = ( n5120 & ~n5133 ) | ( n5120 & n5125 ) | ( ~n5133 & n5125 ) ;
  assign n5482 = ( n5133 & n5480 ) | ( n5133 & n5481 ) | ( n5480 & n5481 ) ;
  assign n5483 = ( n5120 & ~n5481 ) | ( n5120 & n5480 ) | ( ~n5481 & n5480 ) ;
  assign n5484 = ( n5125 & ~n5482 ) | ( n5125 & n5483 ) | ( ~n5482 & n5483 ) ;
  assign n5466 = ( n5127 & ~n5118 ) | ( n5127 & n5131 ) | ( ~n5118 & n5131 ) ;
  assign n5465 = ( n5131 & ~n5327 ) | ( n5131 & 1'b0 ) | ( ~n5327 & 1'b0 ) ;
  assign n5468 = ( n5131 & ~n5466 ) | ( n5131 & n5465 ) | ( ~n5466 & n5465 ) ;
  assign n5467 = ( n5465 & ~n5127 ) | ( n5465 & n5466 ) | ( ~n5127 & n5466 ) ;
  assign n5469 = ( n5118 & ~n5468 ) | ( n5118 & n5467 ) | ( ~n5468 & n5467 ) ;
  assign n5458 = n5098 | n5327 ;
  assign n5459 = ( n5103 & ~n5098 ) | ( n5103 & n5111 ) | ( ~n5098 & n5111 ) ;
  assign n5461 = ( n5098 & n5458 ) | ( n5098 & n5459 ) | ( n5458 & n5459 ) ;
  assign n5460 = ( n5111 & ~n5459 ) | ( n5111 & n5458 ) | ( ~n5459 & n5458 ) ;
  assign n5462 = ( n5103 & ~n5461 ) | ( n5103 & n5460 ) | ( ~n5461 & n5460 ) ;
  assign n5443 = n5109 | n5327 ;
  assign n5444 = ( n5096 & ~n5105 ) | ( n5096 & n5109 ) | ( ~n5105 & n5109 ) ;
  assign n5445 = ( n5105 & n5443 ) | ( n5105 & n5444 ) | ( n5443 & n5444 ) ;
  assign n5446 = ( n5109 & ~n5444 ) | ( n5109 & n5443 ) | ( ~n5444 & n5443 ) ;
  assign n5447 = ( n5096 & ~n5445 ) | ( n5096 & n5446 ) | ( ~n5445 & n5446 ) ;
  assign n5437 = ( n5076 & ~n5081 ) | ( n5076 & n5327 ) | ( ~n5081 & n5327 ) ;
  assign n5436 = n5089 &  n5327 ;
  assign n5438 = ( n5327 & ~n5437 ) | ( n5327 & n5436 ) | ( ~n5437 & n5436 ) ;
  assign n5439 = ( n5436 & ~n5076 ) | ( n5436 & n5437 ) | ( ~n5076 & n5437 ) ;
  assign n5440 = ( n5081 & ~n5438 ) | ( n5081 & n5439 ) | ( ~n5438 & n5439 ) ;
  assign n5421 = n5087 | n5327 ;
  assign n5422 = ( n5074 & ~n5087 ) | ( n5074 & n5083 ) | ( ~n5087 & n5083 ) ;
  assign n5424 = ( n5087 & n5421 ) | ( n5087 & n5422 ) | ( n5421 & n5422 ) ;
  assign n5423 = ( n5083 & ~n5422 ) | ( n5083 & n5421 ) | ( ~n5422 & n5421 ) ;
  assign n5425 = ( n5074 & ~n5424 ) | ( n5074 & n5423 ) | ( ~n5424 & n5423 ) ;
  assign n5414 = n5054 | n5327 ;
  assign n5415 = ( n5054 & ~n5067 ) | ( n5054 & n5059 ) | ( ~n5067 & n5059 ) ;
  assign n5416 = ( n5067 & n5414 ) | ( n5067 & n5415 ) | ( n5414 & n5415 ) ;
  assign n5417 = ( n5054 & ~n5415 ) | ( n5054 & n5414 ) | ( ~n5415 & n5414 ) ;
  assign n5418 = ( n5059 & ~n5416 ) | ( n5059 & n5417 ) | ( ~n5416 & n5417 ) ;
  assign n5399 = n5065 | n5327 ;
  assign n5400 = ( n5052 & ~n5061 ) | ( n5052 & n5065 ) | ( ~n5061 & n5065 ) ;
  assign n5401 = ( n5061 & n5399 ) | ( n5061 & n5400 ) | ( n5399 & n5400 ) ;
  assign n5402 = ( n5065 & ~n5400 ) | ( n5065 & n5399 ) | ( ~n5400 & n5399 ) ;
  assign n5403 = ( n5052 & ~n5401 ) | ( n5052 & n5402 ) | ( ~n5401 & n5402 ) ;
  assign n5392 = n5032 | n5327 ;
  assign n5393 = ( n5037 & ~n5032 ) | ( n5037 & n5045 ) | ( ~n5032 & n5045 ) ;
  assign n5395 = ( n5032 & n5392 ) | ( n5032 & n5393 ) | ( n5392 & n5393 ) ;
  assign n5394 = ( n5045 & ~n5393 ) | ( n5045 & n5392 ) | ( ~n5393 & n5392 ) ;
  assign n5396 = ( n5037 & ~n5395 ) | ( n5037 & n5394 ) | ( ~n5395 & n5394 ) ;
  assign n5377 = n5043 | n5327 ;
  assign n5378 = ( n5030 & ~n5039 ) | ( n5030 & n5043 ) | ( ~n5039 & n5043 ) ;
  assign n5379 = ( n5039 & n5377 ) | ( n5039 & n5378 ) | ( n5377 & n5378 ) ;
  assign n5380 = ( n5043 & ~n5378 ) | ( n5043 & n5377 ) | ( ~n5378 & n5377 ) ;
  assign n5381 = ( n5030 & ~n5379 ) | ( n5030 & n5380 ) | ( ~n5379 & n5380 ) ;
  assign n5370 = ( n5006 & ~n5008 ) | ( n5006 & 1'b0 ) | ( ~n5008 & 1'b0 ) ;
  assign n5371 = ( n5008 & ~n5370 ) | ( n5008 & n5018 ) | ( ~n5370 & n5018 ) ;
  assign n5373 = ( n5327 & n5370 ) | ( n5327 & n5371 ) | ( n5370 & n5371 ) ;
  assign n5372 = ( n5008 & ~n5371 ) | ( n5008 & n5327 ) | ( ~n5371 & n5327 ) ;
  assign n5374 = ( n5018 & ~n5373 ) | ( n5018 & n5372 ) | ( ~n5373 & n5372 ) ;
  assign n5354 = ~x70 & n4990 ;
  assign n5355 = ( x71 & ~n5354 ) | ( x71 & 1'b0 ) | ( ~n5354 & 1'b0 ) ;
  assign n5356 = n5009 | n5355 ;
  assign n5351 = ( n4990 & ~x70 ) | ( n4990 & n5001 ) | ( ~x70 & n5001 ) ;
  assign n5352 = x70 &  n5351 ;
  assign n5353 = ( n4996 & ~n5352 ) | ( n4996 & n5001 ) | ( ~n5352 & n5001 ) ;
  assign n5357 = ( n5327 & ~n5356 ) | ( n5327 & n5353 ) | ( ~n5356 & n5353 ) ;
  assign n5359 = ( n5327 & ~n5357 ) | ( n5327 & 1'b0 ) | ( ~n5357 & 1'b0 ) ;
  assign n5358 = ~n5353 & n5357 ;
  assign n5360 = ( n5356 & ~n5359 ) | ( n5356 & n5358 ) | ( ~n5359 & n5358 ) ;
  assign n5340 = ( n4990 & ~n5324 ) | ( n4990 & 1'b0 ) | ( ~n5324 & 1'b0 ) ;
  assign n5341 = ( n5315 & ~n5319 ) | ( n5315 & n5340 ) | ( ~n5319 & n5340 ) ;
  assign n5342 = ~n5315 & n5341 ;
  assign n5343 = ~n5307 & n5342 ;
  assign n5339 = ~n4993 & n5327 ;
  assign n5344 = ~n5343 & n5339 ;
  assign n5345 = ( x70 & n5344 ) | ( x70 & n5343 ) | ( n5344 & n5343 ) ;
  assign n5346 = x70 | n5343 ;
  assign n5347 = n5339 | n5346 ;
  assign n5348 = ~n5345 & n5347 ;
  assign n5330 = ( x68 & ~n5327 ) | ( x68 & x69 ) | ( ~n5327 & x69 ) ;
  assign n5336 = ( x68 & ~x69 ) | ( x68 & 1'b0 ) | ( ~x69 & 1'b0 ) ;
  assign n4991 = x66 | x67 ;
  assign n5331 = ~x68 & n4991 ;
  assign n5332 = ( x68 & ~n4988 ) | ( x68 & n5331 ) | ( ~n4988 & n5331 ) ;
  assign n5333 = ( n4970 & ~n5332 ) | ( n4970 & n4978 ) | ( ~n5332 & n4978 ) ;
  assign n5334 = ( n4970 & ~n5333 ) | ( n4970 & 1'b0 ) | ( ~n5333 & 1'b0 ) ;
  assign n5335 = ( n5327 & ~x69 ) | ( n5327 & n5334 ) | ( ~x69 & n5334 ) ;
  assign n5337 = ( n5330 & ~n5336 ) | ( n5330 & n5335 ) | ( ~n5336 & n5335 ) ;
  assign n4992 = x68 | n4991 ;
  assign n5328 = x68 &  n5327 ;
  assign n5329 = ( n4990 & ~n4992 ) | ( n4990 & n5328 ) | ( ~n4992 & n5328 ) ;
  assign n5361 = n4668 | n5329 ;
  assign n5362 = ( n5337 & ~n5361 ) | ( n5337 & 1'b0 ) | ( ~n5361 & 1'b0 ) ;
  assign n5363 = n5348 | n5362 ;
  assign n5364 = n5329 &  n5337 ;
  assign n5365 = ( n4668 & ~n5337 ) | ( n4668 & n5364 ) | ( ~n5337 & n5364 ) ;
  assign n5366 = n4353 | n5365 ;
  assign n5367 = ( n5363 & ~n5366 ) | ( n5363 & 1'b0 ) | ( ~n5366 & 1'b0 ) ;
  assign n5368 = n5360 | n5367 ;
  assign n5338 = ~n5329 & n5337 ;
  assign n5349 = ( n5338 & ~n4668 ) | ( n5338 & n5348 ) | ( ~n4668 & n5348 ) ;
  assign n5350 = ( n4353 & ~n5349 ) | ( n4353 & 1'b0 ) | ( ~n5349 & 1'b0 ) ;
  assign n5382 = n4053 | n5350 ;
  assign n5383 = ( n5368 & ~n5382 ) | ( n5368 & 1'b0 ) | ( ~n5382 & 1'b0 ) ;
  assign n5384 = n5374 | n5383 ;
  assign n5385 = ( n5363 & ~n5365 ) | ( n5363 & 1'b0 ) | ( ~n5365 & 1'b0 ) ;
  assign n5386 = ( n5360 & ~n4353 ) | ( n5360 & n5385 ) | ( ~n4353 & n5385 ) ;
  assign n5387 = ( n4053 & ~n5386 ) | ( n4053 & 1'b0 ) | ( ~n5386 & 1'b0 ) ;
  assign n5388 = n3760 | n5387 ;
  assign n5389 = ( n5384 & ~n5388 ) | ( n5384 & 1'b0 ) | ( ~n5388 & 1'b0 ) ;
  assign n5390 = n5381 | n5389 ;
  assign n5369 = ~n5350 & n5368 ;
  assign n5375 = ( n5369 & ~n4053 ) | ( n5369 & n5374 ) | ( ~n4053 & n5374 ) ;
  assign n5376 = ( n3760 & ~n5375 ) | ( n3760 & 1'b0 ) | ( ~n5375 & 1'b0 ) ;
  assign n5404 = n3482 | n5376 ;
  assign n5405 = ( n5390 & ~n5404 ) | ( n5390 & 1'b0 ) | ( ~n5404 & 1'b0 ) ;
  assign n5406 = n5396 | n5405 ;
  assign n5407 = ( n5384 & ~n5387 ) | ( n5384 & 1'b0 ) | ( ~n5387 & 1'b0 ) ;
  assign n5408 = ( n5381 & ~n3760 ) | ( n5381 & n5407 ) | ( ~n3760 & n5407 ) ;
  assign n5409 = ( n3482 & ~n5408 ) | ( n3482 & 1'b0 ) | ( ~n5408 & 1'b0 ) ;
  assign n5410 = n3211 | n5409 ;
  assign n5411 = ( n5406 & ~n5410 ) | ( n5406 & 1'b0 ) | ( ~n5410 & 1'b0 ) ;
  assign n5412 = n5403 | n5411 ;
  assign n5391 = ~n5376 & n5390 ;
  assign n5397 = ( n5391 & ~n3482 ) | ( n5391 & n5396 ) | ( ~n3482 & n5396 ) ;
  assign n5398 = ( n3211 & ~n5397 ) | ( n3211 & 1'b0 ) | ( ~n5397 & 1'b0 ) ;
  assign n5426 = n2955 | n5398 ;
  assign n5427 = ( n5412 & ~n5426 ) | ( n5412 & 1'b0 ) | ( ~n5426 & 1'b0 ) ;
  assign n5428 = n5418 | n5427 ;
  assign n5429 = ( n5406 & ~n5409 ) | ( n5406 & 1'b0 ) | ( ~n5409 & 1'b0 ) ;
  assign n5430 = ( n5403 & ~n3211 ) | ( n5403 & n5429 ) | ( ~n3211 & n5429 ) ;
  assign n5431 = ( n2955 & ~n5430 ) | ( n2955 & 1'b0 ) | ( ~n5430 & 1'b0 ) ;
  assign n5432 = n2706 | n5431 ;
  assign n5433 = ( n5428 & ~n5432 ) | ( n5428 & 1'b0 ) | ( ~n5432 & 1'b0 ) ;
  assign n5434 = n5425 | n5433 ;
  assign n5413 = ~n5398 & n5412 ;
  assign n5419 = ( n5413 & ~n2955 ) | ( n5413 & n5418 ) | ( ~n2955 & n5418 ) ;
  assign n5420 = ( n2706 & ~n5419 ) | ( n2706 & 1'b0 ) | ( ~n5419 & 1'b0 ) ;
  assign n5448 = n2472 | n5420 ;
  assign n5449 = ( n5434 & ~n5448 ) | ( n5434 & 1'b0 ) | ( ~n5448 & 1'b0 ) ;
  assign n5450 = n5440 | n5449 ;
  assign n5451 = ( n5428 & ~n5431 ) | ( n5428 & 1'b0 ) | ( ~n5431 & 1'b0 ) ;
  assign n5452 = ( n5425 & ~n2706 ) | ( n5425 & n5451 ) | ( ~n2706 & n5451 ) ;
  assign n5453 = ( n2472 & ~n5452 ) | ( n2472 & 1'b0 ) | ( ~n5452 & 1'b0 ) ;
  assign n5454 = n2245 | n5453 ;
  assign n5455 = ( n5450 & ~n5454 ) | ( n5450 & 1'b0 ) | ( ~n5454 & 1'b0 ) ;
  assign n5456 = n5447 | n5455 ;
  assign n5435 = ~n5420 & n5434 ;
  assign n5441 = ( n5435 & ~n2472 ) | ( n5435 & n5440 ) | ( ~n2472 & n5440 ) ;
  assign n5442 = ( n2245 & ~n5441 ) | ( n2245 & 1'b0 ) | ( ~n5441 & 1'b0 ) ;
  assign n5470 = ( n2033 & ~n5442 ) | ( n2033 & 1'b0 ) | ( ~n5442 & 1'b0 ) ;
  assign n5471 = n5456 &  n5470 ;
  assign n5472 = n5462 | n5471 ;
  assign n5473 = ( n5450 & ~n5453 ) | ( n5450 & 1'b0 ) | ( ~n5453 & 1'b0 ) ;
  assign n5474 = ( n5447 & ~n2245 ) | ( n5447 & n5473 ) | ( ~n2245 & n5473 ) ;
  assign n5475 = n2033 | n5474 ;
  assign n5476 = ~n1827 & n5475 ;
  assign n5477 = n5472 &  n5476 ;
  assign n5478 = n5469 | n5477 ;
  assign n5457 = ~n5442 & n5456 ;
  assign n5463 = ( n2033 & n5457 ) | ( n2033 & n5462 ) | ( n5457 & n5462 ) ;
  assign n5464 = ( n1827 & ~n5463 ) | ( n1827 & 1'b0 ) | ( ~n5463 & 1'b0 ) ;
  assign n5492 = ( n1636 & ~n5464 ) | ( n1636 & 1'b0 ) | ( ~n5464 & 1'b0 ) ;
  assign n5493 = n5478 &  n5492 ;
  assign n5494 = n5484 | n5493 ;
  assign n5495 = n5472 &  n5475 ;
  assign n5496 = ( n5469 & ~n1827 ) | ( n5469 & n5495 ) | ( ~n1827 & n5495 ) ;
  assign n5497 = n1636 | n5496 ;
  assign n5517 = n5494 &  n5497 ;
  assign n5518 = ( n1452 & n5491 ) | ( n1452 & n5517 ) | ( n5491 & n5517 ) ;
  assign n5519 = ( n1283 & ~n5518 ) | ( n1283 & 1'b0 ) | ( ~n5518 & 1'b0 ) ;
  assign n5640 = ( n5293 & ~n5312 ) | ( n5293 & 1'b0 ) | ( ~n5312 & 1'b0 ) ;
  assign n5641 = ( n5309 & n5327 ) | ( n5309 & n5640 ) | ( n5327 & n5640 ) ;
  assign n5642 = ~n5309 & n5641 ;
  assign n5643 = n5309 | n5312 ;
  assign n5644 = n5327 | n5643 ;
  assign n5645 = ( n5293 & ~n5643 ) | ( n5293 & n5644 ) | ( ~n5643 & n5644 ) ;
  assign n5646 = ~n5642 & n5645 ;
  assign n5647 = n5294 | n5301 ;
  assign n5648 = n5327 | n5647 ;
  assign n5649 = ( n5315 & ~n5647 ) | ( n5315 & n5648 ) | ( ~n5647 & n5648 ) ;
  assign n5650 = n5646 | n5649 ;
  assign n5479 = ~n5464 & n5478 ;
  assign n5485 = ( n1636 & n5479 ) | ( n1636 & n5484 ) | ( n5479 & n5484 ) ;
  assign n5486 = n1452 | n5485 ;
  assign n5498 = n1452 &  n5497 ;
  assign n5499 = n5494 &  n5498 ;
  assign n5500 = n5491 | n5499 ;
  assign n5501 = n5486 &  n5500 ;
  assign n5502 = n5155 &  n5327 ;
  assign n5503 = ( n5142 & ~n5327 ) | ( n5142 & n5147 ) | ( ~n5327 & n5147 ) ;
  assign n5504 = ( n5327 & n5502 ) | ( n5327 & n5503 ) | ( n5502 & n5503 ) ;
  assign n5505 = ( n5142 & ~n5503 ) | ( n5142 & n5502 ) | ( ~n5503 & n5502 ) ;
  assign n5506 = ( n5147 & ~n5504 ) | ( n5147 & n5505 ) | ( ~n5504 & n5505 ) ;
  assign n5507 = ( n5501 & ~n1283 ) | ( n5501 & n5506 ) | ( ~n1283 & n5506 ) ;
  assign n5508 = n1122 | n5507 ;
  assign n5509 = n5175 | n5327 ;
  assign n5510 = ( n5162 & ~n5171 ) | ( n5162 & n5175 ) | ( ~n5171 & n5175 ) ;
  assign n5511 = ( n5171 & n5509 ) | ( n5171 & n5510 ) | ( n5509 & n5510 ) ;
  assign n5512 = ( n5175 & ~n5510 ) | ( n5175 & n5509 ) | ( ~n5510 & n5509 ) ;
  assign n5513 = ( n5162 & ~n5511 ) | ( n5162 & n5512 ) | ( ~n5511 & n5512 ) ;
  assign n5514 = ~n1283 & n5486 ;
  assign n5515 = n5500 &  n5514 ;
  assign n5516 = n5506 | n5515 ;
  assign n5520 = ( n1122 & ~n5519 ) | ( n1122 & 1'b0 ) | ( ~n5519 & 1'b0 ) ;
  assign n5521 = n5516 &  n5520 ;
  assign n5522 = n5513 | n5521 ;
  assign n5523 = n5508 &  n5522 ;
  assign n5524 = ( n5164 & ~n5327 ) | ( n5164 & 1'b0 ) | ( ~n5327 & 1'b0 ) ;
  assign n5525 = ( n5164 & n5169 ) | ( n5164 & n5177 ) | ( n5169 & n5177 ) ;
  assign n5526 = ( n5524 & ~n5177 ) | ( n5524 & n5525 ) | ( ~n5177 & n5525 ) ;
  assign n5527 = ( n5164 & ~n5525 ) | ( n5164 & n5524 ) | ( ~n5525 & n5524 ) ;
  assign n5528 = ( n5169 & ~n5526 ) | ( n5169 & n5527 ) | ( ~n5526 & n5527 ) ;
  assign n5529 = ( n976 & n5523 ) | ( n976 & n5528 ) | ( n5523 & n5528 ) ;
  assign n5530 = ( n837 & ~n5529 ) | ( n837 & 1'b0 ) | ( ~n5529 & 1'b0 ) ;
  assign n5532 = ( n5193 & ~n5184 ) | ( n5193 & n5197 ) | ( ~n5184 & n5197 ) ;
  assign n5531 = ( n5197 & ~n5327 ) | ( n5197 & 1'b0 ) | ( ~n5327 & 1'b0 ) ;
  assign n5534 = ( n5197 & ~n5532 ) | ( n5197 & n5531 ) | ( ~n5532 & n5531 ) ;
  assign n5533 = ( n5531 & ~n5193 ) | ( n5531 & n5532 ) | ( ~n5193 & n5532 ) ;
  assign n5535 = ( n5184 & ~n5534 ) | ( n5184 & n5533 ) | ( ~n5534 & n5533 ) ;
  assign n5536 = n976 &  n5508 ;
  assign n5537 = n5522 &  n5536 ;
  assign n5538 = n5528 | n5537 ;
  assign n5539 = ( n5516 & ~n5519 ) | ( n5516 & 1'b0 ) | ( ~n5519 & 1'b0 ) ;
  assign n5540 = ( n1122 & n5513 ) | ( n1122 & n5539 ) | ( n5513 & n5539 ) ;
  assign n5541 = n976 | n5540 ;
  assign n5542 = ~n837 & n5541 ;
  assign n5543 = n5538 &  n5542 ;
  assign n5544 = n5535 | n5543 ;
  assign n5545 = ~n5530 & n5544 ;
  assign n5546 = n5186 | n5327 ;
  assign n5547 = ( n5186 & ~n5199 ) | ( n5186 & n5191 ) | ( ~n5199 & n5191 ) ;
  assign n5548 = ( n5199 & n5546 ) | ( n5199 & n5547 ) | ( n5546 & n5547 ) ;
  assign n5549 = ( n5186 & ~n5547 ) | ( n5186 & n5546 ) | ( ~n5547 & n5546 ) ;
  assign n5550 = ( n5191 & ~n5548 ) | ( n5191 & n5549 ) | ( ~n5548 & n5549 ) ;
  assign n5551 = ( n5545 & ~n713 ) | ( n5545 & n5550 ) | ( ~n713 & n5550 ) ;
  assign n5552 = ( n595 & ~n5551 ) | ( n595 & 1'b0 ) | ( ~n5551 & 1'b0 ) ;
  assign n5553 = n5219 | n5327 ;
  assign n5554 = ( n5206 & ~n5219 ) | ( n5206 & n5215 ) | ( ~n5219 & n5215 ) ;
  assign n5556 = ( n5219 & n5553 ) | ( n5219 & n5554 ) | ( n5553 & n5554 ) ;
  assign n5555 = ( n5215 & ~n5554 ) | ( n5215 & n5553 ) | ( ~n5554 & n5553 ) ;
  assign n5557 = ( n5206 & ~n5556 ) | ( n5206 & n5555 ) | ( ~n5556 & n5555 ) ;
  assign n5558 = n713 | n5530 ;
  assign n5559 = ( n5544 & ~n5558 ) | ( n5544 & 1'b0 ) | ( ~n5558 & 1'b0 ) ;
  assign n5560 = n5550 | n5559 ;
  assign n5561 = n5538 &  n5541 ;
  assign n5562 = ( n5535 & ~n837 ) | ( n5535 & n5561 ) | ( ~n837 & n5561 ) ;
  assign n5563 = ( n713 & ~n5562 ) | ( n713 & 1'b0 ) | ( ~n5562 & 1'b0 ) ;
  assign n5564 = n595 | n5563 ;
  assign n5565 = ( n5560 & ~n5564 ) | ( n5560 & 1'b0 ) | ( ~n5564 & 1'b0 ) ;
  assign n5566 = n5557 | n5565 ;
  assign n5567 = ~n5552 & n5566 ;
  assign n5569 = ( n5208 & ~n5213 ) | ( n5208 & n5327 ) | ( ~n5213 & n5327 ) ;
  assign n5568 = n5221 &  n5327 ;
  assign n5570 = ( n5327 & ~n5569 ) | ( n5327 & n5568 ) | ( ~n5569 & n5568 ) ;
  assign n5571 = ( n5568 & ~n5208 ) | ( n5568 & n5569 ) | ( ~n5208 & n5569 ) ;
  assign n5572 = ( n5213 & ~n5570 ) | ( n5213 & n5571 ) | ( ~n5570 & n5571 ) ;
  assign n5573 = ( n5567 & ~n492 ) | ( n5567 & n5572 ) | ( ~n492 & n5572 ) ;
  assign n5574 = ( n396 & ~n5573 ) | ( n396 & 1'b0 ) | ( ~n5573 & 1'b0 ) ;
  assign n5575 = n5241 | n5327 ;
  assign n5576 = ( n5228 & ~n5237 ) | ( n5228 & n5241 ) | ( ~n5237 & n5241 ) ;
  assign n5577 = ( n5237 & n5575 ) | ( n5237 & n5576 ) | ( n5575 & n5576 ) ;
  assign n5578 = ( n5241 & ~n5576 ) | ( n5241 & n5575 ) | ( ~n5576 & n5575 ) ;
  assign n5579 = ( n5228 & ~n5577 ) | ( n5228 & n5578 ) | ( ~n5577 & n5578 ) ;
  assign n5580 = n492 | n5552 ;
  assign n5581 = ( n5566 & ~n5580 ) | ( n5566 & 1'b0 ) | ( ~n5580 & 1'b0 ) ;
  assign n5582 = n5572 | n5581 ;
  assign n5583 = ( n5560 & ~n5563 ) | ( n5560 & 1'b0 ) | ( ~n5563 & 1'b0 ) ;
  assign n5584 = ( n5557 & ~n595 ) | ( n5557 & n5583 ) | ( ~n595 & n5583 ) ;
  assign n5585 = ( n492 & ~n5584 ) | ( n492 & 1'b0 ) | ( ~n5584 & 1'b0 ) ;
  assign n5586 = n396 | n5585 ;
  assign n5587 = ( n5582 & ~n5586 ) | ( n5582 & 1'b0 ) | ( ~n5586 & 1'b0 ) ;
  assign n5588 = n5579 | n5587 ;
  assign n5589 = ~n5574 & n5588 ;
  assign n5590 = n5230 | n5327 ;
  assign n5591 = ( n5235 & ~n5230 ) | ( n5235 & n5243 ) | ( ~n5230 & n5243 ) ;
  assign n5593 = ( n5230 & n5590 ) | ( n5230 & n5591 ) | ( n5590 & n5591 ) ;
  assign n5592 = ( n5243 & ~n5591 ) | ( n5243 & n5590 ) | ( ~n5591 & n5590 ) ;
  assign n5594 = ( n5235 & ~n5593 ) | ( n5235 & n5592 ) | ( ~n5593 & n5592 ) ;
  assign n5595 = ( n5589 & ~n315 ) | ( n5589 & n5594 ) | ( ~n315 & n5594 ) ;
  assign n5596 = ( n240 & ~n5595 ) | ( n240 & 1'b0 ) | ( ~n5595 & 1'b0 ) ;
  assign n5597 = n5263 | n5327 ;
  assign n5598 = ( n5250 & ~n5263 ) | ( n5250 & n5259 ) | ( ~n5263 & n5259 ) ;
  assign n5600 = ( n5263 & n5597 ) | ( n5263 & n5598 ) | ( n5597 & n5598 ) ;
  assign n5599 = ( n5259 & ~n5598 ) | ( n5259 & n5597 ) | ( ~n5598 & n5597 ) ;
  assign n5601 = ( n5250 & ~n5600 ) | ( n5250 & n5599 ) | ( ~n5600 & n5599 ) ;
  assign n5602 = n315 | n5574 ;
  assign n5603 = ( n5588 & ~n5602 ) | ( n5588 & 1'b0 ) | ( ~n5602 & 1'b0 ) ;
  assign n5604 = n5594 | n5603 ;
  assign n5605 = ( n5582 & ~n5585 ) | ( n5582 & 1'b0 ) | ( ~n5585 & 1'b0 ) ;
  assign n5606 = ( n5579 & ~n396 ) | ( n5579 & n5605 ) | ( ~n396 & n5605 ) ;
  assign n5607 = ( n315 & ~n5606 ) | ( n315 & 1'b0 ) | ( ~n5606 & 1'b0 ) ;
  assign n5608 = n240 | n5607 ;
  assign n5609 = ( n5604 & ~n5608 ) | ( n5604 & 1'b0 ) | ( ~n5608 & 1'b0 ) ;
  assign n5610 = ( n5601 & ~n5609 ) | ( n5601 & 1'b0 ) | ( ~n5609 & 1'b0 ) ;
  assign n5611 = n5596 | n5610 ;
  assign n5613 = ( n5252 & ~n5257 ) | ( n5252 & n5265 ) | ( ~n5257 & n5265 ) ;
  assign n5612 = n5252 | n5327 ;
  assign n5615 = ( n5252 & ~n5613 ) | ( n5252 & n5612 ) | ( ~n5613 & n5612 ) ;
  assign n5614 = ( n5612 & ~n5265 ) | ( n5612 & n5613 ) | ( ~n5265 & n5613 ) ;
  assign n5616 = ( n5257 & ~n5615 ) | ( n5257 & n5614 ) | ( ~n5615 & n5614 ) ;
  assign n5617 = ( n181 & n5611 ) | ( n181 & n5616 ) | ( n5611 & n5616 ) ;
  assign n5618 = ~n145 & n5617 ;
  assign n5620 = ( n5281 & ~n5272 ) | ( n5281 & n5285 ) | ( ~n5272 & n5285 ) ;
  assign n5619 = n5285 | n5327 ;
  assign n5622 = ( n5285 & ~n5620 ) | ( n5285 & n5619 ) | ( ~n5620 & n5619 ) ;
  assign n5621 = ( n5619 & ~n5281 ) | ( n5619 & n5620 ) | ( ~n5281 & n5620 ) ;
  assign n5623 = ( n5272 & ~n5622 ) | ( n5272 & n5621 ) | ( ~n5622 & n5621 ) ;
  assign n5624 = n181 | n5596 ;
  assign n5625 = n5610 | n5624 ;
  assign n5626 = n5616 &  n5625 ;
  assign n5627 = ( n5604 & ~n5607 ) | ( n5604 & 1'b0 ) | ( ~n5607 & 1'b0 ) ;
  assign n5628 = ( n240 & ~n5627 ) | ( n240 & n5601 ) | ( ~n5627 & n5601 ) ;
  assign n5629 = n181 &  n5628 ;
  assign n5630 = ( n145 & ~n5629 ) | ( n145 & 1'b0 ) | ( ~n5629 & 1'b0 ) ;
  assign n5631 = ~n5626 & n5630 ;
  assign n5632 = n5623 | n5631 ;
  assign n5633 = ~n5618 & n5632 ;
  assign n5634 = n5274 | n5327 ;
  assign n5635 = ( n5274 & ~n5287 ) | ( n5274 & n5279 ) | ( ~n5287 & n5279 ) ;
  assign n5636 = ( n5287 & n5634 ) | ( n5287 & n5635 ) | ( n5634 & n5635 ) ;
  assign n5637 = ( n5274 & ~n5635 ) | ( n5274 & n5634 ) | ( ~n5635 & n5634 ) ;
  assign n5638 = ( n5279 & ~n5636 ) | ( n5279 & n5637 ) | ( ~n5636 & n5637 ) ;
  assign n5639 = ( n5633 & ~n150 ) | ( n5633 & n5638 ) | ( ~n150 & n5638 ) ;
  assign n5651 = ~n5650 & n5639 ;
  assign n5652 = ( n5651 & ~n133 ) | ( n5651 & n5650 ) | ( ~n133 & n5650 ) ;
  assign n5655 = n5626 | n5629 ;
  assign n5656 = ( n145 & ~n5655 ) | ( n145 & n5623 ) | ( ~n5655 & n5623 ) ;
  assign n5657 = ( n150 & ~n5656 ) | ( n150 & 1'b0 ) | ( ~n5656 & 1'b0 ) ;
  assign n5658 = ( n5646 & ~n5657 ) | ( n5646 & 1'b0 ) | ( ~n5657 & 1'b0 ) ;
  assign n5653 = n150 | n5618 ;
  assign n5654 = ( n5632 & ~n5653 ) | ( n5632 & 1'b0 ) | ( ~n5653 & 1'b0 ) ;
  assign n5659 = ~n5638 & n5654 ;
  assign n5660 = ( n5638 & n5658 ) | ( n5638 & n5659 ) | ( n5658 & n5659 ) ;
  assign n5662 = ( n5294 & ~n133 ) | ( n5294 & n5301 ) | ( ~n133 & n5301 ) ;
  assign n5661 = ( n5294 & n5301 ) | ( n5294 & n5327 ) | ( n5301 & n5327 ) ;
  assign n5663 = ~n5301 & n5661 ;
  assign n5664 = ( n5301 & ~n5662 ) | ( n5301 & n5663 ) | ( ~n5662 & n5663 ) ;
  assign n5665 = n5297 | n5324 ;
  assign n5666 = ( n5300 & n5319 ) | ( n5300 & n5665 ) | ( n5319 & n5665 ) ;
  assign n5667 = ( n5300 & ~n5666 ) | ( n5300 & 1'b0 ) | ( ~n5666 & 1'b0 ) ;
  assign n5668 = ( n5307 & ~n5315 ) | ( n5307 & n5667 ) | ( ~n5315 & n5667 ) ;
  assign n5669 = ~n5307 & n5668 ;
  assign n5670 = n5664 | n5669 ;
  assign n5671 = n5660 | n5670 ;
  assign n5672 = ~n5652 &  ~n5671 ;
  assign n5869 = ~n5519 & n5672 ;
  assign n5870 = ( n5506 & ~n5519 ) | ( n5506 & n5515 ) | ( ~n5519 & n5515 ) ;
  assign n5871 = ( n5869 & ~n5515 ) | ( n5869 & n5870 ) | ( ~n5515 & n5870 ) ;
  assign n5872 = ( n5519 & ~n5869 ) | ( n5519 & n5870 ) | ( ~n5869 & n5870 ) ;
  assign n5873 = ( n5871 & ~n5506 ) | ( n5871 & n5872 ) | ( ~n5506 & n5872 ) ;
  assign n5675 = x64 | x65 ;
  assign n5680 = ~x66 & n5675 ;
  assign n5681 = ( x66 & ~n5325 ) | ( x66 & n5680 ) | ( ~n5325 & n5680 ) ;
  assign n5682 = ( n5307 & ~n5315 ) | ( n5307 & n5681 ) | ( ~n5315 & n5681 ) ;
  assign n5683 = ~n5307 & n5682 ;
  assign n5684 = ( x67 & ~n5683 ) | ( x67 & n5672 ) | ( ~n5683 & n5672 ) ;
  assign n5679 = ( x66 & x67 ) | ( x66 & n5672 ) | ( x67 & n5672 ) ;
  assign n5685 = ( x66 & ~x67 ) | ( x66 & 1'b0 ) | ( ~x67 & 1'b0 ) ;
  assign n5686 = ( n5684 & ~n5679 ) | ( n5684 & n5685 ) | ( ~n5679 & n5685 ) ;
  assign n5676 = x66 | n5675 ;
  assign n5677 = ( x66 & ~n5672 ) | ( x66 & 1'b0 ) | ( ~n5672 & 1'b0 ) ;
  assign n5678 = ( n5327 & ~n5676 ) | ( n5327 & n5677 ) | ( ~n5676 & n5677 ) ;
  assign n5687 = ( n5678 & ~n5686 ) | ( n5678 & 1'b0 ) | ( ~n5686 & 1'b0 ) ;
  assign n5688 = ( n4990 & n5686 ) | ( n4990 & n5687 ) | ( n5686 & n5687 ) ;
  assign n5689 = n4990 | n5678 ;
  assign n5690 = n5686 | n5689 ;
  assign n5691 = n4991 | n5672 ;
  assign n5692 = ( n5327 & ~n5669 ) | ( n5327 & 1'b0 ) | ( ~n5669 & 1'b0 ) ;
  assign n5693 = ( n5660 & ~n5664 ) | ( n5660 & n5692 ) | ( ~n5664 & n5692 ) ;
  assign n5694 = ~n5660 & n5693 ;
  assign n5695 = ~n5652 & n5694 ;
  assign n5696 = n5691 | n5695 ;
  assign n5697 = ( x68 & ~n5696 ) | ( x68 & n5695 ) | ( ~n5696 & n5695 ) ;
  assign n5698 = x68 | n5695 ;
  assign n5699 = ( n5691 & ~n5698 ) | ( n5691 & 1'b0 ) | ( ~n5698 & 1'b0 ) ;
  assign n5700 = n5697 | n5699 ;
  assign n5701 = n5690 &  n5700 ;
  assign n5702 = n5688 | n5701 ;
  assign n5703 = ( n5327 & ~x68 ) | ( n5327 & n5334 ) | ( ~x68 & n5334 ) ;
  assign n5704 = x68 &  n5703 ;
  assign n5705 = ( n5329 & ~n5704 ) | ( n5329 & n5334 ) | ( ~n5704 & n5334 ) ;
  assign n5706 = ~x68 & n5327 ;
  assign n5707 = ( x69 & ~n5706 ) | ( x69 & 1'b0 ) | ( ~n5706 & 1'b0 ) ;
  assign n5708 = n5339 | n5707 ;
  assign n5709 = ( n5672 & ~n5705 ) | ( n5672 & n5708 ) | ( ~n5705 & n5708 ) ;
  assign n5710 = n5705 | n5709 ;
  assign n5711 = ~n5672 & n5709 ;
  assign n5712 = ( n5710 & ~n5708 ) | ( n5710 & n5711 ) | ( ~n5708 & n5711 ) ;
  assign n5713 = ( n4668 & n5702 ) | ( n4668 & n5712 ) | ( n5702 & n5712 ) ;
  assign n5714 = n4353 &  n5713 ;
  assign n5715 = ~n5362 & n5365 ;
  assign n5716 = ( n5348 & ~n5362 ) | ( n5348 & n5715 ) | ( ~n5362 & n5715 ) ;
  assign n5717 = ( n5672 & ~n5715 ) | ( n5672 & n5716 ) | ( ~n5715 & n5716 ) ;
  assign n5718 = ( n5362 & ~n5672 ) | ( n5362 & n5716 ) | ( ~n5672 & n5716 ) ;
  assign n5719 = ( n5717 & ~n5348 ) | ( n5717 & n5718 ) | ( ~n5348 & n5718 ) ;
  assign n5720 = n4668 | n5688 ;
  assign n5721 = n5701 | n5720 ;
  assign n5722 = n5712 &  n5721 ;
  assign n5723 = n5678 | n5686 ;
  assign n5724 = ( n4990 & n5700 ) | ( n4990 & n5723 ) | ( n5700 & n5723 ) ;
  assign n5725 = n4668 &  n5724 ;
  assign n5726 = n4353 | n5725 ;
  assign n5727 = n5722 | n5726 ;
  assign n5728 = n5719 &  n5727 ;
  assign n5729 = n5714 | n5728 ;
  assign n5730 = ( n5367 & ~n5672 ) | ( n5367 & 1'b0 ) | ( ~n5672 & 1'b0 ) ;
  assign n5731 = ( n5350 & ~n5672 ) | ( n5350 & n5360 ) | ( ~n5672 & n5360 ) ;
  assign n5732 = ( n5672 & ~n5730 ) | ( n5672 & n5731 ) | ( ~n5730 & n5731 ) ;
  assign n5733 = ( n5730 & ~n5350 ) | ( n5730 & n5731 ) | ( ~n5350 & n5731 ) ;
  assign n5734 = ( n5732 & ~n5360 ) | ( n5732 & n5733 ) | ( ~n5360 & n5733 ) ;
  assign n5735 = ( n4053 & n5729 ) | ( n4053 & n5734 ) | ( n5729 & n5734 ) ;
  assign n5736 = n3760 &  n5735 ;
  assign n5737 = ~n5387 & n5672 ;
  assign n5738 = ( n5374 & ~n5387 ) | ( n5374 & n5383 ) | ( ~n5387 & n5383 ) ;
  assign n5739 = ( n5737 & ~n5383 ) | ( n5737 & n5738 ) | ( ~n5383 & n5738 ) ;
  assign n5740 = ( n5387 & ~n5737 ) | ( n5387 & n5738 ) | ( ~n5737 & n5738 ) ;
  assign n5741 = ( n5739 & ~n5374 ) | ( n5739 & n5740 ) | ( ~n5374 & n5740 ) ;
  assign n5742 = n4053 | n5714 ;
  assign n5743 = n5728 | n5742 ;
  assign n5744 = n5734 &  n5743 ;
  assign n5745 = n5722 | n5725 ;
  assign n5746 = ( n4353 & n5719 ) | ( n4353 & n5745 ) | ( n5719 & n5745 ) ;
  assign n5747 = n4053 &  n5746 ;
  assign n5748 = n3760 | n5747 ;
  assign n5749 = n5744 | n5748 ;
  assign n5750 = n5741 &  n5749 ;
  assign n5751 = n5736 | n5750 ;
  assign n5752 = ( n5389 & ~n5672 ) | ( n5389 & 1'b0 ) | ( ~n5672 & 1'b0 ) ;
  assign n5753 = ( n5672 & ~n5376 ) | ( n5672 & n5752 ) | ( ~n5376 & n5752 ) ;
  assign n5755 = ( n5376 & n5381 ) | ( n5376 & n5753 ) | ( n5381 & n5753 ) ;
  assign n5754 = ( n5376 & ~n5381 ) | ( n5376 & n5753 ) | ( ~n5381 & n5753 ) ;
  assign n5756 = ( n5381 & ~n5755 ) | ( n5381 & n5754 ) | ( ~n5755 & n5754 ) ;
  assign n5757 = ( n3482 & n5751 ) | ( n3482 & n5756 ) | ( n5751 & n5756 ) ;
  assign n5758 = n3211 &  n5757 ;
  assign n5759 = ~n5409 & n5672 ;
  assign n5760 = ( n5396 & ~n5405 ) | ( n5396 & n5409 ) | ( ~n5405 & n5409 ) ;
  assign n5761 = ( n5405 & ~n5759 ) | ( n5405 & n5760 ) | ( ~n5759 & n5760 ) ;
  assign n5762 = ( n5759 & ~n5409 ) | ( n5759 & n5760 ) | ( ~n5409 & n5760 ) ;
  assign n5763 = ( n5761 & ~n5396 ) | ( n5761 & n5762 ) | ( ~n5396 & n5762 ) ;
  assign n5764 = n3482 | n5736 ;
  assign n5765 = n5750 | n5764 ;
  assign n5766 = n5756 &  n5765 ;
  assign n5767 = n5744 | n5747 ;
  assign n5768 = ( n3760 & n5741 ) | ( n3760 & n5767 ) | ( n5741 & n5767 ) ;
  assign n5769 = n3482 &  n5768 ;
  assign n5770 = n3211 | n5769 ;
  assign n5771 = n5766 | n5770 ;
  assign n5772 = n5763 &  n5771 ;
  assign n5773 = n5758 | n5772 ;
  assign n5774 = ~n5398 & n5672 ;
  assign n5775 = ( n5403 & ~n5398 ) | ( n5403 & n5411 ) | ( ~n5398 & n5411 ) ;
  assign n5776 = ( n5774 & ~n5411 ) | ( n5774 & n5775 ) | ( ~n5411 & n5775 ) ;
  assign n5777 = ( n5398 & ~n5774 ) | ( n5398 & n5775 ) | ( ~n5774 & n5775 ) ;
  assign n5778 = ( n5776 & ~n5403 ) | ( n5776 & n5777 ) | ( ~n5403 & n5777 ) ;
  assign n5779 = ( n2955 & n5773 ) | ( n2955 & n5778 ) | ( n5773 & n5778 ) ;
  assign n5780 = n2706 &  n5779 ;
  assign n5781 = ~n5431 & n5672 ;
  assign n5782 = ( n5418 & ~n5427 ) | ( n5418 & n5431 ) | ( ~n5427 & n5431 ) ;
  assign n5783 = ( n5427 & ~n5781 ) | ( n5427 & n5782 ) | ( ~n5781 & n5782 ) ;
  assign n5784 = ( n5781 & ~n5431 ) | ( n5781 & n5782 ) | ( ~n5431 & n5782 ) ;
  assign n5785 = ( n5783 & ~n5418 ) | ( n5783 & n5784 ) | ( ~n5418 & n5784 ) ;
  assign n5786 = n2955 | n5758 ;
  assign n5787 = n5772 | n5786 ;
  assign n5788 = n5778 &  n5787 ;
  assign n5789 = n5766 | n5769 ;
  assign n5790 = ( n3211 & n5763 ) | ( n3211 & n5789 ) | ( n5763 & n5789 ) ;
  assign n5791 = n2955 &  n5790 ;
  assign n5792 = n2706 | n5791 ;
  assign n5793 = n5788 | n5792 ;
  assign n5794 = n5785 &  n5793 ;
  assign n5795 = n5780 | n5794 ;
  assign n5796 = ~n5420 & n5672 ;
  assign n5797 = ( n5420 & ~n5433 ) | ( n5420 & n5425 ) | ( ~n5433 & n5425 ) ;
  assign n5798 = ( n5433 & ~n5796 ) | ( n5433 & n5797 ) | ( ~n5796 & n5797 ) ;
  assign n5799 = ( n5796 & ~n5420 ) | ( n5796 & n5797 ) | ( ~n5420 & n5797 ) ;
  assign n5800 = ( n5798 & ~n5425 ) | ( n5798 & n5799 ) | ( ~n5425 & n5799 ) ;
  assign n5801 = ( n2472 & n5795 ) | ( n2472 & n5800 ) | ( n5795 & n5800 ) ;
  assign n5802 = n2245 &  n5801 ;
  assign n5803 = ~n5453 & n5672 ;
  assign n5804 = ( n5440 & ~n5453 ) | ( n5440 & n5449 ) | ( ~n5453 & n5449 ) ;
  assign n5805 = ( n5803 & ~n5449 ) | ( n5803 & n5804 ) | ( ~n5449 & n5804 ) ;
  assign n5806 = ( n5453 & ~n5803 ) | ( n5453 & n5804 ) | ( ~n5803 & n5804 ) ;
  assign n5807 = ( n5805 & ~n5440 ) | ( n5805 & n5806 ) | ( ~n5440 & n5806 ) ;
  assign n5808 = n2472 | n5780 ;
  assign n5809 = n5794 | n5808 ;
  assign n5810 = n5800 &  n5809 ;
  assign n5811 = n5788 | n5791 ;
  assign n5812 = ( n2706 & n5785 ) | ( n2706 & n5811 ) | ( n5785 & n5811 ) ;
  assign n5813 = n2472 &  n5812 ;
  assign n5814 = n2245 | n5813 ;
  assign n5815 = n5810 | n5814 ;
  assign n5816 = n5807 &  n5815 ;
  assign n5817 = n5802 | n5816 ;
  assign n5818 = ( n5455 & ~n5672 ) | ( n5455 & 1'b0 ) | ( ~n5672 & 1'b0 ) ;
  assign n5819 = ( n5672 & ~n5442 ) | ( n5672 & n5818 ) | ( ~n5442 & n5818 ) ;
  assign n5821 = ( n5442 & n5447 ) | ( n5442 & n5819 ) | ( n5447 & n5819 ) ;
  assign n5820 = ( n5442 & ~n5447 ) | ( n5442 & n5819 ) | ( ~n5447 & n5819 ) ;
  assign n5822 = ( n5447 & ~n5821 ) | ( n5447 & n5820 ) | ( ~n5821 & n5820 ) ;
  assign n5823 = ( n5817 & ~n2033 ) | ( n5817 & n5822 ) | ( ~n2033 & n5822 ) ;
  assign n5824 = n1827 &  n5823 ;
  assign n5826 = ( n5471 & ~n5462 ) | ( n5471 & n5475 ) | ( ~n5462 & n5475 ) ;
  assign n5825 = n5475 &  n5672 ;
  assign n5828 = ( n5475 & ~n5826 ) | ( n5475 & n5825 ) | ( ~n5826 & n5825 ) ;
  assign n5827 = ( n5825 & ~n5471 ) | ( n5825 & n5826 ) | ( ~n5471 & n5826 ) ;
  assign n5829 = ( n5462 & ~n5828 ) | ( n5462 & n5827 ) | ( ~n5828 & n5827 ) ;
  assign n5830 = ( n2033 & ~n5802 ) | ( n2033 & 1'b0 ) | ( ~n5802 & 1'b0 ) ;
  assign n5831 = ~n5816 & n5830 ;
  assign n5832 = ( n5822 & ~n5831 ) | ( n5822 & 1'b0 ) | ( ~n5831 & 1'b0 ) ;
  assign n5833 = n5810 | n5813 ;
  assign n5834 = ( n2245 & n5807 ) | ( n2245 & n5833 ) | ( n5807 & n5833 ) ;
  assign n5835 = ~n2033 & n5834 ;
  assign n5836 = n1827 | n5835 ;
  assign n5837 = n5832 | n5836 ;
  assign n5838 = ~n5829 & n5837 ;
  assign n5839 = n5824 | n5838 ;
  assign n5840 = ~n5464 & n5672 ;
  assign n5841 = ( n5469 & ~n5464 ) | ( n5469 & n5477 ) | ( ~n5464 & n5477 ) ;
  assign n5842 = ( n5840 & ~n5477 ) | ( n5840 & n5841 ) | ( ~n5477 & n5841 ) ;
  assign n5843 = ( n5464 & ~n5840 ) | ( n5464 & n5841 ) | ( ~n5840 & n5841 ) ;
  assign n5844 = ( n5842 & ~n5469 ) | ( n5842 & n5843 ) | ( ~n5469 & n5843 ) ;
  assign n5845 = ( n5839 & ~n1636 ) | ( n5839 & n5844 ) | ( ~n1636 & n5844 ) ;
  assign n5846 = ~n1452 & n5845 ;
  assign n5848 = ( n5493 & ~n5484 ) | ( n5493 & n5497 ) | ( ~n5484 & n5497 ) ;
  assign n5847 = n5497 &  n5672 ;
  assign n5850 = ( n5497 & ~n5848 ) | ( n5497 & n5847 ) | ( ~n5848 & n5847 ) ;
  assign n5849 = ( n5847 & ~n5493 ) | ( n5847 & n5848 ) | ( ~n5493 & n5848 ) ;
  assign n5851 = ( n5484 & ~n5850 ) | ( n5484 & n5849 ) | ( ~n5850 & n5849 ) ;
  assign n5852 = ( n1636 & ~n5824 ) | ( n1636 & 1'b0 ) | ( ~n5824 & 1'b0 ) ;
  assign n5853 = ~n5838 & n5852 ;
  assign n5854 = ( n5844 & ~n5853 ) | ( n5844 & 1'b0 ) | ( ~n5853 & 1'b0 ) ;
  assign n5855 = n5832 | n5835 ;
  assign n5856 = ( n1827 & ~n5829 ) | ( n1827 & n5855 ) | ( ~n5829 & n5855 ) ;
  assign n5857 = ~n1636 & n5856 ;
  assign n5858 = ( n1452 & ~n5857 ) | ( n1452 & 1'b0 ) | ( ~n5857 & 1'b0 ) ;
  assign n5859 = ~n5854 & n5858 ;
  assign n5860 = n5851 | n5859 ;
  assign n5861 = ~n5846 & n5860 ;
  assign n5863 = ( n5486 & ~n5491 ) | ( n5486 & n5499 ) | ( ~n5491 & n5499 ) ;
  assign n5862 = n5486 &  n5672 ;
  assign n5865 = ( n5486 & ~n5863 ) | ( n5486 & n5862 ) | ( ~n5863 & n5862 ) ;
  assign n5864 = ( n5862 & ~n5499 ) | ( n5862 & n5863 ) | ( ~n5499 & n5863 ) ;
  assign n5866 = ( n5491 & ~n5865 ) | ( n5491 & n5864 ) | ( ~n5865 & n5864 ) ;
  assign n5867 = ( n5861 & ~n1283 ) | ( n5861 & n5866 ) | ( ~n1283 & n5866 ) ;
  assign n5868 = n1122 | n5867 ;
  assign n5972 = ~n5596 & n5672 ;
  assign n5973 = ( n5596 & ~n5609 ) | ( n5596 & n5601 ) | ( ~n5609 & n5601 ) ;
  assign n5974 = ( n5609 & ~n5972 ) | ( n5609 & n5973 ) | ( ~n5972 & n5973 ) ;
  assign n5975 = ( n5972 & ~n5596 ) | ( n5972 & n5973 ) | ( ~n5596 & n5973 ) ;
  assign n5976 = ( n5974 & ~n5601 ) | ( n5974 & n5975 ) | ( ~n5601 & n5975 ) ;
  assign n5874 = n1283 | n5846 ;
  assign n5875 = ( n5860 & ~n5874 ) | ( n5860 & 1'b0 ) | ( ~n5874 & 1'b0 ) ;
  assign n5876 = n5866 | n5875 ;
  assign n5877 = n5854 | n5857 ;
  assign n5878 = ( n1452 & ~n5877 ) | ( n1452 & n5851 ) | ( ~n5877 & n5851 ) ;
  assign n5879 = ( n1283 & ~n5878 ) | ( n1283 & 1'b0 ) | ( ~n5878 & 1'b0 ) ;
  assign n5880 = ( n1122 & ~n5879 ) | ( n1122 & 1'b0 ) | ( ~n5879 & 1'b0 ) ;
  assign n5881 = n5876 &  n5880 ;
  assign n5882 = ( n5873 & ~n5881 ) | ( n5873 & 1'b0 ) | ( ~n5881 & 1'b0 ) ;
  assign n5883 = ( n5868 & ~n5882 ) | ( n5868 & 1'b0 ) | ( ~n5882 & 1'b0 ) ;
  assign n5884 = ( n5521 & ~n5672 ) | ( n5521 & 1'b0 ) | ( ~n5672 & 1'b0 ) ;
  assign n5885 = ( n5508 & n5672 ) | ( n5508 & n5884 ) | ( n5672 & n5884 ) ;
  assign n5886 = ( n5508 & ~n5885 ) | ( n5508 & n5513 ) | ( ~n5885 & n5513 ) ;
  assign n5887 = ( n5513 & ~n5508 ) | ( n5513 & n5885 ) | ( ~n5508 & n5885 ) ;
  assign n5888 = ( n5886 & ~n5513 ) | ( n5886 & n5887 ) | ( ~n5513 & n5887 ) ;
  assign n5889 = ( n976 & n5883 ) | ( n976 & n5888 ) | ( n5883 & n5888 ) ;
  assign n5890 = ( n837 & ~n5889 ) | ( n837 & 1'b0 ) | ( ~n5889 & 1'b0 ) ;
  assign n5892 = ( n5537 & ~n5528 ) | ( n5537 & n5541 ) | ( ~n5528 & n5541 ) ;
  assign n5891 = n5541 &  n5672 ;
  assign n5894 = ( n5541 & ~n5892 ) | ( n5541 & n5891 ) | ( ~n5892 & n5891 ) ;
  assign n5893 = ( n5891 & ~n5537 ) | ( n5891 & n5892 ) | ( ~n5537 & n5892 ) ;
  assign n5895 = ( n5528 & ~n5894 ) | ( n5528 & n5893 ) | ( ~n5894 & n5893 ) ;
  assign n5896 = n976 &  n5868 ;
  assign n5897 = ~n5882 & n5896 ;
  assign n5898 = n5888 | n5897 ;
  assign n5899 = ( n5876 & ~n5879 ) | ( n5876 & 1'b0 ) | ( ~n5879 & 1'b0 ) ;
  assign n5900 = ( n1122 & ~n5873 ) | ( n1122 & n5899 ) | ( ~n5873 & n5899 ) ;
  assign n5901 = n976 | n5900 ;
  assign n5902 = ~n837 & n5901 ;
  assign n5903 = n5898 &  n5902 ;
  assign n5904 = n5895 | n5903 ;
  assign n5905 = ~n5890 & n5904 ;
  assign n5906 = ~n5530 & n5672 ;
  assign n5907 = ( n5535 & ~n5530 ) | ( n5535 & n5543 ) | ( ~n5530 & n5543 ) ;
  assign n5908 = ( n5906 & ~n5543 ) | ( n5906 & n5907 ) | ( ~n5543 & n5907 ) ;
  assign n5909 = ( n5530 & ~n5906 ) | ( n5530 & n5907 ) | ( ~n5906 & n5907 ) ;
  assign n5910 = ( n5908 & ~n5535 ) | ( n5908 & n5909 ) | ( ~n5535 & n5909 ) ;
  assign n5911 = ( n713 & ~n5905 ) | ( n713 & n5910 ) | ( ~n5905 & n5910 ) ;
  assign n5912 = n595 &  n5911 ;
  assign n5913 = ~n5563 & n5672 ;
  assign n5914 = ( n5550 & ~n5559 ) | ( n5550 & n5563 ) | ( ~n5559 & n5563 ) ;
  assign n5915 = ( n5559 & ~n5913 ) | ( n5559 & n5914 ) | ( ~n5913 & n5914 ) ;
  assign n5916 = ( n5913 & ~n5563 ) | ( n5913 & n5914 ) | ( ~n5563 & n5914 ) ;
  assign n5917 = ( n5915 & ~n5550 ) | ( n5915 & n5916 ) | ( ~n5550 & n5916 ) ;
  assign n5918 = n713 | n5890 ;
  assign n5919 = ( n5904 & ~n5918 ) | ( n5904 & 1'b0 ) | ( ~n5918 & 1'b0 ) ;
  assign n5920 = ( n5910 & ~n5919 ) | ( n5910 & 1'b0 ) | ( ~n5919 & 1'b0 ) ;
  assign n5921 = n5898 &  n5901 ;
  assign n5922 = ( n5895 & ~n837 ) | ( n5895 & n5921 ) | ( ~n837 & n5921 ) ;
  assign n5923 = ( n713 & ~n5922 ) | ( n713 & 1'b0 ) | ( ~n5922 & 1'b0 ) ;
  assign n5924 = n595 | n5923 ;
  assign n5925 = n5920 | n5924 ;
  assign n5926 = n5917 &  n5925 ;
  assign n5927 = n5912 | n5926 ;
  assign n5928 = ~n5552 & n5672 ;
  assign n5929 = ( n5552 & ~n5565 ) | ( n5552 & n5557 ) | ( ~n5565 & n5557 ) ;
  assign n5930 = ( n5565 & ~n5928 ) | ( n5565 & n5929 ) | ( ~n5928 & n5929 ) ;
  assign n5931 = ( n5928 & ~n5552 ) | ( n5928 & n5929 ) | ( ~n5552 & n5929 ) ;
  assign n5932 = ( n5930 & ~n5557 ) | ( n5930 & n5931 ) | ( ~n5557 & n5931 ) ;
  assign n5933 = ( n492 & n5927 ) | ( n492 & n5932 ) | ( n5927 & n5932 ) ;
  assign n5934 = n396 &  n5933 ;
  assign n5935 = ~n5585 & n5672 ;
  assign n5936 = ( n5572 & ~n5585 ) | ( n5572 & n5581 ) | ( ~n5585 & n5581 ) ;
  assign n5937 = ( n5935 & ~n5581 ) | ( n5935 & n5936 ) | ( ~n5581 & n5936 ) ;
  assign n5938 = ( n5585 & ~n5935 ) | ( n5585 & n5936 ) | ( ~n5935 & n5936 ) ;
  assign n5939 = ( n5937 & ~n5572 ) | ( n5937 & n5938 ) | ( ~n5572 & n5938 ) ;
  assign n5940 = n492 | n5912 ;
  assign n5941 = n5926 | n5940 ;
  assign n5942 = n5932 &  n5941 ;
  assign n5943 = n5920 | n5923 ;
  assign n5944 = ( n595 & n5917 ) | ( n595 & n5943 ) | ( n5917 & n5943 ) ;
  assign n5945 = n492 &  n5944 ;
  assign n5946 = n396 | n5945 ;
  assign n5947 = n5942 | n5946 ;
  assign n5948 = n5939 &  n5947 ;
  assign n5949 = n5934 | n5948 ;
  assign n5950 = ( n5587 & ~n5672 ) | ( n5587 & 1'b0 ) | ( ~n5672 & 1'b0 ) ;
  assign n5951 = ( n5579 & ~n5574 ) | ( n5579 & n5672 ) | ( ~n5574 & n5672 ) ;
  assign n5952 = ( n5950 & ~n5672 ) | ( n5950 & n5951 ) | ( ~n5672 & n5951 ) ;
  assign n5953 = ( n5574 & ~n5950 ) | ( n5574 & n5951 ) | ( ~n5950 & n5951 ) ;
  assign n5954 = ( n5952 & ~n5579 ) | ( n5952 & n5953 ) | ( ~n5579 & n5953 ) ;
  assign n5955 = ( n315 & n5949 ) | ( n315 & n5954 ) | ( n5949 & n5954 ) ;
  assign n5956 = n240 &  n5955 ;
  assign n5957 = ~n5607 & n5672 ;
  assign n5958 = ( n5594 & ~n5603 ) | ( n5594 & n5607 ) | ( ~n5603 & n5607 ) ;
  assign n5959 = ( n5603 & ~n5957 ) | ( n5603 & n5958 ) | ( ~n5957 & n5958 ) ;
  assign n5960 = ( n5957 & ~n5607 ) | ( n5957 & n5958 ) | ( ~n5607 & n5958 ) ;
  assign n5961 = ( n5959 & ~n5594 ) | ( n5959 & n5960 ) | ( ~n5594 & n5960 ) ;
  assign n5962 = n315 | n5934 ;
  assign n5963 = n5948 | n5962 ;
  assign n5964 = n5954 &  n5963 ;
  assign n5965 = n5942 | n5945 ;
  assign n5966 = ( n396 & n5939 ) | ( n396 & n5965 ) | ( n5939 & n5965 ) ;
  assign n5967 = n315 &  n5966 ;
  assign n5968 = n240 | n5967 ;
  assign n5969 = n5964 | n5968 ;
  assign n5970 = n5961 &  n5969 ;
  assign n5971 = n5956 | n5970 ;
  assign n5977 = ( n181 & ~n5976 ) | ( n181 & n5971 ) | ( ~n5976 & n5971 ) ;
  assign n5978 = ~n145 & n5977 ;
  assign n5980 = ( n5625 & ~n5616 ) | ( n5625 & n5629 ) | ( ~n5616 & n5629 ) ;
  assign n5979 = ~n5629 & n5672 ;
  assign n5981 = ( n5625 & ~n5980 ) | ( n5625 & n5979 ) | ( ~n5980 & n5979 ) ;
  assign n5982 = ( n5979 & ~n5629 ) | ( n5979 & n5980 ) | ( ~n5629 & n5980 ) ;
  assign n5983 = ( n5616 & ~n5981 ) | ( n5616 & n5982 ) | ( ~n5981 & n5982 ) ;
  assign n5984 = n181 | n5956 ;
  assign n5985 = n5970 | n5984 ;
  assign n5986 = ~n5976 & n5985 ;
  assign n5987 = n5964 | n5967 ;
  assign n5988 = ( n240 & n5961 ) | ( n240 & n5987 ) | ( n5961 & n5987 ) ;
  assign n5989 = n181 &  n5988 ;
  assign n5990 = ( n145 & ~n5989 ) | ( n145 & 1'b0 ) | ( ~n5989 & 1'b0 ) ;
  assign n5991 = ~n5986 & n5990 ;
  assign n5992 = ( n5983 & ~n5991 ) | ( n5983 & 1'b0 ) | ( ~n5991 & 1'b0 ) ;
  assign n5993 = n5978 | n5992 ;
  assign n5994 = ( n5631 & ~n5672 ) | ( n5631 & 1'b0 ) | ( ~n5672 & 1'b0 ) ;
  assign n5995 = ( n5618 & ~n5672 ) | ( n5618 & n5623 ) | ( ~n5672 & n5623 ) ;
  assign n5996 = ( n5672 & ~n5994 ) | ( n5672 & n5995 ) | ( ~n5994 & n5995 ) ;
  assign n5997 = ( n5994 & ~n5618 ) | ( n5994 & n5995 ) | ( ~n5618 & n5995 ) ;
  assign n5998 = ( n5996 & ~n5623 ) | ( n5996 & n5997 ) | ( ~n5623 & n5997 ) ;
  assign n5999 = ( n150 & n5993 ) | ( n150 & n5998 ) | ( n5993 & n5998 ) ;
  assign n6000 = ( n5638 & ~n5654 ) | ( n5638 & 1'b0 ) | ( ~n5654 & 1'b0 ) ;
  assign n6001 = ( n5657 & ~n5672 ) | ( n5657 & n6000 ) | ( ~n5672 & n6000 ) ;
  assign n6002 = ~n5657 & n6001 ;
  assign n6003 = n5654 | n5657 ;
  assign n6004 = ~n6003 & n5672 ;
  assign n6005 = ( n6004 & ~n5638 ) | ( n6004 & n6003 ) | ( ~n5638 & n6003 ) ;
  assign n6006 = n6002 | n6005 ;
  assign n6007 = n5639 | n5646 ;
  assign n6008 = ~n6007 & n5672 ;
  assign n6009 = ( n6008 & ~n5660 ) | ( n6008 & n6007 ) | ( ~n5660 & n6007 ) ;
  assign n6010 = n6006 &  n6009 ;
  assign n6011 = ~n5999 & n6010 ;
  assign n6012 = ( n133 & ~n6011 ) | ( n133 & n6010 ) | ( ~n6011 & n6010 ) ;
  assign n6013 = n150 | n5978 ;
  assign n6014 = n5992 | n6013 ;
  assign n6019 = ( n5998 & ~n6014 ) | ( n5998 & 1'b0 ) | ( ~n6014 & 1'b0 ) ;
  assign n6015 = n5986 | n5989 ;
  assign n6016 = ( n5983 & ~n145 ) | ( n5983 & n6015 ) | ( ~n145 & n6015 ) ;
  assign n6017 = n150 &  n6016 ;
  assign n6018 = n6006 | n6017 ;
  assign n6020 = ( n5998 & ~n6019 ) | ( n5998 & n6018 ) | ( ~n6019 & n6018 ) ;
  assign n6022 = ( n5639 & ~n133 ) | ( n5639 & n5646 ) | ( ~n133 & n5646 ) ;
  assign n6021 = ( n5639 & ~n5672 ) | ( n5639 & n5646 ) | ( ~n5672 & n5646 ) ;
  assign n6023 = ~n5646 & n6021 ;
  assign n6024 = ( n5646 & ~n6022 ) | ( n5646 & n6023 ) | ( ~n6022 & n6023 ) ;
  assign n6025 = n5642 | n5669 ;
  assign n6026 = ( n5645 & n5664 ) | ( n5645 & n6025 ) | ( n5664 & n6025 ) ;
  assign n6027 = ( n5645 & ~n6026 ) | ( n5645 & 1'b0 ) | ( ~n6026 & 1'b0 ) ;
  assign n6028 = ( n5652 & ~n5660 ) | ( n5652 & n6027 ) | ( ~n5660 & n6027 ) ;
  assign n6029 = ~n5652 & n6028 ;
  assign n6030 = n6024 | n6029 ;
  assign n6031 = ( n6020 & ~n6030 ) | ( n6020 & 1'b0 ) | ( ~n6030 & 1'b0 ) ;
  assign n6032 = ~n6012 | ~n6031 ;
  assign n6251 = ( n5868 & ~n6032 ) | ( n5868 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n6252 = ( n5868 & n5873 ) | ( n5868 & n5881 ) | ( n5873 & n5881 ) ;
  assign n6253 = ( n6251 & ~n5881 ) | ( n6251 & n6252 ) | ( ~n5881 & n6252 ) ;
  assign n6254 = ( n5868 & ~n6252 ) | ( n5868 & n6251 ) | ( ~n6252 & n6251 ) ;
  assign n6255 = ( n5873 & ~n6253 ) | ( n5873 & n6254 ) | ( ~n6253 & n6254 ) ;
  assign n6033 = x64 &  n6032 ;
  assign n5674 = x64 | n5673 ;
  assign n6034 = ( n5672 & ~n6033 ) | ( n5672 & n5674 ) | ( ~n6033 & n5674 ) ;
  assign n6035 = ( x64 & ~n6032 ) | ( x64 & x65 ) | ( ~n6032 & x65 ) ;
  assign n6041 = ( x64 & ~x65 ) | ( x64 & 1'b0 ) | ( ~x65 & 1'b0 ) ;
  assign n6036 = ~x64 & n5673 ;
  assign n6037 = ( x64 & ~n5670 ) | ( x64 & n6036 ) | ( ~n5670 & n6036 ) ;
  assign n6038 = ( n5652 & ~n5660 ) | ( n5652 & n6037 ) | ( ~n5660 & n6037 ) ;
  assign n6039 = ~n5652 & n6038 ;
  assign n6040 = ( n6032 & ~x65 ) | ( n6032 & n6039 ) | ( ~x65 & n6039 ) ;
  assign n6042 = ( n6035 & ~n6041 ) | ( n6035 & n6040 ) | ( ~n6041 & n6040 ) ;
  assign n6043 = n6034 &  n6042 ;
  assign n6045 = n5672 | n6029 ;
  assign n6046 = ( n6020 & n6024 ) | ( n6020 & n6045 ) | ( n6024 & n6045 ) ;
  assign n6047 = ( n6020 & ~n6046 ) | ( n6020 & 1'b0 ) | ( ~n6046 & 1'b0 ) ;
  assign n6048 = n6012 &  n6047 ;
  assign n6044 = ~n5675 & n6032 ;
  assign n6049 = ~n6048 & n6044 ;
  assign n6050 = ( x66 & n6049 ) | ( x66 & n6048 ) | ( n6049 & n6048 ) ;
  assign n6051 = x66 | n6048 ;
  assign n6052 = n6044 | n6051 ;
  assign n6053 = ~n6050 & n6052 ;
  assign n6054 = ( n6043 & ~n5327 ) | ( n6043 & n6053 ) | ( ~n5327 & n6053 ) ;
  assign n6055 = ( n4990 & ~n6054 ) | ( n4990 & 1'b0 ) | ( ~n6054 & 1'b0 ) ;
  assign n6059 = x66 | n5672 ;
  assign n6060 = x67 &  n6059 ;
  assign n6061 = ( n5691 & ~n6060 ) | ( n5691 & 1'b0 ) | ( ~n6060 & 1'b0 ) ;
  assign n6056 = ( x66 & ~n5683 ) | ( x66 & n5672 ) | ( ~n5683 & n5672 ) ;
  assign n6057 = ( x66 & ~n6056 ) | ( x66 & 1'b0 ) | ( ~n6056 & 1'b0 ) ;
  assign n6058 = ( n5678 & ~n6057 ) | ( n5678 & n5683 ) | ( ~n6057 & n5683 ) ;
  assign n6062 = ( n6032 & n6058 ) | ( n6032 & n6061 ) | ( n6058 & n6061 ) ;
  assign n6063 = ~n6058 & n6062 ;
  assign n6064 = ( n6032 & ~n6062 ) | ( n6032 & 1'b0 ) | ( ~n6062 & 1'b0 ) ;
  assign n6065 = ( n6061 & ~n6063 ) | ( n6061 & n6064 ) | ( ~n6063 & n6064 ) ;
  assign n6066 = ~n5327 & n6034 ;
  assign n6067 = n6042 &  n6066 ;
  assign n6068 = n6053 | n6067 ;
  assign n6069 = ~n6034 & n6042 ;
  assign n6070 = ( n5327 & ~n6042 ) | ( n5327 & n6069 ) | ( ~n6042 & n6069 ) ;
  assign n6071 = n4990 | n6070 ;
  assign n6072 = ( n6068 & ~n6071 ) | ( n6068 & 1'b0 ) | ( ~n6071 & 1'b0 ) ;
  assign n6073 = ( n6065 & ~n6072 ) | ( n6065 & 1'b0 ) | ( ~n6072 & 1'b0 ) ;
  assign n6074 = n6055 | n6073 ;
  assign n6075 = n5688 &  n5690 ;
  assign n6076 = ( n5690 & n5700 ) | ( n5690 & n6075 ) | ( n5700 & n6075 ) ;
  assign n6077 = ( n6076 & ~n5690 ) | ( n6076 & n6032 ) | ( ~n5690 & n6032 ) ;
  assign n6078 = ( n6032 & ~n6076 ) | ( n6032 & n6075 ) | ( ~n6076 & n6075 ) ;
  assign n6079 = ( n5700 & ~n6077 ) | ( n5700 & n6078 ) | ( ~n6077 & n6078 ) ;
  assign n6080 = ( n4668 & n6074 ) | ( n4668 & n6079 ) | ( n6074 & n6079 ) ;
  assign n6081 = n4353 &  n6080 ;
  assign n6083 = ( n5721 & ~n5712 ) | ( n5721 & n5725 ) | ( ~n5712 & n5725 ) ;
  assign n6082 = n5725 | n6032 ;
  assign n6085 = ( n5725 & ~n6083 ) | ( n5725 & n6082 ) | ( ~n6083 & n6082 ) ;
  assign n6084 = ( n6082 & ~n5721 ) | ( n6082 & n6083 ) | ( ~n5721 & n6083 ) ;
  assign n6086 = ( n5712 & ~n6085 ) | ( n5712 & n6084 ) | ( ~n6085 & n6084 ) ;
  assign n6087 = n4668 | n6055 ;
  assign n6088 = n6073 | n6087 ;
  assign n6089 = n6079 &  n6088 ;
  assign n6090 = ( n6068 & ~n6070 ) | ( n6068 & 1'b0 ) | ( ~n6070 & 1'b0 ) ;
  assign n6091 = ( n4990 & ~n6090 ) | ( n4990 & n6065 ) | ( ~n6090 & n6065 ) ;
  assign n6092 = n4668 &  n6091 ;
  assign n6093 = n4353 | n6092 ;
  assign n6094 = n6089 | n6093 ;
  assign n6095 = n6086 &  n6094 ;
  assign n6096 = n6081 | n6095 ;
  assign n6097 = n5714 | n6032 ;
  assign n6098 = ( n5714 & n5719 ) | ( n5714 & n5727 ) | ( n5719 & n5727 ) ;
  assign n6099 = ( n6097 & ~n5727 ) | ( n6097 & n6098 ) | ( ~n5727 & n6098 ) ;
  assign n6100 = ( n5714 & ~n6098 ) | ( n5714 & n6097 ) | ( ~n6098 & n6097 ) ;
  assign n6101 = ( n5719 & ~n6099 ) | ( n5719 & n6100 ) | ( ~n6099 & n6100 ) ;
  assign n6102 = ( n4053 & n6096 ) | ( n4053 & n6101 ) | ( n6096 & n6101 ) ;
  assign n6103 = n3760 &  n6102 ;
  assign n6104 = n5747 | n6032 ;
  assign n6105 = ( n5734 & n5743 ) | ( n5734 & n5747 ) | ( n5743 & n5747 ) ;
  assign n6106 = ( n6104 & ~n5743 ) | ( n6104 & n6105 ) | ( ~n5743 & n6105 ) ;
  assign n6107 = ( n5747 & ~n6105 ) | ( n5747 & n6104 ) | ( ~n6105 & n6104 ) ;
  assign n6108 = ( n5734 & ~n6106 ) | ( n5734 & n6107 ) | ( ~n6106 & n6107 ) ;
  assign n6109 = n4053 | n6081 ;
  assign n6110 = n6095 | n6109 ;
  assign n6111 = n6101 &  n6110 ;
  assign n6112 = n6089 | n6092 ;
  assign n6113 = ( n4353 & n6086 ) | ( n4353 & n6112 ) | ( n6086 & n6112 ) ;
  assign n6114 = n4053 &  n6113 ;
  assign n6115 = n3760 | n6114 ;
  assign n6116 = n6111 | n6115 ;
  assign n6117 = n6108 &  n6116 ;
  assign n6118 = n6103 | n6117 ;
  assign n6119 = ~n5749 & n6032 ;
  assign n6120 = ( n5736 & n5741 ) | ( n5736 & n6032 ) | ( n5741 & n6032 ) ;
  assign n6122 = ( n6119 & ~n5736 ) | ( n6119 & n6120 ) | ( ~n5736 & n6120 ) ;
  assign n6121 = ( n6032 & ~n6120 ) | ( n6032 & n6119 ) | ( ~n6120 & n6119 ) ;
  assign n6123 = ( n5741 & ~n6122 ) | ( n5741 & n6121 ) | ( ~n6122 & n6121 ) ;
  assign n6124 = ( n3482 & n6118 ) | ( n3482 & n6123 ) | ( n6118 & n6123 ) ;
  assign n6125 = n3211 &  n6124 ;
  assign n6126 = n5769 | n6032 ;
  assign n6127 = ( n5756 & n5765 ) | ( n5756 & n5769 ) | ( n5765 & n5769 ) ;
  assign n6128 = ( n6126 & ~n5765 ) | ( n6126 & n6127 ) | ( ~n5765 & n6127 ) ;
  assign n6129 = ( n5769 & ~n6127 ) | ( n5769 & n6126 ) | ( ~n6127 & n6126 ) ;
  assign n6130 = ( n5756 & ~n6128 ) | ( n5756 & n6129 ) | ( ~n6128 & n6129 ) ;
  assign n6131 = n3482 | n6103 ;
  assign n6132 = n6117 | n6131 ;
  assign n6133 = n6123 &  n6132 ;
  assign n6134 = n6111 | n6114 ;
  assign n6135 = ( n3760 & n6108 ) | ( n3760 & n6134 ) | ( n6108 & n6134 ) ;
  assign n6136 = n3482 &  n6135 ;
  assign n6137 = n3211 | n6136 ;
  assign n6138 = n6133 | n6137 ;
  assign n6139 = n6130 &  n6138 ;
  assign n6140 = n6125 | n6139 ;
  assign n6141 = ~n5771 & n6032 ;
  assign n6142 = ( n5758 & ~n6141 ) | ( n5758 & n6032 ) | ( ~n6141 & n6032 ) ;
  assign n6143 = ( n5758 & ~n6142 ) | ( n5758 & n5763 ) | ( ~n6142 & n5763 ) ;
  assign n6144 = ( n5763 & ~n5758 ) | ( n5763 & n6142 ) | ( ~n5758 & n6142 ) ;
  assign n6145 = ( n6143 & ~n5763 ) | ( n6143 & n6144 ) | ( ~n5763 & n6144 ) ;
  assign n6146 = ( n2955 & n6140 ) | ( n2955 & n6145 ) | ( n6140 & n6145 ) ;
  assign n6147 = n2706 &  n6146 ;
  assign n6149 = ( n5787 & ~n5778 ) | ( n5787 & n5791 ) | ( ~n5778 & n5791 ) ;
  assign n6148 = n5791 | n6032 ;
  assign n6151 = ( n5791 & ~n6149 ) | ( n5791 & n6148 ) | ( ~n6149 & n6148 ) ;
  assign n6150 = ( n6148 & ~n5787 ) | ( n6148 & n6149 ) | ( ~n5787 & n6149 ) ;
  assign n6152 = ( n5778 & ~n6151 ) | ( n5778 & n6150 ) | ( ~n6151 & n6150 ) ;
  assign n6153 = n2955 | n6125 ;
  assign n6154 = n6139 | n6153 ;
  assign n6155 = n6145 &  n6154 ;
  assign n6156 = n6133 | n6136 ;
  assign n6157 = ( n3211 & n6130 ) | ( n3211 & n6156 ) | ( n6130 & n6156 ) ;
  assign n6158 = n2955 &  n6157 ;
  assign n6159 = n2706 | n6158 ;
  assign n6160 = n6155 | n6159 ;
  assign n6161 = n6152 &  n6160 ;
  assign n6162 = n6147 | n6161 ;
  assign n6164 = ( n5780 & ~n5785 ) | ( n5780 & n6032 ) | ( ~n5785 & n6032 ) ;
  assign n6163 = ~n5793 & n6032 ;
  assign n6165 = ( n6032 & ~n6164 ) | ( n6032 & n6163 ) | ( ~n6164 & n6163 ) ;
  assign n6166 = ( n6163 & ~n5780 ) | ( n6163 & n6164 ) | ( ~n5780 & n6164 ) ;
  assign n6167 = ( n5785 & ~n6165 ) | ( n5785 & n6166 ) | ( ~n6165 & n6166 ) ;
  assign n6168 = ( n2472 & n6162 ) | ( n2472 & n6167 ) | ( n6162 & n6167 ) ;
  assign n6169 = n2245 &  n6168 ;
  assign n6171 = ( n5809 & ~n5800 ) | ( n5809 & n5813 ) | ( ~n5800 & n5813 ) ;
  assign n6170 = n5813 | n6032 ;
  assign n6173 = ( n5813 & ~n6171 ) | ( n5813 & n6170 ) | ( ~n6171 & n6170 ) ;
  assign n6172 = ( n6170 & ~n5809 ) | ( n6170 & n6171 ) | ( ~n5809 & n6171 ) ;
  assign n6174 = ( n5800 & ~n6173 ) | ( n5800 & n6172 ) | ( ~n6173 & n6172 ) ;
  assign n6175 = n2472 | n6147 ;
  assign n6176 = n6161 | n6175 ;
  assign n6177 = n6167 &  n6176 ;
  assign n6178 = n6155 | n6158 ;
  assign n6179 = ( n2706 & n6152 ) | ( n2706 & n6178 ) | ( n6152 & n6178 ) ;
  assign n6180 = n2472 &  n6179 ;
  assign n6181 = n2245 | n6180 ;
  assign n6182 = n6177 | n6181 ;
  assign n6183 = n6174 &  n6182 ;
  assign n6184 = n6169 | n6183 ;
  assign n6185 = ~n5815 & n6032 ;
  assign n6186 = ( n5802 & n5807 ) | ( n5802 & n6032 ) | ( n5807 & n6032 ) ;
  assign n6188 = ( n6185 & ~n5802 ) | ( n6185 & n6186 ) | ( ~n5802 & n6186 ) ;
  assign n6187 = ( n6032 & ~n6186 ) | ( n6032 & n6185 ) | ( ~n6186 & n6185 ) ;
  assign n6189 = ( n5807 & ~n6188 ) | ( n5807 & n6187 ) | ( ~n6188 & n6187 ) ;
  assign n6190 = ( n6184 & ~n2033 ) | ( n6184 & n6189 ) | ( ~n2033 & n6189 ) ;
  assign n6191 = n1827 &  n6190 ;
  assign n6192 = n5835 | n6032 ;
  assign n6193 = ( n5822 & ~n5831 ) | ( n5822 & n5835 ) | ( ~n5831 & n5835 ) ;
  assign n6194 = ( n5831 & n6192 ) | ( n5831 & n6193 ) | ( n6192 & n6193 ) ;
  assign n6195 = ( n5835 & ~n6193 ) | ( n5835 & n6192 ) | ( ~n6193 & n6192 ) ;
  assign n6196 = ( n5822 & ~n6194 ) | ( n5822 & n6195 ) | ( ~n6194 & n6195 ) ;
  assign n6197 = ( n2033 & ~n6169 ) | ( n2033 & 1'b0 ) | ( ~n6169 & 1'b0 ) ;
  assign n6198 = ~n6183 & n6197 ;
  assign n6199 = ( n6189 & ~n6198 ) | ( n6189 & 1'b0 ) | ( ~n6198 & 1'b0 ) ;
  assign n6200 = n6177 | n6180 ;
  assign n6201 = ( n2245 & n6174 ) | ( n2245 & n6200 ) | ( n6174 & n6200 ) ;
  assign n6202 = ~n2033 & n6201 ;
  assign n6203 = n1827 | n6202 ;
  assign n6204 = n6199 | n6203 ;
  assign n6205 = n6196 &  n6204 ;
  assign n6206 = n6191 | n6205 ;
  assign n6207 = ~n5837 & n6032 ;
  assign n6208 = ( n5824 & ~n6207 ) | ( n5824 & n6032 ) | ( ~n6207 & n6032 ) ;
  assign n6209 = ( n5829 & ~n5824 ) | ( n5829 & n6208 ) | ( ~n5824 & n6208 ) ;
  assign n6210 = ( n5824 & ~n6208 ) | ( n5824 & n5829 ) | ( ~n6208 & n5829 ) ;
  assign n6211 = ( n6209 & ~n5829 ) | ( n6209 & n6210 ) | ( ~n5829 & n6210 ) ;
  assign n6212 = ( n1636 & ~n6206 ) | ( n1636 & n6211 ) | ( ~n6206 & n6211 ) ;
  assign n6213 = n1452 | n6212 ;
  assign n6214 = n5857 | n6032 ;
  assign n6215 = ( n5844 & ~n5857 ) | ( n5844 & n5853 ) | ( ~n5857 & n5853 ) ;
  assign n6217 = ( n5857 & n6214 ) | ( n5857 & n6215 ) | ( n6214 & n6215 ) ;
  assign n6216 = ( n5853 & ~n6215 ) | ( n5853 & n6214 ) | ( ~n6215 & n6214 ) ;
  assign n6218 = ( n5844 & ~n6217 ) | ( n5844 & n6216 ) | ( ~n6217 & n6216 ) ;
  assign n6219 = ( n1636 & ~n6191 ) | ( n1636 & 1'b0 ) | ( ~n6191 & 1'b0 ) ;
  assign n6220 = ~n6205 & n6219 ;
  assign n6221 = n6211 | n6220 ;
  assign n6222 = n6199 | n6202 ;
  assign n6223 = ( n1827 & n6196 ) | ( n1827 & n6222 ) | ( n6196 & n6222 ) ;
  assign n6224 = ~n1636 & n6223 ;
  assign n6225 = ( n1452 & ~n6224 ) | ( n1452 & 1'b0 ) | ( ~n6224 & 1'b0 ) ;
  assign n6226 = n6221 &  n6225 ;
  assign n6227 = ( n6218 & ~n6226 ) | ( n6218 & 1'b0 ) | ( ~n6226 & 1'b0 ) ;
  assign n6228 = ( n6213 & ~n6227 ) | ( n6213 & 1'b0 ) | ( ~n6227 & 1'b0 ) ;
  assign n6229 = n5846 | n6032 ;
  assign n6230 = ( n5851 & ~n5846 ) | ( n5851 & n5859 ) | ( ~n5846 & n5859 ) ;
  assign n6232 = ( n5846 & n6229 ) | ( n5846 & n6230 ) | ( n6229 & n6230 ) ;
  assign n6231 = ( n5859 & ~n6230 ) | ( n5859 & n6229 ) | ( ~n6230 & n6229 ) ;
  assign n6233 = ( n5851 & ~n6232 ) | ( n5851 & n6231 ) | ( ~n6232 & n6231 ) ;
  assign n6234 = ( n6228 & ~n1283 ) | ( n6228 & n6233 ) | ( ~n1283 & n6233 ) ;
  assign n6235 = n1122 | n6234 ;
  assign n6236 = n5879 | n6032 ;
  assign n6237 = ( n5866 & ~n5875 ) | ( n5866 & n5879 ) | ( ~n5875 & n5879 ) ;
  assign n6238 = ( n5875 & n6236 ) | ( n5875 & n6237 ) | ( n6236 & n6237 ) ;
  assign n6239 = ( n5879 & ~n6237 ) | ( n5879 & n6236 ) | ( ~n6237 & n6236 ) ;
  assign n6240 = ( n5866 & ~n6238 ) | ( n5866 & n6239 ) | ( ~n6238 & n6239 ) ;
  assign n6241 = ~n1283 & n6213 ;
  assign n6242 = ~n6227 & n6241 ;
  assign n6243 = n6233 | n6242 ;
  assign n6244 = ( n6221 & ~n6224 ) | ( n6221 & 1'b0 ) | ( ~n6224 & 1'b0 ) ;
  assign n6245 = ( n1452 & ~n6218 ) | ( n1452 & n6244 ) | ( ~n6218 & n6244 ) ;
  assign n6246 = ( n1283 & ~n6245 ) | ( n1283 & 1'b0 ) | ( ~n6245 & 1'b0 ) ;
  assign n6247 = ( n1122 & ~n6246 ) | ( n1122 & 1'b0 ) | ( ~n6246 & 1'b0 ) ;
  assign n6248 = n6243 &  n6247 ;
  assign n6249 = n6240 | n6248 ;
  assign n6250 = n6235 &  n6249 ;
  assign n6256 = ( n976 & ~n6255 ) | ( n976 & n6250 ) | ( ~n6255 & n6250 ) ;
  assign n6257 = ( n837 & ~n6256 ) | ( n837 & 1'b0 ) | ( ~n6256 & 1'b0 ) ;
  assign n6258 = ( n5901 & ~n6032 ) | ( n5901 & 1'b0 ) | ( ~n6032 & 1'b0 ) ;
  assign n6259 = ( n5888 & n5897 ) | ( n5888 & n5901 ) | ( n5897 & n5901 ) ;
  assign n6260 = ( n6258 & ~n5897 ) | ( n6258 & n6259 ) | ( ~n5897 & n6259 ) ;
  assign n6261 = ( n5901 & ~n6259 ) | ( n5901 & n6258 ) | ( ~n6259 & n6258 ) ;
  assign n6262 = ( n5888 & ~n6260 ) | ( n5888 & n6261 ) | ( ~n6260 & n6261 ) ;
  assign n6263 = n976 &  n6235 ;
  assign n6264 = n6249 &  n6263 ;
  assign n6265 = ( n6255 & ~n6264 ) | ( n6255 & 1'b0 ) | ( ~n6264 & 1'b0 ) ;
  assign n6266 = ( n6243 & ~n6246 ) | ( n6243 & 1'b0 ) | ( ~n6246 & 1'b0 ) ;
  assign n6267 = ( n1122 & n6240 ) | ( n1122 & n6266 ) | ( n6240 & n6266 ) ;
  assign n6268 = n976 | n6267 ;
  assign n6269 = ~n837 & n6268 ;
  assign n6270 = ~n6265 & n6269 ;
  assign n6271 = n6262 | n6270 ;
  assign n6272 = ~n6257 & n6271 ;
  assign n6273 = n5903 &  n6032 ;
  assign n6274 = ( n5890 & ~n6273 ) | ( n5890 & n6032 ) | ( ~n6273 & n6032 ) ;
  assign n6275 = ( n5895 & ~n5890 ) | ( n5895 & n6274 ) | ( ~n5890 & n6274 ) ;
  assign n6276 = ( n5890 & ~n6274 ) | ( n5890 & n5895 ) | ( ~n6274 & n5895 ) ;
  assign n6277 = ( n6275 & ~n5895 ) | ( n6275 & n6276 ) | ( ~n5895 & n6276 ) ;
  assign n6278 = ( n6272 & ~n713 ) | ( n6272 & n6277 ) | ( ~n713 & n6277 ) ;
  assign n6279 = ( n595 & ~n6278 ) | ( n595 & 1'b0 ) | ( ~n6278 & 1'b0 ) ;
  assign n6280 = n5923 | n6032 ;
  assign n6281 = ( n5910 & ~n5923 ) | ( n5910 & n5919 ) | ( ~n5923 & n5919 ) ;
  assign n6283 = ( n5923 & n6280 ) | ( n5923 & n6281 ) | ( n6280 & n6281 ) ;
  assign n6282 = ( n5919 & ~n6281 ) | ( n5919 & n6280 ) | ( ~n6281 & n6280 ) ;
  assign n6284 = ( n5910 & ~n6283 ) | ( n5910 & n6282 ) | ( ~n6283 & n6282 ) ;
  assign n6285 = n713 | n6257 ;
  assign n6286 = ( n6271 & ~n6285 ) | ( n6271 & 1'b0 ) | ( ~n6285 & 1'b0 ) ;
  assign n6287 = n6277 | n6286 ;
  assign n6288 = ~n6265 & n6268 ;
  assign n6289 = ( n6262 & ~n837 ) | ( n6262 & n6288 ) | ( ~n837 & n6288 ) ;
  assign n6290 = ( n713 & ~n6289 ) | ( n713 & 1'b0 ) | ( ~n6289 & 1'b0 ) ;
  assign n6291 = n595 | n6290 ;
  assign n6292 = ( n6287 & ~n6291 ) | ( n6287 & 1'b0 ) | ( ~n6291 & 1'b0 ) ;
  assign n6293 = ( n6284 & ~n6292 ) | ( n6284 & 1'b0 ) | ( ~n6292 & 1'b0 ) ;
  assign n6294 = n6279 | n6293 ;
  assign n6295 = n5912 | n6032 ;
  assign n6296 = ( n5912 & n5917 ) | ( n5912 & n5925 ) | ( n5917 & n5925 ) ;
  assign n6297 = ( n6295 & ~n5925 ) | ( n6295 & n6296 ) | ( ~n5925 & n6296 ) ;
  assign n6298 = ( n5912 & ~n6296 ) | ( n5912 & n6295 ) | ( ~n6296 & n6295 ) ;
  assign n6299 = ( n5917 & ~n6297 ) | ( n5917 & n6298 ) | ( ~n6297 & n6298 ) ;
  assign n6300 = ( n492 & n6294 ) | ( n492 & n6299 ) | ( n6294 & n6299 ) ;
  assign n6301 = n396 &  n6300 ;
  assign n6303 = ( n5941 & ~n5932 ) | ( n5941 & n5945 ) | ( ~n5932 & n5945 ) ;
  assign n6302 = n5945 | n6032 ;
  assign n6305 = ( n5945 & ~n6303 ) | ( n5945 & n6302 ) | ( ~n6303 & n6302 ) ;
  assign n6304 = ( n6302 & ~n5941 ) | ( n6302 & n6303 ) | ( ~n5941 & n6303 ) ;
  assign n6306 = ( n5932 & ~n6305 ) | ( n5932 & n6304 ) | ( ~n6305 & n6304 ) ;
  assign n6307 = n492 | n6279 ;
  assign n6308 = n6293 | n6307 ;
  assign n6309 = n6299 &  n6308 ;
  assign n6310 = ( n6287 & ~n6290 ) | ( n6287 & 1'b0 ) | ( ~n6290 & 1'b0 ) ;
  assign n6311 = ( n595 & ~n6310 ) | ( n595 & n6284 ) | ( ~n6310 & n6284 ) ;
  assign n6312 = n492 &  n6311 ;
  assign n6313 = n396 | n6312 ;
  assign n6314 = n6309 | n6313 ;
  assign n6315 = n6306 &  n6314 ;
  assign n6316 = n6301 | n6315 ;
  assign n6318 = ( n5934 & ~n5939 ) | ( n5934 & n5947 ) | ( ~n5939 & n5947 ) ;
  assign n6317 = n5934 | n6032 ;
  assign n6320 = ( n5934 & ~n6318 ) | ( n5934 & n6317 ) | ( ~n6318 & n6317 ) ;
  assign n6319 = ( n6317 & ~n5947 ) | ( n6317 & n6318 ) | ( ~n5947 & n6318 ) ;
  assign n6321 = ( n5939 & ~n6320 ) | ( n5939 & n6319 ) | ( ~n6320 & n6319 ) ;
  assign n6322 = ( n315 & n6316 ) | ( n315 & n6321 ) | ( n6316 & n6321 ) ;
  assign n6323 = n240 &  n6322 ;
  assign n6324 = n5967 | n6032 ;
  assign n6325 = ( n5954 & n5963 ) | ( n5954 & n5967 ) | ( n5963 & n5967 ) ;
  assign n6326 = ( n6324 & ~n5963 ) | ( n6324 & n6325 ) | ( ~n5963 & n6325 ) ;
  assign n6327 = ( n5967 & ~n6325 ) | ( n5967 & n6324 ) | ( ~n6325 & n6324 ) ;
  assign n6328 = ( n5954 & ~n6326 ) | ( n5954 & n6327 ) | ( ~n6326 & n6327 ) ;
  assign n6329 = n315 | n6301 ;
  assign n6330 = n6315 | n6329 ;
  assign n6331 = n6321 &  n6330 ;
  assign n6332 = n6309 | n6312 ;
  assign n6333 = ( n396 & n6306 ) | ( n396 & n6332 ) | ( n6306 & n6332 ) ;
  assign n6334 = n315 &  n6333 ;
  assign n6335 = n240 | n6334 ;
  assign n6336 = n6331 | n6335 ;
  assign n6337 = n6328 &  n6336 ;
  assign n6338 = n6323 | n6337 ;
  assign n6340 = ( n5956 & ~n5961 ) | ( n5956 & n6032 ) | ( ~n5961 & n6032 ) ;
  assign n6339 = ~n5969 & n6032 ;
  assign n6341 = ( n6032 & ~n6340 ) | ( n6032 & n6339 ) | ( ~n6340 & n6339 ) ;
  assign n6342 = ( n6339 & ~n5956 ) | ( n6339 & n6340 ) | ( ~n5956 & n6340 ) ;
  assign n6343 = ( n5961 & ~n6341 ) | ( n5961 & n6342 ) | ( ~n6341 & n6342 ) ;
  assign n6344 = ( n181 & n6338 ) | ( n181 & n6343 ) | ( n6338 & n6343 ) ;
  assign n6345 = ~n145 & n6344 ;
  assign n6346 = n5989 | n6032 ;
  assign n6347 = ( n5976 & n5985 ) | ( n5976 & n5989 ) | ( n5985 & n5989 ) ;
  assign n6348 = ( n6346 & ~n5985 ) | ( n6346 & n6347 ) | ( ~n5985 & n6347 ) ;
  assign n6349 = ( n5989 & ~n6347 ) | ( n5989 & n6346 ) | ( ~n6347 & n6346 ) ;
  assign n6350 = ( n5976 & ~n6348 ) | ( n5976 & n6349 ) | ( ~n6348 & n6349 ) ;
  assign n6351 = n181 | n6323 ;
  assign n6352 = n6337 | n6351 ;
  assign n6353 = n6343 &  n6352 ;
  assign n6354 = n6331 | n6334 ;
  assign n6355 = ( n240 & n6328 ) | ( n240 & n6354 ) | ( n6328 & n6354 ) ;
  assign n6356 = n181 &  n6355 ;
  assign n6357 = ( n145 & ~n6356 ) | ( n145 & 1'b0 ) | ( ~n6356 & 1'b0 ) ;
  assign n6358 = ~n6353 & n6357 ;
  assign n6359 = n6350 | n6358 ;
  assign n6360 = ~n6345 & n6359 ;
  assign n6361 = n5991 &  n6032 ;
  assign n6362 = ( n5978 & ~n6361 ) | ( n5978 & n6032 ) | ( ~n6361 & n6032 ) ;
  assign n6363 = ( n5978 & ~n6362 ) | ( n5978 & n5983 ) | ( ~n6362 & n5983 ) ;
  assign n6364 = ( n5983 & ~n5978 ) | ( n5983 & n6362 ) | ( ~n5978 & n6362 ) ;
  assign n6365 = ( n6363 & ~n5983 ) | ( n6363 & n6364 ) | ( ~n5983 & n6364 ) ;
  assign n6366 = ( n150 & ~n6360 ) | ( n150 & n6365 ) | ( ~n6360 & n6365 ) ;
  assign n6367 = n5998 | n6017 ;
  assign n6368 = ( n6014 & ~n6032 ) | ( n6014 & n6367 ) | ( ~n6032 & n6367 ) ;
  assign n6369 = ( n6014 & ~n6368 ) | ( n6014 & 1'b0 ) | ( ~n6368 & 1'b0 ) ;
  assign n6370 = ( n6014 & ~n6017 ) | ( n6014 & 1'b0 ) | ( ~n6017 & 1'b0 ) ;
  assign n6371 = ~n6032 & n6370 ;
  assign n6372 = ( n5998 & ~n6370 ) | ( n5998 & n6371 ) | ( ~n6370 & n6371 ) ;
  assign n6373 = n6369 | n6372 ;
  assign n6374 = n5999 &  n6006 ;
  assign n6375 = ~n6032 & n6374 ;
  assign n6376 = ( n6020 & ~n6374 ) | ( n6020 & n6375 ) | ( ~n6374 & n6375 ) ;
  assign n6377 = n6373 &  n6376 ;
  assign n6378 = ~n6366 & n6377 ;
  assign n6379 = ( n133 & ~n6378 ) | ( n133 & n6377 ) | ( ~n6378 & n6377 ) ;
  assign n6380 = n150 | n6345 ;
  assign n6381 = ( n6359 & ~n6380 ) | ( n6359 & 1'b0 ) | ( ~n6380 & 1'b0 ) ;
  assign n6386 = n6381 &  n6365 ;
  assign n6382 = n6353 | n6356 ;
  assign n6383 = ( n145 & ~n6382 ) | ( n145 & n6350 ) | ( ~n6382 & n6350 ) ;
  assign n6384 = ( n150 & ~n6383 ) | ( n150 & 1'b0 ) | ( ~n6383 & 1'b0 ) ;
  assign n6385 = n6373 | n6384 ;
  assign n6387 = ( n6365 & ~n6386 ) | ( n6365 & n6385 ) | ( ~n6386 & n6385 ) ;
  assign n6389 = ( n133 & n5999 ) | ( n133 & n6006 ) | ( n5999 & n6006 ) ;
  assign n6388 = ( n5999 & ~n6032 ) | ( n5999 & n6006 ) | ( ~n6032 & n6006 ) ;
  assign n6390 = ( n6006 & ~n6388 ) | ( n6006 & 1'b0 ) | ( ~n6388 & 1'b0 ) ;
  assign n6391 = ( n6389 & ~n6006 ) | ( n6389 & n6390 ) | ( ~n6006 & n6390 ) ;
  assign n6392 = n6002 | n6029 ;
  assign n6393 = ( n6024 & ~n6005 ) | ( n6024 & n6392 ) | ( ~n6005 & n6392 ) ;
  assign n6394 = n6005 | n6393 ;
  assign n6395 = ( n6012 & ~n6020 ) | ( n6012 & n6394 ) | ( ~n6020 & n6394 ) ;
  assign n6396 = ( n6012 & ~n6395 ) | ( n6012 & 1'b0 ) | ( ~n6395 & 1'b0 ) ;
  assign n6397 = n6391 | n6396 ;
  assign n6398 = ( n6387 & ~n6397 ) | ( n6387 & 1'b0 ) | ( ~n6397 & 1'b0 ) ;
  assign n6399 = n6379 &  n6398 ;
  assign n6418 = n5673 | n6399 ;
  assign n6808 = x62 | n6399 ;
  assign n6809 = x63 &  n6808 ;
  assign n6810 = ( n6418 & ~n6809 ) | ( n6418 & 1'b0 ) | ( ~n6809 & 1'b0 ) ;
  assign n6402 = x60 | x61 ;
  assign n6403 = x62 | n6402 ;
  assign n6404 = ( x62 & ~n6399 ) | ( x62 & 1'b0 ) | ( ~n6399 & 1'b0 ) ;
  assign n6405 = ( n6032 & ~n6403 ) | ( n6032 & n6404 ) | ( ~n6403 & n6404 ) ;
  assign n6407 = ~x62 & n6402 ;
  assign n6408 = ( x62 & ~n6030 ) | ( x62 & n6407 ) | ( ~n6030 & n6407 ) ;
  assign n6409 = ( n6020 & ~n6012 ) | ( n6020 & n6408 ) | ( ~n6012 & n6408 ) ;
  assign n6410 = n6012 &  n6409 ;
  assign n6805 = ( x62 & ~n6410 ) | ( x62 & n6399 ) | ( ~n6410 & n6399 ) ;
  assign n6806 = ( x62 & ~n6805 ) | ( x62 & 1'b0 ) | ( ~n6805 & 1'b0 ) ;
  assign n6807 = ( n6405 & ~n6806 ) | ( n6405 & n6410 ) | ( ~n6806 & n6410 ) ;
  assign n6677 = ( n6292 & ~n6399 ) | ( n6292 & 1'b0 ) | ( ~n6399 & 1'b0 ) ;
  assign n6678 = ( n6284 & ~n6279 ) | ( n6284 & n6399 ) | ( ~n6279 & n6399 ) ;
  assign n6679 = ( n6677 & ~n6399 ) | ( n6677 & n6678 ) | ( ~n6399 & n6678 ) ;
  assign n6680 = ( n6279 & ~n6677 ) | ( n6279 & n6678 ) | ( ~n6677 & n6678 ) ;
  assign n6681 = ( n6679 & ~n6284 ) | ( n6679 & n6680 ) | ( ~n6284 & n6680 ) ;
  assign n6457 = ( n6072 & ~n6399 ) | ( n6072 & 1'b0 ) | ( ~n6399 & 1'b0 ) ;
  assign n6458 = ( n6399 & ~n6055 ) | ( n6399 & n6457 ) | ( ~n6055 & n6457 ) ;
  assign n6459 = ( n6055 & n6065 ) | ( n6055 & n6458 ) | ( n6065 & n6458 ) ;
  assign n6460 = ( n6055 & ~n6065 ) | ( n6055 & n6458 ) | ( ~n6065 & n6458 ) ;
  assign n6461 = ( n6065 & ~n6459 ) | ( n6065 & n6460 ) | ( ~n6459 & n6460 ) ;
  assign n6430 = ~x64 & n6032 ;
  assign n6431 = ~x65 & n6430 ;
  assign n6432 = ( x65 & ~n6430 ) | ( x65 & 1'b0 ) | ( ~n6430 & 1'b0 ) ;
  assign n6433 = n6431 | n6432 ;
  assign n6434 = ~n6033 & n6039 ;
  assign n6436 = ( n6034 & ~n6433 ) | ( n6034 & n6434 ) | ( ~n6433 & n6434 ) ;
  assign n6435 = n6034 &  n6399 ;
  assign n6438 = ( n6034 & ~n6436 ) | ( n6034 & n6435 ) | ( ~n6436 & n6435 ) ;
  assign n6437 = ( n6435 & ~n6434 ) | ( n6435 & n6436 ) | ( ~n6434 & n6436 ) ;
  assign n6439 = ( n6433 & ~n6438 ) | ( n6433 & n6437 ) | ( ~n6438 & n6437 ) ;
  assign n6411 = ( x63 & ~n6410 ) | ( x63 & n6399 ) | ( ~n6410 & n6399 ) ;
  assign n6406 = ( x62 & x63 ) | ( x62 & n6399 ) | ( x63 & n6399 ) ;
  assign n6412 = ( x62 & ~x63 ) | ( x62 & 1'b0 ) | ( ~x63 & 1'b0 ) ;
  assign n6413 = ( n6411 & ~n6406 ) | ( n6411 & n6412 ) | ( ~n6406 & n6412 ) ;
  assign n6414 = ( n6405 & ~n6413 ) | ( n6405 & 1'b0 ) | ( ~n6413 & 1'b0 ) ;
  assign n6415 = ( n6413 & ~n5672 ) | ( n6413 & n6414 ) | ( ~n5672 & n6414 ) ;
  assign n6416 = ( n5672 & ~n6405 ) | ( n5672 & 1'b0 ) | ( ~n6405 & 1'b0 ) ;
  assign n6417 = ~n6413 & n6416 ;
  assign n6419 = ( n6032 & ~n6396 ) | ( n6032 & 1'b0 ) | ( ~n6396 & 1'b0 ) ;
  assign n6420 = ( n6387 & ~n6419 ) | ( n6387 & n6391 ) | ( ~n6419 & n6391 ) ;
  assign n6421 = ( n6387 & ~n6420 ) | ( n6387 & 1'b0 ) | ( ~n6420 & 1'b0 ) ;
  assign n6422 = n6379 &  n6421 ;
  assign n6423 = n6418 | n6422 ;
  assign n6424 = ( x64 & ~n6423 ) | ( x64 & n6422 ) | ( ~n6423 & n6422 ) ;
  assign n6425 = x64 | n6422 ;
  assign n6426 = ( n6418 & ~n6425 ) | ( n6418 & 1'b0 ) | ( ~n6425 & 1'b0 ) ;
  assign n6427 = n6424 | n6426 ;
  assign n6428 = ~n6417 & n6427 ;
  assign n6429 = n6415 | n6428 ;
  assign n6440 = ( n5327 & ~n6439 ) | ( n5327 & n6429 ) | ( ~n6439 & n6429 ) ;
  assign n6441 = n4990 &  n6440 ;
  assign n6442 = ~n6067 & n6070 ;
  assign n6443 = ( n6067 & ~n6442 ) | ( n6067 & n6053 ) | ( ~n6442 & n6053 ) ;
  assign n6444 = ( n6443 & ~n6399 ) | ( n6443 & n6442 ) | ( ~n6399 & n6442 ) ;
  assign n6445 = ( n6399 & ~n6067 ) | ( n6399 & n6443 ) | ( ~n6067 & n6443 ) ;
  assign n6446 = ( n6444 & ~n6053 ) | ( n6444 & n6445 ) | ( ~n6053 & n6445 ) ;
  assign n6447 = n5327 | n6415 ;
  assign n6448 = n6428 | n6447 ;
  assign n6449 = ~n6439 & n6448 ;
  assign n6450 = n6405 | n6413 ;
  assign n6451 = ( n6427 & ~n5672 ) | ( n6427 & n6450 ) | ( ~n5672 & n6450 ) ;
  assign n6452 = n5327 &  n6451 ;
  assign n6453 = n4990 | n6452 ;
  assign n6454 = n6449 | n6453 ;
  assign n6455 = n6446 &  n6454 ;
  assign n6456 = n6441 | n6455 ;
  assign n6462 = ( n4668 & ~n6461 ) | ( n4668 & n6456 ) | ( ~n6461 & n6456 ) ;
  assign n6463 = n4353 &  n6462 ;
  assign n6464 = ~n6092 & n6399 ;
  assign n6465 = ( n6079 & n6088 ) | ( n6079 & n6092 ) | ( n6088 & n6092 ) ;
  assign n6467 = ( n6464 & ~n6092 ) | ( n6464 & n6465 ) | ( ~n6092 & n6465 ) ;
  assign n6466 = ( n6088 & ~n6465 ) | ( n6088 & n6464 ) | ( ~n6465 & n6464 ) ;
  assign n6468 = ( n6079 & ~n6467 ) | ( n6079 & n6466 ) | ( ~n6467 & n6466 ) ;
  assign n6469 = n4668 | n6441 ;
  assign n6470 = n6455 | n6469 ;
  assign n6471 = ~n6461 & n6470 ;
  assign n6472 = n6449 | n6452 ;
  assign n6473 = ( n4990 & n6446 ) | ( n4990 & n6472 ) | ( n6446 & n6472 ) ;
  assign n6474 = n4668 &  n6473 ;
  assign n6475 = n4353 | n6474 ;
  assign n6476 = n6471 | n6475 ;
  assign n6477 = n6468 &  n6476 ;
  assign n6478 = n6463 | n6477 ;
  assign n6479 = n6094 | n6399 ;
  assign n6480 = ( n6086 & ~n6081 ) | ( n6086 & n6399 ) | ( ~n6081 & n6399 ) ;
  assign n6482 = ( n6081 & n6479 ) | ( n6081 & n6480 ) | ( n6479 & n6480 ) ;
  assign n6481 = ( n6399 & ~n6480 ) | ( n6399 & n6479 ) | ( ~n6480 & n6479 ) ;
  assign n6483 = ( n6086 & ~n6482 ) | ( n6086 & n6481 ) | ( ~n6482 & n6481 ) ;
  assign n6484 = ( n4053 & n6478 ) | ( n4053 & n6483 ) | ( n6478 & n6483 ) ;
  assign n6485 = n3760 &  n6484 ;
  assign n6487 = ( n6110 & ~n6101 ) | ( n6110 & n6114 ) | ( ~n6101 & n6114 ) ;
  assign n6486 = ~n6114 & n6399 ;
  assign n6488 = ( n6110 & ~n6487 ) | ( n6110 & n6486 ) | ( ~n6487 & n6486 ) ;
  assign n6489 = ( n6486 & ~n6114 ) | ( n6486 & n6487 ) | ( ~n6114 & n6487 ) ;
  assign n6490 = ( n6101 & ~n6488 ) | ( n6101 & n6489 ) | ( ~n6488 & n6489 ) ;
  assign n6491 = n4053 | n6463 ;
  assign n6492 = n6477 | n6491 ;
  assign n6493 = n6483 &  n6492 ;
  assign n6494 = n6471 | n6474 ;
  assign n6495 = ( n4353 & n6468 ) | ( n4353 & n6494 ) | ( n6468 & n6494 ) ;
  assign n6496 = n4053 &  n6495 ;
  assign n6497 = n3760 | n6496 ;
  assign n6498 = n6493 | n6497 ;
  assign n6499 = n6490 &  n6498 ;
  assign n6500 = n6485 | n6499 ;
  assign n6501 = ~n6103 & n6399 ;
  assign n6502 = ( n6103 & n6108 ) | ( n6103 & n6116 ) | ( n6108 & n6116 ) ;
  assign n6504 = ( n6501 & ~n6103 ) | ( n6501 & n6502 ) | ( ~n6103 & n6502 ) ;
  assign n6503 = ( n6116 & ~n6502 ) | ( n6116 & n6501 ) | ( ~n6502 & n6501 ) ;
  assign n6505 = ( n6108 & ~n6504 ) | ( n6108 & n6503 ) | ( ~n6504 & n6503 ) ;
  assign n6506 = ( n3482 & n6500 ) | ( n3482 & n6505 ) | ( n6500 & n6505 ) ;
  assign n6507 = n3211 &  n6506 ;
  assign n6508 = ~n6136 & n6399 ;
  assign n6509 = ( n6123 & n6132 ) | ( n6123 & n6136 ) | ( n6132 & n6136 ) ;
  assign n6511 = ( n6508 & ~n6136 ) | ( n6508 & n6509 ) | ( ~n6136 & n6509 ) ;
  assign n6510 = ( n6132 & ~n6509 ) | ( n6132 & n6508 ) | ( ~n6509 & n6508 ) ;
  assign n6512 = ( n6123 & ~n6511 ) | ( n6123 & n6510 ) | ( ~n6511 & n6510 ) ;
  assign n6513 = n3482 | n6485 ;
  assign n6514 = n6499 | n6513 ;
  assign n6515 = n6505 &  n6514 ;
  assign n6516 = n6493 | n6496 ;
  assign n6517 = ( n3760 & n6490 ) | ( n3760 & n6516 ) | ( n6490 & n6516 ) ;
  assign n6518 = n3482 &  n6517 ;
  assign n6519 = n3211 | n6518 ;
  assign n6520 = n6515 | n6519 ;
  assign n6521 = n6512 &  n6520 ;
  assign n6522 = n6507 | n6521 ;
  assign n6523 = n6138 | n6399 ;
  assign n6524 = ( n6125 & ~n6399 ) | ( n6125 & n6523 ) | ( ~n6399 & n6523 ) ;
  assign n6525 = ( n6125 & ~n6524 ) | ( n6125 & n6130 ) | ( ~n6524 & n6130 ) ;
  assign n6526 = ( n6130 & ~n6125 ) | ( n6130 & n6524 ) | ( ~n6125 & n6524 ) ;
  assign n6527 = ( n6525 & ~n6130 ) | ( n6525 & n6526 ) | ( ~n6130 & n6526 ) ;
  assign n6528 = ( n2955 & n6522 ) | ( n2955 & n6527 ) | ( n6522 & n6527 ) ;
  assign n6529 = n2706 &  n6528 ;
  assign n6530 = ~n6158 & n6399 ;
  assign n6531 = ( n6145 & n6154 ) | ( n6145 & n6158 ) | ( n6154 & n6158 ) ;
  assign n6533 = ( n6530 & ~n6158 ) | ( n6530 & n6531 ) | ( ~n6158 & n6531 ) ;
  assign n6532 = ( n6154 & ~n6531 ) | ( n6154 & n6530 ) | ( ~n6531 & n6530 ) ;
  assign n6534 = ( n6145 & ~n6533 ) | ( n6145 & n6532 ) | ( ~n6533 & n6532 ) ;
  assign n6535 = n2955 | n6507 ;
  assign n6536 = n6521 | n6535 ;
  assign n6537 = n6527 &  n6536 ;
  assign n6538 = n6515 | n6518 ;
  assign n6539 = ( n3211 & n6512 ) | ( n3211 & n6538 ) | ( n6512 & n6538 ) ;
  assign n6540 = n2955 &  n6539 ;
  assign n6541 = n2706 | n6540 ;
  assign n6542 = n6537 | n6541 ;
  assign n6543 = n6534 &  n6542 ;
  assign n6544 = n6529 | n6543 ;
  assign n6545 = n6160 | n6399 ;
  assign n6546 = ( n6147 & ~n6399 ) | ( n6147 & n6545 ) | ( ~n6399 & n6545 ) ;
  assign n6547 = ( n6147 & ~n6546 ) | ( n6147 & n6152 ) | ( ~n6546 & n6152 ) ;
  assign n6548 = ( n6152 & ~n6147 ) | ( n6152 & n6546 ) | ( ~n6147 & n6546 ) ;
  assign n6549 = ( n6547 & ~n6152 ) | ( n6547 & n6548 ) | ( ~n6152 & n6548 ) ;
  assign n6550 = ( n2472 & n6544 ) | ( n2472 & n6549 ) | ( n6544 & n6549 ) ;
  assign n6551 = n2245 &  n6550 ;
  assign n6552 = ~n6180 & n6399 ;
  assign n6553 = ( n6167 & n6176 ) | ( n6167 & n6180 ) | ( n6176 & n6180 ) ;
  assign n6555 = ( n6552 & ~n6180 ) | ( n6552 & n6553 ) | ( ~n6180 & n6553 ) ;
  assign n6554 = ( n6176 & ~n6553 ) | ( n6176 & n6552 ) | ( ~n6553 & n6552 ) ;
  assign n6556 = ( n6167 & ~n6555 ) | ( n6167 & n6554 ) | ( ~n6555 & n6554 ) ;
  assign n6557 = n2472 | n6529 ;
  assign n6558 = n6543 | n6557 ;
  assign n6559 = n6549 &  n6558 ;
  assign n6560 = n6537 | n6540 ;
  assign n6561 = ( n2706 & n6534 ) | ( n2706 & n6560 ) | ( n6534 & n6560 ) ;
  assign n6562 = n2472 &  n6561 ;
  assign n6563 = n2245 | n6562 ;
  assign n6564 = n6559 | n6563 ;
  assign n6565 = n6556 &  n6564 ;
  assign n6566 = n6551 | n6565 ;
  assign n6567 = n6182 | n6399 ;
  assign n6568 = ( n6169 & ~n6399 ) | ( n6169 & n6174 ) | ( ~n6399 & n6174 ) ;
  assign n6569 = ( n6399 & n6567 ) | ( n6399 & n6568 ) | ( n6567 & n6568 ) ;
  assign n6570 = ( n6169 & ~n6568 ) | ( n6169 & n6567 ) | ( ~n6568 & n6567 ) ;
  assign n6571 = ( n6174 & ~n6569 ) | ( n6174 & n6570 ) | ( ~n6569 & n6570 ) ;
  assign n6572 = ( n6566 & ~n2033 ) | ( n6566 & n6571 ) | ( ~n2033 & n6571 ) ;
  assign n6573 = n1827 &  n6572 ;
  assign n6574 = ~n6202 & n6399 ;
  assign n6575 = ( n6189 & ~n6198 ) | ( n6189 & n6202 ) | ( ~n6198 & n6202 ) ;
  assign n6576 = ( n6198 & ~n6574 ) | ( n6198 & n6575 ) | ( ~n6574 & n6575 ) ;
  assign n6577 = ( n6574 & ~n6202 ) | ( n6574 & n6575 ) | ( ~n6202 & n6575 ) ;
  assign n6578 = ( n6576 & ~n6189 ) | ( n6576 & n6577 ) | ( ~n6189 & n6577 ) ;
  assign n6579 = ( n2033 & ~n6551 ) | ( n2033 & 1'b0 ) | ( ~n6551 & 1'b0 ) ;
  assign n6580 = ~n6565 & n6579 ;
  assign n6581 = ( n6571 & ~n6580 ) | ( n6571 & 1'b0 ) | ( ~n6580 & 1'b0 ) ;
  assign n6582 = n6559 | n6562 ;
  assign n6583 = ( n2245 & n6556 ) | ( n2245 & n6582 ) | ( n6556 & n6582 ) ;
  assign n6584 = ~n2033 & n6583 ;
  assign n6585 = n1827 | n6584 ;
  assign n6586 = n6581 | n6585 ;
  assign n6587 = ~n6578 & n6586 ;
  assign n6588 = n6573 | n6587 ;
  assign n6589 = n6204 | n6399 ;
  assign n6590 = ( n6191 & ~n6399 ) | ( n6191 & n6589 ) | ( ~n6399 & n6589 ) ;
  assign n6591 = ( n6191 & ~n6590 ) | ( n6191 & n6196 ) | ( ~n6590 & n6196 ) ;
  assign n6592 = ( n6196 & ~n6191 ) | ( n6196 & n6590 ) | ( ~n6191 & n6590 ) ;
  assign n6593 = ( n6591 & ~n6196 ) | ( n6591 & n6592 ) | ( ~n6196 & n6592 ) ;
  assign n6594 = ( n6588 & ~n1636 ) | ( n6588 & n6593 ) | ( ~n1636 & n6593 ) ;
  assign n6595 = ~n1452 & n6594 ;
  assign n6596 = ~n6224 & n6399 ;
  assign n6597 = ( n6211 & ~n6224 ) | ( n6211 & n6220 ) | ( ~n6224 & n6220 ) ;
  assign n6598 = ( n6596 & ~n6220 ) | ( n6596 & n6597 ) | ( ~n6220 & n6597 ) ;
  assign n6599 = ( n6224 & ~n6596 ) | ( n6224 & n6597 ) | ( ~n6596 & n6597 ) ;
  assign n6600 = ( n6598 & ~n6211 ) | ( n6598 & n6599 ) | ( ~n6211 & n6599 ) ;
  assign n6601 = ( n1636 & ~n6573 ) | ( n1636 & 1'b0 ) | ( ~n6573 & 1'b0 ) ;
  assign n6602 = ~n6587 & n6601 ;
  assign n6603 = ( n6593 & ~n6602 ) | ( n6593 & 1'b0 ) | ( ~n6602 & 1'b0 ) ;
  assign n6604 = n6581 | n6584 ;
  assign n6605 = ( n1827 & ~n6578 ) | ( n1827 & n6604 ) | ( ~n6578 & n6604 ) ;
  assign n6606 = ~n1636 & n6605 ;
  assign n6607 = ( n1452 & ~n6606 ) | ( n1452 & 1'b0 ) | ( ~n6606 & 1'b0 ) ;
  assign n6608 = ~n6603 & n6607 ;
  assign n6609 = ( n6600 & ~n6608 ) | ( n6600 & 1'b0 ) | ( ~n6608 & 1'b0 ) ;
  assign n6610 = n6595 | n6609 ;
  assign n6611 = ~n6399 & n6226 ;
  assign n6612 = ( n6213 & n6611 ) | ( n6213 & n6399 ) | ( n6611 & n6399 ) ;
  assign n6613 = ( n6218 & ~n6213 ) | ( n6218 & n6612 ) | ( ~n6213 & n6612 ) ;
  assign n6614 = ( n6213 & ~n6612 ) | ( n6213 & n6218 ) | ( ~n6612 & n6218 ) ;
  assign n6615 = ( n6613 & ~n6218 ) | ( n6613 & n6614 ) | ( ~n6218 & n6614 ) ;
  assign n6616 = ( n1283 & n6610 ) | ( n1283 & n6615 ) | ( n6610 & n6615 ) ;
  assign n6617 = ~n1122 & n6616 ;
  assign n6618 = ~n6246 & n6399 ;
  assign n6619 = ( n6233 & ~n6242 ) | ( n6233 & n6246 ) | ( ~n6242 & n6246 ) ;
  assign n6620 = ( n6242 & ~n6618 ) | ( n6242 & n6619 ) | ( ~n6618 & n6619 ) ;
  assign n6621 = ( n6618 & ~n6246 ) | ( n6618 & n6619 ) | ( ~n6246 & n6619 ) ;
  assign n6622 = ( n6620 & ~n6233 ) | ( n6620 & n6621 ) | ( ~n6233 & n6621 ) ;
  assign n6623 = n1283 | n6595 ;
  assign n6624 = n6609 | n6623 ;
  assign n6625 = n6615 &  n6624 ;
  assign n6626 = n6603 | n6606 ;
  assign n6627 = ( n6600 & ~n1452 ) | ( n6600 & n6626 ) | ( ~n1452 & n6626 ) ;
  assign n6628 = n1283 &  n6627 ;
  assign n6629 = ( n1122 & ~n6628 ) | ( n1122 & 1'b0 ) | ( ~n6628 & 1'b0 ) ;
  assign n6630 = ~n6625 & n6629 ;
  assign n6631 = ( n6622 & ~n6630 ) | ( n6622 & 1'b0 ) | ( ~n6630 & 1'b0 ) ;
  assign n6632 = n6617 | n6631 ;
  assign n6633 = n6235 &  n6399 ;
  assign n6634 = ( n6235 & n6240 ) | ( n6235 & n6248 ) | ( n6240 & n6248 ) ;
  assign n6635 = ( n6633 & ~n6248 ) | ( n6633 & n6634 ) | ( ~n6248 & n6634 ) ;
  assign n6636 = ( n6235 & ~n6634 ) | ( n6235 & n6633 ) | ( ~n6634 & n6633 ) ;
  assign n6637 = ( n6240 & ~n6635 ) | ( n6240 & n6636 ) | ( ~n6635 & n6636 ) ;
  assign n6638 = ( n976 & ~n6632 ) | ( n976 & n6637 ) | ( ~n6632 & n6637 ) ;
  assign n6639 = ( n837 & ~n6638 ) | ( n837 & 1'b0 ) | ( ~n6638 & 1'b0 ) ;
  assign n6640 = n6268 &  n6399 ;
  assign n6641 = ( n6255 & n6264 ) | ( n6255 & n6268 ) | ( n6264 & n6268 ) ;
  assign n6642 = ( n6640 & ~n6264 ) | ( n6640 & n6641 ) | ( ~n6264 & n6641 ) ;
  assign n6643 = ( n6268 & ~n6641 ) | ( n6268 & n6640 ) | ( ~n6641 & n6640 ) ;
  assign n6644 = ( n6255 & ~n6642 ) | ( n6255 & n6643 ) | ( ~n6642 & n6643 ) ;
  assign n6645 = ( n976 & ~n6617 ) | ( n976 & 1'b0 ) | ( ~n6617 & 1'b0 ) ;
  assign n6646 = ~n6631 & n6645 ;
  assign n6647 = n6637 | n6646 ;
  assign n6648 = n6625 | n6628 ;
  assign n6649 = ( n6622 & ~n1122 ) | ( n6622 & n6648 ) | ( ~n1122 & n6648 ) ;
  assign n6650 = ~n976 & n6649 ;
  assign n6651 = n837 | n6650 ;
  assign n6652 = ( n6647 & ~n6651 ) | ( n6647 & 1'b0 ) | ( ~n6651 & 1'b0 ) ;
  assign n6653 = ( n6644 & ~n6652 ) | ( n6644 & 1'b0 ) | ( ~n6652 & 1'b0 ) ;
  assign n6654 = n6639 | n6653 ;
  assign n6655 = ~n6257 & n6399 ;
  assign n6656 = ( n6257 & ~n6270 ) | ( n6257 & n6262 ) | ( ~n6270 & n6262 ) ;
  assign n6657 = ( n6270 & ~n6655 ) | ( n6270 & n6656 ) | ( ~n6655 & n6656 ) ;
  assign n6658 = ( n6655 & ~n6257 ) | ( n6655 & n6656 ) | ( ~n6257 & n6656 ) ;
  assign n6659 = ( n6657 & ~n6262 ) | ( n6657 & n6658 ) | ( ~n6262 & n6658 ) ;
  assign n6660 = ( n713 & n6654 ) | ( n713 & n6659 ) | ( n6654 & n6659 ) ;
  assign n6661 = n595 &  n6660 ;
  assign n6662 = ~n6290 & n6399 ;
  assign n6663 = ( n6277 & ~n6290 ) | ( n6277 & n6286 ) | ( ~n6290 & n6286 ) ;
  assign n6664 = ( n6662 & ~n6286 ) | ( n6662 & n6663 ) | ( ~n6286 & n6663 ) ;
  assign n6665 = ( n6290 & ~n6662 ) | ( n6290 & n6663 ) | ( ~n6662 & n6663 ) ;
  assign n6666 = ( n6664 & ~n6277 ) | ( n6664 & n6665 ) | ( ~n6277 & n6665 ) ;
  assign n6667 = n713 | n6639 ;
  assign n6668 = n6653 | n6667 ;
  assign n6669 = n6659 &  n6668 ;
  assign n6670 = ( n6647 & ~n6650 ) | ( n6647 & 1'b0 ) | ( ~n6650 & 1'b0 ) ;
  assign n6671 = ( n837 & ~n6670 ) | ( n837 & n6644 ) | ( ~n6670 & n6644 ) ;
  assign n6672 = n713 &  n6671 ;
  assign n6673 = n595 | n6672 ;
  assign n6674 = n6669 | n6673 ;
  assign n6675 = n6666 &  n6674 ;
  assign n6676 = n6661 | n6675 ;
  assign n6682 = ( n492 & ~n6681 ) | ( n492 & n6676 ) | ( ~n6681 & n6676 ) ;
  assign n6683 = n396 &  n6682 ;
  assign n6685 = ( n6308 & ~n6299 ) | ( n6308 & n6312 ) | ( ~n6299 & n6312 ) ;
  assign n6684 = ~n6312 & n6399 ;
  assign n6686 = ( n6308 & ~n6685 ) | ( n6308 & n6684 ) | ( ~n6685 & n6684 ) ;
  assign n6687 = ( n6684 & ~n6312 ) | ( n6684 & n6685 ) | ( ~n6312 & n6685 ) ;
  assign n6688 = ( n6299 & ~n6686 ) | ( n6299 & n6687 ) | ( ~n6686 & n6687 ) ;
  assign n6689 = n492 | n6661 ;
  assign n6690 = n6675 | n6689 ;
  assign n6691 = ~n6681 & n6690 ;
  assign n6692 = n6669 | n6672 ;
  assign n6693 = ( n595 & n6666 ) | ( n595 & n6692 ) | ( n6666 & n6692 ) ;
  assign n6694 = n492 &  n6693 ;
  assign n6695 = n396 | n6694 ;
  assign n6696 = n6691 | n6695 ;
  assign n6697 = n6688 &  n6696 ;
  assign n6698 = n6683 | n6697 ;
  assign n6699 = ~n6301 & n6399 ;
  assign n6700 = ( n6301 & n6306 ) | ( n6301 & n6314 ) | ( n6306 & n6314 ) ;
  assign n6702 = ( n6699 & ~n6301 ) | ( n6699 & n6700 ) | ( ~n6301 & n6700 ) ;
  assign n6701 = ( n6314 & ~n6700 ) | ( n6314 & n6699 ) | ( ~n6700 & n6699 ) ;
  assign n6703 = ( n6306 & ~n6702 ) | ( n6306 & n6701 ) | ( ~n6702 & n6701 ) ;
  assign n6704 = ( n315 & n6698 ) | ( n315 & n6703 ) | ( n6698 & n6703 ) ;
  assign n6705 = n240 &  n6704 ;
  assign n6707 = ( n6330 & ~n6321 ) | ( n6330 & n6334 ) | ( ~n6321 & n6334 ) ;
  assign n6706 = ~n6334 & n6399 ;
  assign n6708 = ( n6330 & ~n6707 ) | ( n6330 & n6706 ) | ( ~n6707 & n6706 ) ;
  assign n6709 = ( n6706 & ~n6334 ) | ( n6706 & n6707 ) | ( ~n6334 & n6707 ) ;
  assign n6710 = ( n6321 & ~n6708 ) | ( n6321 & n6709 ) | ( ~n6708 & n6709 ) ;
  assign n6711 = n315 | n6683 ;
  assign n6712 = n6697 | n6711 ;
  assign n6713 = n6703 &  n6712 ;
  assign n6714 = n6691 | n6694 ;
  assign n6715 = ( n396 & n6688 ) | ( n396 & n6714 ) | ( n6688 & n6714 ) ;
  assign n6716 = n315 &  n6715 ;
  assign n6717 = n240 | n6716 ;
  assign n6718 = n6713 | n6717 ;
  assign n6719 = n6710 &  n6718 ;
  assign n6720 = n6705 | n6719 ;
  assign n6722 = ( n6323 & ~n6328 ) | ( n6323 & n6336 ) | ( ~n6328 & n6336 ) ;
  assign n6721 = ~n6323 & n6399 ;
  assign n6723 = ( n6336 & ~n6722 ) | ( n6336 & n6721 ) | ( ~n6722 & n6721 ) ;
  assign n6724 = ( n6721 & ~n6323 ) | ( n6721 & n6722 ) | ( ~n6323 & n6722 ) ;
  assign n6725 = ( n6328 & ~n6723 ) | ( n6328 & n6724 ) | ( ~n6723 & n6724 ) ;
  assign n6726 = ( n181 & n6720 ) | ( n181 & n6725 ) | ( n6720 & n6725 ) ;
  assign n6727 = ~n145 & n6726 ;
  assign n6728 = ~n6356 & n6399 ;
  assign n6729 = ( n6343 & n6352 ) | ( n6343 & n6356 ) | ( n6352 & n6356 ) ;
  assign n6731 = ( n6728 & ~n6356 ) | ( n6728 & n6729 ) | ( ~n6356 & n6729 ) ;
  assign n6730 = ( n6352 & ~n6729 ) | ( n6352 & n6728 ) | ( ~n6729 & n6728 ) ;
  assign n6732 = ( n6343 & ~n6731 ) | ( n6343 & n6730 ) | ( ~n6731 & n6730 ) ;
  assign n6733 = n181 | n6705 ;
  assign n6734 = n6719 | n6733 ;
  assign n6735 = n6725 &  n6734 ;
  assign n6736 = n6713 | n6716 ;
  assign n6737 = ( n240 & n6710 ) | ( n240 & n6736 ) | ( n6710 & n6736 ) ;
  assign n6738 = n181 &  n6737 ;
  assign n6739 = ( n145 & ~n6738 ) | ( n145 & 1'b0 ) | ( ~n6738 & 1'b0 ) ;
  assign n6740 = ~n6735 & n6739 ;
  assign n6741 = ( n6732 & ~n6740 ) | ( n6732 & 1'b0 ) | ( ~n6740 & 1'b0 ) ;
  assign n6742 = n6727 | n6741 ;
  assign n6743 = ~n6345 & n6399 ;
  assign n6744 = ( n6345 & ~n6358 ) | ( n6345 & n6350 ) | ( ~n6358 & n6350 ) ;
  assign n6745 = ( n6358 & ~n6743 ) | ( n6358 & n6744 ) | ( ~n6743 & n6744 ) ;
  assign n6746 = ( n6743 & ~n6345 ) | ( n6743 & n6744 ) | ( ~n6345 & n6744 ) ;
  assign n6747 = ( n6745 & ~n6350 ) | ( n6745 & n6746 ) | ( ~n6350 & n6746 ) ;
  assign n6748 = ( n150 & n6742 ) | ( n150 & n6747 ) | ( n6742 & n6747 ) ;
  assign n6749 = n6365 | n6381 ;
  assign n6750 = ( n6399 & ~n6384 ) | ( n6399 & n6749 ) | ( ~n6384 & n6749 ) ;
  assign n6751 = n6384 | n6750 ;
  assign n6752 = n6381 | n6384 ;
  assign n6753 = ~n6752 & n6399 ;
  assign n6754 = ( n6365 & n6753 ) | ( n6365 & n6752 ) | ( n6753 & n6752 ) ;
  assign n6755 = ( n6751 & ~n6754 ) | ( n6751 & 1'b0 ) | ( ~n6754 & 1'b0 ) ;
  assign n6756 = n6366 &  n6373 ;
  assign n6757 = n6399 &  n6756 ;
  assign n6758 = ( n6387 & ~n6756 ) | ( n6387 & n6757 ) | ( ~n6756 & n6757 ) ;
  assign n6759 = ~n6755 & n6758 ;
  assign n6760 = ~n6748 & n6759 ;
  assign n6761 = ( n133 & ~n6760 ) | ( n133 & n6759 ) | ( ~n6760 & n6759 ) ;
  assign n6764 = n6735 | n6738 ;
  assign n6765 = ( n6732 & ~n145 ) | ( n6732 & n6764 ) | ( ~n145 & n6764 ) ;
  assign n6766 = n150 &  n6765 ;
  assign n6767 = ( n6755 & ~n6766 ) | ( n6755 & 1'b0 ) | ( ~n6766 & 1'b0 ) ;
  assign n6762 = n150 | n6727 ;
  assign n6763 = n6741 | n6762 ;
  assign n6768 = ( n6747 & ~n6763 ) | ( n6747 & 1'b0 ) | ( ~n6763 & 1'b0 ) ;
  assign n6769 = ( n6767 & ~n6747 ) | ( n6767 & n6768 ) | ( ~n6747 & n6768 ) ;
  assign n6771 = ( n133 & n6366 ) | ( n133 & n6373 ) | ( n6366 & n6373 ) ;
  assign n6770 = ( n6366 & n6373 ) | ( n6366 & n6399 ) | ( n6373 & n6399 ) ;
  assign n6772 = ( n6373 & ~n6770 ) | ( n6373 & 1'b0 ) | ( ~n6770 & 1'b0 ) ;
  assign n6773 = ( n6771 & ~n6373 ) | ( n6771 & n6772 ) | ( ~n6373 & n6772 ) ;
  assign n6774 = n6369 | n6396 ;
  assign n6775 = ( n6391 & ~n6372 ) | ( n6391 & n6774 ) | ( ~n6372 & n6774 ) ;
  assign n6776 = n6372 | n6775 ;
  assign n6777 = ( n6379 & ~n6387 ) | ( n6379 & n6776 ) | ( ~n6387 & n6776 ) ;
  assign n6778 = ( n6379 & ~n6777 ) | ( n6379 & 1'b0 ) | ( ~n6777 & 1'b0 ) ;
  assign n6779 = n6773 | n6778 ;
  assign n6780 = n6769 | n6779 ;
  assign n6781 = ~n6761 |  n6780 ;
  assign n6811 = ( n6781 & n6807 ) | ( n6781 & n6810 ) | ( n6807 & n6810 ) ;
  assign n6812 = ~n6807 & n6811 ;
  assign n6813 = ( n6781 & ~n6811 ) | ( n6781 & 1'b0 ) | ( ~n6811 & 1'b0 ) ;
  assign n6814 = ( n6810 & ~n6812 ) | ( n6810 & n6813 ) | ( ~n6812 & n6813 ) ;
  assign n6782 = x60 &  n6781 ;
  assign n6400 = x58 | x59 ;
  assign n6401 = x60 | n6400 ;
  assign n6783 = ( n6399 & ~n6782 ) | ( n6399 & n6401 ) | ( ~n6782 & n6401 ) ;
  assign n6784 = ( x60 & ~n6781 ) | ( x60 & x61 ) | ( ~n6781 & x61 ) ;
  assign n6790 = ( x60 & ~x61 ) | ( x60 & 1'b0 ) | ( ~x61 & 1'b0 ) ;
  assign n6785 = ~x60 & n6400 ;
  assign n6786 = ( x60 & ~n6397 ) | ( x60 & n6785 ) | ( ~n6397 & n6785 ) ;
  assign n6787 = ( n6387 & ~n6379 ) | ( n6387 & n6786 ) | ( ~n6379 & n6786 ) ;
  assign n6788 = n6379 &  n6787 ;
  assign n6789 = ( n6781 & ~x61 ) | ( n6781 & n6788 ) | ( ~x61 & n6788 ) ;
  assign n6791 = ( n6784 & ~n6790 ) | ( n6784 & n6789 ) | ( ~n6790 & n6789 ) ;
  assign n6792 = n6783 &  n6791 ;
  assign n6794 = n6399 | n6778 ;
  assign n6795 = ( n6773 & ~n6769 ) | ( n6773 & n6794 ) | ( ~n6769 & n6794 ) ;
  assign n6796 = n6769 | n6795 ;
  assign n6797 = ( n6761 & ~n6796 ) | ( n6761 & 1'b0 ) | ( ~n6796 & 1'b0 ) ;
  assign n6793 = ~n6402 & n6781 ;
  assign n6798 = ( n6793 & ~n6797 ) | ( n6793 & 1'b0 ) | ( ~n6797 & 1'b0 ) ;
  assign n6799 = ( x62 & n6797 ) | ( x62 & n6798 ) | ( n6797 & n6798 ) ;
  assign n6800 = x62 | n6797 ;
  assign n6801 = n6793 | n6800 ;
  assign n6802 = ~n6799 & n6801 ;
  assign n6803 = ( n6792 & ~n6032 ) | ( n6792 & n6802 ) | ( ~n6032 & n6802 ) ;
  assign n6804 = n5672 | n6803 ;
  assign n6815 = ~n6032 & n6783 ;
  assign n6816 = n6791 &  n6815 ;
  assign n6817 = n6802 | n6816 ;
  assign n6818 = ~n6783 & n6791 ;
  assign n6819 = ( n6032 & ~n6791 ) | ( n6032 & n6818 ) | ( ~n6791 & n6818 ) ;
  assign n6820 = ( n5672 & ~n6819 ) | ( n5672 & 1'b0 ) | ( ~n6819 & 1'b0 ) ;
  assign n6821 = n6817 &  n6820 ;
  assign n7228 = ( n6804 & ~n6814 ) | ( n6804 & n6821 ) | ( ~n6814 & n6821 ) ;
  assign n6822 = ( n6814 & ~n6821 ) | ( n6814 & 1'b0 ) | ( ~n6821 & 1'b0 ) ;
  assign n6823 = ( n6804 & ~n6822 ) | ( n6804 & 1'b0 ) | ( ~n6822 & 1'b0 ) ;
  assign n6824 = ( n6415 & ~n6417 ) | ( n6415 & 1'b0 ) | ( ~n6417 & 1'b0 ) ;
  assign n6825 = ( n6417 & ~n6824 ) | ( n6417 & n6781 ) | ( ~n6824 & n6781 ) ;
  assign n6826 = ( n6417 & ~n6825 ) | ( n6417 & n6427 ) | ( ~n6825 & n6427 ) ;
  assign n6827 = ( n6427 & ~n6417 ) | ( n6427 & n6825 ) | ( ~n6417 & n6825 ) ;
  assign n6828 = ( n6826 & ~n6427 ) | ( n6826 & n6827 ) | ( ~n6427 & n6827 ) ;
  assign n6829 = ( n5327 & ~n6823 ) | ( n5327 & n6828 ) | ( ~n6823 & n6828 ) ;
  assign n6830 = n4990 &  n6829 ;
  assign n6831 = ~n5327 & n6804 ;
  assign n6832 = ~n6822 & n6831 ;
  assign n6833 = ( n6828 & ~n6832 ) | ( n6828 & 1'b0 ) | ( ~n6832 & 1'b0 ) ;
  assign n6834 = ( n6817 & ~n6819 ) | ( n6817 & 1'b0 ) | ( ~n6819 & 1'b0 ) ;
  assign n6835 = ( n5672 & ~n6814 ) | ( n5672 & n6834 ) | ( ~n6814 & n6834 ) ;
  assign n6836 = ( n5327 & ~n6835 ) | ( n5327 & 1'b0 ) | ( ~n6835 & 1'b0 ) ;
  assign n6837 = n4990 | n6836 ;
  assign n6838 = n6833 | n6837 ;
  assign n6839 = ( n6448 & ~n6439 ) | ( n6448 & n6452 ) | ( ~n6439 & n6452 ) ;
  assign n6840 = ( n6452 & ~n6839 ) | ( n6452 & n6781 ) | ( ~n6839 & n6781 ) ;
  assign n6841 = ( n6781 & ~n6448 ) | ( n6781 & n6839 ) | ( ~n6448 & n6839 ) ;
  assign n6842 = ( n6439 & ~n6840 ) | ( n6439 & n6841 ) | ( ~n6840 & n6841 ) ;
  assign n6843 = ( n6838 & ~n6842 ) | ( n6838 & 1'b0 ) | ( ~n6842 & 1'b0 ) ;
  assign n6844 = n6830 | n6843 ;
  assign n6846 = ( n6441 & ~n6446 ) | ( n6441 & n6781 ) | ( ~n6446 & n6781 ) ;
  assign n6845 = ~n6454 & n6781 ;
  assign n6847 = ( n6781 & ~n6846 ) | ( n6781 & n6845 ) | ( ~n6846 & n6845 ) ;
  assign n6848 = ( n6845 & ~n6441 ) | ( n6845 & n6846 ) | ( ~n6441 & n6846 ) ;
  assign n6849 = ( n6446 & ~n6847 ) | ( n6446 & n6848 ) | ( ~n6847 & n6848 ) ;
  assign n6850 = ( n4668 & n6844 ) | ( n4668 & n6849 ) | ( n6844 & n6849 ) ;
  assign n6851 = n4353 &  n6850 ;
  assign n6853 = ( n6470 & ~n6461 ) | ( n6470 & n6474 ) | ( ~n6461 & n6474 ) ;
  assign n6852 = n6474 | n6781 ;
  assign n6855 = ( n6474 & ~n6853 ) | ( n6474 & n6852 ) | ( ~n6853 & n6852 ) ;
  assign n6854 = ( n6852 & ~n6470 ) | ( n6852 & n6853 ) | ( ~n6470 & n6853 ) ;
  assign n6856 = ( n6461 & ~n6855 ) | ( n6461 & n6854 ) | ( ~n6855 & n6854 ) ;
  assign n6857 = n4668 | n6830 ;
  assign n6858 = n6843 | n6857 ;
  assign n6859 = n6849 &  n6858 ;
  assign n6860 = n6833 | n6836 ;
  assign n6861 = ( n4990 & ~n6842 ) | ( n4990 & n6860 ) | ( ~n6842 & n6860 ) ;
  assign n6862 = n4668 &  n6861 ;
  assign n6863 = n4353 | n6862 ;
  assign n6864 = n6859 | n6863 ;
  assign n6865 = ~n6856 & n6864 ;
  assign n6866 = n6851 | n6865 ;
  assign n6867 = ~n6476 & n6781 ;
  assign n6868 = ( n6463 & n6468 ) | ( n6463 & n6781 ) | ( n6468 & n6781 ) ;
  assign n6870 = ( n6867 & ~n6463 ) | ( n6867 & n6868 ) | ( ~n6463 & n6868 ) ;
  assign n6869 = ( n6781 & ~n6868 ) | ( n6781 & n6867 ) | ( ~n6868 & n6867 ) ;
  assign n6871 = ( n6468 & ~n6870 ) | ( n6468 & n6869 ) | ( ~n6870 & n6869 ) ;
  assign n6872 = ( n4053 & n6866 ) | ( n4053 & n6871 ) | ( n6866 & n6871 ) ;
  assign n6873 = n3760 &  n6872 ;
  assign n6874 = n6496 | n6781 ;
  assign n6875 = ( n6483 & n6492 ) | ( n6483 & n6496 ) | ( n6492 & n6496 ) ;
  assign n6876 = ( n6874 & ~n6492 ) | ( n6874 & n6875 ) | ( ~n6492 & n6875 ) ;
  assign n6877 = ( n6496 & ~n6875 ) | ( n6496 & n6874 ) | ( ~n6875 & n6874 ) ;
  assign n6878 = ( n6483 & ~n6876 ) | ( n6483 & n6877 ) | ( ~n6876 & n6877 ) ;
  assign n6879 = n4053 | n6851 ;
  assign n6880 = n6865 | n6879 ;
  assign n6881 = n6871 &  n6880 ;
  assign n6882 = n6859 | n6862 ;
  assign n6883 = ( n4353 & ~n6856 ) | ( n4353 & n6882 ) | ( ~n6856 & n6882 ) ;
  assign n6884 = n4053 &  n6883 ;
  assign n6885 = n3760 | n6884 ;
  assign n6886 = n6881 | n6885 ;
  assign n6887 = n6878 &  n6886 ;
  assign n6888 = n6873 | n6887 ;
  assign n6890 = ( n6485 & ~n6490 ) | ( n6485 & n6781 ) | ( ~n6490 & n6781 ) ;
  assign n6889 = ~n6498 & n6781 ;
  assign n6891 = ( n6781 & ~n6890 ) | ( n6781 & n6889 ) | ( ~n6890 & n6889 ) ;
  assign n6892 = ( n6889 & ~n6485 ) | ( n6889 & n6890 ) | ( ~n6485 & n6890 ) ;
  assign n6893 = ( n6490 & ~n6891 ) | ( n6490 & n6892 ) | ( ~n6891 & n6892 ) ;
  assign n6894 = ( n3482 & n6888 ) | ( n3482 & n6893 ) | ( n6888 & n6893 ) ;
  assign n6895 = n3211 &  n6894 ;
  assign n6897 = ( n6514 & ~n6505 ) | ( n6514 & n6518 ) | ( ~n6505 & n6518 ) ;
  assign n6896 = n6518 | n6781 ;
  assign n6899 = ( n6518 & ~n6897 ) | ( n6518 & n6896 ) | ( ~n6897 & n6896 ) ;
  assign n6898 = ( n6896 & ~n6514 ) | ( n6896 & n6897 ) | ( ~n6514 & n6897 ) ;
  assign n6900 = ( n6505 & ~n6899 ) | ( n6505 & n6898 ) | ( ~n6899 & n6898 ) ;
  assign n6901 = n3482 | n6873 ;
  assign n6902 = n6887 | n6901 ;
  assign n6903 = n6893 &  n6902 ;
  assign n6904 = n6881 | n6884 ;
  assign n6905 = ( n3760 & n6878 ) | ( n3760 & n6904 ) | ( n6878 & n6904 ) ;
  assign n6906 = n3482 &  n6905 ;
  assign n6907 = n3211 | n6906 ;
  assign n6908 = n6903 | n6907 ;
  assign n6909 = n6900 &  n6908 ;
  assign n6910 = n6895 | n6909 ;
  assign n6912 = ( n6507 & ~n6512 ) | ( n6507 & n6781 ) | ( ~n6512 & n6781 ) ;
  assign n6911 = ~n6520 & n6781 ;
  assign n6913 = ( n6781 & ~n6912 ) | ( n6781 & n6911 ) | ( ~n6912 & n6911 ) ;
  assign n6914 = ( n6911 & ~n6507 ) | ( n6911 & n6912 ) | ( ~n6507 & n6912 ) ;
  assign n6915 = ( n6512 & ~n6913 ) | ( n6512 & n6914 ) | ( ~n6913 & n6914 ) ;
  assign n6916 = ( n2955 & n6910 ) | ( n2955 & n6915 ) | ( n6910 & n6915 ) ;
  assign n6917 = n2706 &  n6916 ;
  assign n6918 = n6540 | n6781 ;
  assign n6919 = ( n6527 & n6536 ) | ( n6527 & n6540 ) | ( n6536 & n6540 ) ;
  assign n6920 = ( n6918 & ~n6536 ) | ( n6918 & n6919 ) | ( ~n6536 & n6919 ) ;
  assign n6921 = ( n6540 & ~n6919 ) | ( n6540 & n6918 ) | ( ~n6919 & n6918 ) ;
  assign n6922 = ( n6527 & ~n6920 ) | ( n6527 & n6921 ) | ( ~n6920 & n6921 ) ;
  assign n6923 = n2955 | n6895 ;
  assign n6924 = n6909 | n6923 ;
  assign n6925 = n6915 &  n6924 ;
  assign n6926 = n6903 | n6906 ;
  assign n6927 = ( n3211 & n6900 ) | ( n3211 & n6926 ) | ( n6900 & n6926 ) ;
  assign n6928 = n2955 &  n6927 ;
  assign n6929 = n2706 | n6928 ;
  assign n6930 = n6925 | n6929 ;
  assign n6931 = n6922 &  n6930 ;
  assign n6932 = n6917 | n6931 ;
  assign n6933 = ~n6542 & n6781 ;
  assign n6934 = ( n6529 & n6534 ) | ( n6529 & n6781 ) | ( n6534 & n6781 ) ;
  assign n6936 = ( n6933 & ~n6529 ) | ( n6933 & n6934 ) | ( ~n6529 & n6934 ) ;
  assign n6935 = ( n6781 & ~n6934 ) | ( n6781 & n6933 ) | ( ~n6934 & n6933 ) ;
  assign n6937 = ( n6534 & ~n6936 ) | ( n6534 & n6935 ) | ( ~n6936 & n6935 ) ;
  assign n6938 = ( n2472 & n6932 ) | ( n2472 & n6937 ) | ( n6932 & n6937 ) ;
  assign n6939 = n2245 &  n6938 ;
  assign n6940 = n6562 | n6781 ;
  assign n6941 = ( n6549 & n6558 ) | ( n6549 & n6562 ) | ( n6558 & n6562 ) ;
  assign n6942 = ( n6940 & ~n6558 ) | ( n6940 & n6941 ) | ( ~n6558 & n6941 ) ;
  assign n6943 = ( n6562 & ~n6941 ) | ( n6562 & n6940 ) | ( ~n6941 & n6940 ) ;
  assign n6944 = ( n6549 & ~n6942 ) | ( n6549 & n6943 ) | ( ~n6942 & n6943 ) ;
  assign n6945 = n2472 | n6917 ;
  assign n6946 = n6931 | n6945 ;
  assign n6947 = n6937 &  n6946 ;
  assign n6948 = n6925 | n6928 ;
  assign n6949 = ( n2706 & n6922 ) | ( n2706 & n6948 ) | ( n6922 & n6948 ) ;
  assign n6950 = n2472 &  n6949 ;
  assign n6951 = n2245 | n6950 ;
  assign n6952 = n6947 | n6951 ;
  assign n6953 = n6944 &  n6952 ;
  assign n6954 = n6939 | n6953 ;
  assign n6955 = ~n6564 & n6781 ;
  assign n6956 = ( n6551 & n6556 ) | ( n6551 & n6781 ) | ( n6556 & n6781 ) ;
  assign n6958 = ( n6955 & ~n6551 ) | ( n6955 & n6956 ) | ( ~n6551 & n6956 ) ;
  assign n6957 = ( n6781 & ~n6956 ) | ( n6781 & n6955 ) | ( ~n6956 & n6955 ) ;
  assign n6959 = ( n6556 & ~n6958 ) | ( n6556 & n6957 ) | ( ~n6958 & n6957 ) ;
  assign n6960 = ( n6954 & ~n2033 ) | ( n6954 & n6959 ) | ( ~n2033 & n6959 ) ;
  assign n6961 = n1827 &  n6960 ;
  assign n6962 = n6584 | n6781 ;
  assign n6963 = ( n6571 & ~n6580 ) | ( n6571 & n6584 ) | ( ~n6580 & n6584 ) ;
  assign n6964 = ( n6580 & n6962 ) | ( n6580 & n6963 ) | ( n6962 & n6963 ) ;
  assign n6965 = ( n6584 & ~n6963 ) | ( n6584 & n6962 ) | ( ~n6963 & n6962 ) ;
  assign n6966 = ( n6571 & ~n6964 ) | ( n6571 & n6965 ) | ( ~n6964 & n6965 ) ;
  assign n6967 = ( n2033 & ~n6939 ) | ( n2033 & 1'b0 ) | ( ~n6939 & 1'b0 ) ;
  assign n6968 = ~n6953 & n6967 ;
  assign n6969 = ( n6959 & ~n6968 ) | ( n6959 & 1'b0 ) | ( ~n6968 & 1'b0 ) ;
  assign n6970 = n6947 | n6950 ;
  assign n6971 = ( n2245 & n6944 ) | ( n2245 & n6970 ) | ( n6944 & n6970 ) ;
  assign n6972 = ~n2033 & n6971 ;
  assign n6973 = n1827 | n6972 ;
  assign n6974 = n6969 | n6973 ;
  assign n6975 = n6966 &  n6974 ;
  assign n6976 = n6961 | n6975 ;
  assign n6977 = ~n6586 & n6781 ;
  assign n6978 = ( n6573 & n6578 ) | ( n6573 & n6781 ) | ( n6578 & n6781 ) ;
  assign n6980 = ( n6977 & ~n6573 ) | ( n6977 & n6978 ) | ( ~n6573 & n6978 ) ;
  assign n6979 = ( n6781 & ~n6978 ) | ( n6781 & n6977 ) | ( ~n6978 & n6977 ) ;
  assign n6981 = ( n6578 & ~n6980 ) | ( n6578 & n6979 ) | ( ~n6980 & n6979 ) ;
  assign n6982 = ( n1636 & ~n6976 ) | ( n1636 & n6981 ) | ( ~n6976 & n6981 ) ;
  assign n6983 = n1452 | n6982 ;
  assign n6984 = n6606 | n6781 ;
  assign n6985 = ( n6593 & ~n6602 ) | ( n6593 & n6606 ) | ( ~n6602 & n6606 ) ;
  assign n6986 = ( n6602 & n6984 ) | ( n6602 & n6985 ) | ( n6984 & n6985 ) ;
  assign n6987 = ( n6606 & ~n6985 ) | ( n6606 & n6984 ) | ( ~n6985 & n6984 ) ;
  assign n6988 = ( n6593 & ~n6986 ) | ( n6593 & n6987 ) | ( ~n6986 & n6987 ) ;
  assign n6989 = ( n1636 & ~n6961 ) | ( n1636 & 1'b0 ) | ( ~n6961 & 1'b0 ) ;
  assign n6990 = ~n6975 & n6989 ;
  assign n6991 = n6981 | n6990 ;
  assign n6992 = n6969 | n6972 ;
  assign n6993 = ( n1827 & n6966 ) | ( n1827 & n6992 ) | ( n6966 & n6992 ) ;
  assign n6994 = ~n1636 & n6993 ;
  assign n6995 = ( n1452 & ~n6994 ) | ( n1452 & 1'b0 ) | ( ~n6994 & 1'b0 ) ;
  assign n6996 = n6991 &  n6995 ;
  assign n6997 = ( n6988 & ~n6996 ) | ( n6988 & 1'b0 ) | ( ~n6996 & 1'b0 ) ;
  assign n6998 = ( n6983 & ~n6997 ) | ( n6983 & 1'b0 ) | ( ~n6997 & 1'b0 ) ;
  assign n6999 = n6608 &  n6781 ;
  assign n7000 = ( n6595 & n6600 ) | ( n6595 & n6781 ) | ( n6600 & n6781 ) ;
  assign n7002 = ( n6999 & ~n6595 ) | ( n6999 & n7000 ) | ( ~n6595 & n7000 ) ;
  assign n7001 = ( n6781 & ~n7000 ) | ( n6781 & n6999 ) | ( ~n7000 & n6999 ) ;
  assign n7003 = ( n6600 & ~n7002 ) | ( n6600 & n7001 ) | ( ~n7002 & n7001 ) ;
  assign n7004 = ( n1283 & ~n6998 ) | ( n1283 & n7003 ) | ( ~n6998 & n7003 ) ;
  assign n7005 = ~n1122 & n7004 ;
  assign n7006 = n6628 | n6781 ;
  assign n7007 = ( n6615 & n6624 ) | ( n6615 & n6628 ) | ( n6624 & n6628 ) ;
  assign n7008 = ( n7006 & ~n6624 ) | ( n7006 & n7007 ) | ( ~n6624 & n7007 ) ;
  assign n7009 = ( n6628 & ~n7007 ) | ( n6628 & n7006 ) | ( ~n7007 & n7006 ) ;
  assign n7010 = ( n6615 & ~n7008 ) | ( n6615 & n7009 ) | ( ~n7008 & n7009 ) ;
  assign n7011 = ~n1283 & n6983 ;
  assign n7012 = ~n6997 & n7011 ;
  assign n7013 = ( n7003 & ~n7012 ) | ( n7003 & 1'b0 ) | ( ~n7012 & 1'b0 ) ;
  assign n7014 = ( n6991 & ~n6994 ) | ( n6991 & 1'b0 ) | ( ~n6994 & 1'b0 ) ;
  assign n7015 = ( n1452 & ~n6988 ) | ( n1452 & n7014 ) | ( ~n6988 & n7014 ) ;
  assign n7016 = ( n1283 & ~n7015 ) | ( n1283 & 1'b0 ) | ( ~n7015 & 1'b0 ) ;
  assign n7017 = ( n1122 & ~n7016 ) | ( n1122 & 1'b0 ) | ( ~n7016 & 1'b0 ) ;
  assign n7018 = ~n7013 & n7017 ;
  assign n7019 = ( n7010 & ~n7018 ) | ( n7010 & 1'b0 ) | ( ~n7018 & 1'b0 ) ;
  assign n7020 = n7005 | n7019 ;
  assign n7021 = n6630 &  n6781 ;
  assign n7022 = ( n6617 & n6622 ) | ( n6617 & n6781 ) | ( n6622 & n6781 ) ;
  assign n7024 = ( n7021 & ~n6617 ) | ( n7021 & n7022 ) | ( ~n6617 & n7022 ) ;
  assign n7023 = ( n6781 & ~n7022 ) | ( n6781 & n7021 ) | ( ~n7022 & n7021 ) ;
  assign n7025 = ( n6622 & ~n7024 ) | ( n6622 & n7023 ) | ( ~n7024 & n7023 ) ;
  assign n7026 = ( n7020 & ~n976 ) | ( n7020 & n7025 ) | ( ~n976 & n7025 ) ;
  assign n7027 = n837 &  n7026 ;
  assign n7028 = n6650 | n6781 ;
  assign n7029 = ( n6637 & ~n6646 ) | ( n6637 & n6650 ) | ( ~n6646 & n6650 ) ;
  assign n7030 = ( n6646 & n7028 ) | ( n6646 & n7029 ) | ( n7028 & n7029 ) ;
  assign n7031 = ( n6650 & ~n7029 ) | ( n6650 & n7028 ) | ( ~n7029 & n7028 ) ;
  assign n7032 = ( n6637 & ~n7030 ) | ( n6637 & n7031 ) | ( ~n7030 & n7031 ) ;
  assign n7033 = ( n976 & ~n7005 ) | ( n976 & 1'b0 ) | ( ~n7005 & 1'b0 ) ;
  assign n7034 = ~n7019 & n7033 ;
  assign n7035 = ( n7025 & ~n7034 ) | ( n7025 & 1'b0 ) | ( ~n7034 & 1'b0 ) ;
  assign n7036 = n7013 | n7016 ;
  assign n7037 = ( n7010 & ~n1122 ) | ( n7010 & n7036 ) | ( ~n1122 & n7036 ) ;
  assign n7038 = ~n976 & n7037 ;
  assign n7039 = n837 | n7038 ;
  assign n7040 = n7035 | n7039 ;
  assign n7041 = ~n7032 & n7040 ;
  assign n7042 = n7027 | n7041 ;
  assign n7044 = ( n6639 & ~n6644 ) | ( n6639 & n6781 ) | ( ~n6644 & n6781 ) ;
  assign n7043 = n6652 &  n6781 ;
  assign n7045 = ( n6781 & ~n7044 ) | ( n6781 & n7043 ) | ( ~n7044 & n7043 ) ;
  assign n7046 = ( n7043 & ~n6639 ) | ( n7043 & n7044 ) | ( ~n6639 & n7044 ) ;
  assign n7047 = ( n6644 & ~n7045 ) | ( n6644 & n7046 ) | ( ~n7045 & n7046 ) ;
  assign n7048 = ( n713 & n7042 ) | ( n713 & n7047 ) | ( n7042 & n7047 ) ;
  assign n7049 = n595 &  n7048 ;
  assign n7051 = ( n6668 & ~n6659 ) | ( n6668 & n6672 ) | ( ~n6659 & n6672 ) ;
  assign n7050 = n6672 | n6781 ;
  assign n7053 = ( n6672 & ~n7051 ) | ( n6672 & n7050 ) | ( ~n7051 & n7050 ) ;
  assign n7052 = ( n7050 & ~n6668 ) | ( n7050 & n7051 ) | ( ~n6668 & n7051 ) ;
  assign n7054 = ( n6659 & ~n7053 ) | ( n6659 & n7052 ) | ( ~n7053 & n7052 ) ;
  assign n7055 = n713 | n7027 ;
  assign n7056 = n7041 | n7055 ;
  assign n7057 = n7047 &  n7056 ;
  assign n7058 = n7035 | n7038 ;
  assign n7059 = ( n837 & ~n7032 ) | ( n837 & n7058 ) | ( ~n7032 & n7058 ) ;
  assign n7060 = n713 &  n7059 ;
  assign n7061 = n595 | n7060 ;
  assign n7062 = n7057 | n7061 ;
  assign n7063 = n7054 &  n7062 ;
  assign n7064 = n7049 | n7063 ;
  assign n7065 = ~n6674 & n6781 ;
  assign n7066 = ( n6661 & ~n7065 ) | ( n6661 & n6781 ) | ( ~n7065 & n6781 ) ;
  assign n7067 = ( n6661 & ~n7066 ) | ( n6661 & n6666 ) | ( ~n7066 & n6666 ) ;
  assign n7068 = ( n6666 & ~n6661 ) | ( n6666 & n7066 ) | ( ~n6661 & n7066 ) ;
  assign n7069 = ( n7067 & ~n6666 ) | ( n7067 & n7068 ) | ( ~n6666 & n7068 ) ;
  assign n7070 = ( n492 & n7064 ) | ( n492 & n7069 ) | ( n7064 & n7069 ) ;
  assign n7071 = n396 &  n7070 ;
  assign n7073 = ( n6690 & ~n6681 ) | ( n6690 & n6694 ) | ( ~n6681 & n6694 ) ;
  assign n7072 = n6694 | n6781 ;
  assign n7075 = ( n6694 & ~n7073 ) | ( n6694 & n7072 ) | ( ~n7073 & n7072 ) ;
  assign n7074 = ( n7072 & ~n6690 ) | ( n7072 & n7073 ) | ( ~n6690 & n7073 ) ;
  assign n7076 = ( n6681 & ~n7075 ) | ( n6681 & n7074 ) | ( ~n7075 & n7074 ) ;
  assign n7077 = n492 | n7049 ;
  assign n7078 = n7063 | n7077 ;
  assign n7079 = n7069 &  n7078 ;
  assign n7080 = n7057 | n7060 ;
  assign n7081 = ( n595 & n7054 ) | ( n595 & n7080 ) | ( n7054 & n7080 ) ;
  assign n7082 = n492 &  n7081 ;
  assign n7083 = n396 | n7082 ;
  assign n7084 = n7079 | n7083 ;
  assign n7085 = ~n7076 & n7084 ;
  assign n7086 = n7071 | n7085 ;
  assign n7087 = ~n6696 & n6781 ;
  assign n7088 = ( n6683 & ~n7087 ) | ( n6683 & n6781 ) | ( ~n7087 & n6781 ) ;
  assign n7089 = ( n6683 & ~n7088 ) | ( n6683 & n6688 ) | ( ~n7088 & n6688 ) ;
  assign n7090 = ( n6688 & ~n6683 ) | ( n6688 & n7088 ) | ( ~n6683 & n7088 ) ;
  assign n7091 = ( n7089 & ~n6688 ) | ( n7089 & n7090 ) | ( ~n6688 & n7090 ) ;
  assign n7092 = ( n315 & n7086 ) | ( n315 & n7091 ) | ( n7086 & n7091 ) ;
  assign n7093 = n240 &  n7092 ;
  assign n7095 = ( n6712 & ~n6703 ) | ( n6712 & n6716 ) | ( ~n6703 & n6716 ) ;
  assign n7094 = n6716 | n6781 ;
  assign n7097 = ( n6716 & ~n7095 ) | ( n6716 & n7094 ) | ( ~n7095 & n7094 ) ;
  assign n7096 = ( n7094 & ~n6712 ) | ( n7094 & n7095 ) | ( ~n6712 & n7095 ) ;
  assign n7098 = ( n6703 & ~n7097 ) | ( n6703 & n7096 ) | ( ~n7097 & n7096 ) ;
  assign n7099 = n315 | n7071 ;
  assign n7100 = n7085 | n7099 ;
  assign n7101 = n7091 &  n7100 ;
  assign n7102 = n7079 | n7082 ;
  assign n7103 = ( n396 & ~n7076 ) | ( n396 & n7102 ) | ( ~n7076 & n7102 ) ;
  assign n7104 = n315 &  n7103 ;
  assign n7105 = n240 | n7104 ;
  assign n7106 = n7101 | n7105 ;
  assign n7107 = n7098 &  n7106 ;
  assign n7108 = n7093 | n7107 ;
  assign n7109 = n6705 | n6781 ;
  assign n7110 = ( n6705 & n6710 ) | ( n6705 & n6718 ) | ( n6710 & n6718 ) ;
  assign n7111 = ( n7109 & ~n6718 ) | ( n7109 & n7110 ) | ( ~n6718 & n7110 ) ;
  assign n7112 = ( n6705 & ~n7110 ) | ( n6705 & n7109 ) | ( ~n7110 & n7109 ) ;
  assign n7113 = ( n6710 & ~n7111 ) | ( n6710 & n7112 ) | ( ~n7111 & n7112 ) ;
  assign n7114 = ( n181 & n7108 ) | ( n181 & n7113 ) | ( n7108 & n7113 ) ;
  assign n7115 = ~n145 & n7114 ;
  assign n7117 = ( n6734 & ~n6725 ) | ( n6734 & n6738 ) | ( ~n6725 & n6738 ) ;
  assign n7116 = n6738 | n6781 ;
  assign n7119 = ( n6738 & ~n7117 ) | ( n6738 & n7116 ) | ( ~n7117 & n7116 ) ;
  assign n7118 = ( n7116 & ~n6734 ) | ( n7116 & n7117 ) | ( ~n6734 & n7117 ) ;
  assign n7120 = ( n6725 & ~n7119 ) | ( n6725 & n7118 ) | ( ~n7119 & n7118 ) ;
  assign n7121 = n181 | n7093 ;
  assign n7122 = n7107 | n7121 ;
  assign n7123 = n7113 &  n7122 ;
  assign n7124 = n7101 | n7104 ;
  assign n7125 = ( n240 & n7098 ) | ( n240 & n7124 ) | ( n7098 & n7124 ) ;
  assign n7126 = n181 &  n7125 ;
  assign n7127 = ( n145 & ~n7126 ) | ( n145 & 1'b0 ) | ( ~n7126 & 1'b0 ) ;
  assign n7128 = ~n7123 & n7127 ;
  assign n7129 = ( n7120 & ~n7128 ) | ( n7120 & 1'b0 ) | ( ~n7128 & 1'b0 ) ;
  assign n7130 = n7115 | n7129 ;
  assign n7132 = ( n6727 & ~n6732 ) | ( n6727 & n6781 ) | ( ~n6732 & n6781 ) ;
  assign n7131 = n6740 &  n6781 ;
  assign n7133 = ( n6781 & ~n7132 ) | ( n6781 & n7131 ) | ( ~n7132 & n7131 ) ;
  assign n7134 = ( n7131 & ~n6727 ) | ( n7131 & n7132 ) | ( ~n6727 & n7132 ) ;
  assign n7135 = ( n6732 & ~n7133 ) | ( n6732 & n7134 ) | ( ~n7133 & n7134 ) ;
  assign n7136 = ( n150 & n7130 ) | ( n150 & n7135 ) | ( n7130 & n7135 ) ;
  assign n7137 = n6747 | n6766 ;
  assign n7138 = ( n6763 & ~n6781 ) | ( n6763 & n7137 ) | ( ~n6781 & n7137 ) ;
  assign n7139 = ( n6763 & ~n7138 ) | ( n6763 & 1'b0 ) | ( ~n7138 & 1'b0 ) ;
  assign n7140 = ( n6763 & ~n6766 ) | ( n6763 & 1'b0 ) | ( ~n6766 & 1'b0 ) ;
  assign n7141 = ~n6781 & n7140 ;
  assign n7142 = ( n6747 & ~n7140 ) | ( n6747 & n7141 ) | ( ~n7140 & n7141 ) ;
  assign n7143 = n7139 | n7142 ;
  assign n7144 = ( n6748 & ~n6755 ) | ( n6748 & 1'b0 ) | ( ~n6755 & 1'b0 ) ;
  assign n7145 = ~n6781 & n7144 ;
  assign n7146 = ( n6769 & ~n7145 ) | ( n6769 & n7144 ) | ( ~n7145 & n7144 ) ;
  assign n7147 = ( n7143 & ~n7146 ) | ( n7143 & 1'b0 ) | ( ~n7146 & 1'b0 ) ;
  assign n7148 = ~n7136 & n7147 ;
  assign n7149 = ( n133 & ~n7148 ) | ( n133 & n7147 ) | ( ~n7148 & n7147 ) ;
  assign n7150 = n150 | n7115 ;
  assign n7151 = n7129 | n7150 ;
  assign n7156 = ( n7135 & ~n7151 ) | ( n7135 & 1'b0 ) | ( ~n7151 & 1'b0 ) ;
  assign n7152 = n7123 | n7126 ;
  assign n7153 = ( n7120 & ~n145 ) | ( n7120 & n7152 ) | ( ~n145 & n7152 ) ;
  assign n7154 = n150 &  n7153 ;
  assign n7155 = n7143 | n7154 ;
  assign n7157 = ( n7135 & ~n7156 ) | ( n7135 & n7155 ) | ( ~n7156 & n7155 ) ;
  assign n7159 = ( n133 & ~n6755 ) | ( n133 & n6748 ) | ( ~n6755 & n6748 ) ;
  assign n7158 = ( n6755 & ~n6748 ) | ( n6755 & n6781 ) | ( ~n6748 & n6781 ) ;
  assign n7160 = ~n6755 & n7158 ;
  assign n7161 = ( n6755 & n7159 ) | ( n6755 & n7160 ) | ( n7159 & n7160 ) ;
  assign n7162 = ( n6751 & ~n6778 ) | ( n6751 & 1'b0 ) | ( ~n6778 & 1'b0 ) ;
  assign n7163 = ( n6754 & ~n6773 ) | ( n6754 & n7162 ) | ( ~n6773 & n7162 ) ;
  assign n7164 = ~n6754 & n7163 ;
  assign n7165 = ( n6761 & ~n7164 ) | ( n6761 & n6769 ) | ( ~n7164 & n6769 ) ;
  assign n7166 = ( n6761 & ~n7165 ) | ( n6761 & 1'b0 ) | ( ~n7165 & 1'b0 ) ;
  assign n7167 = n7161 | n7166 ;
  assign n7168 = ( n7157 & ~n7167 ) | ( n7157 & 1'b0 ) | ( ~n7167 & 1'b0 ) ;
  assign n7169 = n7149 &  n7168 ;
  assign n7227 = n6804 &  n7169 ;
  assign n7230 = ( n6804 & ~n7228 ) | ( n6804 & n7227 ) | ( ~n7228 & n7227 ) ;
  assign n7229 = ( n7227 & ~n6821 ) | ( n7227 & n7228 ) | ( ~n6821 & n7228 ) ;
  assign n7231 = ( n6814 & ~n7230 ) | ( n6814 & n7229 ) | ( ~n7230 & n7229 ) ;
  assign n7212 = ~n6816 & n6819 ;
  assign n7213 = ( n6802 & ~n6816 ) | ( n6802 & n7212 ) | ( ~n6816 & n7212 ) ;
  assign n7214 = ( n7169 & ~n7212 ) | ( n7169 & n7213 ) | ( ~n7212 & n7213 ) ;
  assign n7215 = ( n6816 & ~n7169 ) | ( n6816 & n7213 ) | ( ~n7169 & n7213 ) ;
  assign n7216 = ( n7214 & ~n6802 ) | ( n7214 & n7215 ) | ( ~n6802 & n7215 ) ;
  assign n7203 = ~x60 & n6781 ;
  assign n7204 = ( x61 & ~n7203 ) | ( x61 & 1'b0 ) | ( ~n7203 & 1'b0 ) ;
  assign n7205 = n6793 | n7204 ;
  assign n7200 = ( n6781 & ~x60 ) | ( n6781 & n6788 ) | ( ~x60 & n6788 ) ;
  assign n7201 = x60 &  n7200 ;
  assign n7202 = ( n6783 & ~n6788 ) | ( n6783 & n7201 ) | ( ~n6788 & n7201 ) ;
  assign n7206 = ( n7169 & n7202 ) | ( n7169 & n7205 ) | ( n7202 & n7205 ) ;
  assign n7208 = ~n7169 & n7206 ;
  assign n7207 = ( n7202 & ~n7206 ) | ( n7202 & 1'b0 ) | ( ~n7206 & 1'b0 ) ;
  assign n7209 = ( n7205 & ~n7208 ) | ( n7205 & n7207 ) | ( ~n7208 & n7207 ) ;
  assign n7172 = x56 | x57 ;
  assign n7177 = ~x58 & n7172 ;
  assign n7178 = ( x58 & ~n6779 ) | ( x58 & n7177 ) | ( ~n6779 & n7177 ) ;
  assign n7179 = ( n6761 & ~n7178 ) | ( n6761 & n6769 ) | ( ~n7178 & n6769 ) ;
  assign n7180 = ( n6761 & ~n7179 ) | ( n6761 & 1'b0 ) | ( ~n7179 & 1'b0 ) ;
  assign n7181 = ( x59 & ~n7180 ) | ( x59 & n7169 ) | ( ~n7180 & n7169 ) ;
  assign n7176 = ( x58 & x59 ) | ( x58 & n7169 ) | ( x59 & n7169 ) ;
  assign n7182 = ( x58 & ~x59 ) | ( x58 & 1'b0 ) | ( ~x59 & 1'b0 ) ;
  assign n7183 = ( n7181 & ~n7176 ) | ( n7181 & n7182 ) | ( ~n7176 & n7182 ) ;
  assign n7173 = x58 | n7172 ;
  assign n7174 = ( x58 & ~n7169 ) | ( x58 & 1'b0 ) | ( ~n7169 & 1'b0 ) ;
  assign n7175 = ( n6781 & ~n7173 ) | ( n6781 & n7174 ) | ( ~n7173 & n7174 ) ;
  assign n7186 = ( n6399 & ~n7175 ) | ( n6399 & 1'b0 ) | ( ~n7175 & 1'b0 ) ;
  assign n7187 = ~n7183 & n7186 ;
  assign n7188 = n6400 | n7169 ;
  assign n7189 = ( n6781 & ~n7166 ) | ( n6781 & 1'b0 ) | ( ~n7166 & 1'b0 ) ;
  assign n7190 = ( n7157 & ~n7189 ) | ( n7157 & n7161 ) | ( ~n7189 & n7161 ) ;
  assign n7191 = ( n7157 & ~n7190 ) | ( n7157 & 1'b0 ) | ( ~n7190 & 1'b0 ) ;
  assign n7192 = n7149 &  n7191 ;
  assign n7193 = n7188 | n7192 ;
  assign n7194 = ( x60 & ~n7193 ) | ( x60 & n7192 ) | ( ~n7193 & n7192 ) ;
  assign n7195 = x60 | n7192 ;
  assign n7196 = ( n7188 & ~n7195 ) | ( n7188 & 1'b0 ) | ( ~n7195 & 1'b0 ) ;
  assign n7197 = n7194 | n7196 ;
  assign n7198 = ~n7187 & n7197 ;
  assign n7184 = ~n7183 & n7175 ;
  assign n7185 = ( n7184 & ~n6399 ) | ( n7184 & n7183 ) | ( ~n6399 & n7183 ) ;
  assign n7217 = n6032 | n7185 ;
  assign n7218 = n7198 | n7217 ;
  assign n7219 = ~n7209 & n7218 ;
  assign n7220 = n7175 | n7183 ;
  assign n7221 = ( n7197 & ~n6399 ) | ( n7197 & n7220 ) | ( ~n6399 & n7220 ) ;
  assign n7222 = n6032 &  n7221 ;
  assign n7223 = ( n5672 & ~n7222 ) | ( n5672 & 1'b0 ) | ( ~n7222 & 1'b0 ) ;
  assign n7224 = ~n7219 & n7223 ;
  assign n7225 = ( n7216 & ~n7224 ) | ( n7216 & 1'b0 ) | ( ~n7224 & 1'b0 ) ;
  assign n7199 = n7185 | n7198 ;
  assign n7210 = ( n6032 & ~n7209 ) | ( n6032 & n7199 ) | ( ~n7209 & n7199 ) ;
  assign n7211 = ~n5672 & n7210 ;
  assign n7239 = n5327 | n7211 ;
  assign n7240 = n7225 | n7239 ;
  assign n7242 = n7219 | n7222 ;
  assign n7243 = ( n7216 & ~n5672 ) | ( n7216 & n7242 ) | ( ~n5672 & n7242 ) ;
  assign n7244 = n5327 &  n7243 ;
  assign n7645 = ( n7240 & ~n7231 ) | ( n7240 & n7244 ) | ( ~n7231 & n7244 ) ;
  assign n7534 = ~n7169 & n7128 ;
  assign n7535 = ( n7534 & ~n7115 ) | ( n7534 & n7169 ) | ( ~n7115 & n7169 ) ;
  assign n7536 = ( n7115 & n7120 ) | ( n7115 & n7535 ) | ( n7120 & n7535 ) ;
  assign n7537 = ( n7115 & ~n7120 ) | ( n7115 & n7535 ) | ( ~n7120 & n7535 ) ;
  assign n7538 = ( n7120 & ~n7536 ) | ( n7120 & n7537 ) | ( ~n7536 & n7537 ) ;
  assign n7490 = n7084 | n7169 ;
  assign n7491 = ( n7071 & ~n7169 ) | ( n7071 & n7490 ) | ( ~n7169 & n7490 ) ;
  assign n7492 = ( n7076 & ~n7071 ) | ( n7076 & n7491 ) | ( ~n7071 & n7491 ) ;
  assign n7493 = ( n7071 & ~n7491 ) | ( n7071 & n7076 ) | ( ~n7491 & n7076 ) ;
  assign n7494 = ( n7492 & ~n7076 ) | ( n7492 & n7493 ) | ( ~n7076 & n7493 ) ;
  assign n7270 = n6864 | n7169 ;
  assign n7271 = ( n6856 & ~n6851 ) | ( n6856 & n7169 ) | ( ~n6851 & n7169 ) ;
  assign n7273 = ( n6851 & n7270 ) | ( n6851 & n7271 ) | ( n7270 & n7271 ) ;
  assign n7272 = ( n7169 & ~n7271 ) | ( n7169 & n7270 ) | ( ~n7271 & n7270 ) ;
  assign n7274 = ( n6856 & ~n7273 ) | ( n6856 & n7272 ) | ( ~n7273 & n7272 ) ;
  assign n7249 = ( n6830 & n6838 ) | ( n6830 & n6842 ) | ( n6838 & n6842 ) ;
  assign n7251 = ( n7169 & ~n6830 ) | ( n7169 & n7249 ) | ( ~n6830 & n7249 ) ;
  assign n7250 = ( n6838 & ~n7249 ) | ( n6838 & n7169 ) | ( ~n7249 & n7169 ) ;
  assign n7252 = ( n6842 & ~n7251 ) | ( n6842 & n7250 ) | ( ~n7251 & n7250 ) ;
  assign n7226 = n7211 | n7225 ;
  assign n7232 = ( n5327 & n7226 ) | ( n5327 & n7231 ) | ( n7226 & n7231 ) ;
  assign n7233 = n4990 &  n7232 ;
  assign n7234 = ~n6836 & n7169 ;
  assign n7235 = ( n6828 & ~n6832 ) | ( n6828 & n6836 ) | ( ~n6832 & n6836 ) ;
  assign n7236 = ( n6832 & ~n7234 ) | ( n6832 & n7235 ) | ( ~n7234 & n7235 ) ;
  assign n7237 = ( n7234 & ~n6836 ) | ( n7234 & n7235 ) | ( ~n6836 & n7235 ) ;
  assign n7238 = ( n7236 & ~n6828 ) | ( n7236 & n7237 ) | ( ~n6828 & n7237 ) ;
  assign n7241 = n7231 &  n7240 ;
  assign n7245 = n4990 | n7244 ;
  assign n7246 = n7241 | n7245 ;
  assign n7247 = ~n7238 & n7246 ;
  assign n7248 = n7233 | n7247 ;
  assign n7253 = ( n4668 & ~n7252 ) | ( n4668 & n7248 ) | ( ~n7252 & n7248 ) ;
  assign n7254 = n4353 &  n7253 ;
  assign n7255 = ~n6862 & n7169 ;
  assign n7256 = ( n6849 & n6858 ) | ( n6849 & n6862 ) | ( n6858 & n6862 ) ;
  assign n7258 = ( n7255 & ~n6862 ) | ( n7255 & n7256 ) | ( ~n6862 & n7256 ) ;
  assign n7257 = ( n6858 & ~n7256 ) | ( n6858 & n7255 ) | ( ~n7256 & n7255 ) ;
  assign n7259 = ( n6849 & ~n7258 ) | ( n6849 & n7257 ) | ( ~n7258 & n7257 ) ;
  assign n7260 = n4668 | n7233 ;
  assign n7261 = n7247 | n7260 ;
  assign n7262 = ~n7252 & n7261 ;
  assign n7263 = n7241 | n7244 ;
  assign n7264 = ( n4990 & ~n7238 ) | ( n4990 & n7263 ) | ( ~n7238 & n7263 ) ;
  assign n7265 = n4668 &  n7264 ;
  assign n7266 = n4353 | n7265 ;
  assign n7267 = n7262 | n7266 ;
  assign n7268 = n7259 &  n7267 ;
  assign n7269 = n7254 | n7268 ;
  assign n7275 = ( n4053 & ~n7274 ) | ( n4053 & n7269 ) | ( ~n7274 & n7269 ) ;
  assign n7276 = n3760 &  n7275 ;
  assign n7277 = ~n6884 & n7169 ;
  assign n7278 = ( n6871 & n6880 ) | ( n6871 & n6884 ) | ( n6880 & n6884 ) ;
  assign n7280 = ( n7277 & ~n6884 ) | ( n7277 & n7278 ) | ( ~n6884 & n7278 ) ;
  assign n7279 = ( n6880 & ~n7278 ) | ( n6880 & n7277 ) | ( ~n7278 & n7277 ) ;
  assign n7281 = ( n6871 & ~n7280 ) | ( n6871 & n7279 ) | ( ~n7280 & n7279 ) ;
  assign n7282 = n4053 | n7254 ;
  assign n7283 = n7268 | n7282 ;
  assign n7284 = ~n7274 & n7283 ;
  assign n7285 = n7262 | n7265 ;
  assign n7286 = ( n4353 & n7259 ) | ( n4353 & n7285 ) | ( n7259 & n7285 ) ;
  assign n7287 = n4053 &  n7286 ;
  assign n7288 = n3760 | n7287 ;
  assign n7289 = n7284 | n7288 ;
  assign n7290 = n7281 &  n7289 ;
  assign n7291 = n7276 | n7290 ;
  assign n7292 = n6886 | n7169 ;
  assign n7293 = ( n6873 & ~n7169 ) | ( n6873 & n6878 ) | ( ~n7169 & n6878 ) ;
  assign n7294 = ( n7169 & n7292 ) | ( n7169 & n7293 ) | ( n7292 & n7293 ) ;
  assign n7295 = ( n6873 & ~n7293 ) | ( n6873 & n7292 ) | ( ~n7293 & n7292 ) ;
  assign n7296 = ( n6878 & ~n7294 ) | ( n6878 & n7295 ) | ( ~n7294 & n7295 ) ;
  assign n7297 = ( n3482 & n7291 ) | ( n3482 & n7296 ) | ( n7291 & n7296 ) ;
  assign n7298 = n3211 &  n7297 ;
  assign n7299 = ~n6906 & n7169 ;
  assign n7300 = ( n6893 & n6902 ) | ( n6893 & n6906 ) | ( n6902 & n6906 ) ;
  assign n7302 = ( n7299 & ~n6906 ) | ( n7299 & n7300 ) | ( ~n6906 & n7300 ) ;
  assign n7301 = ( n6902 & ~n7300 ) | ( n6902 & n7299 ) | ( ~n7300 & n7299 ) ;
  assign n7303 = ( n6893 & ~n7302 ) | ( n6893 & n7301 ) | ( ~n7302 & n7301 ) ;
  assign n7304 = n3482 | n7276 ;
  assign n7305 = n7290 | n7304 ;
  assign n7306 = n7296 &  n7305 ;
  assign n7307 = n7284 | n7287 ;
  assign n7308 = ( n3760 & n7281 ) | ( n3760 & n7307 ) | ( n7281 & n7307 ) ;
  assign n7309 = n3482 &  n7308 ;
  assign n7310 = n3211 | n7309 ;
  assign n7311 = n7306 | n7310 ;
  assign n7312 = n7303 &  n7311 ;
  assign n7313 = n7298 | n7312 ;
  assign n7314 = n6908 | n7169 ;
  assign n7315 = ( n6895 & ~n7169 ) | ( n6895 & n7314 ) | ( ~n7169 & n7314 ) ;
  assign n7316 = ( n6895 & ~n7315 ) | ( n6895 & n6900 ) | ( ~n7315 & n6900 ) ;
  assign n7317 = ( n6900 & ~n6895 ) | ( n6900 & n7315 ) | ( ~n6895 & n7315 ) ;
  assign n7318 = ( n7316 & ~n6900 ) | ( n7316 & n7317 ) | ( ~n6900 & n7317 ) ;
  assign n7319 = ( n2955 & n7313 ) | ( n2955 & n7318 ) | ( n7313 & n7318 ) ;
  assign n7320 = n2706 &  n7319 ;
  assign n7321 = ~n6928 & n7169 ;
  assign n7322 = ( n6915 & n6924 ) | ( n6915 & n6928 ) | ( n6924 & n6928 ) ;
  assign n7324 = ( n7321 & ~n6928 ) | ( n7321 & n7322 ) | ( ~n6928 & n7322 ) ;
  assign n7323 = ( n6924 & ~n7322 ) | ( n6924 & n7321 ) | ( ~n7322 & n7321 ) ;
  assign n7325 = ( n6915 & ~n7324 ) | ( n6915 & n7323 ) | ( ~n7324 & n7323 ) ;
  assign n7326 = n2955 | n7298 ;
  assign n7327 = n7312 | n7326 ;
  assign n7328 = n7318 &  n7327 ;
  assign n7329 = n7306 | n7309 ;
  assign n7330 = ( n3211 & n7303 ) | ( n3211 & n7329 ) | ( n7303 & n7329 ) ;
  assign n7331 = n2955 &  n7330 ;
  assign n7332 = n2706 | n7331 ;
  assign n7333 = n7328 | n7332 ;
  assign n7334 = n7325 &  n7333 ;
  assign n7335 = n7320 | n7334 ;
  assign n7336 = n6930 | n7169 ;
  assign n7337 = ( n6917 & ~n7169 ) | ( n6917 & n6922 ) | ( ~n7169 & n6922 ) ;
  assign n7338 = ( n7169 & n7336 ) | ( n7169 & n7337 ) | ( n7336 & n7337 ) ;
  assign n7339 = ( n6917 & ~n7337 ) | ( n6917 & n7336 ) | ( ~n7337 & n7336 ) ;
  assign n7340 = ( n6922 & ~n7338 ) | ( n6922 & n7339 ) | ( ~n7338 & n7339 ) ;
  assign n7341 = ( n2472 & n7335 ) | ( n2472 & n7340 ) | ( n7335 & n7340 ) ;
  assign n7342 = n2245 &  n7341 ;
  assign n7343 = ~n6950 & n7169 ;
  assign n7344 = ( n6937 & n6946 ) | ( n6937 & n6950 ) | ( n6946 & n6950 ) ;
  assign n7346 = ( n7343 & ~n6950 ) | ( n7343 & n7344 ) | ( ~n6950 & n7344 ) ;
  assign n7345 = ( n6946 & ~n7344 ) | ( n6946 & n7343 ) | ( ~n7344 & n7343 ) ;
  assign n7347 = ( n6937 & ~n7346 ) | ( n6937 & n7345 ) | ( ~n7346 & n7345 ) ;
  assign n7348 = n2472 | n7320 ;
  assign n7349 = n7334 | n7348 ;
  assign n7350 = n7340 &  n7349 ;
  assign n7351 = n7328 | n7331 ;
  assign n7352 = ( n2706 & n7325 ) | ( n2706 & n7351 ) | ( n7325 & n7351 ) ;
  assign n7353 = n2472 &  n7352 ;
  assign n7354 = n2245 | n7353 ;
  assign n7355 = n7350 | n7354 ;
  assign n7356 = n7347 &  n7355 ;
  assign n7357 = n7342 | n7356 ;
  assign n7358 = n6952 | n7169 ;
  assign n7359 = ( n6939 & ~n7169 ) | ( n6939 & n6944 ) | ( ~n7169 & n6944 ) ;
  assign n7360 = ( n7169 & n7358 ) | ( n7169 & n7359 ) | ( n7358 & n7359 ) ;
  assign n7361 = ( n6939 & ~n7359 ) | ( n6939 & n7358 ) | ( ~n7359 & n7358 ) ;
  assign n7362 = ( n6944 & ~n7360 ) | ( n6944 & n7361 ) | ( ~n7360 & n7361 ) ;
  assign n7363 = ( n7357 & ~n2033 ) | ( n7357 & n7362 ) | ( ~n2033 & n7362 ) ;
  assign n7364 = n1827 &  n7363 ;
  assign n7365 = ~n6972 & n7169 ;
  assign n7366 = ( n6959 & ~n6968 ) | ( n6959 & n6972 ) | ( ~n6968 & n6972 ) ;
  assign n7367 = ( n6968 & ~n7365 ) | ( n6968 & n7366 ) | ( ~n7365 & n7366 ) ;
  assign n7368 = ( n7365 & ~n6972 ) | ( n7365 & n7366 ) | ( ~n6972 & n7366 ) ;
  assign n7369 = ( n7367 & ~n6959 ) | ( n7367 & n7368 ) | ( ~n6959 & n7368 ) ;
  assign n7370 = ( n2033 & ~n7342 ) | ( n2033 & 1'b0 ) | ( ~n7342 & 1'b0 ) ;
  assign n7371 = ~n7356 & n7370 ;
  assign n7372 = ( n7362 & ~n7371 ) | ( n7362 & 1'b0 ) | ( ~n7371 & 1'b0 ) ;
  assign n7373 = n7350 | n7353 ;
  assign n7374 = ( n2245 & n7347 ) | ( n2245 & n7373 ) | ( n7347 & n7373 ) ;
  assign n7375 = ~n2033 & n7374 ;
  assign n7376 = n1827 | n7375 ;
  assign n7377 = n7372 | n7376 ;
  assign n7378 = ~n7369 & n7377 ;
  assign n7379 = n7364 | n7378 ;
  assign n7380 = n6974 | n7169 ;
  assign n7381 = ( n6961 & ~n7169 ) | ( n6961 & n7380 ) | ( ~n7169 & n7380 ) ;
  assign n7382 = ( n6961 & ~n7381 ) | ( n6961 & n6966 ) | ( ~n7381 & n6966 ) ;
  assign n7383 = ( n6966 & ~n6961 ) | ( n6966 & n7381 ) | ( ~n6961 & n7381 ) ;
  assign n7384 = ( n7382 & ~n6966 ) | ( n7382 & n7383 ) | ( ~n6966 & n7383 ) ;
  assign n7385 = ( n7379 & ~n1636 ) | ( n7379 & n7384 ) | ( ~n1636 & n7384 ) ;
  assign n7386 = ~n1452 & n7385 ;
  assign n7387 = ~n6994 & n7169 ;
  assign n7388 = ( n6981 & ~n6994 ) | ( n6981 & n6990 ) | ( ~n6994 & n6990 ) ;
  assign n7389 = ( n7387 & ~n6990 ) | ( n7387 & n7388 ) | ( ~n6990 & n7388 ) ;
  assign n7390 = ( n6994 & ~n7387 ) | ( n6994 & n7388 ) | ( ~n7387 & n7388 ) ;
  assign n7391 = ( n7389 & ~n6981 ) | ( n7389 & n7390 ) | ( ~n6981 & n7390 ) ;
  assign n7392 = ( n1636 & ~n7364 ) | ( n1636 & 1'b0 ) | ( ~n7364 & 1'b0 ) ;
  assign n7393 = ~n7378 & n7392 ;
  assign n7394 = ( n7384 & ~n7393 ) | ( n7384 & 1'b0 ) | ( ~n7393 & 1'b0 ) ;
  assign n7395 = n7372 | n7375 ;
  assign n7396 = ( n1827 & ~n7369 ) | ( n1827 & n7395 ) | ( ~n7369 & n7395 ) ;
  assign n7397 = ~n1636 & n7396 ;
  assign n7398 = ( n1452 & ~n7397 ) | ( n1452 & 1'b0 ) | ( ~n7397 & 1'b0 ) ;
  assign n7399 = ~n7394 & n7398 ;
  assign n7400 = ( n7391 & ~n7399 ) | ( n7391 & 1'b0 ) | ( ~n7399 & 1'b0 ) ;
  assign n7401 = n7386 | n7400 ;
  assign n7402 = ( n6996 & ~n7169 ) | ( n6996 & 1'b0 ) | ( ~n7169 & 1'b0 ) ;
  assign n7403 = ( n6983 & n6988 ) | ( n6983 & n7169 ) | ( n6988 & n7169 ) ;
  assign n7404 = ( n7402 & ~n7169 ) | ( n7402 & n7403 ) | ( ~n7169 & n7403 ) ;
  assign n7405 = ( n6983 & ~n7403 ) | ( n6983 & n7402 ) | ( ~n7403 & n7402 ) ;
  assign n7406 = ( n6988 & ~n7404 ) | ( n6988 & n7405 ) | ( ~n7404 & n7405 ) ;
  assign n7407 = ( n1283 & n7401 ) | ( n1283 & n7406 ) | ( n7401 & n7406 ) ;
  assign n7408 = ~n1122 & n7407 ;
  assign n7409 = ~n7016 & n7169 ;
  assign n7410 = ( n7003 & ~n7012 ) | ( n7003 & n7016 ) | ( ~n7012 & n7016 ) ;
  assign n7411 = ( n7012 & ~n7409 ) | ( n7012 & n7410 ) | ( ~n7409 & n7410 ) ;
  assign n7412 = ( n7409 & ~n7016 ) | ( n7409 & n7410 ) | ( ~n7016 & n7410 ) ;
  assign n7413 = ( n7411 & ~n7003 ) | ( n7411 & n7412 ) | ( ~n7003 & n7412 ) ;
  assign n7414 = n1283 | n7386 ;
  assign n7415 = n7400 | n7414 ;
  assign n7416 = n7406 &  n7415 ;
  assign n7417 = n7394 | n7397 ;
  assign n7418 = ( n7391 & ~n1452 ) | ( n7391 & n7417 ) | ( ~n1452 & n7417 ) ;
  assign n7419 = n1283 &  n7418 ;
  assign n7420 = ( n1122 & ~n7419 ) | ( n1122 & 1'b0 ) | ( ~n7419 & 1'b0 ) ;
  assign n7421 = ~n7416 & n7420 ;
  assign n7422 = n7413 | n7421 ;
  assign n7423 = ~n7408 & n7422 ;
  assign n7424 = ( n7018 & ~n7169 ) | ( n7018 & 1'b0 ) | ( ~n7169 & 1'b0 ) ;
  assign n7425 = ( n7010 & ~n7005 ) | ( n7010 & n7169 ) | ( ~n7005 & n7169 ) ;
  assign n7426 = ( n7424 & ~n7169 ) | ( n7424 & n7425 ) | ( ~n7169 & n7425 ) ;
  assign n7427 = ( n7005 & ~n7424 ) | ( n7005 & n7425 ) | ( ~n7424 & n7425 ) ;
  assign n7428 = ( n7426 & ~n7010 ) | ( n7426 & n7427 ) | ( ~n7010 & n7427 ) ;
  assign n7429 = ( n976 & n7423 ) | ( n976 & n7428 ) | ( n7423 & n7428 ) ;
  assign n7430 = ( n837 & ~n7429 ) | ( n837 & 1'b0 ) | ( ~n7429 & 1'b0 ) ;
  assign n7431 = ~n7038 & n7169 ;
  assign n7432 = ( n7025 & ~n7034 ) | ( n7025 & n7038 ) | ( ~n7034 & n7038 ) ;
  assign n7433 = ( n7034 & ~n7431 ) | ( n7034 & n7432 ) | ( ~n7431 & n7432 ) ;
  assign n7434 = ( n7431 & ~n7038 ) | ( n7431 & n7432 ) | ( ~n7038 & n7432 ) ;
  assign n7435 = ( n7433 & ~n7025 ) | ( n7433 & n7434 ) | ( ~n7025 & n7434 ) ;
  assign n7436 = ( n976 & ~n7408 ) | ( n976 & 1'b0 ) | ( ~n7408 & 1'b0 ) ;
  assign n7437 = n7422 &  n7436 ;
  assign n7438 = n7428 | n7437 ;
  assign n7439 = n7416 | n7419 ;
  assign n7440 = ( n1122 & ~n7439 ) | ( n1122 & n7413 ) | ( ~n7439 & n7413 ) ;
  assign n7441 = n976 | n7440 ;
  assign n7442 = ~n837 & n7441 ;
  assign n7443 = n7438 &  n7442 ;
  assign n7444 = n7435 | n7443 ;
  assign n7445 = ~n7430 & n7444 ;
  assign n7446 = n7040 | n7169 ;
  assign n7447 = ( n7032 & ~n7027 ) | ( n7032 & n7169 ) | ( ~n7027 & n7169 ) ;
  assign n7449 = ( n7027 & n7446 ) | ( n7027 & n7447 ) | ( n7446 & n7447 ) ;
  assign n7448 = ( n7169 & ~n7447 ) | ( n7169 & n7446 ) | ( ~n7447 & n7446 ) ;
  assign n7450 = ( n7032 & ~n7449 ) | ( n7032 & n7448 ) | ( ~n7449 & n7448 ) ;
  assign n7451 = ( n7445 & ~n713 ) | ( n7445 & n7450 ) | ( ~n713 & n7450 ) ;
  assign n7452 = ( n595 & ~n7451 ) | ( n595 & 1'b0 ) | ( ~n7451 & 1'b0 ) ;
  assign n7453 = ~n7060 & n7169 ;
  assign n7454 = ( n7047 & n7056 ) | ( n7047 & n7060 ) | ( n7056 & n7060 ) ;
  assign n7456 = ( n7453 & ~n7060 ) | ( n7453 & n7454 ) | ( ~n7060 & n7454 ) ;
  assign n7455 = ( n7056 & ~n7454 ) | ( n7056 & n7453 ) | ( ~n7454 & n7453 ) ;
  assign n7457 = ( n7047 & ~n7456 ) | ( n7047 & n7455 ) | ( ~n7456 & n7455 ) ;
  assign n7458 = n713 | n7430 ;
  assign n7459 = ( n7444 & ~n7458 ) | ( n7444 & 1'b0 ) | ( ~n7458 & 1'b0 ) ;
  assign n7460 = n7450 | n7459 ;
  assign n7461 = n7438 &  n7441 ;
  assign n7462 = ( n7435 & ~n837 ) | ( n7435 & n7461 ) | ( ~n837 & n7461 ) ;
  assign n7463 = ( n713 & ~n7462 ) | ( n713 & 1'b0 ) | ( ~n7462 & 1'b0 ) ;
  assign n7464 = n595 | n7463 ;
  assign n7465 = ( n7460 & ~n7464 ) | ( n7460 & 1'b0 ) | ( ~n7464 & 1'b0 ) ;
  assign n7466 = ( n7457 & ~n7465 ) | ( n7457 & 1'b0 ) | ( ~n7465 & 1'b0 ) ;
  assign n7467 = n7452 | n7466 ;
  assign n7468 = n7062 | n7169 ;
  assign n7469 = ( n7049 & ~n7169 ) | ( n7049 & n7054 ) | ( ~n7169 & n7054 ) ;
  assign n7470 = ( n7169 & n7468 ) | ( n7169 & n7469 ) | ( n7468 & n7469 ) ;
  assign n7471 = ( n7049 & ~n7469 ) | ( n7049 & n7468 ) | ( ~n7469 & n7468 ) ;
  assign n7472 = ( n7054 & ~n7470 ) | ( n7054 & n7471 ) | ( ~n7470 & n7471 ) ;
  assign n7473 = ( n492 & n7467 ) | ( n492 & n7472 ) | ( n7467 & n7472 ) ;
  assign n7474 = n396 &  n7473 ;
  assign n7475 = ~n7082 & n7169 ;
  assign n7476 = ( n7069 & n7078 ) | ( n7069 & n7082 ) | ( n7078 & n7082 ) ;
  assign n7478 = ( n7475 & ~n7082 ) | ( n7475 & n7476 ) | ( ~n7082 & n7476 ) ;
  assign n7477 = ( n7078 & ~n7476 ) | ( n7078 & n7475 ) | ( ~n7476 & n7475 ) ;
  assign n7479 = ( n7069 & ~n7478 ) | ( n7069 & n7477 ) | ( ~n7478 & n7477 ) ;
  assign n7480 = n492 | n7452 ;
  assign n7481 = n7466 | n7480 ;
  assign n7482 = n7472 &  n7481 ;
  assign n7483 = ( n7460 & ~n7463 ) | ( n7460 & 1'b0 ) | ( ~n7463 & 1'b0 ) ;
  assign n7484 = ( n595 & ~n7483 ) | ( n595 & n7457 ) | ( ~n7483 & n7457 ) ;
  assign n7485 = n492 &  n7484 ;
  assign n7486 = n396 | n7485 ;
  assign n7487 = n7482 | n7486 ;
  assign n7488 = n7479 &  n7487 ;
  assign n7489 = n7474 | n7488 ;
  assign n7495 = ( n315 & ~n7494 ) | ( n315 & n7489 ) | ( ~n7494 & n7489 ) ;
  assign n7496 = n240 &  n7495 ;
  assign n7497 = ~n7104 & n7169 ;
  assign n7498 = ( n7091 & n7100 ) | ( n7091 & n7104 ) | ( n7100 & n7104 ) ;
  assign n7500 = ( n7497 & ~n7104 ) | ( n7497 & n7498 ) | ( ~n7104 & n7498 ) ;
  assign n7499 = ( n7100 & ~n7498 ) | ( n7100 & n7497 ) | ( ~n7498 & n7497 ) ;
  assign n7501 = ( n7091 & ~n7500 ) | ( n7091 & n7499 ) | ( ~n7500 & n7499 ) ;
  assign n7502 = n315 | n7474 ;
  assign n7503 = n7488 | n7502 ;
  assign n7504 = ~n7494 & n7503 ;
  assign n7505 = n7482 | n7485 ;
  assign n7506 = ( n396 & n7479 ) | ( n396 & n7505 ) | ( n7479 & n7505 ) ;
  assign n7507 = n315 &  n7506 ;
  assign n7508 = n240 | n7507 ;
  assign n7509 = n7504 | n7508 ;
  assign n7510 = n7501 &  n7509 ;
  assign n7511 = n7496 | n7510 ;
  assign n7512 = n7106 | n7169 ;
  assign n7513 = ( n7098 & ~n7093 ) | ( n7098 & n7169 ) | ( ~n7093 & n7169 ) ;
  assign n7515 = ( n7093 & n7512 ) | ( n7093 & n7513 ) | ( n7512 & n7513 ) ;
  assign n7514 = ( n7169 & ~n7513 ) | ( n7169 & n7512 ) | ( ~n7513 & n7512 ) ;
  assign n7516 = ( n7098 & ~n7515 ) | ( n7098 & n7514 ) | ( ~n7515 & n7514 ) ;
  assign n7517 = ( n181 & n7511 ) | ( n181 & n7516 ) | ( n7511 & n7516 ) ;
  assign n7518 = ~n145 & n7517 ;
  assign n7520 = ( n7122 & ~n7113 ) | ( n7122 & n7126 ) | ( ~n7113 & n7126 ) ;
  assign n7519 = ~n7126 & n7169 ;
  assign n7521 = ( n7122 & ~n7520 ) | ( n7122 & n7519 ) | ( ~n7520 & n7519 ) ;
  assign n7522 = ( n7519 & ~n7126 ) | ( n7519 & n7520 ) | ( ~n7126 & n7520 ) ;
  assign n7523 = ( n7113 & ~n7521 ) | ( n7113 & n7522 ) | ( ~n7521 & n7522 ) ;
  assign n7524 = n181 | n7496 ;
  assign n7525 = n7510 | n7524 ;
  assign n7526 = n7516 &  n7525 ;
  assign n7527 = n7504 | n7507 ;
  assign n7528 = ( n240 & n7501 ) | ( n240 & n7527 ) | ( n7501 & n7527 ) ;
  assign n7529 = n181 &  n7528 ;
  assign n7530 = ( n145 & ~n7529 ) | ( n145 & 1'b0 ) | ( ~n7529 & 1'b0 ) ;
  assign n7531 = ~n7526 & n7530 ;
  assign n7532 = ( n7523 & ~n7531 ) | ( n7523 & 1'b0 ) | ( ~n7531 & 1'b0 ) ;
  assign n7533 = n7518 | n7532 ;
  assign n7539 = ( n150 & ~n7538 ) | ( n150 & n7533 ) | ( ~n7538 & n7533 ) ;
  assign n7540 = ~n7135 & n7151 ;
  assign n7541 = ( n7154 & ~n7169 ) | ( n7154 & n7540 ) | ( ~n7169 & n7540 ) ;
  assign n7542 = ~n7154 & n7541 ;
  assign n7543 = ( n7151 & ~n7154 ) | ( n7151 & 1'b0 ) | ( ~n7154 & 1'b0 ) ;
  assign n7544 = n7169 &  n7543 ;
  assign n7545 = ( n7135 & ~n7543 ) | ( n7135 & n7544 ) | ( ~n7543 & n7544 ) ;
  assign n7546 = n7542 | n7545 ;
  assign n7547 = n7136 &  n7143 ;
  assign n7548 = n7169 &  n7547 ;
  assign n7549 = ( n7157 & ~n7547 ) | ( n7157 & n7548 ) | ( ~n7547 & n7548 ) ;
  assign n7550 = n7546 &  n7549 ;
  assign n7551 = ~n7539 & n7550 ;
  assign n7552 = ( n133 & ~n7551 ) | ( n133 & n7550 ) | ( ~n7551 & n7550 ) ;
  assign n7555 = n7526 | n7529 ;
  assign n7556 = ( n7523 & ~n145 ) | ( n7523 & n7555 ) | ( ~n145 & n7555 ) ;
  assign n7557 = n150 &  n7556 ;
  assign n7558 = n7546 | n7557 ;
  assign n7553 = n150 | n7518 ;
  assign n7554 = n7532 | n7553 ;
  assign n7559 = n7538 | n7554 ;
  assign n7560 = ( n7558 & ~n7538 ) | ( n7558 & n7559 ) | ( ~n7538 & n7559 ) ;
  assign n7562 = ( n133 & n7136 ) | ( n133 & n7143 ) | ( n7136 & n7143 ) ;
  assign n7561 = ( n7136 & n7143 ) | ( n7136 & n7169 ) | ( n7143 & n7169 ) ;
  assign n7563 = ( n7143 & ~n7561 ) | ( n7143 & 1'b0 ) | ( ~n7561 & 1'b0 ) ;
  assign n7564 = ( n7562 & ~n7143 ) | ( n7562 & n7563 ) | ( ~n7143 & n7563 ) ;
  assign n7565 = n7139 | n7166 ;
  assign n7566 = ( n7161 & ~n7142 ) | ( n7161 & n7565 ) | ( ~n7142 & n7565 ) ;
  assign n7567 = n7142 | n7566 ;
  assign n7568 = ( n7149 & ~n7157 ) | ( n7149 & n7567 ) | ( ~n7157 & n7567 ) ;
  assign n7569 = ( n7149 & ~n7568 ) | ( n7149 & 1'b0 ) | ( ~n7568 & 1'b0 ) ;
  assign n7570 = n7564 | n7569 ;
  assign n7571 = ( n7560 & ~n7570 ) | ( n7560 & 1'b0 ) | ( ~n7570 & 1'b0 ) ;
  assign n7572 = n7552 &  n7571 ;
  assign n7644 = ~n7244 & n7572 ;
  assign n7646 = ( n7240 & ~n7645 ) | ( n7240 & n7644 ) | ( ~n7645 & n7644 ) ;
  assign n7647 = ( n7644 & ~n7244 ) | ( n7644 & n7645 ) | ( ~n7244 & n7645 ) ;
  assign n7648 = ( n7231 & ~n7646 ) | ( n7231 & n7647 ) | ( ~n7646 & n7647 ) ;
  assign n7637 = ~n7211 & n7572 ;
  assign n7638 = ( n7211 & ~n7224 ) | ( n7211 & n7216 ) | ( ~n7224 & n7216 ) ;
  assign n7639 = ( n7224 & ~n7637 ) | ( n7224 & n7638 ) | ( ~n7637 & n7638 ) ;
  assign n7640 = ( n7637 & ~n7211 ) | ( n7637 & n7638 ) | ( ~n7211 & n7638 ) ;
  assign n7641 = ( n7639 & ~n7216 ) | ( n7639 & n7640 ) | ( ~n7216 & n7640 ) ;
  assign n7622 = ~n7222 & n7572 ;
  assign n7623 = ( n7209 & n7218 ) | ( n7209 & n7222 ) | ( n7218 & n7222 ) ;
  assign n7625 = ( n7622 & ~n7222 ) | ( n7622 & n7623 ) | ( ~n7222 & n7623 ) ;
  assign n7624 = ( n7218 & ~n7623 ) | ( n7218 & n7622 ) | ( ~n7623 & n7622 ) ;
  assign n7626 = ( n7209 & ~n7625 ) | ( n7209 & n7624 ) | ( ~n7625 & n7624 ) ;
  assign n7615 = ( n7185 & ~n7187 ) | ( n7185 & 1'b0 ) | ( ~n7187 & 1'b0 ) ;
  assign n7616 = ( n7197 & ~n7187 ) | ( n7197 & n7615 ) | ( ~n7187 & n7615 ) ;
  assign n7617 = ( n7187 & ~n7572 ) | ( n7187 & n7616 ) | ( ~n7572 & n7616 ) ;
  assign n7618 = ( n7572 & ~n7615 ) | ( n7572 & n7616 ) | ( ~n7615 & n7616 ) ;
  assign n7619 = ( n7617 & ~n7197 ) | ( n7617 & n7618 ) | ( ~n7197 & n7618 ) ;
  assign n7596 = ( x58 & ~n7180 ) | ( x58 & n7169 ) | ( ~n7180 & n7169 ) ;
  assign n7597 = ( x58 & ~n7596 ) | ( x58 & 1'b0 ) | ( ~n7596 & 1'b0 ) ;
  assign n7598 = ( n7175 & ~n7597 ) | ( n7175 & n7180 ) | ( ~n7597 & n7180 ) ;
  assign n7599 = x58 | n7169 ;
  assign n7600 = x59 &  n7599 ;
  assign n7601 = ( n7188 & ~n7600 ) | ( n7188 & 1'b0 ) | ( ~n7600 & 1'b0 ) ;
  assign n7602 = ( n7598 & ~n7572 ) | ( n7598 & n7601 ) | ( ~n7572 & n7601 ) ;
  assign n7603 = ~n7598 & n7602 ;
  assign n7604 = n7572 | n7602 ;
  assign n7605 = ( n7603 & ~n7601 ) | ( n7603 & n7604 ) | ( ~n7601 & n7604 ) ;
  assign n7584 = n7172 | n7572 ;
  assign n7585 = n7169 | n7569 ;
  assign n7586 = ( n7560 & n7564 ) | ( n7560 & n7585 ) | ( n7564 & n7585 ) ;
  assign n7587 = ( n7560 & ~n7586 ) | ( n7560 & 1'b0 ) | ( ~n7586 & 1'b0 ) ;
  assign n7588 = n7552 &  n7587 ;
  assign n7589 = n7584 | n7588 ;
  assign n7590 = ( x58 & ~n7589 ) | ( x58 & n7588 ) | ( ~n7589 & n7588 ) ;
  assign n7591 = x58 | n7588 ;
  assign n7592 = ( n7584 & ~n7591 ) | ( n7584 & 1'b0 ) | ( ~n7591 & 1'b0 ) ;
  assign n7593 = n7590 | n7592 ;
  assign n7170 = x54 | x55 ;
  assign n7576 = ~x56 & n7170 ;
  assign n7577 = ( x56 & ~n7167 ) | ( x56 & n7576 ) | ( ~n7167 & n7576 ) ;
  assign n7578 = ( n7157 & ~n7149 ) | ( n7157 & n7577 ) | ( ~n7149 & n7577 ) ;
  assign n7579 = n7149 &  n7578 ;
  assign n7580 = ( x57 & ~n7579 ) | ( x57 & n7572 ) | ( ~n7579 & n7572 ) ;
  assign n7575 = ( x56 & x57 ) | ( x56 & n7572 ) | ( x57 & n7572 ) ;
  assign n7581 = ( x56 & ~x57 ) | ( x56 & 1'b0 ) | ( ~x57 & 1'b0 ) ;
  assign n7582 = ( n7580 & ~n7575 ) | ( n7580 & n7581 ) | ( ~n7575 & n7581 ) ;
  assign n7573 = ( x56 & ~n7572 ) | ( x56 & 1'b0 ) | ( ~n7572 & 1'b0 ) ;
  assign n7171 = x56 | n7170 ;
  assign n7574 = ( n7169 & ~n7573 ) | ( n7169 & n7171 ) | ( ~n7573 & n7171 ) ;
  assign n7606 = ~n6781 & n7574 ;
  assign n7607 = ~n7582 & n7606 ;
  assign n7608 = ( n7593 & ~n7607 ) | ( n7593 & 1'b0 ) | ( ~n7607 & 1'b0 ) ;
  assign n7609 = n7574 | n7582 ;
  assign n7610 = ( n6781 & ~n7609 ) | ( n6781 & n7582 ) | ( ~n7609 & n7582 ) ;
  assign n7611 = ( n6399 & ~n7610 ) | ( n6399 & 1'b0 ) | ( ~n7610 & 1'b0 ) ;
  assign n7612 = ~n7608 & n7611 ;
  assign n7613 = n7605 | n7612 ;
  assign n7583 = ( n7574 & ~n7582 ) | ( n7574 & 1'b0 ) | ( ~n7582 & 1'b0 ) ;
  assign n7594 = ( n6781 & ~n7583 ) | ( n6781 & n7593 ) | ( ~n7583 & n7593 ) ;
  assign n7595 = ~n6399 & n7594 ;
  assign n7627 = n6032 | n7595 ;
  assign n7628 = ( n7613 & ~n7627 ) | ( n7613 & 1'b0 ) | ( ~n7627 & 1'b0 ) ;
  assign n7629 = n7619 | n7628 ;
  assign n7630 = n7608 | n7610 ;
  assign n7631 = ( n6399 & ~n7630 ) | ( n6399 & n7605 ) | ( ~n7630 & n7605 ) ;
  assign n7632 = ( n6032 & ~n7631 ) | ( n6032 & 1'b0 ) | ( ~n7631 & 1'b0 ) ;
  assign n7633 = ( n5672 & ~n7632 ) | ( n5672 & 1'b0 ) | ( ~n7632 & 1'b0 ) ;
  assign n7634 = n7629 &  n7633 ;
  assign n7635 = n7626 | n7634 ;
  assign n7614 = ~n7595 & n7613 ;
  assign n7620 = ( n7614 & ~n6032 ) | ( n7614 & n7619 ) | ( ~n6032 & n7619 ) ;
  assign n7621 = n5672 | n7620 ;
  assign n7649 = ~n5327 & n7621 ;
  assign n7650 = n7635 &  n7649 ;
  assign n7651 = n7641 | n7650 ;
  assign n7652 = ( n7629 & ~n7632 ) | ( n7629 & 1'b0 ) | ( ~n7632 & 1'b0 ) ;
  assign n7653 = ( n5672 & n7626 ) | ( n5672 & n7652 ) | ( n7626 & n7652 ) ;
  assign n7654 = ( n5327 & ~n7653 ) | ( n5327 & 1'b0 ) | ( ~n7653 & 1'b0 ) ;
  assign n7655 = n4990 | n7654 ;
  assign n7656 = ( n7651 & ~n7655 ) | ( n7651 & 1'b0 ) | ( ~n7655 & 1'b0 ) ;
  assign n7636 = n7621 &  n7635 ;
  assign n7642 = ( n7636 & ~n5327 ) | ( n7636 & n7641 ) | ( ~n5327 & n7641 ) ;
  assign n7643 = ( n4990 & ~n7642 ) | ( n4990 & 1'b0 ) | ( ~n7642 & 1'b0 ) ;
  assign n7944 = ~n7518 & n7572 ;
  assign n7945 = ( n7523 & ~n7518 ) | ( n7523 & n7531 ) | ( ~n7518 & n7531 ) ;
  assign n7946 = ( n7944 & ~n7531 ) | ( n7944 & n7945 ) | ( ~n7531 & n7945 ) ;
  assign n7947 = ( n7518 & ~n7944 ) | ( n7518 & n7945 ) | ( ~n7944 & n7945 ) ;
  assign n7948 = ( n7946 & ~n7523 ) | ( n7946 & n7947 ) | ( ~n7523 & n7947 ) ;
  assign n7878 = ( n7465 & ~n7572 ) | ( n7465 & 1'b0 ) | ( ~n7572 & 1'b0 ) ;
  assign n7879 = ( n7452 & ~n7572 ) | ( n7452 & n7457 ) | ( ~n7572 & n7457 ) ;
  assign n7880 = ( n7572 & ~n7878 ) | ( n7572 & n7879 ) | ( ~n7878 & n7879 ) ;
  assign n7881 = ( n7878 & ~n7452 ) | ( n7878 & n7879 ) | ( ~n7452 & n7879 ) ;
  assign n7882 = ( n7880 & ~n7457 ) | ( n7880 & n7881 ) | ( ~n7457 & n7881 ) ;
  assign n7834 = ~n7572 & n7421 ;
  assign n7835 = ( n7834 & ~n7408 ) | ( n7834 & n7572 ) | ( ~n7408 & n7572 ) ;
  assign n7837 = ( n7408 & n7413 ) | ( n7408 & n7835 ) | ( n7413 & n7835 ) ;
  assign n7836 = ( n7408 & ~n7413 ) | ( n7408 & n7835 ) | ( ~n7413 & n7835 ) ;
  assign n7838 = ( n7413 & ~n7837 ) | ( n7413 & n7836 ) | ( ~n7837 & n7836 ) ;
  assign n7660 = ( n7233 & ~n7238 ) | ( n7233 & n7246 ) | ( ~n7238 & n7246 ) ;
  assign n7659 = ~n7233 & n7572 ;
  assign n7661 = ( n7246 & ~n7660 ) | ( n7246 & n7659 ) | ( ~n7660 & n7659 ) ;
  assign n7662 = ( n7659 & ~n7233 ) | ( n7659 & n7660 ) | ( ~n7233 & n7660 ) ;
  assign n7663 = ( n7238 & ~n7661 ) | ( n7238 & n7662 ) | ( ~n7661 & n7662 ) ;
  assign n7657 = ( n7648 & ~n7656 ) | ( n7648 & 1'b0 ) | ( ~n7656 & 1'b0 ) ;
  assign n7658 = n7643 | n7657 ;
  assign n7664 = ( n4668 & ~n7663 ) | ( n4668 & n7658 ) | ( ~n7663 & n7658 ) ;
  assign n7665 = n4353 &  n7664 ;
  assign n7666 = n4668 | n7643 ;
  assign n7667 = n7657 | n7666 ;
  assign n7668 = ~n7663 & n7667 ;
  assign n7669 = ( n7651 & ~n7654 ) | ( n7651 & 1'b0 ) | ( ~n7654 & 1'b0 ) ;
  assign n7670 = ( n4990 & ~n7669 ) | ( n4990 & n7648 ) | ( ~n7669 & n7648 ) ;
  assign n7671 = n4668 &  n7670 ;
  assign n7672 = n4353 | n7671 ;
  assign n7673 = n7668 | n7672 ;
  assign n7674 = ( n7252 & n7261 ) | ( n7252 & n7265 ) | ( n7261 & n7265 ) ;
  assign n7676 = ( n7572 & ~n7265 ) | ( n7572 & n7674 ) | ( ~n7265 & n7674 ) ;
  assign n7675 = ( n7261 & ~n7674 ) | ( n7261 & n7572 ) | ( ~n7674 & n7572 ) ;
  assign n7677 = ( n7252 & ~n7676 ) | ( n7252 & n7675 ) | ( ~n7676 & n7675 ) ;
  assign n7678 = ( n7673 & ~n7677 ) | ( n7673 & 1'b0 ) | ( ~n7677 & 1'b0 ) ;
  assign n7679 = n7665 | n7678 ;
  assign n7680 = n7267 | n7572 ;
  assign n7681 = ( n7254 & ~n7572 ) | ( n7254 & n7259 ) | ( ~n7572 & n7259 ) ;
  assign n7682 = ( n7572 & n7680 ) | ( n7572 & n7681 ) | ( n7680 & n7681 ) ;
  assign n7683 = ( n7254 & ~n7681 ) | ( n7254 & n7680 ) | ( ~n7681 & n7680 ) ;
  assign n7684 = ( n7259 & ~n7682 ) | ( n7259 & n7683 ) | ( ~n7682 & n7683 ) ;
  assign n7685 = ( n4053 & n7679 ) | ( n4053 & n7684 ) | ( n7679 & n7684 ) ;
  assign n7686 = n3760 &  n7685 ;
  assign n7688 = ( n7283 & ~n7274 ) | ( n7283 & n7287 ) | ( ~n7274 & n7287 ) ;
  assign n7687 = ~n7287 & n7572 ;
  assign n7689 = ( n7283 & ~n7688 ) | ( n7283 & n7687 ) | ( ~n7688 & n7687 ) ;
  assign n7690 = ( n7687 & ~n7287 ) | ( n7687 & n7688 ) | ( ~n7287 & n7688 ) ;
  assign n7691 = ( n7274 & ~n7689 ) | ( n7274 & n7690 ) | ( ~n7689 & n7690 ) ;
  assign n7692 = n4053 | n7665 ;
  assign n7693 = n7678 | n7692 ;
  assign n7694 = n7684 &  n7693 ;
  assign n7695 = n7668 | n7671 ;
  assign n7696 = ( n4353 & ~n7677 ) | ( n4353 & n7695 ) | ( ~n7677 & n7695 ) ;
  assign n7697 = n4053 &  n7696 ;
  assign n7698 = n3760 | n7697 ;
  assign n7699 = n7694 | n7698 ;
  assign n7700 = ~n7691 & n7699 ;
  assign n7701 = n7686 | n7700 ;
  assign n7702 = n7289 | n7572 ;
  assign n7703 = ( n7276 & ~n7572 ) | ( n7276 & n7281 ) | ( ~n7572 & n7281 ) ;
  assign n7704 = ( n7572 & n7702 ) | ( n7572 & n7703 ) | ( n7702 & n7703 ) ;
  assign n7705 = ( n7276 & ~n7703 ) | ( n7276 & n7702 ) | ( ~n7703 & n7702 ) ;
  assign n7706 = ( n7281 & ~n7704 ) | ( n7281 & n7705 ) | ( ~n7704 & n7705 ) ;
  assign n7707 = ( n3482 & n7701 ) | ( n3482 & n7706 ) | ( n7701 & n7706 ) ;
  assign n7708 = n3211 &  n7707 ;
  assign n7709 = ~n7309 & n7572 ;
  assign n7710 = ( n7296 & n7305 ) | ( n7296 & n7309 ) | ( n7305 & n7309 ) ;
  assign n7712 = ( n7709 & ~n7309 ) | ( n7709 & n7710 ) | ( ~n7309 & n7710 ) ;
  assign n7711 = ( n7305 & ~n7710 ) | ( n7305 & n7709 ) | ( ~n7710 & n7709 ) ;
  assign n7713 = ( n7296 & ~n7712 ) | ( n7296 & n7711 ) | ( ~n7712 & n7711 ) ;
  assign n7714 = n3482 | n7686 ;
  assign n7715 = n7700 | n7714 ;
  assign n7716 = n7706 &  n7715 ;
  assign n7717 = n7694 | n7697 ;
  assign n7718 = ( n3760 & ~n7691 ) | ( n3760 & n7717 ) | ( ~n7691 & n7717 ) ;
  assign n7719 = n3482 &  n7718 ;
  assign n7720 = n3211 | n7719 ;
  assign n7721 = n7716 | n7720 ;
  assign n7722 = n7713 &  n7721 ;
  assign n7723 = n7708 | n7722 ;
  assign n7725 = ( n7298 & ~n7572 ) | ( n7298 & n7303 ) | ( ~n7572 & n7303 ) ;
  assign n7724 = n7311 | n7572 ;
  assign n7726 = ( n7572 & n7725 ) | ( n7572 & n7724 ) | ( n7725 & n7724 ) ;
  assign n7727 = ( n7724 & ~n7725 ) | ( n7724 & n7298 ) | ( ~n7725 & n7298 ) ;
  assign n7728 = ( n7303 & ~n7726 ) | ( n7303 & n7727 ) | ( ~n7726 & n7727 ) ;
  assign n7729 = ( n2955 & n7723 ) | ( n2955 & n7728 ) | ( n7723 & n7728 ) ;
  assign n7730 = n2706 &  n7729 ;
  assign n7731 = ~n7331 & n7572 ;
  assign n7732 = ( n7318 & n7327 ) | ( n7318 & n7331 ) | ( n7327 & n7331 ) ;
  assign n7734 = ( n7731 & ~n7331 ) | ( n7731 & n7732 ) | ( ~n7331 & n7732 ) ;
  assign n7733 = ( n7327 & ~n7732 ) | ( n7327 & n7731 ) | ( ~n7732 & n7731 ) ;
  assign n7735 = ( n7318 & ~n7734 ) | ( n7318 & n7733 ) | ( ~n7734 & n7733 ) ;
  assign n7736 = n2955 | n7708 ;
  assign n7737 = n7722 | n7736 ;
  assign n7738 = n7728 &  n7737 ;
  assign n7739 = n7716 | n7719 ;
  assign n7740 = ( n3211 & n7713 ) | ( n3211 & n7739 ) | ( n7713 & n7739 ) ;
  assign n7741 = n2955 &  n7740 ;
  assign n7742 = n2706 | n7741 ;
  assign n7743 = n7738 | n7742 ;
  assign n7744 = n7735 &  n7743 ;
  assign n7745 = n7730 | n7744 ;
  assign n7746 = n7333 | n7572 ;
  assign n7747 = ( n7320 & ~n7572 ) | ( n7320 & n7746 ) | ( ~n7572 & n7746 ) ;
  assign n7748 = ( n7320 & ~n7747 ) | ( n7320 & n7325 ) | ( ~n7747 & n7325 ) ;
  assign n7749 = ( n7325 & ~n7320 ) | ( n7325 & n7747 ) | ( ~n7320 & n7747 ) ;
  assign n7750 = ( n7748 & ~n7325 ) | ( n7748 & n7749 ) | ( ~n7325 & n7749 ) ;
  assign n7751 = ( n2472 & n7745 ) | ( n2472 & n7750 ) | ( n7745 & n7750 ) ;
  assign n7752 = n2245 &  n7751 ;
  assign n7753 = ~n7353 & n7572 ;
  assign n7754 = ( n7340 & n7349 ) | ( n7340 & n7353 ) | ( n7349 & n7353 ) ;
  assign n7756 = ( n7753 & ~n7353 ) | ( n7753 & n7754 ) | ( ~n7353 & n7754 ) ;
  assign n7755 = ( n7349 & ~n7754 ) | ( n7349 & n7753 ) | ( ~n7754 & n7753 ) ;
  assign n7757 = ( n7340 & ~n7756 ) | ( n7340 & n7755 ) | ( ~n7756 & n7755 ) ;
  assign n7758 = n2472 | n7730 ;
  assign n7759 = n7744 | n7758 ;
  assign n7760 = n7750 &  n7759 ;
  assign n7761 = n7738 | n7741 ;
  assign n7762 = ( n2706 & n7735 ) | ( n2706 & n7761 ) | ( n7735 & n7761 ) ;
  assign n7763 = n2472 &  n7762 ;
  assign n7764 = n2245 | n7763 ;
  assign n7765 = n7760 | n7764 ;
  assign n7766 = n7757 &  n7765 ;
  assign n7767 = n7752 | n7766 ;
  assign n7768 = n7355 | n7572 ;
  assign n7769 = ( n7347 & ~n7342 ) | ( n7347 & n7572 ) | ( ~n7342 & n7572 ) ;
  assign n7771 = ( n7768 & n7342 ) | ( n7768 & n7769 ) | ( n7342 & n7769 ) ;
  assign n7770 = ( n7572 & ~n7769 ) | ( n7572 & n7768 ) | ( ~n7769 & n7768 ) ;
  assign n7772 = ( n7347 & ~n7771 ) | ( n7347 & n7770 ) | ( ~n7771 & n7770 ) ;
  assign n7773 = ( n7767 & ~n2033 ) | ( n7767 & n7772 ) | ( ~n2033 & n7772 ) ;
  assign n7774 = n1827 &  n7773 ;
  assign n7775 = ~n7375 & n7572 ;
  assign n7776 = ( n7362 & ~n7371 ) | ( n7362 & n7375 ) | ( ~n7371 & n7375 ) ;
  assign n7777 = ( n7371 & ~n7775 ) | ( n7371 & n7776 ) | ( ~n7775 & n7776 ) ;
  assign n7778 = ( n7775 & ~n7375 ) | ( n7775 & n7776 ) | ( ~n7375 & n7776 ) ;
  assign n7779 = ( n7777 & ~n7362 ) | ( n7777 & n7778 ) | ( ~n7362 & n7778 ) ;
  assign n7780 = ( n2033 & ~n7752 ) | ( n2033 & 1'b0 ) | ( ~n7752 & 1'b0 ) ;
  assign n7781 = ~n7766 & n7780 ;
  assign n7782 = ( n7772 & ~n7781 ) | ( n7772 & 1'b0 ) | ( ~n7781 & 1'b0 ) ;
  assign n7783 = n7760 | n7763 ;
  assign n7784 = ( n2245 & n7757 ) | ( n2245 & n7783 ) | ( n7757 & n7783 ) ;
  assign n7785 = ~n2033 & n7784 ;
  assign n7786 = n1827 | n7785 ;
  assign n7787 = n7782 | n7786 ;
  assign n7788 = ~n7779 & n7787 ;
  assign n7789 = n7774 | n7788 ;
  assign n7790 = n7377 | n7572 ;
  assign n7791 = ( n7364 & ~n7572 ) | ( n7364 & n7790 ) | ( ~n7572 & n7790 ) ;
  assign n7792 = ( n7369 & ~n7364 ) | ( n7369 & n7791 ) | ( ~n7364 & n7791 ) ;
  assign n7793 = ( n7364 & ~n7791 ) | ( n7364 & n7369 ) | ( ~n7791 & n7369 ) ;
  assign n7794 = ( n7792 & ~n7369 ) | ( n7792 & n7793 ) | ( ~n7369 & n7793 ) ;
  assign n7795 = ( n1636 & ~n7789 ) | ( n1636 & n7794 ) | ( ~n7789 & n7794 ) ;
  assign n7796 = n1452 | n7795 ;
  assign n7797 = ~n7397 & n7572 ;
  assign n7798 = ( n7384 & ~n7393 ) | ( n7384 & n7397 ) | ( ~n7393 & n7397 ) ;
  assign n7799 = ( n7393 & ~n7797 ) | ( n7393 & n7798 ) | ( ~n7797 & n7798 ) ;
  assign n7800 = ( n7797 & ~n7397 ) | ( n7797 & n7798 ) | ( ~n7397 & n7798 ) ;
  assign n7801 = ( n7799 & ~n7384 ) | ( n7799 & n7800 ) | ( ~n7384 & n7800 ) ;
  assign n7802 = ( n1636 & ~n7774 ) | ( n1636 & 1'b0 ) | ( ~n7774 & 1'b0 ) ;
  assign n7803 = ~n7788 & n7802 ;
  assign n7804 = n7794 | n7803 ;
  assign n7805 = n7782 | n7785 ;
  assign n7806 = ( n1827 & ~n7779 ) | ( n1827 & n7805 ) | ( ~n7779 & n7805 ) ;
  assign n7807 = ~n1636 & n7806 ;
  assign n7808 = ( n1452 & ~n7807 ) | ( n1452 & 1'b0 ) | ( ~n7807 & 1'b0 ) ;
  assign n7809 = n7804 &  n7808 ;
  assign n7810 = n7801 | n7809 ;
  assign n7811 = n7796 &  n7810 ;
  assign n7812 = ( n7399 & ~n7572 ) | ( n7399 & 1'b0 ) | ( ~n7572 & 1'b0 ) ;
  assign n7813 = ( n7391 & ~n7386 ) | ( n7391 & n7572 ) | ( ~n7386 & n7572 ) ;
  assign n7814 = ( n7812 & ~n7572 ) | ( n7812 & n7813 ) | ( ~n7572 & n7813 ) ;
  assign n7815 = ( n7386 & ~n7812 ) | ( n7386 & n7813 ) | ( ~n7812 & n7813 ) ;
  assign n7816 = ( n7814 & ~n7391 ) | ( n7814 & n7815 ) | ( ~n7391 & n7815 ) ;
  assign n7817 = ( n7811 & ~n1283 ) | ( n7811 & n7816 ) | ( ~n1283 & n7816 ) ;
  assign n7818 = n1122 | n7817 ;
  assign n7819 = ~n7419 & n7572 ;
  assign n7820 = ( n7406 & n7415 ) | ( n7406 & n7419 ) | ( n7415 & n7419 ) ;
  assign n7822 = ( n7819 & ~n7419 ) | ( n7819 & n7820 ) | ( ~n7419 & n7820 ) ;
  assign n7821 = ( n7415 & ~n7820 ) | ( n7415 & n7819 ) | ( ~n7820 & n7819 ) ;
  assign n7823 = ( n7406 & ~n7822 ) | ( n7406 & n7821 ) | ( ~n7822 & n7821 ) ;
  assign n7824 = ~n1283 & n7796 ;
  assign n7825 = n7810 &  n7824 ;
  assign n7826 = n7816 | n7825 ;
  assign n7827 = ( n7804 & ~n7807 ) | ( n7804 & 1'b0 ) | ( ~n7807 & 1'b0 ) ;
  assign n7828 = ( n1452 & n7801 ) | ( n1452 & n7827 ) | ( n7801 & n7827 ) ;
  assign n7829 = ( n1283 & ~n7828 ) | ( n1283 & 1'b0 ) | ( ~n7828 & 1'b0 ) ;
  assign n7830 = ( n1122 & ~n7829 ) | ( n1122 & 1'b0 ) | ( ~n7829 & 1'b0 ) ;
  assign n7831 = n7826 &  n7830 ;
  assign n7832 = ( n7823 & ~n7831 ) | ( n7823 & 1'b0 ) | ( ~n7831 & 1'b0 ) ;
  assign n7833 = ( n7818 & ~n7832 ) | ( n7818 & 1'b0 ) | ( ~n7832 & 1'b0 ) ;
  assign n7839 = ( n976 & ~n7838 ) | ( n976 & n7833 ) | ( ~n7838 & n7833 ) ;
  assign n7840 = ( n837 & ~n7839 ) | ( n837 & 1'b0 ) | ( ~n7839 & 1'b0 ) ;
  assign n7841 = n7441 &  n7572 ;
  assign n7842 = ( n7428 & n7437 ) | ( n7428 & n7441 ) | ( n7437 & n7441 ) ;
  assign n7843 = ( n7841 & ~n7437 ) | ( n7841 & n7842 ) | ( ~n7437 & n7842 ) ;
  assign n7844 = ( n7441 & ~n7842 ) | ( n7441 & n7841 ) | ( ~n7842 & n7841 ) ;
  assign n7845 = ( n7428 & ~n7843 ) | ( n7428 & n7844 ) | ( ~n7843 & n7844 ) ;
  assign n7846 = n976 &  n7818 ;
  assign n7847 = ~n7832 & n7846 ;
  assign n7848 = ( n7838 & ~n7847 ) | ( n7838 & 1'b0 ) | ( ~n7847 & 1'b0 ) ;
  assign n7849 = ( n7826 & ~n7829 ) | ( n7826 & 1'b0 ) | ( ~n7829 & 1'b0 ) ;
  assign n7850 = ( n1122 & ~n7823 ) | ( n1122 & n7849 ) | ( ~n7823 & n7849 ) ;
  assign n7851 = n976 | n7850 ;
  assign n7852 = ~n837 & n7851 ;
  assign n7853 = ~n7848 & n7852 ;
  assign n7854 = n7845 | n7853 ;
  assign n7855 = ~n7840 & n7854 ;
  assign n7856 = ( n7443 & ~n7572 ) | ( n7443 & 1'b0 ) | ( ~n7572 & 1'b0 ) ;
  assign n7857 = ( n7430 & ~n7572 ) | ( n7430 & n7435 ) | ( ~n7572 & n7435 ) ;
  assign n7858 = ( n7572 & ~n7856 ) | ( n7572 & n7857 ) | ( ~n7856 & n7857 ) ;
  assign n7859 = ( n7856 & ~n7430 ) | ( n7856 & n7857 ) | ( ~n7430 & n7857 ) ;
  assign n7860 = ( n7858 & ~n7435 ) | ( n7858 & n7859 ) | ( ~n7435 & n7859 ) ;
  assign n7861 = ( n713 & ~n7855 ) | ( n713 & n7860 ) | ( ~n7855 & n7860 ) ;
  assign n7862 = n595 &  n7861 ;
  assign n7863 = ~n7463 & n7572 ;
  assign n7864 = ( n7450 & ~n7463 ) | ( n7450 & n7459 ) | ( ~n7463 & n7459 ) ;
  assign n7865 = ( n7863 & ~n7459 ) | ( n7863 & n7864 ) | ( ~n7459 & n7864 ) ;
  assign n7866 = ( n7463 & ~n7863 ) | ( n7463 & n7864 ) | ( ~n7863 & n7864 ) ;
  assign n7867 = ( n7865 & ~n7450 ) | ( n7865 & n7866 ) | ( ~n7450 & n7866 ) ;
  assign n7868 = n713 | n7840 ;
  assign n7869 = ( n7854 & ~n7868 ) | ( n7854 & 1'b0 ) | ( ~n7868 & 1'b0 ) ;
  assign n7870 = ( n7860 & ~n7869 ) | ( n7860 & 1'b0 ) | ( ~n7869 & 1'b0 ) ;
  assign n7871 = ~n7848 & n7851 ;
  assign n7872 = ( n7845 & ~n837 ) | ( n7845 & n7871 ) | ( ~n837 & n7871 ) ;
  assign n7873 = ( n713 & ~n7872 ) | ( n713 & 1'b0 ) | ( ~n7872 & 1'b0 ) ;
  assign n7874 = n595 | n7873 ;
  assign n7875 = n7870 | n7874 ;
  assign n7876 = n7867 &  n7875 ;
  assign n7877 = n7862 | n7876 ;
  assign n7883 = ( n492 & ~n7882 ) | ( n492 & n7877 ) | ( ~n7882 & n7877 ) ;
  assign n7884 = n396 &  n7883 ;
  assign n7885 = ~n7485 & n7572 ;
  assign n7886 = ( n7472 & n7481 ) | ( n7472 & n7485 ) | ( n7481 & n7485 ) ;
  assign n7888 = ( n7885 & ~n7485 ) | ( n7885 & n7886 ) | ( ~n7485 & n7886 ) ;
  assign n7887 = ( n7481 & ~n7886 ) | ( n7481 & n7885 ) | ( ~n7886 & n7885 ) ;
  assign n7889 = ( n7472 & ~n7888 ) | ( n7472 & n7887 ) | ( ~n7888 & n7887 ) ;
  assign n7890 = n492 | n7862 ;
  assign n7891 = n7876 | n7890 ;
  assign n7892 = ~n7882 & n7891 ;
  assign n7893 = n7870 | n7873 ;
  assign n7894 = ( n595 & n7867 ) | ( n595 & n7893 ) | ( n7867 & n7893 ) ;
  assign n7895 = n492 &  n7894 ;
  assign n7896 = n396 | n7895 ;
  assign n7897 = n7892 | n7896 ;
  assign n7898 = n7889 &  n7897 ;
  assign n7899 = n7884 | n7898 ;
  assign n7900 = n7487 | n7572 ;
  assign n7901 = ( n7479 & ~n7474 ) | ( n7479 & n7572 ) | ( ~n7474 & n7572 ) ;
  assign n7903 = ( n7900 & n7474 ) | ( n7900 & n7901 ) | ( n7474 & n7901 ) ;
  assign n7902 = ( n7572 & ~n7901 ) | ( n7572 & n7900 ) | ( ~n7901 & n7900 ) ;
  assign n7904 = ( n7479 & ~n7903 ) | ( n7479 & n7902 ) | ( ~n7903 & n7902 ) ;
  assign n7905 = ( n315 & n7899 ) | ( n315 & n7904 ) | ( n7899 & n7904 ) ;
  assign n7906 = n240 &  n7905 ;
  assign n7908 = ( n7503 & ~n7494 ) | ( n7503 & n7507 ) | ( ~n7494 & n7507 ) ;
  assign n7907 = ~n7507 & n7572 ;
  assign n7909 = ( n7503 & ~n7908 ) | ( n7503 & n7907 ) | ( ~n7908 & n7907 ) ;
  assign n7910 = ( n7907 & ~n7507 ) | ( n7907 & n7908 ) | ( ~n7507 & n7908 ) ;
  assign n7911 = ( n7494 & ~n7909 ) | ( n7494 & n7910 ) | ( ~n7909 & n7910 ) ;
  assign n7912 = n315 | n7884 ;
  assign n7913 = n7898 | n7912 ;
  assign n7914 = n7904 &  n7913 ;
  assign n7915 = n7892 | n7895 ;
  assign n7916 = ( n396 & n7889 ) | ( n396 & n7915 ) | ( n7889 & n7915 ) ;
  assign n7917 = n315 &  n7916 ;
  assign n7918 = n240 | n7917 ;
  assign n7919 = n7914 | n7918 ;
  assign n7920 = ~n7911 & n7919 ;
  assign n7921 = n7906 | n7920 ;
  assign n7922 = n7509 | n7572 ;
  assign n7923 = ( n7496 & ~n7572 ) | ( n7496 & n7501 ) | ( ~n7572 & n7501 ) ;
  assign n7924 = ( n7572 & n7922 ) | ( n7572 & n7923 ) | ( n7922 & n7923 ) ;
  assign n7925 = ( n7496 & ~n7923 ) | ( n7496 & n7922 ) | ( ~n7923 & n7922 ) ;
  assign n7926 = ( n7501 & ~n7924 ) | ( n7501 & n7925 ) | ( ~n7924 & n7925 ) ;
  assign n7927 = ( n181 & n7921 ) | ( n181 & n7926 ) | ( n7921 & n7926 ) ;
  assign n7928 = ~n145 & n7927 ;
  assign n7930 = ( n7525 & ~n7516 ) | ( n7525 & n7529 ) | ( ~n7516 & n7529 ) ;
  assign n7929 = ~n7529 & n7572 ;
  assign n7931 = ( n7525 & ~n7930 ) | ( n7525 & n7929 ) | ( ~n7930 & n7929 ) ;
  assign n7932 = ( n7929 & ~n7529 ) | ( n7929 & n7930 ) | ( ~n7529 & n7930 ) ;
  assign n7933 = ( n7516 & ~n7931 ) | ( n7516 & n7932 ) | ( ~n7931 & n7932 ) ;
  assign n7934 = n181 | n7906 ;
  assign n7935 = n7920 | n7934 ;
  assign n7936 = n7926 &  n7935 ;
  assign n7937 = n7914 | n7917 ;
  assign n7938 = ( n240 & ~n7911 ) | ( n240 & n7937 ) | ( ~n7911 & n7937 ) ;
  assign n7939 = n181 &  n7938 ;
  assign n7940 = ( n145 & ~n7939 ) | ( n145 & 1'b0 ) | ( ~n7939 & 1'b0 ) ;
  assign n7941 = ~n7936 & n7940 ;
  assign n7942 = ( n7933 & ~n7941 ) | ( n7933 & 1'b0 ) | ( ~n7941 & 1'b0 ) ;
  assign n7943 = n7928 | n7942 ;
  assign n7949 = ( n150 & ~n7948 ) | ( n150 & n7943 ) | ( ~n7948 & n7943 ) ;
  assign n7950 = ( n7538 & ~n7557 ) | ( n7538 & 1'b0 ) | ( ~n7557 & 1'b0 ) ;
  assign n7951 = ( n7554 & ~n7950 ) | ( n7554 & n7572 ) | ( ~n7950 & n7572 ) ;
  assign n7952 = ( n7554 & ~n7951 ) | ( n7554 & 1'b0 ) | ( ~n7951 & 1'b0 ) ;
  assign n7953 = ( n7554 & ~n7557 ) | ( n7554 & 1'b0 ) | ( ~n7557 & 1'b0 ) ;
  assign n7954 = n7572 &  n7953 ;
  assign n7955 = ( n7538 & ~n7954 ) | ( n7538 & n7953 ) | ( ~n7954 & n7953 ) ;
  assign n7956 = ~n7952 & n7955 ;
  assign n7957 = n7539 &  n7546 ;
  assign n7958 = n7572 &  n7957 ;
  assign n7959 = ( n7560 & ~n7957 ) | ( n7560 & n7958 ) | ( ~n7957 & n7958 ) ;
  assign n7960 = ~n7956 & n7959 ;
  assign n7961 = ~n7949 & n7960 ;
  assign n7962 = ( n133 & ~n7961 ) | ( n133 & n7960 ) | ( ~n7961 & n7960 ) ;
  assign n7963 = n150 | n7928 ;
  assign n7964 = n7942 | n7963 ;
  assign n7969 = n7948 | n7964 ;
  assign n7965 = n7936 | n7939 ;
  assign n7966 = ( n7933 & ~n145 ) | ( n7933 & n7965 ) | ( ~n145 & n7965 ) ;
  assign n7967 = n150 &  n7966 ;
  assign n7968 = ( n7956 & ~n7967 ) | ( n7956 & 1'b0 ) | ( ~n7967 & 1'b0 ) ;
  assign n7970 = ( n7948 & ~n7969 ) | ( n7948 & n7968 ) | ( ~n7969 & n7968 ) ;
  assign n7972 = ( n133 & n7539 ) | ( n133 & n7546 ) | ( n7539 & n7546 ) ;
  assign n7971 = ( n7539 & n7546 ) | ( n7539 & n7572 ) | ( n7546 & n7572 ) ;
  assign n7973 = ( n7546 & ~n7971 ) | ( n7546 & 1'b0 ) | ( ~n7971 & 1'b0 ) ;
  assign n7974 = ( n7972 & ~n7546 ) | ( n7972 & n7973 ) | ( ~n7546 & n7973 ) ;
  assign n7975 = n7542 | n7569 ;
  assign n7976 = ( n7564 & ~n7545 ) | ( n7564 & n7975 ) | ( ~n7545 & n7975 ) ;
  assign n7977 = n7545 | n7976 ;
  assign n7978 = ( n7552 & ~n7560 ) | ( n7552 & n7977 ) | ( ~n7560 & n7977 ) ;
  assign n7979 = ( n7552 & ~n7978 ) | ( n7552 & 1'b0 ) | ( ~n7978 & 1'b0 ) ;
  assign n7980 = n7974 | n7979 ;
  assign n7981 = n7970 | n7980 ;
  assign n7982 = ~n7962 |  n7981 ;
  assign n8084 = n7643 | n7982 ;
  assign n8085 = ( n7643 & ~n7656 ) | ( n7643 & n7648 ) | ( ~n7656 & n7648 ) ;
  assign n8086 = ( n7656 & n8084 ) | ( n7656 & n8085 ) | ( n8084 & n8085 ) ;
  assign n8087 = ( n7643 & ~n8085 ) | ( n7643 & n8084 ) | ( ~n8085 & n8084 ) ;
  assign n8088 = ( n7648 & ~n8086 ) | ( n7648 & n8087 ) | ( ~n8086 & n8087 ) ;
  assign n8069 = n7654 | n7982 ;
  assign n8070 = ( n7641 & ~n7650 ) | ( n7641 & n7654 ) | ( ~n7650 & n7654 ) ;
  assign n8071 = ( n7650 & n8069 ) | ( n7650 & n8070 ) | ( n8069 & n8070 ) ;
  assign n8072 = ( n7654 & ~n8070 ) | ( n7654 & n8069 ) | ( ~n8070 & n8069 ) ;
  assign n8073 = ( n7641 & ~n8071 ) | ( n7641 & n8072 ) | ( ~n8071 & n8072 ) ;
  assign n8062 = n7634 &  n7982 ;
  assign n8063 = ( n7621 & ~n7982 ) | ( n7621 & n8062 ) | ( ~n7982 & n8062 ) ;
  assign n8064 = ( n7621 & ~n8063 ) | ( n7621 & n7626 ) | ( ~n8063 & n7626 ) ;
  assign n8065 = ( n7626 & ~n7621 ) | ( n7626 & n8063 ) | ( ~n7621 & n8063 ) ;
  assign n8066 = ( n8064 & ~n7626 ) | ( n8064 & n8065 ) | ( ~n7626 & n8065 ) ;
  assign n8047 = n7632 | n7982 ;
  assign n8048 = ( n7619 & ~n7632 ) | ( n7619 & n7628 ) | ( ~n7632 & n7628 ) ;
  assign n8050 = ( n7632 & n8047 ) | ( n7632 & n8048 ) | ( n8047 & n8048 ) ;
  assign n8049 = ( n7628 & ~n8048 ) | ( n7628 & n8047 ) | ( ~n8048 & n8047 ) ;
  assign n8051 = ( n7619 & ~n8050 ) | ( n7619 & n8049 ) | ( ~n8050 & n8049 ) ;
  assign n8040 = n7612 &  n7982 ;
  assign n8041 = ( n7595 & n7605 ) | ( n7595 & n7982 ) | ( n7605 & n7982 ) ;
  assign n8043 = ( n8040 & ~n7595 ) | ( n8040 & n8041 ) | ( ~n7595 & n8041 ) ;
  assign n8042 = ( n7982 & ~n8041 ) | ( n7982 & n8040 ) | ( ~n8041 & n8040 ) ;
  assign n8044 = ( n7605 & ~n8043 ) | ( n7605 & n8042 ) | ( ~n8043 & n8042 ) ;
  assign n8025 = ~n7607 & n7610 ;
  assign n8026 = ( n7593 & ~n7607 ) | ( n7593 & n8025 ) | ( ~n7607 & n8025 ) ;
  assign n8028 = ( n7607 & n7982 ) | ( n7607 & n8026 ) | ( n7982 & n8026 ) ;
  assign n8027 = ( n7982 & ~n8026 ) | ( n7982 & n8025 ) | ( ~n8026 & n8025 ) ;
  assign n8029 = ( n7593 & ~n8028 ) | ( n7593 & n8027 ) | ( ~n8028 & n8027 ) ;
  assign n8016 = x56 | n7572 ;
  assign n8017 = x57 &  n8016 ;
  assign n8018 = ( n7584 & ~n8017 ) | ( n7584 & 1'b0 ) | ( ~n8017 & 1'b0 ) ;
  assign n8013 = ( x56 & ~n7579 ) | ( x56 & n7572 ) | ( ~n7579 & n7572 ) ;
  assign n8014 = ( x56 & ~n8013 ) | ( x56 & 1'b0 ) | ( ~n8013 & 1'b0 ) ;
  assign n8015 = ( n7574 & ~n7579 ) | ( n7574 & n8014 ) | ( ~n7579 & n8014 ) ;
  assign n8019 = ( n7982 & ~n8015 ) | ( n7982 & n8018 ) | ( ~n8015 & n8018 ) ;
  assign n8020 = n8015 &  n8019 ;
  assign n8021 = ( n7982 & ~n8019 ) | ( n7982 & 1'b0 ) | ( ~n8019 & 1'b0 ) ;
  assign n8022 = ( n8018 & ~n8020 ) | ( n8018 & n8021 ) | ( ~n8020 & n8021 ) ;
  assign n7989 = ( x54 & ~n7982 ) | ( x54 & x55 ) | ( ~n7982 & x55 ) ;
  assign n7995 = ( x54 & ~x55 ) | ( x54 & 1'b0 ) | ( ~x55 & 1'b0 ) ;
  assign n7985 = x52 | x53 ;
  assign n7990 = ~x54 & n7985 ;
  assign n7991 = ( x54 & ~n7570 ) | ( x54 & n7990 ) | ( ~n7570 & n7990 ) ;
  assign n7992 = ( n7560 & ~n7552 ) | ( n7560 & n7991 ) | ( ~n7552 & n7991 ) ;
  assign n7993 = n7552 &  n7992 ;
  assign n7994 = ( n7982 & ~x55 ) | ( n7982 & n7993 ) | ( ~x55 & n7993 ) ;
  assign n7996 = ( n7989 & ~n7995 ) | ( n7989 & n7994 ) | ( ~n7995 & n7994 ) ;
  assign n7987 = x54 &  n7982 ;
  assign n7986 = x54 | n7985 ;
  assign n7988 = ( n7572 & ~n7987 ) | ( n7572 & n7986 ) | ( ~n7987 & n7986 ) ;
  assign n7999 = n7169 &  n7988 ;
  assign n8000 = n7996 &  n7999 ;
  assign n8002 = n7572 | n7979 ;
  assign n8003 = ( n7974 & ~n7970 ) | ( n7974 & n8002 ) | ( ~n7970 & n8002 ) ;
  assign n8004 = n7970 | n8003 ;
  assign n8005 = ( n7962 & ~n8004 ) | ( n7962 & 1'b0 ) | ( ~n8004 & 1'b0 ) ;
  assign n8001 = ~n7170 & n7982 ;
  assign n8006 = ~n8005 & n8001 ;
  assign n8007 = ( x56 & n8006 ) | ( x56 & n8005 ) | ( n8006 & n8005 ) ;
  assign n8008 = x56 | n8005 ;
  assign n8009 = n8001 | n8008 ;
  assign n8010 = ~n8007 & n8009 ;
  assign n8011 = n8000 | n8010 ;
  assign n7997 = ~n7988 & n7996 ;
  assign n7998 = ( n7169 & ~n7997 ) | ( n7169 & n7996 ) | ( ~n7997 & n7996 ) ;
  assign n8030 = ~n6781 & n7998 ;
  assign n8031 = n8011 &  n8030 ;
  assign n8032 = ( n8022 & ~n8031 ) | ( n8022 & 1'b0 ) | ( ~n8031 & 1'b0 ) ;
  assign n8033 = n7988 &  n7996 ;
  assign n8034 = ( n7169 & n8010 ) | ( n7169 & n8033 ) | ( n8010 & n8033 ) ;
  assign n8035 = ( n6781 & ~n8034 ) | ( n6781 & 1'b0 ) | ( ~n8034 & 1'b0 ) ;
  assign n8036 = ( n6399 & ~n8035 ) | ( n6399 & 1'b0 ) | ( ~n8035 & 1'b0 ) ;
  assign n8037 = ~n8032 & n8036 ;
  assign n8038 = ( n8029 & ~n8037 ) | ( n8029 & 1'b0 ) | ( ~n8037 & 1'b0 ) ;
  assign n8012 = n7998 &  n8011 ;
  assign n8023 = ( n6781 & ~n8012 ) | ( n6781 & n8022 ) | ( ~n8012 & n8022 ) ;
  assign n8024 = ~n6399 & n8023 ;
  assign n8052 = n6032 | n8024 ;
  assign n8053 = n8038 | n8052 ;
  assign n8054 = ~n8044 & n8053 ;
  assign n8055 = n8032 | n8035 ;
  assign n8056 = ( n8029 & ~n6399 ) | ( n8029 & n8055 ) | ( ~n6399 & n8055 ) ;
  assign n8057 = n6032 &  n8056 ;
  assign n8058 = ( n5672 & ~n8057 ) | ( n5672 & 1'b0 ) | ( ~n8057 & 1'b0 ) ;
  assign n8059 = ~n8054 & n8058 ;
  assign n8060 = n8051 | n8059 ;
  assign n8039 = n8024 | n8038 ;
  assign n8045 = ( n6032 & ~n8044 ) | ( n6032 & n8039 ) | ( ~n8044 & n8039 ) ;
  assign n8046 = ~n5672 & n8045 ;
  assign n8074 = n5327 | n8046 ;
  assign n8075 = ( n8060 & ~n8074 ) | ( n8060 & 1'b0 ) | ( ~n8074 & 1'b0 ) ;
  assign n8076 = n8066 | n8075 ;
  assign n8077 = n8054 | n8057 ;
  assign n8078 = ( n5672 & ~n8077 ) | ( n5672 & n8051 ) | ( ~n8077 & n8051 ) ;
  assign n8079 = ( n5327 & ~n8078 ) | ( n5327 & 1'b0 ) | ( ~n8078 & 1'b0 ) ;
  assign n8080 = n4990 | n8079 ;
  assign n8081 = ( n8076 & ~n8080 ) | ( n8076 & 1'b0 ) | ( ~n8080 & 1'b0 ) ;
  assign n8082 = n8073 | n8081 ;
  assign n8061 = ~n8046 & n8060 ;
  assign n8067 = ( n8061 & ~n5327 ) | ( n8061 & n8066 ) | ( ~n5327 & n8066 ) ;
  assign n8068 = ( n4990 & ~n8067 ) | ( n4990 & 1'b0 ) | ( ~n8067 & 1'b0 ) ;
  assign n8096 = n4668 | n8068 ;
  assign n8097 = ( n8082 & ~n8096 ) | ( n8082 & 1'b0 ) | ( ~n8096 & 1'b0 ) ;
  assign n8099 = ( n8076 & ~n8079 ) | ( n8076 & 1'b0 ) | ( ~n8079 & 1'b0 ) ;
  assign n8100 = ( n8073 & ~n4990 ) | ( n8073 & n8099 ) | ( ~n4990 & n8099 ) ;
  assign n8101 = ( n4668 & ~n8100 ) | ( n4668 & 1'b0 ) | ( ~n8100 & 1'b0 ) ;
  assign n8375 = n7948 &  n7964 ;
  assign n8376 = ( n7967 & n7982 ) | ( n7967 & n8375 ) | ( n7982 & n8375 ) ;
  assign n8377 = ~n7967 & n8376 ;
  assign n8378 = ( n7964 & ~n7967 ) | ( n7964 & 1'b0 ) | ( ~n7967 & 1'b0 ) ;
  assign n8379 = ~n7982 & n8378 ;
  assign n8380 = ( n7948 & ~n8379 ) | ( n7948 & n8378 ) | ( ~n8379 & n8378 ) ;
  assign n8381 = ~n8377 & n8380 ;
  assign n8382 = ( n7949 & ~n7956 ) | ( n7949 & 1'b0 ) | ( ~n7956 & 1'b0 ) ;
  assign n8383 = ~n7982 & n8382 ;
  assign n8384 = ( n7970 & ~n8383 ) | ( n7970 & n8382 ) | ( ~n8383 & n8382 ) ;
  assign n8385 = n8381 | n8384 ;
  assign n8347 = ~n7919 & n7982 ;
  assign n8348 = ( n7906 & n7911 ) | ( n7906 & n7982 ) | ( n7911 & n7982 ) ;
  assign n8350 = ( n8347 & ~n7906 ) | ( n8347 & n8348 ) | ( ~n7906 & n8348 ) ;
  assign n8349 = ( n7982 & ~n8348 ) | ( n7982 & n8347 ) | ( ~n8348 & n8347 ) ;
  assign n8351 = ( n7911 & ~n8350 ) | ( n7911 & n8349 ) | ( ~n8350 & n8349 ) ;
  assign n8281 = n7853 &  n7982 ;
  assign n8282 = ( n7840 & n7845 ) | ( n7840 & n7982 ) | ( n7845 & n7982 ) ;
  assign n8284 = ( n8281 & ~n7840 ) | ( n8281 & n8282 ) | ( ~n7840 & n8282 ) ;
  assign n8283 = ( n7982 & ~n8282 ) | ( n7982 & n8281 ) | ( ~n8282 & n8281 ) ;
  assign n8285 = ( n7845 & ~n8284 ) | ( n7845 & n8283 ) | ( ~n8284 & n8283 ) ;
  assign n8260 = ( n7818 & ~n7982 ) | ( n7818 & n7823 ) | ( ~n7982 & n7823 ) ;
  assign n8259 = n7831 &  n7982 ;
  assign n8261 = ( n7982 & n8260 ) | ( n7982 & n8259 ) | ( n8260 & n8259 ) ;
  assign n8262 = ( n8259 & ~n8260 ) | ( n8259 & n7818 ) | ( ~n8260 & n7818 ) ;
  assign n8263 = ( n7823 & ~n8261 ) | ( n7823 & n8262 ) | ( ~n8261 & n8262 ) ;
  assign n8128 = ( n7686 & ~n7691 ) | ( n7686 & n7982 ) | ( ~n7691 & n7982 ) ;
  assign n8127 = ~n7699 & n7982 ;
  assign n8129 = ( n7982 & ~n8128 ) | ( n7982 & n8127 ) | ( ~n8128 & n8127 ) ;
  assign n8130 = ( n8127 & ~n7686 ) | ( n8127 & n8128 ) | ( ~n7686 & n8128 ) ;
  assign n8131 = ( n7691 & ~n8129 ) | ( n7691 & n8130 ) | ( ~n8129 & n8130 ) ;
  assign n8106 = ( n7665 & ~n7677 ) | ( n7665 & n7673 ) | ( ~n7677 & n7673 ) ;
  assign n8107 = ( n7665 & ~n8106 ) | ( n7665 & n7982 ) | ( ~n8106 & n7982 ) ;
  assign n8108 = ( n7982 & ~n7673 ) | ( n7982 & n8106 ) | ( ~n7673 & n8106 ) ;
  assign n8109 = ( n7677 & ~n8107 ) | ( n7677 & n8108 ) | ( ~n8107 & n8108 ) ;
  assign n8083 = ~n8068 & n8082 ;
  assign n8089 = ( n4668 & ~n8083 ) | ( n4668 & n8088 ) | ( ~n8083 & n8088 ) ;
  assign n8090 = n4353 &  n8089 ;
  assign n8091 = n7671 | n7982 ;
  assign n8092 = ( n7663 & n7667 ) | ( n7663 & n7671 ) | ( n7667 & n7671 ) ;
  assign n8093 = ( n8091 & ~n7667 ) | ( n8091 & n8092 ) | ( ~n7667 & n8092 ) ;
  assign n8094 = ( n7671 & ~n8092 ) | ( n7671 & n8091 ) | ( ~n8092 & n8091 ) ;
  assign n8095 = ( n7663 & ~n8093 ) | ( n7663 & n8094 ) | ( ~n8093 & n8094 ) ;
  assign n8098 = ( n8088 & ~n8097 ) | ( n8088 & 1'b0 ) | ( ~n8097 & 1'b0 ) ;
  assign n8102 = n4353 | n8101 ;
  assign n8103 = n8098 | n8102 ;
  assign n8104 = ~n8095 & n8103 ;
  assign n8105 = n8090 | n8104 ;
  assign n8110 = ( n4053 & ~n8109 ) | ( n4053 & n8105 ) | ( ~n8109 & n8105 ) ;
  assign n8111 = n3760 &  n8110 ;
  assign n8112 = n7697 | n7982 ;
  assign n8113 = ( n7684 & n7693 ) | ( n7684 & n7697 ) | ( n7693 & n7697 ) ;
  assign n8114 = ( n8112 & ~n7693 ) | ( n8112 & n8113 ) | ( ~n7693 & n8113 ) ;
  assign n8115 = ( n7697 & ~n8113 ) | ( n7697 & n8112 ) | ( ~n8113 & n8112 ) ;
  assign n8116 = ( n7684 & ~n8114 ) | ( n7684 & n8115 ) | ( ~n8114 & n8115 ) ;
  assign n8117 = n4053 | n8090 ;
  assign n8118 = n8104 | n8117 ;
  assign n8119 = ~n8109 & n8118 ;
  assign n8120 = n8098 | n8101 ;
  assign n8121 = ( n4353 & ~n8095 ) | ( n4353 & n8120 ) | ( ~n8095 & n8120 ) ;
  assign n8122 = n4053 &  n8121 ;
  assign n8123 = n3760 | n8122 ;
  assign n8124 = n8119 | n8123 ;
  assign n8125 = n8116 &  n8124 ;
  assign n8126 = n8111 | n8125 ;
  assign n8132 = ( n3482 & ~n8131 ) | ( n3482 & n8126 ) | ( ~n8131 & n8126 ) ;
  assign n8133 = n3211 &  n8132 ;
  assign n8134 = n7719 | n7982 ;
  assign n8135 = ( n7706 & n7715 ) | ( n7706 & n7719 ) | ( n7715 & n7719 ) ;
  assign n8136 = ( n8134 & ~n7715 ) | ( n8134 & n8135 ) | ( ~n7715 & n8135 ) ;
  assign n8137 = ( n7719 & ~n8135 ) | ( n7719 & n8134 ) | ( ~n8135 & n8134 ) ;
  assign n8138 = ( n7706 & ~n8136 ) | ( n7706 & n8137 ) | ( ~n8136 & n8137 ) ;
  assign n8139 = n3482 | n8111 ;
  assign n8140 = n8125 | n8139 ;
  assign n8141 = ~n8131 & n8140 ;
  assign n8142 = n8119 | n8122 ;
  assign n8143 = ( n3760 & n8116 ) | ( n3760 & n8142 ) | ( n8116 & n8142 ) ;
  assign n8144 = n3482 &  n8143 ;
  assign n8145 = n3211 | n8144 ;
  assign n8146 = n8141 | n8145 ;
  assign n8147 = n8138 &  n8146 ;
  assign n8148 = n8133 | n8147 ;
  assign n8149 = ~n7721 & n7982 ;
  assign n8150 = ( n7708 & n7713 ) | ( n7708 & n7982 ) | ( n7713 & n7982 ) ;
  assign n8152 = ( n8149 & ~n7708 ) | ( n8149 & n8150 ) | ( ~n7708 & n8150 ) ;
  assign n8151 = ( n7982 & ~n8150 ) | ( n7982 & n8149 ) | ( ~n8150 & n8149 ) ;
  assign n8153 = ( n7713 & ~n8152 ) | ( n7713 & n8151 ) | ( ~n8152 & n8151 ) ;
  assign n8154 = ( n2955 & n8148 ) | ( n2955 & n8153 ) | ( n8148 & n8153 ) ;
  assign n8155 = n2706 &  n8154 ;
  assign n8156 = n7741 | n7982 ;
  assign n8157 = ( n7728 & n7737 ) | ( n7728 & n7741 ) | ( n7737 & n7741 ) ;
  assign n8158 = ( n8156 & ~n7737 ) | ( n8156 & n8157 ) | ( ~n7737 & n8157 ) ;
  assign n8159 = ( n7741 & ~n8157 ) | ( n7741 & n8156 ) | ( ~n8157 & n8156 ) ;
  assign n8160 = ( n7728 & ~n8158 ) | ( n7728 & n8159 ) | ( ~n8158 & n8159 ) ;
  assign n8161 = n2955 | n8133 ;
  assign n8162 = n8147 | n8161 ;
  assign n8163 = n8153 &  n8162 ;
  assign n8164 = n8141 | n8144 ;
  assign n8165 = ( n3211 & n8138 ) | ( n3211 & n8164 ) | ( n8138 & n8164 ) ;
  assign n8166 = n2955 &  n8165 ;
  assign n8167 = n2706 | n8166 ;
  assign n8168 = n8163 | n8167 ;
  assign n8169 = n8160 &  n8168 ;
  assign n8170 = n8155 | n8169 ;
  assign n8171 = ~n7743 & n7982 ;
  assign n8172 = ( n7730 & n7735 ) | ( n7730 & n7982 ) | ( n7735 & n7982 ) ;
  assign n8174 = ( n8171 & ~n7730 ) | ( n8171 & n8172 ) | ( ~n7730 & n8172 ) ;
  assign n8173 = ( n7982 & ~n8172 ) | ( n7982 & n8171 ) | ( ~n8172 & n8171 ) ;
  assign n8175 = ( n7735 & ~n8174 ) | ( n7735 & n8173 ) | ( ~n8174 & n8173 ) ;
  assign n8176 = ( n2472 & n8170 ) | ( n2472 & n8175 ) | ( n8170 & n8175 ) ;
  assign n8177 = n2245 &  n8176 ;
  assign n8178 = n7763 | n7982 ;
  assign n8179 = ( n7750 & n7759 ) | ( n7750 & n7763 ) | ( n7759 & n7763 ) ;
  assign n8180 = ( n8178 & ~n7759 ) | ( n8178 & n8179 ) | ( ~n7759 & n8179 ) ;
  assign n8181 = ( n7763 & ~n8179 ) | ( n7763 & n8178 ) | ( ~n8179 & n8178 ) ;
  assign n8182 = ( n7750 & ~n8180 ) | ( n7750 & n8181 ) | ( ~n8180 & n8181 ) ;
  assign n8183 = n2472 | n8155 ;
  assign n8184 = n8169 | n8183 ;
  assign n8185 = n8175 &  n8184 ;
  assign n8186 = n8163 | n8166 ;
  assign n8187 = ( n2706 & n8160 ) | ( n2706 & n8186 ) | ( n8160 & n8186 ) ;
  assign n8188 = n2472 &  n8187 ;
  assign n8189 = n2245 | n8188 ;
  assign n8190 = n8185 | n8189 ;
  assign n8191 = n8182 &  n8190 ;
  assign n8192 = n8177 | n8191 ;
  assign n8193 = ~n7765 & n7982 ;
  assign n8194 = ( n7752 & n7757 ) | ( n7752 & n7982 ) | ( n7757 & n7982 ) ;
  assign n8196 = ( n8193 & ~n7752 ) | ( n8193 & n8194 ) | ( ~n7752 & n8194 ) ;
  assign n8195 = ( n7982 & ~n8194 ) | ( n7982 & n8193 ) | ( ~n8194 & n8193 ) ;
  assign n8197 = ( n7757 & ~n8196 ) | ( n7757 & n8195 ) | ( ~n8196 & n8195 ) ;
  assign n8198 = ( n8192 & ~n2033 ) | ( n8192 & n8197 ) | ( ~n2033 & n8197 ) ;
  assign n8199 = n1827 &  n8198 ;
  assign n8200 = n7785 | n7982 ;
  assign n8201 = ( n7772 & ~n7781 ) | ( n7772 & n7785 ) | ( ~n7781 & n7785 ) ;
  assign n8202 = ( n7781 & n8200 ) | ( n7781 & n8201 ) | ( n8200 & n8201 ) ;
  assign n8203 = ( n7785 & ~n8201 ) | ( n7785 & n8200 ) | ( ~n8201 & n8200 ) ;
  assign n8204 = ( n7772 & ~n8202 ) | ( n7772 & n8203 ) | ( ~n8202 & n8203 ) ;
  assign n8205 = ( n2033 & ~n8177 ) | ( n2033 & 1'b0 ) | ( ~n8177 & 1'b0 ) ;
  assign n8206 = ~n8191 & n8205 ;
  assign n8207 = ( n8197 & ~n8206 ) | ( n8197 & 1'b0 ) | ( ~n8206 & 1'b0 ) ;
  assign n8208 = n8185 | n8188 ;
  assign n8209 = ( n2245 & n8182 ) | ( n2245 & n8208 ) | ( n8182 & n8208 ) ;
  assign n8210 = ~n2033 & n8209 ;
  assign n8211 = n1827 | n8210 ;
  assign n8212 = n8207 | n8211 ;
  assign n8213 = n8204 &  n8212 ;
  assign n8214 = n8199 | n8213 ;
  assign n8215 = ~n7787 & n7982 ;
  assign n8216 = ( n7774 & n7779 ) | ( n7774 & n7982 ) | ( n7779 & n7982 ) ;
  assign n8218 = ( n8215 & ~n7774 ) | ( n8215 & n8216 ) | ( ~n7774 & n8216 ) ;
  assign n8217 = ( n7982 & ~n8216 ) | ( n7982 & n8215 ) | ( ~n8216 & n8215 ) ;
  assign n8219 = ( n7779 & ~n8218 ) | ( n7779 & n8217 ) | ( ~n8218 & n8217 ) ;
  assign n8220 = ( n1636 & ~n8214 ) | ( n1636 & n8219 ) | ( ~n8214 & n8219 ) ;
  assign n8221 = n1452 | n8220 ;
  assign n8222 = n7807 | n7982 ;
  assign n8223 = ( n7794 & ~n7807 ) | ( n7794 & n7803 ) | ( ~n7807 & n7803 ) ;
  assign n8225 = ( n7807 & n8222 ) | ( n7807 & n8223 ) | ( n8222 & n8223 ) ;
  assign n8224 = ( n7803 & ~n8223 ) | ( n7803 & n8222 ) | ( ~n8223 & n8222 ) ;
  assign n8226 = ( n7794 & ~n8225 ) | ( n7794 & n8224 ) | ( ~n8225 & n8224 ) ;
  assign n8227 = ( n1636 & ~n8199 ) | ( n1636 & 1'b0 ) | ( ~n8199 & 1'b0 ) ;
  assign n8228 = ~n8213 & n8227 ;
  assign n8229 = n8219 | n8228 ;
  assign n8230 = n8207 | n8210 ;
  assign n8231 = ( n1827 & n8204 ) | ( n1827 & n8230 ) | ( n8204 & n8230 ) ;
  assign n8232 = ~n1636 & n8231 ;
  assign n8233 = ( n1452 & ~n8232 ) | ( n1452 & 1'b0 ) | ( ~n8232 & 1'b0 ) ;
  assign n8234 = n8229 &  n8233 ;
  assign n8235 = n8226 | n8234 ;
  assign n8236 = n8221 &  n8235 ;
  assign n8237 = n7809 &  n7982 ;
  assign n8238 = ( n7801 & ~n7796 ) | ( n7801 & n7982 ) | ( ~n7796 & n7982 ) ;
  assign n8240 = ( n7796 & n8237 ) | ( n7796 & n8238 ) | ( n8237 & n8238 ) ;
  assign n8239 = ( n7982 & ~n8238 ) | ( n7982 & n8237 ) | ( ~n8238 & n8237 ) ;
  assign n8241 = ( n7801 & ~n8240 ) | ( n7801 & n8239 ) | ( ~n8240 & n8239 ) ;
  assign n8242 = ( n8236 & ~n1283 ) | ( n8236 & n8241 ) | ( ~n1283 & n8241 ) ;
  assign n8243 = n1122 | n8242 ;
  assign n8244 = n7829 | n7982 ;
  assign n8245 = ( n7816 & ~n7829 ) | ( n7816 & n7825 ) | ( ~n7829 & n7825 ) ;
  assign n8247 = ( n7829 & n8244 ) | ( n7829 & n8245 ) | ( n8244 & n8245 ) ;
  assign n8246 = ( n7825 & ~n8245 ) | ( n7825 & n8244 ) | ( ~n8245 & n8244 ) ;
  assign n8248 = ( n7816 & ~n8247 ) | ( n7816 & n8246 ) | ( ~n8247 & n8246 ) ;
  assign n8249 = ~n1283 & n8221 ;
  assign n8250 = n8235 &  n8249 ;
  assign n8251 = n8241 | n8250 ;
  assign n8252 = ( n8229 & ~n8232 ) | ( n8229 & 1'b0 ) | ( ~n8232 & 1'b0 ) ;
  assign n8253 = ( n1452 & n8226 ) | ( n1452 & n8252 ) | ( n8226 & n8252 ) ;
  assign n8254 = ( n1283 & ~n8253 ) | ( n1283 & 1'b0 ) | ( ~n8253 & 1'b0 ) ;
  assign n8255 = ( n1122 & ~n8254 ) | ( n1122 & 1'b0 ) | ( ~n8254 & 1'b0 ) ;
  assign n8256 = n8251 &  n8255 ;
  assign n8257 = n8248 | n8256 ;
  assign n8258 = n8243 &  n8257 ;
  assign n8264 = ( n976 & ~n8263 ) | ( n976 & n8258 ) | ( ~n8263 & n8258 ) ;
  assign n8265 = ( n837 & ~n8264 ) | ( n837 & 1'b0 ) | ( ~n8264 & 1'b0 ) ;
  assign n8267 = ( n7847 & ~n7838 ) | ( n7847 & n7851 ) | ( ~n7838 & n7851 ) ;
  assign n8266 = ( n7851 & ~n7982 ) | ( n7851 & 1'b0 ) | ( ~n7982 & 1'b0 ) ;
  assign n8269 = ( n7851 & ~n8267 ) | ( n7851 & n8266 ) | ( ~n8267 & n8266 ) ;
  assign n8268 = ( n8266 & ~n7847 ) | ( n8266 & n8267 ) | ( ~n7847 & n8267 ) ;
  assign n8270 = ( n7838 & ~n8269 ) | ( n7838 & n8268 ) | ( ~n8269 & n8268 ) ;
  assign n8271 = n976 &  n8243 ;
  assign n8272 = n8257 &  n8271 ;
  assign n8273 = ( n8263 & ~n8272 ) | ( n8263 & 1'b0 ) | ( ~n8272 & 1'b0 ) ;
  assign n8274 = ( n8251 & ~n8254 ) | ( n8251 & 1'b0 ) | ( ~n8254 & 1'b0 ) ;
  assign n8275 = ( n1122 & n8248 ) | ( n1122 & n8274 ) | ( n8248 & n8274 ) ;
  assign n8276 = n976 | n8275 ;
  assign n8277 = ~n837 & n8276 ;
  assign n8278 = ~n8273 & n8277 ;
  assign n8279 = ( n8270 & ~n8278 ) | ( n8270 & 1'b0 ) | ( ~n8278 & 1'b0 ) ;
  assign n8280 = n8265 | n8279 ;
  assign n8286 = ( n713 & ~n8285 ) | ( n713 & n8280 ) | ( ~n8285 & n8280 ) ;
  assign n8287 = n595 &  n8286 ;
  assign n8288 = n7873 | n7982 ;
  assign n8289 = ( n7860 & ~n7869 ) | ( n7860 & n7873 ) | ( ~n7869 & n7873 ) ;
  assign n8290 = ( n7869 & n8288 ) | ( n7869 & n8289 ) | ( n8288 & n8289 ) ;
  assign n8291 = ( n7873 & ~n8289 ) | ( n7873 & n8288 ) | ( ~n8289 & n8288 ) ;
  assign n8292 = ( n7860 & ~n8290 ) | ( n7860 & n8291 ) | ( ~n8290 & n8291 ) ;
  assign n8293 = n713 | n8265 ;
  assign n8294 = n8279 | n8293 ;
  assign n8295 = ~n8285 & n8294 ;
  assign n8296 = ~n8273 & n8276 ;
  assign n8297 = ( n837 & ~n8296 ) | ( n837 & n8270 ) | ( ~n8296 & n8270 ) ;
  assign n8298 = n713 &  n8297 ;
  assign n8299 = n595 | n8298 ;
  assign n8300 = n8295 | n8299 ;
  assign n8301 = n8292 &  n8300 ;
  assign n8302 = n8287 | n8301 ;
  assign n8303 = ~n7875 & n7982 ;
  assign n8304 = ( n7862 & n7867 ) | ( n7862 & n7982 ) | ( n7867 & n7982 ) ;
  assign n8306 = ( n8303 & ~n7862 ) | ( n8303 & n8304 ) | ( ~n7862 & n8304 ) ;
  assign n8305 = ( n7982 & ~n8304 ) | ( n7982 & n8303 ) | ( ~n8304 & n8303 ) ;
  assign n8307 = ( n7867 & ~n8306 ) | ( n7867 & n8305 ) | ( ~n8306 & n8305 ) ;
  assign n8308 = ( n492 & n8302 ) | ( n492 & n8307 ) | ( n8302 & n8307 ) ;
  assign n8309 = n396 &  n8308 ;
  assign n8311 = ( n7891 & ~n7882 ) | ( n7891 & n7895 ) | ( ~n7882 & n7895 ) ;
  assign n8310 = n7895 | n7982 ;
  assign n8313 = ( n7895 & ~n8311 ) | ( n7895 & n8310 ) | ( ~n8311 & n8310 ) ;
  assign n8312 = ( n8310 & ~n7891 ) | ( n8310 & n8311 ) | ( ~n7891 & n8311 ) ;
  assign n8314 = ( n7882 & ~n8313 ) | ( n7882 & n8312 ) | ( ~n8313 & n8312 ) ;
  assign n8315 = n492 | n8287 ;
  assign n8316 = n8301 | n8315 ;
  assign n8317 = n8307 &  n8316 ;
  assign n8318 = n8295 | n8298 ;
  assign n8319 = ( n595 & n8292 ) | ( n595 & n8318 ) | ( n8292 & n8318 ) ;
  assign n8320 = n492 &  n8319 ;
  assign n8321 = n396 | n8320 ;
  assign n8322 = n8317 | n8321 ;
  assign n8323 = ~n8314 & n8322 ;
  assign n8324 = n8309 | n8323 ;
  assign n8325 = ~n7897 & n7982 ;
  assign n8326 = ( n7884 & n7889 ) | ( n7884 & n7982 ) | ( n7889 & n7982 ) ;
  assign n8328 = ( n8325 & ~n7884 ) | ( n8325 & n8326 ) | ( ~n7884 & n8326 ) ;
  assign n8327 = ( n7982 & ~n8326 ) | ( n7982 & n8325 ) | ( ~n8326 & n8325 ) ;
  assign n8329 = ( n7889 & ~n8328 ) | ( n7889 & n8327 ) | ( ~n8328 & n8327 ) ;
  assign n8330 = ( n315 & n8324 ) | ( n315 & n8329 ) | ( n8324 & n8329 ) ;
  assign n8331 = n240 &  n8330 ;
  assign n8332 = n7917 | n7982 ;
  assign n8333 = ( n7904 & n7913 ) | ( n7904 & n7917 ) | ( n7913 & n7917 ) ;
  assign n8334 = ( n8332 & ~n7913 ) | ( n8332 & n8333 ) | ( ~n7913 & n8333 ) ;
  assign n8335 = ( n7917 & ~n8333 ) | ( n7917 & n8332 ) | ( ~n8333 & n8332 ) ;
  assign n8336 = ( n7904 & ~n8334 ) | ( n7904 & n8335 ) | ( ~n8334 & n8335 ) ;
  assign n8337 = n315 | n8309 ;
  assign n8338 = n8323 | n8337 ;
  assign n8339 = n8329 &  n8338 ;
  assign n8340 = n8317 | n8320 ;
  assign n8341 = ( n396 & ~n8314 ) | ( n396 & n8340 ) | ( ~n8314 & n8340 ) ;
  assign n8342 = n315 &  n8341 ;
  assign n8343 = n240 | n8342 ;
  assign n8344 = n8339 | n8343 ;
  assign n8345 = n8336 &  n8344 ;
  assign n8346 = n8331 | n8345 ;
  assign n8352 = ( n181 & ~n8351 ) | ( n181 & n8346 ) | ( ~n8351 & n8346 ) ;
  assign n8353 = ~n145 & n8352 ;
  assign n8355 = ( n7935 & ~n7926 ) | ( n7935 & n7939 ) | ( ~n7926 & n7939 ) ;
  assign n8354 = n7939 | n7982 ;
  assign n8357 = ( n7939 & ~n8355 ) | ( n7939 & n8354 ) | ( ~n8355 & n8354 ) ;
  assign n8356 = ( n8354 & ~n7935 ) | ( n8354 & n8355 ) | ( ~n7935 & n8355 ) ;
  assign n8358 = ( n7926 & ~n8357 ) | ( n7926 & n8356 ) | ( ~n8357 & n8356 ) ;
  assign n8359 = n181 | n8331 ;
  assign n8360 = n8345 | n8359 ;
  assign n8361 = ~n8351 & n8360 ;
  assign n8362 = n8339 | n8342 ;
  assign n8363 = ( n240 & n8336 ) | ( n240 & n8362 ) | ( n8336 & n8362 ) ;
  assign n8364 = n181 &  n8363 ;
  assign n8365 = ( n145 & ~n8364 ) | ( n145 & 1'b0 ) | ( ~n8364 & 1'b0 ) ;
  assign n8366 = ~n8361 & n8365 ;
  assign n8367 = ( n8358 & ~n8366 ) | ( n8358 & 1'b0 ) | ( ~n8366 & 1'b0 ) ;
  assign n8368 = n8353 | n8367 ;
  assign n8369 = n7928 | n7982 ;
  assign n8370 = ( n7933 & ~n7928 ) | ( n7933 & n7941 ) | ( ~n7928 & n7941 ) ;
  assign n8372 = ( n7928 & n8369 ) | ( n7928 & n8370 ) | ( n8369 & n8370 ) ;
  assign n8371 = ( n7941 & ~n8370 ) | ( n7941 & n8369 ) | ( ~n8370 & n8369 ) ;
  assign n8373 = ( n7933 & ~n8372 ) | ( n7933 & n8371 ) | ( ~n8372 & n8371 ) ;
  assign n8374 = ( n150 & n8368 ) | ( n150 & n8373 ) | ( n8368 & n8373 ) ;
  assign n8386 = n8374 | n8385 ;
  assign n8387 = ( n133 & ~n8385 ) | ( n133 & n8386 ) | ( ~n8385 & n8386 ) ;
  assign n8390 = n8361 | n8364 ;
  assign n8391 = ( n8358 & ~n145 ) | ( n8358 & n8390 ) | ( ~n145 & n8390 ) ;
  assign n8392 = n150 &  n8391 ;
  assign n8393 = ( n8381 & ~n8392 ) | ( n8381 & 1'b0 ) | ( ~n8392 & 1'b0 ) ;
  assign n8388 = n150 | n8353 ;
  assign n8389 = n8367 | n8388 ;
  assign n8394 = ( n8373 & ~n8389 ) | ( n8373 & 1'b0 ) | ( ~n8389 & 1'b0 ) ;
  assign n8395 = ( n8393 & ~n8373 ) | ( n8393 & n8394 ) | ( ~n8373 & n8394 ) ;
  assign n8397 = ( n133 & ~n7956 ) | ( n133 & n7949 ) | ( ~n7956 & n7949 ) ;
  assign n8396 = ( n7956 & ~n7949 ) | ( n7956 & n7982 ) | ( ~n7949 & n7982 ) ;
  assign n8398 = ~n7956 & n8396 ;
  assign n8399 = ( n7956 & n8397 ) | ( n7956 & n8398 ) | ( n8397 & n8398 ) ;
  assign n8400 = n7952 | n7979 ;
  assign n8401 = ( n7955 & n7974 ) | ( n7955 & n8400 ) | ( n7974 & n8400 ) ;
  assign n8402 = ( n7955 & ~n8401 ) | ( n7955 & 1'b0 ) | ( ~n8401 & 1'b0 ) ;
  assign n8403 = ( n7962 & ~n8402 ) | ( n7962 & n7970 ) | ( ~n8402 & n7970 ) ;
  assign n8404 = ( n7962 & ~n8403 ) | ( n7962 & 1'b0 ) | ( ~n8403 & 1'b0 ) ;
  assign n8405 = n8399 | n8404 ;
  assign n8406 = n8395 | n8405 ;
  assign n8407 = ~n8387 |  n8406 ;
  assign n8523 = n8101 | n8407 ;
  assign n8524 = ( n8088 & ~n8097 ) | ( n8088 & n8101 ) | ( ~n8097 & n8101 ) ;
  assign n8525 = ( n8097 & n8523 ) | ( n8097 & n8524 ) | ( n8523 & n8524 ) ;
  assign n8526 = ( n8101 & ~n8524 ) | ( n8101 & n8523 ) | ( ~n8524 & n8523 ) ;
  assign n8527 = ( n8088 & ~n8525 ) | ( n8088 & n8526 ) | ( ~n8525 & n8526 ) ;
  assign n8517 = ( n8068 & ~n8073 ) | ( n8068 & n8407 ) | ( ~n8073 & n8407 ) ;
  assign n8516 = n8081 &  n8407 ;
  assign n8518 = ( n8407 & ~n8517 ) | ( n8407 & n8516 ) | ( ~n8517 & n8516 ) ;
  assign n8519 = ( n8516 & ~n8068 ) | ( n8516 & n8517 ) | ( ~n8068 & n8517 ) ;
  assign n8520 = ( n8073 & ~n8518 ) | ( n8073 & n8519 ) | ( ~n8518 & n8519 ) ;
  assign n8501 = n8079 | n8407 ;
  assign n8502 = ( n8066 & ~n8075 ) | ( n8066 & n8079 ) | ( ~n8075 & n8079 ) ;
  assign n8503 = ( n8075 & n8501 ) | ( n8075 & n8502 ) | ( n8501 & n8502 ) ;
  assign n8504 = ( n8079 & ~n8502 ) | ( n8079 & n8501 ) | ( ~n8502 & n8501 ) ;
  assign n8505 = ( n8066 & ~n8503 ) | ( n8066 & n8504 ) | ( ~n8503 & n8504 ) ;
  assign n8494 = n8059 &  n8407 ;
  assign n8495 = ( n8046 & ~n8494 ) | ( n8046 & n8407 ) | ( ~n8494 & n8407 ) ;
  assign n8496 = ( n8051 & ~n8046 ) | ( n8051 & n8495 ) | ( ~n8046 & n8495 ) ;
  assign n8497 = ( n8046 & ~n8495 ) | ( n8046 & n8051 ) | ( ~n8495 & n8051 ) ;
  assign n8498 = ( n8496 & ~n8051 ) | ( n8496 & n8497 ) | ( ~n8051 & n8497 ) ;
  assign n8480 = ( n8053 & ~n8044 ) | ( n8053 & n8057 ) | ( ~n8044 & n8057 ) ;
  assign n8479 = ( n8053 & ~n8407 ) | ( n8053 & 1'b0 ) | ( ~n8407 & 1'b0 ) ;
  assign n8481 = ( n8053 & ~n8480 ) | ( n8053 & n8479 ) | ( ~n8480 & n8479 ) ;
  assign n8482 = ( n8479 & ~n8057 ) | ( n8479 & n8480 ) | ( ~n8057 & n8480 ) ;
  assign n8483 = ( n8044 & ~n8481 ) | ( n8044 & n8482 ) | ( ~n8481 & n8482 ) ;
  assign n8472 = n8024 | n8407 ;
  assign n8473 = ( n8024 & ~n8037 ) | ( n8024 & n8029 ) | ( ~n8037 & n8029 ) ;
  assign n8474 = ( n8037 & n8472 ) | ( n8037 & n8473 ) | ( n8472 & n8473 ) ;
  assign n8475 = ( n8024 & ~n8473 ) | ( n8024 & n8472 ) | ( ~n8473 & n8472 ) ;
  assign n8476 = ( n8029 & ~n8474 ) | ( n8029 & n8475 ) | ( ~n8474 & n8475 ) ;
  assign n8457 = n8031 | n8407 ;
  assign n8458 = ( n8022 & ~n8031 ) | ( n8022 & n8035 ) | ( ~n8031 & n8035 ) ;
  assign n8459 = ( n8031 & n8457 ) | ( n8031 & n8458 ) | ( n8457 & n8458 ) ;
  assign n8460 = ( n8035 & ~n8458 ) | ( n8035 & n8457 ) | ( ~n8458 & n8457 ) ;
  assign n8461 = ( n8022 & ~n8459 ) | ( n8022 & n8460 ) | ( ~n8459 & n8460 ) ;
  assign n8450 = n7998 | n8000 ;
  assign n8451 = ( n8000 & n8010 ) | ( n8000 & n8450 ) | ( n8010 & n8450 ) ;
  assign n8453 = ( n8407 & ~n8450 ) | ( n8407 & n8451 ) | ( ~n8450 & n8451 ) ;
  assign n8452 = ( n8000 & ~n8451 ) | ( n8000 & n8407 ) | ( ~n8451 & n8407 ) ;
  assign n8454 = ( n8010 & ~n8453 ) | ( n8010 & n8452 ) | ( ~n8453 & n8452 ) ;
  assign n8434 = ~x54 & n7982 ;
  assign n8435 = ( x55 & ~n8434 ) | ( x55 & 1'b0 ) | ( ~n8434 & 1'b0 ) ;
  assign n8436 = n8001 | n8435 ;
  assign n8431 = ( n7982 & ~x54 ) | ( n7982 & n7993 ) | ( ~x54 & n7993 ) ;
  assign n8432 = x54 &  n8431 ;
  assign n8433 = ( n7988 & ~n7993 ) | ( n7988 & n8432 ) | ( ~n7993 & n8432 ) ;
  assign n8437 = ( n8433 & ~n8407 ) | ( n8433 & n8436 ) | ( ~n8407 & n8436 ) ;
  assign n8439 = n8407 &  n8437 ;
  assign n8438 = ( n8433 & ~n8437 ) | ( n8433 & 1'b0 ) | ( ~n8437 & 1'b0 ) ;
  assign n8440 = ( n8436 & ~n8439 ) | ( n8436 & n8438 ) | ( ~n8439 & n8438 ) ;
  assign n8420 = ( n7982 & ~n8404 ) | ( n7982 & 1'b0 ) | ( ~n8404 & 1'b0 ) ;
  assign n8421 = ( n8395 & ~n8399 ) | ( n8395 & n8420 ) | ( ~n8399 & n8420 ) ;
  assign n8422 = ~n8395 & n8421 ;
  assign n8423 = n8387 &  n8422 ;
  assign n8419 = ~n7985 & n8407 ;
  assign n8424 = ( n8419 & ~n8423 ) | ( n8419 & 1'b0 ) | ( ~n8423 & 1'b0 ) ;
  assign n8425 = ( x54 & n8423 ) | ( x54 & n8424 ) | ( n8423 & n8424 ) ;
  assign n8426 = x54 | n8423 ;
  assign n8427 = n8419 | n8426 ;
  assign n8428 = ~n8425 & n8427 ;
  assign n8410 = ( x52 & ~n8407 ) | ( x52 & x53 ) | ( ~n8407 & x53 ) ;
  assign n8416 = ( x52 & ~x53 ) | ( x52 & 1'b0 ) | ( ~x53 & 1'b0 ) ;
  assign n7983 = x50 | x51 ;
  assign n8411 = ~x52 & n7983 ;
  assign n8412 = ( x52 & ~n7980 ) | ( x52 & n8411 ) | ( ~n7980 & n8411 ) ;
  assign n8413 = ( n7962 & ~n8412 ) | ( n7962 & n7970 ) | ( ~n8412 & n7970 ) ;
  assign n8414 = ( n7962 & ~n8413 ) | ( n7962 & 1'b0 ) | ( ~n8413 & 1'b0 ) ;
  assign n8415 = ( n8407 & ~x53 ) | ( n8407 & n8414 ) | ( ~x53 & n8414 ) ;
  assign n8417 = ( n8410 & ~n8416 ) | ( n8410 & n8415 ) | ( ~n8416 & n8415 ) ;
  assign n7984 = x52 | n7983 ;
  assign n8408 = x52 &  n8407 ;
  assign n8409 = ( n7982 & ~n7984 ) | ( n7982 & n8408 ) | ( ~n7984 & n8408 ) ;
  assign n8441 = ( n7572 & ~n8409 ) | ( n7572 & 1'b0 ) | ( ~n8409 & 1'b0 ) ;
  assign n8442 = n8417 &  n8441 ;
  assign n8443 = n8428 | n8442 ;
  assign n8444 = n8409 &  n8417 ;
  assign n8445 = ( n7572 & ~n8444 ) | ( n7572 & n8417 ) | ( ~n8444 & n8417 ) ;
  assign n8446 = n7169 &  n8445 ;
  assign n8447 = n8443 &  n8446 ;
  assign n8448 = n8440 | n8447 ;
  assign n8418 = ~n8409 & n8417 ;
  assign n8429 = ( n7572 & n8418 ) | ( n7572 & n8428 ) | ( n8418 & n8428 ) ;
  assign n8430 = n7169 | n8429 ;
  assign n8462 = ~n6781 & n8430 ;
  assign n8463 = n8448 &  n8462 ;
  assign n8464 = n8454 | n8463 ;
  assign n8465 = n8443 &  n8445 ;
  assign n8466 = ( n7169 & n8440 ) | ( n7169 & n8465 ) | ( n8440 & n8465 ) ;
  assign n8467 = ( n6781 & ~n8466 ) | ( n6781 & 1'b0 ) | ( ~n8466 & 1'b0 ) ;
  assign n8468 = ( n6399 & ~n8467 ) | ( n6399 & 1'b0 ) | ( ~n8467 & 1'b0 ) ;
  assign n8469 = n8464 &  n8468 ;
  assign n8470 = ( n8461 & ~n8469 ) | ( n8461 & 1'b0 ) | ( ~n8469 & 1'b0 ) ;
  assign n8449 = n8430 &  n8448 ;
  assign n8455 = ( n8449 & ~n6781 ) | ( n8449 & n8454 ) | ( ~n6781 & n8454 ) ;
  assign n8456 = n6399 | n8455 ;
  assign n8484 = ~n6032 & n8456 ;
  assign n8485 = ~n8470 & n8484 ;
  assign n8486 = ( n8476 & ~n8485 ) | ( n8476 & 1'b0 ) | ( ~n8485 & 1'b0 ) ;
  assign n8487 = ( n8464 & ~n8467 ) | ( n8464 & 1'b0 ) | ( ~n8467 & 1'b0 ) ;
  assign n8488 = ( n6399 & ~n8461 ) | ( n6399 & n8487 ) | ( ~n8461 & n8487 ) ;
  assign n8489 = ( n6032 & ~n8488 ) | ( n6032 & 1'b0 ) | ( ~n8488 & 1'b0 ) ;
  assign n8490 = ( n5672 & ~n8489 ) | ( n5672 & 1'b0 ) | ( ~n8489 & 1'b0 ) ;
  assign n8491 = ~n8486 & n8490 ;
  assign n8492 = n8483 | n8491 ;
  assign n8471 = ( n8456 & ~n8470 ) | ( n8456 & 1'b0 ) | ( ~n8470 & 1'b0 ) ;
  assign n8477 = ( n6032 & ~n8471 ) | ( n6032 & n8476 ) | ( ~n8471 & n8476 ) ;
  assign n8478 = ~n5672 & n8477 ;
  assign n8506 = n5327 | n8478 ;
  assign n8507 = ( n8492 & ~n8506 ) | ( n8492 & 1'b0 ) | ( ~n8506 & 1'b0 ) ;
  assign n8508 = n8498 | n8507 ;
  assign n8509 = n8486 | n8489 ;
  assign n8510 = ( n5672 & ~n8509 ) | ( n5672 & n8483 ) | ( ~n8509 & n8483 ) ;
  assign n8511 = ( n5327 & ~n8510 ) | ( n5327 & 1'b0 ) | ( ~n8510 & 1'b0 ) ;
  assign n8512 = n4990 | n8511 ;
  assign n8513 = ( n8508 & ~n8512 ) | ( n8508 & 1'b0 ) | ( ~n8512 & 1'b0 ) ;
  assign n8514 = n8505 | n8513 ;
  assign n8493 = ~n8478 & n8492 ;
  assign n8499 = ( n8493 & ~n5327 ) | ( n8493 & n8498 ) | ( ~n5327 & n8498 ) ;
  assign n8500 = ( n4990 & ~n8499 ) | ( n4990 & 1'b0 ) | ( ~n8499 & 1'b0 ) ;
  assign n8528 = n4668 | n8500 ;
  assign n8529 = ( n8514 & ~n8528 ) | ( n8514 & 1'b0 ) | ( ~n8528 & 1'b0 ) ;
  assign n8530 = n8520 | n8529 ;
  assign n8531 = ( n8508 & ~n8511 ) | ( n8508 & 1'b0 ) | ( ~n8511 & 1'b0 ) ;
  assign n8532 = ( n8505 & ~n4990 ) | ( n8505 & n8531 ) | ( ~n4990 & n8531 ) ;
  assign n8533 = ( n4668 & ~n8532 ) | ( n4668 & 1'b0 ) | ( ~n8532 & 1'b0 ) ;
  assign n8534 = n4353 | n8533 ;
  assign n8535 = ( n8530 & ~n8534 ) | ( n8530 & 1'b0 ) | ( ~n8534 & 1'b0 ) ;
  assign n8758 = ( n8309 & ~n8314 ) | ( n8309 & n8407 ) | ( ~n8314 & n8407 ) ;
  assign n8757 = ~n8322 & n8407 ;
  assign n8759 = ( n8407 & ~n8758 ) | ( n8407 & n8757 ) | ( ~n8758 & n8757 ) ;
  assign n8760 = ( n8757 & ~n8309 ) | ( n8757 & n8758 ) | ( ~n8309 & n8758 ) ;
  assign n8761 = ( n8314 & ~n8759 ) | ( n8314 & n8760 ) | ( ~n8759 & n8760 ) ;
  assign n8538 = ~n8103 & n8407 ;
  assign n8539 = ( n8090 & n8095 ) | ( n8090 & n8407 ) | ( n8095 & n8407 ) ;
  assign n8541 = ( n8538 & ~n8090 ) | ( n8538 & n8539 ) | ( ~n8090 & n8539 ) ;
  assign n8540 = ( n8407 & ~n8539 ) | ( n8407 & n8538 ) | ( ~n8539 & n8538 ) ;
  assign n8542 = ( n8095 & ~n8541 ) | ( n8095 & n8540 ) | ( ~n8541 & n8540 ) ;
  assign n8515 = ~n8500 & n8514 ;
  assign n8521 = ( n8515 & ~n4668 ) | ( n8515 & n8520 ) | ( ~n4668 & n8520 ) ;
  assign n8522 = ( n4353 & ~n8521 ) | ( n4353 & 1'b0 ) | ( ~n8521 & 1'b0 ) ;
  assign n8536 = ( n8527 & ~n8535 ) | ( n8527 & 1'b0 ) | ( ~n8535 & 1'b0 ) ;
  assign n8537 = n8522 | n8536 ;
  assign n8543 = ( n4053 & ~n8542 ) | ( n4053 & n8537 ) | ( ~n8542 & n8537 ) ;
  assign n8544 = n3760 &  n8543 ;
  assign n8545 = n4053 | n8522 ;
  assign n8546 = n8536 | n8545 ;
  assign n8547 = ~n8542 & n8546 ;
  assign n8548 = ( n8530 & ~n8533 ) | ( n8530 & 1'b0 ) | ( ~n8533 & 1'b0 ) ;
  assign n8549 = ( n4353 & ~n8548 ) | ( n4353 & n8527 ) | ( ~n8548 & n8527 ) ;
  assign n8550 = n4053 &  n8549 ;
  assign n8551 = n3760 | n8550 ;
  assign n8552 = n8547 | n8551 ;
  assign n8553 = ( n8118 & ~n8109 ) | ( n8118 & n8122 ) | ( ~n8109 & n8122 ) ;
  assign n8555 = ( n8122 & ~n8553 ) | ( n8122 & n8407 ) | ( ~n8553 & n8407 ) ;
  assign n8554 = ( n8407 & ~n8118 ) | ( n8407 & n8553 ) | ( ~n8118 & n8553 ) ;
  assign n8556 = ( n8109 & ~n8555 ) | ( n8109 & n8554 ) | ( ~n8555 & n8554 ) ;
  assign n8557 = ( n8552 & ~n8556 ) | ( n8552 & 1'b0 ) | ( ~n8556 & 1'b0 ) ;
  assign n8558 = n8544 | n8557 ;
  assign n8559 = ~n8124 & n8407 ;
  assign n8560 = ( n8111 & n8116 ) | ( n8111 & n8407 ) | ( n8116 & n8407 ) ;
  assign n8562 = ( n8559 & ~n8111 ) | ( n8559 & n8560 ) | ( ~n8111 & n8560 ) ;
  assign n8561 = ( n8407 & ~n8560 ) | ( n8407 & n8559 ) | ( ~n8560 & n8559 ) ;
  assign n8563 = ( n8116 & ~n8562 ) | ( n8116 & n8561 ) | ( ~n8562 & n8561 ) ;
  assign n8564 = ( n3482 & n8558 ) | ( n3482 & n8563 ) | ( n8558 & n8563 ) ;
  assign n8565 = n3211 &  n8564 ;
  assign n8566 = ( n8140 & ~n8407 ) | ( n8140 & 1'b0 ) | ( ~n8407 & 1'b0 ) ;
  assign n8567 = ( n8140 & n8131 ) | ( n8140 & n8144 ) | ( n8131 & n8144 ) ;
  assign n8569 = ( n8566 & ~n8144 ) | ( n8566 & n8567 ) | ( ~n8144 & n8567 ) ;
  assign n8568 = ( n8140 & ~n8567 ) | ( n8140 & n8566 ) | ( ~n8567 & n8566 ) ;
  assign n8570 = ( n8131 & ~n8569 ) | ( n8131 & n8568 ) | ( ~n8569 & n8568 ) ;
  assign n8571 = n3482 | n8544 ;
  assign n8572 = n8557 | n8571 ;
  assign n8573 = n8563 &  n8572 ;
  assign n8574 = n8547 | n8550 ;
  assign n8575 = ( n3760 & ~n8556 ) | ( n3760 & n8574 ) | ( ~n8556 & n8574 ) ;
  assign n8576 = n3482 &  n8575 ;
  assign n8577 = n3211 | n8576 ;
  assign n8578 = n8573 | n8577 ;
  assign n8579 = ~n8570 & n8578 ;
  assign n8580 = n8565 | n8579 ;
  assign n8581 = ~n8146 & n8407 ;
  assign n8582 = ( n8133 & n8138 ) | ( n8133 & n8407 ) | ( n8138 & n8407 ) ;
  assign n8584 = ( n8581 & ~n8133 ) | ( n8581 & n8582 ) | ( ~n8133 & n8582 ) ;
  assign n8583 = ( n8407 & ~n8582 ) | ( n8407 & n8581 ) | ( ~n8582 & n8581 ) ;
  assign n8585 = ( n8138 & ~n8584 ) | ( n8138 & n8583 ) | ( ~n8584 & n8583 ) ;
  assign n8586 = ( n2955 & n8580 ) | ( n2955 & n8585 ) | ( n8580 & n8585 ) ;
  assign n8587 = n2706 &  n8586 ;
  assign n8588 = ( n8162 & ~n8407 ) | ( n8162 & 1'b0 ) | ( ~n8407 & 1'b0 ) ;
  assign n8589 = ( n8162 & ~n8588 ) | ( n8162 & n8166 ) | ( ~n8588 & n8166 ) ;
  assign n8590 = ( n8153 & ~n8589 ) | ( n8153 & n8166 ) | ( ~n8589 & n8166 ) ;
  assign n8591 = ( n8153 & ~n8166 ) | ( n8153 & n8589 ) | ( ~n8166 & n8589 ) ;
  assign n8592 = ( n8590 & ~n8153 ) | ( n8590 & n8591 ) | ( ~n8153 & n8591 ) ;
  assign n8593 = n2955 | n8565 ;
  assign n8594 = n8579 | n8593 ;
  assign n8595 = n8585 &  n8594 ;
  assign n8596 = n8573 | n8576 ;
  assign n8597 = ( n3211 & ~n8570 ) | ( n3211 & n8596 ) | ( ~n8570 & n8596 ) ;
  assign n8598 = n2955 &  n8597 ;
  assign n8599 = n2706 | n8598 ;
  assign n8600 = n8595 | n8599 ;
  assign n8601 = n8592 &  n8600 ;
  assign n8602 = n8587 | n8601 ;
  assign n8603 = ~n8168 & n8407 ;
  assign n8604 = ( n8155 & n8160 ) | ( n8155 & n8407 ) | ( n8160 & n8407 ) ;
  assign n8606 = ( n8603 & ~n8155 ) | ( n8603 & n8604 ) | ( ~n8155 & n8604 ) ;
  assign n8605 = ( n8407 & ~n8604 ) | ( n8407 & n8603 ) | ( ~n8604 & n8603 ) ;
  assign n8607 = ( n8160 & ~n8606 ) | ( n8160 & n8605 ) | ( ~n8606 & n8605 ) ;
  assign n8608 = ( n2472 & n8602 ) | ( n2472 & n8607 ) | ( n8602 & n8607 ) ;
  assign n8609 = n2245 &  n8608 ;
  assign n8611 = ( n8184 & ~n8175 ) | ( n8184 & n8188 ) | ( ~n8175 & n8188 ) ;
  assign n8610 = ( n8184 & ~n8407 ) | ( n8184 & 1'b0 ) | ( ~n8407 & 1'b0 ) ;
  assign n8612 = ( n8184 & ~n8611 ) | ( n8184 & n8610 ) | ( ~n8611 & n8610 ) ;
  assign n8613 = ( n8610 & ~n8188 ) | ( n8610 & n8611 ) | ( ~n8188 & n8611 ) ;
  assign n8614 = ( n8175 & ~n8612 ) | ( n8175 & n8613 ) | ( ~n8612 & n8613 ) ;
  assign n8615 = n2472 | n8587 ;
  assign n8616 = n8601 | n8615 ;
  assign n8617 = n8607 &  n8616 ;
  assign n8618 = n8595 | n8598 ;
  assign n8619 = ( n2706 & n8592 ) | ( n2706 & n8618 ) | ( n8592 & n8618 ) ;
  assign n8620 = n2472 &  n8619 ;
  assign n8621 = n2245 | n8620 ;
  assign n8622 = n8617 | n8621 ;
  assign n8623 = n8614 &  n8622 ;
  assign n8624 = n8609 | n8623 ;
  assign n8625 = ~n8190 & n8407 ;
  assign n8626 = ( n8177 & n8182 ) | ( n8177 & n8407 ) | ( n8182 & n8407 ) ;
  assign n8628 = ( n8625 & ~n8177 ) | ( n8625 & n8626 ) | ( ~n8177 & n8626 ) ;
  assign n8627 = ( n8407 & ~n8626 ) | ( n8407 & n8625 ) | ( ~n8626 & n8625 ) ;
  assign n8629 = ( n8182 & ~n8628 ) | ( n8182 & n8627 ) | ( ~n8628 & n8627 ) ;
  assign n8630 = ( n8624 & ~n2033 ) | ( n8624 & n8629 ) | ( ~n2033 & n8629 ) ;
  assign n8631 = n1827 &  n8630 ;
  assign n8632 = n8206 | n8407 ;
  assign n8633 = ( n8210 & ~n8206 ) | ( n8210 & n8632 ) | ( ~n8206 & n8632 ) ;
  assign n8634 = ( n8197 & ~n8633 ) | ( n8197 & n8210 ) | ( ~n8633 & n8210 ) ;
  assign n8635 = ( n8197 & ~n8210 ) | ( n8197 & n8633 ) | ( ~n8210 & n8633 ) ;
  assign n8636 = ( n8634 & ~n8197 ) | ( n8634 & n8635 ) | ( ~n8197 & n8635 ) ;
  assign n8637 = ( n2033 & ~n8609 ) | ( n2033 & 1'b0 ) | ( ~n8609 & 1'b0 ) ;
  assign n8638 = ~n8623 & n8637 ;
  assign n8639 = ( n8629 & ~n8638 ) | ( n8629 & 1'b0 ) | ( ~n8638 & 1'b0 ) ;
  assign n8640 = n8617 | n8620 ;
  assign n8641 = ( n2245 & n8614 ) | ( n2245 & n8640 ) | ( n8614 & n8640 ) ;
  assign n8642 = ~n2033 & n8641 ;
  assign n8643 = n1827 | n8642 ;
  assign n8644 = n8639 | n8643 ;
  assign n8645 = n8636 &  n8644 ;
  assign n8646 = n8631 | n8645 ;
  assign n8648 = ( n8199 & ~n8204 ) | ( n8199 & n8407 ) | ( ~n8204 & n8407 ) ;
  assign n8647 = ~n8212 & n8407 ;
  assign n8649 = ( n8407 & ~n8648 ) | ( n8407 & n8647 ) | ( ~n8648 & n8647 ) ;
  assign n8650 = ( n8647 & ~n8199 ) | ( n8647 & n8648 ) | ( ~n8199 & n8648 ) ;
  assign n8651 = ( n8204 & ~n8649 ) | ( n8204 & n8650 ) | ( ~n8649 & n8650 ) ;
  assign n8652 = ( n8646 & ~n1636 ) | ( n8646 & n8651 ) | ( ~n1636 & n8651 ) ;
  assign n8653 = ~n1452 & n8652 ;
  assign n8654 = n8232 | n8407 ;
  assign n8655 = ( n8219 & ~n8232 ) | ( n8219 & n8228 ) | ( ~n8232 & n8228 ) ;
  assign n8657 = ( n8232 & n8654 ) | ( n8232 & n8655 ) | ( n8654 & n8655 ) ;
  assign n8656 = ( n8228 & ~n8655 ) | ( n8228 & n8654 ) | ( ~n8655 & n8654 ) ;
  assign n8658 = ( n8219 & ~n8657 ) | ( n8219 & n8656 ) | ( ~n8657 & n8656 ) ;
  assign n8659 = ( n1636 & ~n8631 ) | ( n1636 & 1'b0 ) | ( ~n8631 & 1'b0 ) ;
  assign n8660 = ~n8645 & n8659 ;
  assign n8661 = ( n8651 & ~n8660 ) | ( n8651 & 1'b0 ) | ( ~n8660 & 1'b0 ) ;
  assign n8662 = n8639 | n8642 ;
  assign n8663 = ( n1827 & n8636 ) | ( n1827 & n8662 ) | ( n8636 & n8662 ) ;
  assign n8664 = ~n1636 & n8663 ;
  assign n8665 = ( n1452 & ~n8664 ) | ( n1452 & 1'b0 ) | ( ~n8664 & 1'b0 ) ;
  assign n8666 = ~n8661 & n8665 ;
  assign n8667 = n8658 | n8666 ;
  assign n8668 = ~n8653 & n8667 ;
  assign n8669 = n8234 &  n8407 ;
  assign n8670 = ( n8226 & ~n8221 ) | ( n8226 & n8407 ) | ( ~n8221 & n8407 ) ;
  assign n8672 = ( n8221 & n8669 ) | ( n8221 & n8670 ) | ( n8669 & n8670 ) ;
  assign n8671 = ( n8407 & ~n8670 ) | ( n8407 & n8669 ) | ( ~n8670 & n8669 ) ;
  assign n8673 = ( n8226 & ~n8672 ) | ( n8226 & n8671 ) | ( ~n8672 & n8671 ) ;
  assign n8674 = ( n8668 & ~n1283 ) | ( n8668 & n8673 ) | ( ~n1283 & n8673 ) ;
  assign n8675 = n1122 | n8674 ;
  assign n8676 = n8250 | n8407 ;
  assign n8677 = ( n8250 & ~n8254 ) | ( n8250 & n8241 ) | ( ~n8254 & n8241 ) ;
  assign n8679 = ( n8676 & n8254 ) | ( n8676 & n8677 ) | ( n8254 & n8677 ) ;
  assign n8678 = ( n8250 & ~n8677 ) | ( n8250 & n8676 ) | ( ~n8677 & n8676 ) ;
  assign n8680 = ( n8241 & ~n8679 ) | ( n8241 & n8678 ) | ( ~n8679 & n8678 ) ;
  assign n8681 = n1283 | n8653 ;
  assign n8682 = ( n8667 & ~n8681 ) | ( n8667 & 1'b0 ) | ( ~n8681 & 1'b0 ) ;
  assign n8683 = n8673 | n8682 ;
  assign n8684 = n8661 | n8664 ;
  assign n8685 = ( n1452 & ~n8684 ) | ( n1452 & n8658 ) | ( ~n8684 & n8658 ) ;
  assign n8686 = ( n1283 & ~n8685 ) | ( n1283 & 1'b0 ) | ( ~n8685 & 1'b0 ) ;
  assign n8687 = ( n1122 & ~n8686 ) | ( n1122 & 1'b0 ) | ( ~n8686 & 1'b0 ) ;
  assign n8688 = n8683 &  n8687 ;
  assign n8689 = n8680 | n8688 ;
  assign n8690 = n8675 &  n8689 ;
  assign n8691 = n8256 &  n8407 ;
  assign n8692 = ( n8248 & ~n8243 ) | ( n8248 & n8407 ) | ( ~n8243 & n8407 ) ;
  assign n8694 = ( n8691 & n8243 ) | ( n8691 & n8692 ) | ( n8243 & n8692 ) ;
  assign n8693 = ( n8407 & ~n8692 ) | ( n8407 & n8691 ) | ( ~n8692 & n8691 ) ;
  assign n8695 = ( n8248 & ~n8694 ) | ( n8248 & n8693 ) | ( ~n8694 & n8693 ) ;
  assign n8696 = ( n976 & n8690 ) | ( n976 & n8695 ) | ( n8690 & n8695 ) ;
  assign n8697 = ( n837 & ~n8696 ) | ( n837 & 1'b0 ) | ( ~n8696 & 1'b0 ) ;
  assign n8699 = ( n8272 & ~n8263 ) | ( n8272 & n8276 ) | ( ~n8263 & n8276 ) ;
  assign n8698 = n8272 | n8407 ;
  assign n8700 = ( n8272 & ~n8699 ) | ( n8272 & n8698 ) | ( ~n8699 & n8698 ) ;
  assign n8701 = ( n8698 & ~n8276 ) | ( n8698 & n8699 ) | ( ~n8276 & n8699 ) ;
  assign n8702 = ( n8263 & ~n8700 ) | ( n8263 & n8701 ) | ( ~n8700 & n8701 ) ;
  assign n8703 = n976 &  n8675 ;
  assign n8704 = n8689 &  n8703 ;
  assign n8705 = n8695 | n8704 ;
  assign n8706 = ( n8683 & ~n8686 ) | ( n8683 & 1'b0 ) | ( ~n8686 & 1'b0 ) ;
  assign n8707 = ( n1122 & n8680 ) | ( n1122 & n8706 ) | ( n8680 & n8706 ) ;
  assign n8708 = n976 | n8707 ;
  assign n8709 = ~n837 & n8708 ;
  assign n8710 = n8705 &  n8709 ;
  assign n8711 = ( n8702 & ~n8710 ) | ( n8702 & 1'b0 ) | ( ~n8710 & 1'b0 ) ;
  assign n8712 = n8697 | n8711 ;
  assign n8714 = ( n8265 & ~n8270 ) | ( n8265 & n8407 ) | ( ~n8270 & n8407 ) ;
  assign n8713 = n8278 &  n8407 ;
  assign n8715 = ( n8407 & ~n8714 ) | ( n8407 & n8713 ) | ( ~n8714 & n8713 ) ;
  assign n8716 = ( n8713 & ~n8265 ) | ( n8713 & n8714 ) | ( ~n8265 & n8714 ) ;
  assign n8717 = ( n8270 & ~n8715 ) | ( n8270 & n8716 ) | ( ~n8715 & n8716 ) ;
  assign n8718 = ( n713 & n8712 ) | ( n713 & n8717 ) | ( n8712 & n8717 ) ;
  assign n8719 = n595 &  n8718 ;
  assign n8721 = ( n8294 & ~n8285 ) | ( n8294 & n8298 ) | ( ~n8285 & n8298 ) ;
  assign n8720 = n8298 | n8407 ;
  assign n8723 = ( n8298 & ~n8721 ) | ( n8298 & n8720 ) | ( ~n8721 & n8720 ) ;
  assign n8722 = ( n8720 & ~n8294 ) | ( n8720 & n8721 ) | ( ~n8294 & n8721 ) ;
  assign n8724 = ( n8285 & ~n8723 ) | ( n8285 & n8722 ) | ( ~n8723 & n8722 ) ;
  assign n8725 = n713 | n8697 ;
  assign n8726 = n8711 | n8725 ;
  assign n8727 = n8717 &  n8726 ;
  assign n8728 = n8705 &  n8708 ;
  assign n8729 = ( n837 & ~n8728 ) | ( n837 & n8702 ) | ( ~n8728 & n8702 ) ;
  assign n8730 = n713 &  n8729 ;
  assign n8731 = n595 | n8730 ;
  assign n8732 = n8727 | n8731 ;
  assign n8733 = ~n8724 & n8732 ;
  assign n8734 = n8719 | n8733 ;
  assign n8735 = ~n8300 & n8407 ;
  assign n8736 = ( n8287 & ~n8735 ) | ( n8287 & n8407 ) | ( ~n8735 & n8407 ) ;
  assign n8737 = ( n8287 & ~n8736 ) | ( n8287 & n8292 ) | ( ~n8736 & n8292 ) ;
  assign n8738 = ( n8292 & ~n8287 ) | ( n8292 & n8736 ) | ( ~n8287 & n8736 ) ;
  assign n8739 = ( n8737 & ~n8292 ) | ( n8737 & n8738 ) | ( ~n8292 & n8738 ) ;
  assign n8740 = ( n492 & n8734 ) | ( n492 & n8739 ) | ( n8734 & n8739 ) ;
  assign n8741 = n396 &  n8740 ;
  assign n8742 = ( n8316 & ~n8407 ) | ( n8316 & 1'b0 ) | ( ~n8407 & 1'b0 ) ;
  assign n8743 = ( n8316 & ~n8742 ) | ( n8316 & n8320 ) | ( ~n8742 & n8320 ) ;
  assign n8744 = ( n8307 & ~n8743 ) | ( n8307 & n8320 ) | ( ~n8743 & n8320 ) ;
  assign n8745 = ( n8307 & ~n8320 ) | ( n8307 & n8743 ) | ( ~n8320 & n8743 ) ;
  assign n8746 = ( n8744 & ~n8307 ) | ( n8744 & n8745 ) | ( ~n8307 & n8745 ) ;
  assign n8747 = n492 | n8719 ;
  assign n8748 = n8733 | n8747 ;
  assign n8749 = n8739 &  n8748 ;
  assign n8750 = n8727 | n8730 ;
  assign n8751 = ( n595 & ~n8724 ) | ( n595 & n8750 ) | ( ~n8724 & n8750 ) ;
  assign n8752 = n492 &  n8751 ;
  assign n8753 = n396 | n8752 ;
  assign n8754 = n8749 | n8753 ;
  assign n8755 = n8746 &  n8754 ;
  assign n8756 = n8741 | n8755 ;
  assign n8762 = ( n315 & ~n8761 ) | ( n315 & n8756 ) | ( ~n8761 & n8756 ) ;
  assign n8763 = n240 &  n8762 ;
  assign n8764 = ( n8338 & ~n8407 ) | ( n8338 & 1'b0 ) | ( ~n8407 & 1'b0 ) ;
  assign n8765 = ( n8338 & ~n8764 ) | ( n8338 & n8342 ) | ( ~n8764 & n8342 ) ;
  assign n8766 = ( n8329 & ~n8765 ) | ( n8329 & n8342 ) | ( ~n8765 & n8342 ) ;
  assign n8767 = ( n8329 & ~n8342 ) | ( n8329 & n8765 ) | ( ~n8342 & n8765 ) ;
  assign n8768 = ( n8766 & ~n8329 ) | ( n8766 & n8767 ) | ( ~n8329 & n8767 ) ;
  assign n8769 = n315 | n8741 ;
  assign n8770 = n8755 | n8769 ;
  assign n8771 = ~n8761 & n8770 ;
  assign n8772 = n8749 | n8752 ;
  assign n8773 = ( n396 & n8746 ) | ( n396 & n8772 ) | ( n8746 & n8772 ) ;
  assign n8774 = n315 &  n8773 ;
  assign n8775 = n240 | n8774 ;
  assign n8776 = n8771 | n8775 ;
  assign n8777 = n8768 &  n8776 ;
  assign n8778 = n8763 | n8777 ;
  assign n8779 = ~n8344 & n8407 ;
  assign n8780 = ( n8331 & n8336 ) | ( n8331 & n8407 ) | ( n8336 & n8407 ) ;
  assign n8782 = ( n8779 & ~n8331 ) | ( n8779 & n8780 ) | ( ~n8331 & n8780 ) ;
  assign n8781 = ( n8407 & ~n8780 ) | ( n8407 & n8779 ) | ( ~n8780 & n8779 ) ;
  assign n8783 = ( n8336 & ~n8782 ) | ( n8336 & n8781 ) | ( ~n8782 & n8781 ) ;
  assign n8784 = ( n181 & n8778 ) | ( n181 & n8783 ) | ( n8778 & n8783 ) ;
  assign n8785 = ~n145 & n8784 ;
  assign n8786 = ( n8360 & ~n8407 ) | ( n8360 & 1'b0 ) | ( ~n8407 & 1'b0 ) ;
  assign n8787 = ( n8360 & n8351 ) | ( n8360 & n8364 ) | ( n8351 & n8364 ) ;
  assign n8789 = ( n8786 & ~n8364 ) | ( n8786 & n8787 ) | ( ~n8364 & n8787 ) ;
  assign n8788 = ( n8360 & ~n8787 ) | ( n8360 & n8786 ) | ( ~n8787 & n8786 ) ;
  assign n8790 = ( n8351 & ~n8789 ) | ( n8351 & n8788 ) | ( ~n8789 & n8788 ) ;
  assign n8791 = n181 | n8763 ;
  assign n8792 = n8777 | n8791 ;
  assign n8793 = n8783 &  n8792 ;
  assign n8794 = n8771 | n8774 ;
  assign n8795 = ( n240 & n8768 ) | ( n240 & n8794 ) | ( n8768 & n8794 ) ;
  assign n8796 = n181 &  n8795 ;
  assign n8797 = ( n145 & ~n8796 ) | ( n145 & 1'b0 ) | ( ~n8796 & 1'b0 ) ;
  assign n8798 = ~n8793 & n8797 ;
  assign n8799 = n8790 | n8798 ;
  assign n8800 = ~n8785 & n8799 ;
  assign n8801 = n8366 &  n8407 ;
  assign n8802 = ( n8353 & n8358 ) | ( n8353 & n8407 ) | ( n8358 & n8407 ) ;
  assign n8804 = ( n8801 & ~n8353 ) | ( n8801 & n8802 ) | ( ~n8353 & n8802 ) ;
  assign n8803 = ( n8407 & ~n8802 ) | ( n8407 & n8801 ) | ( ~n8802 & n8801 ) ;
  assign n8805 = ( n8358 & ~n8804 ) | ( n8358 & n8803 ) | ( ~n8804 & n8803 ) ;
  assign n8806 = ( n150 & ~n8800 ) | ( n150 & n8805 ) | ( ~n8800 & n8805 ) ;
  assign n8807 = n8373 | n8392 ;
  assign n8808 = ( n8389 & ~n8407 ) | ( n8389 & n8807 ) | ( ~n8407 & n8807 ) ;
  assign n8809 = ( n8389 & ~n8808 ) | ( n8389 & 1'b0 ) | ( ~n8808 & 1'b0 ) ;
  assign n8810 = ( n8389 & ~n8392 ) | ( n8389 & 1'b0 ) | ( ~n8392 & 1'b0 ) ;
  assign n8811 = ~n8407 & n8810 ;
  assign n8812 = ( n8373 & ~n8810 ) | ( n8373 & n8811 ) | ( ~n8810 & n8811 ) ;
  assign n8813 = n8809 | n8812 ;
  assign n8814 = ( n8374 & ~n8381 ) | ( n8374 & 1'b0 ) | ( ~n8381 & 1'b0 ) ;
  assign n8815 = ~n8407 & n8814 ;
  assign n8816 = ( n8395 & ~n8815 ) | ( n8395 & n8814 ) | ( ~n8815 & n8814 ) ;
  assign n8817 = ( n8813 & ~n8816 ) | ( n8813 & 1'b0 ) | ( ~n8816 & 1'b0 ) ;
  assign n8818 = ~n8806 & n8817 ;
  assign n8819 = ( n133 & ~n8818 ) | ( n133 & n8817 ) | ( ~n8818 & n8817 ) ;
  assign n8820 = n150 | n8785 ;
  assign n8821 = ( n8799 & ~n8820 ) | ( n8799 & 1'b0 ) | ( ~n8820 & 1'b0 ) ;
  assign n8826 = n8805 &  n8821 ;
  assign n8822 = n8793 | n8796 ;
  assign n8823 = ( n145 & ~n8822 ) | ( n145 & n8790 ) | ( ~n8822 & n8790 ) ;
  assign n8824 = ( n150 & ~n8823 ) | ( n150 & 1'b0 ) | ( ~n8823 & 1'b0 ) ;
  assign n8825 = n8813 | n8824 ;
  assign n8827 = ( n8805 & ~n8826 ) | ( n8805 & n8825 ) | ( ~n8826 & n8825 ) ;
  assign n8829 = ( n133 & ~n8381 ) | ( n133 & n8374 ) | ( ~n8381 & n8374 ) ;
  assign n8828 = ( n8381 & ~n8374 ) | ( n8381 & n8407 ) | ( ~n8374 & n8407 ) ;
  assign n8830 = ~n8381 & n8828 ;
  assign n8831 = ( n8381 & n8829 ) | ( n8381 & n8830 ) | ( n8829 & n8830 ) ;
  assign n8832 = n8377 | n8404 ;
  assign n8833 = ( n8380 & n8399 ) | ( n8380 & n8832 ) | ( n8399 & n8832 ) ;
  assign n8834 = ( n8380 & ~n8833 ) | ( n8380 & 1'b0 ) | ( ~n8833 & 1'b0 ) ;
  assign n8835 = ( n8387 & ~n8834 ) | ( n8387 & n8395 ) | ( ~n8834 & n8395 ) ;
  assign n8836 = ( n8387 & ~n8835 ) | ( n8387 & 1'b0 ) | ( ~n8835 & 1'b0 ) ;
  assign n8837 = n8831 | n8836 ;
  assign n8838 = ( n8827 & ~n8837 ) | ( n8827 & 1'b0 ) | ( ~n8837 & 1'b0 ) ;
  assign n8839 = ~n8819 | ~n8838 ;
  assign n8985 = n8535 &  n8839 ;
  assign n8986 = ( n8522 & n8527 ) | ( n8522 & n8839 ) | ( n8527 & n8839 ) ;
  assign n8988 = ( n8985 & ~n8522 ) | ( n8985 & n8986 ) | ( ~n8522 & n8986 ) ;
  assign n8987 = ( n8839 & ~n8986 ) | ( n8839 & n8985 ) | ( ~n8986 & n8985 ) ;
  assign n8989 = ( n8527 & ~n8988 ) | ( n8527 & n8987 ) | ( ~n8988 & n8987 ) ;
  assign n8970 = n8533 | n8839 ;
  assign n8971 = ( n8520 & ~n8533 ) | ( n8520 & n8529 ) | ( ~n8533 & n8529 ) ;
  assign n8973 = ( n8533 & n8970 ) | ( n8533 & n8971 ) | ( n8970 & n8971 ) ;
  assign n8972 = ( n8529 & ~n8971 ) | ( n8529 & n8970 ) | ( ~n8971 & n8970 ) ;
  assign n8974 = ( n8520 & ~n8973 ) | ( n8520 & n8972 ) | ( ~n8973 & n8972 ) ;
  assign n8963 = n8513 &  n8839 ;
  assign n8964 = ( n8500 & n8505 ) | ( n8500 & n8839 ) | ( n8505 & n8839 ) ;
  assign n8966 = ( n8963 & ~n8500 ) | ( n8963 & n8964 ) | ( ~n8500 & n8964 ) ;
  assign n8965 = ( n8839 & ~n8964 ) | ( n8839 & n8963 ) | ( ~n8964 & n8963 ) ;
  assign n8967 = ( n8505 & ~n8966 ) | ( n8505 & n8965 ) | ( ~n8966 & n8965 ) ;
  assign n8948 = n8511 | n8839 ;
  assign n8949 = ( n8498 & ~n8511 ) | ( n8498 & n8507 ) | ( ~n8511 & n8507 ) ;
  assign n8951 = ( n8511 & n8948 ) | ( n8511 & n8949 ) | ( n8948 & n8949 ) ;
  assign n8950 = ( n8507 & ~n8949 ) | ( n8507 & n8948 ) | ( ~n8949 & n8948 ) ;
  assign n8952 = ( n8498 & ~n8951 ) | ( n8498 & n8950 ) | ( ~n8951 & n8950 ) ;
  assign n8941 = n8478 | n8839 ;
  assign n8942 = ( n8483 & ~n8478 ) | ( n8483 & n8491 ) | ( ~n8478 & n8491 ) ;
  assign n8944 = ( n8478 & n8941 ) | ( n8478 & n8942 ) | ( n8941 & n8942 ) ;
  assign n8943 = ( n8491 & ~n8942 ) | ( n8491 & n8941 ) | ( ~n8942 & n8941 ) ;
  assign n8945 = ( n8483 & ~n8944 ) | ( n8483 & n8943 ) | ( ~n8944 & n8943 ) ;
  assign n8926 = n8489 | n8839 ;
  assign n8927 = ( n8476 & ~n8489 ) | ( n8476 & n8485 ) | ( ~n8489 & n8485 ) ;
  assign n8929 = ( n8489 & n8926 ) | ( n8489 & n8927 ) | ( n8926 & n8927 ) ;
  assign n8928 = ( n8485 & ~n8927 ) | ( n8485 & n8926 ) | ( ~n8927 & n8926 ) ;
  assign n8930 = ( n8476 & ~n8929 ) | ( n8476 & n8928 ) | ( ~n8929 & n8928 ) ;
  assign n8920 = ( n8456 & ~n8461 ) | ( n8456 & n8469 ) | ( ~n8461 & n8469 ) ;
  assign n8919 = ( n8456 & ~n8839 ) | ( n8456 & 1'b0 ) | ( ~n8839 & 1'b0 ) ;
  assign n8922 = ( n8456 & ~n8920 ) | ( n8456 & n8919 ) | ( ~n8920 & n8919 ) ;
  assign n8921 = ( n8919 & ~n8469 ) | ( n8919 & n8920 ) | ( ~n8469 & n8920 ) ;
  assign n8923 = ( n8461 & ~n8922 ) | ( n8461 & n8921 ) | ( ~n8922 & n8921 ) ;
  assign n8904 = n8467 | n8839 ;
  assign n8905 = ( n8454 & ~n8463 ) | ( n8454 & n8467 ) | ( ~n8463 & n8467 ) ;
  assign n8906 = ( n8463 & n8904 ) | ( n8463 & n8905 ) | ( n8904 & n8905 ) ;
  assign n8907 = ( n8467 & ~n8905 ) | ( n8467 & n8904 ) | ( ~n8905 & n8904 ) ;
  assign n8908 = ( n8454 & ~n8906 ) | ( n8454 & n8907 ) | ( ~n8906 & n8907 ) ;
  assign n8897 = n8447 &  n8839 ;
  assign n8898 = ( n8440 & ~n8430 ) | ( n8440 & n8839 ) | ( ~n8430 & n8839 ) ;
  assign n8900 = ( n8430 & n8897 ) | ( n8430 & n8898 ) | ( n8897 & n8898 ) ;
  assign n8899 = ( n8839 & ~n8898 ) | ( n8839 & n8897 ) | ( ~n8898 & n8897 ) ;
  assign n8901 = ( n8440 & ~n8900 ) | ( n8440 & n8899 ) | ( ~n8900 & n8899 ) ;
  assign n8882 = n8442 | n8445 ;
  assign n8883 = ( n8442 & ~n8428 ) | ( n8442 & n8882 ) | ( ~n8428 & n8882 ) ;
  assign n8885 = ( n8442 & ~n8883 ) | ( n8442 & n8839 ) | ( ~n8883 & n8839 ) ;
  assign n8884 = ( n8839 & ~n8882 ) | ( n8839 & n8883 ) | ( ~n8882 & n8883 ) ;
  assign n8886 = ( n8428 & ~n8885 ) | ( n8428 & n8884 ) | ( ~n8885 & n8884 ) ;
  assign n8873 = ~x52 & n8407 ;
  assign n8874 = ( x53 & ~n8873 ) | ( x53 & 1'b0 ) | ( ~n8873 & 1'b0 ) ;
  assign n8875 = n8419 | n8874 ;
  assign n8870 = ( n8407 & ~x52 ) | ( n8407 & n8414 ) | ( ~x52 & n8414 ) ;
  assign n8871 = x52 &  n8870 ;
  assign n8872 = ( n8409 & ~n8871 ) | ( n8409 & n8414 ) | ( ~n8871 & n8414 ) ;
  assign n8876 = ( n8839 & ~n8875 ) | ( n8839 & n8872 ) | ( ~n8875 & n8872 ) ;
  assign n8878 = ( n8839 & ~n8876 ) | ( n8839 & 1'b0 ) | ( ~n8876 & 1'b0 ) ;
  assign n8877 = ~n8872 & n8876 ;
  assign n8879 = ( n8875 & ~n8878 ) | ( n8875 & n8877 ) | ( ~n8878 & n8877 ) ;
  assign n8846 = ( x50 & ~n8839 ) | ( x50 & x51 ) | ( ~n8839 & x51 ) ;
  assign n8852 = ( x50 & ~x51 ) | ( x50 & 1'b0 ) | ( ~x51 & 1'b0 ) ;
  assign n8842 = x48 | x49 ;
  assign n8847 = ~x50 & n8842 ;
  assign n8848 = ( x50 & ~n8405 ) | ( x50 & n8847 ) | ( ~n8405 & n8847 ) ;
  assign n8849 = ( n8387 & ~n8848 ) | ( n8387 & n8395 ) | ( ~n8848 & n8395 ) ;
  assign n8850 = ( n8387 & ~n8849 ) | ( n8387 & 1'b0 ) | ( ~n8849 & 1'b0 ) ;
  assign n8851 = ( n8839 & ~x51 ) | ( n8839 & n8850 ) | ( ~x51 & n8850 ) ;
  assign n8853 = ( n8846 & ~n8852 ) | ( n8846 & n8851 ) | ( ~n8852 & n8851 ) ;
  assign n8843 = x50 | n8842 ;
  assign n8844 = x50 &  n8839 ;
  assign n8845 = ( n8407 & ~n8843 ) | ( n8407 & n8844 ) | ( ~n8843 & n8844 ) ;
  assign n8856 = n7982 | n8845 ;
  assign n8857 = ( n8853 & ~n8856 ) | ( n8853 & 1'b0 ) | ( ~n8856 & 1'b0 ) ;
  assign n8859 = ( n8407 & ~n8836 ) | ( n8407 & 1'b0 ) | ( ~n8836 & 1'b0 ) ;
  assign n8860 = ( n8827 & ~n8859 ) | ( n8827 & n8831 ) | ( ~n8859 & n8831 ) ;
  assign n8861 = ( n8827 & ~n8860 ) | ( n8827 & 1'b0 ) | ( ~n8860 & 1'b0 ) ;
  assign n8862 = n8819 &  n8861 ;
  assign n8858 = ~n7983 & n8839 ;
  assign n8863 = ( n8858 & ~n8862 ) | ( n8858 & 1'b0 ) | ( ~n8862 & 1'b0 ) ;
  assign n8864 = ( x52 & n8862 ) | ( x52 & n8863 ) | ( n8862 & n8863 ) ;
  assign n8865 = x52 | n8862 ;
  assign n8866 = n8858 | n8865 ;
  assign n8867 = ~n8864 & n8866 ;
  assign n8868 = n8857 | n8867 ;
  assign n8854 = n8845 &  n8853 ;
  assign n8855 = ( n7982 & ~n8853 ) | ( n7982 & n8854 ) | ( ~n8853 & n8854 ) ;
  assign n8887 = ( n7572 & ~n8855 ) | ( n7572 & 1'b0 ) | ( ~n8855 & 1'b0 ) ;
  assign n8888 = n8868 &  n8887 ;
  assign n8889 = n8879 | n8888 ;
  assign n8890 = ~n8845 & n8853 ;
  assign n8891 = ( n8867 & ~n7982 ) | ( n8867 & n8890 ) | ( ~n7982 & n8890 ) ;
  assign n8892 = n7572 | n8891 ;
  assign n8893 = n7169 &  n8892 ;
  assign n8894 = n8889 &  n8893 ;
  assign n8895 = n8886 | n8894 ;
  assign n8869 = ~n8855 & n8868 ;
  assign n8880 = ( n7572 & n8869 ) | ( n7572 & n8879 ) | ( n8869 & n8879 ) ;
  assign n8881 = n7169 | n8880 ;
  assign n8909 = ~n6781 & n8881 ;
  assign n8910 = n8895 &  n8909 ;
  assign n8911 = n8901 | n8910 ;
  assign n8912 = n8889 &  n8892 ;
  assign n8913 = ( n7169 & n8886 ) | ( n7169 & n8912 ) | ( n8886 & n8912 ) ;
  assign n8914 = ( n6781 & ~n8913 ) | ( n6781 & 1'b0 ) | ( ~n8913 & 1'b0 ) ;
  assign n8915 = ( n6399 & ~n8914 ) | ( n6399 & 1'b0 ) | ( ~n8914 & 1'b0 ) ;
  assign n8916 = n8911 &  n8915 ;
  assign n8917 = n8908 | n8916 ;
  assign n8896 = n8881 &  n8895 ;
  assign n8902 = ( n8896 & ~n6781 ) | ( n8896 & n8901 ) | ( ~n6781 & n8901 ) ;
  assign n8903 = n6399 | n8902 ;
  assign n8931 = ~n6032 & n8903 ;
  assign n8932 = n8917 &  n8931 ;
  assign n8933 = ( n8923 & ~n8932 ) | ( n8923 & 1'b0 ) | ( ~n8932 & 1'b0 ) ;
  assign n8934 = ( n8911 & ~n8914 ) | ( n8911 & 1'b0 ) | ( ~n8914 & 1'b0 ) ;
  assign n8935 = ( n6399 & n8908 ) | ( n6399 & n8934 ) | ( n8908 & n8934 ) ;
  assign n8936 = ( n6032 & ~n8935 ) | ( n6032 & 1'b0 ) | ( ~n8935 & 1'b0 ) ;
  assign n8937 = ( n5672 & ~n8936 ) | ( n5672 & 1'b0 ) | ( ~n8936 & 1'b0 ) ;
  assign n8938 = ~n8933 & n8937 ;
  assign n8939 = ( n8930 & ~n8938 ) | ( n8930 & 1'b0 ) | ( ~n8938 & 1'b0 ) ;
  assign n8918 = n8903 &  n8917 ;
  assign n8924 = ( n6032 & ~n8918 ) | ( n6032 & n8923 ) | ( ~n8918 & n8923 ) ;
  assign n8925 = ~n5672 & n8924 ;
  assign n8953 = n5327 | n8925 ;
  assign n8954 = n8939 | n8953 ;
  assign n8955 = ~n8945 & n8954 ;
  assign n8956 = n8933 | n8936 ;
  assign n8957 = ( n8930 & ~n5672 ) | ( n8930 & n8956 ) | ( ~n5672 & n8956 ) ;
  assign n8958 = n5327 &  n8957 ;
  assign n8959 = n4990 | n8958 ;
  assign n8960 = n8955 | n8959 ;
  assign n8961 = ~n8952 & n8960 ;
  assign n8940 = n8925 | n8939 ;
  assign n8946 = ( n5327 & ~n8945 ) | ( n5327 & n8940 ) | ( ~n8945 & n8940 ) ;
  assign n8947 = n4990 &  n8946 ;
  assign n8975 = n4668 | n8947 ;
  assign n8976 = n8961 | n8975 ;
  assign n8977 = ~n8967 & n8976 ;
  assign n8978 = n8955 | n8958 ;
  assign n8979 = ( n4990 & ~n8952 ) | ( n4990 & n8978 ) | ( ~n8952 & n8978 ) ;
  assign n8980 = n4668 &  n8979 ;
  assign n9000 = n8977 | n8980 ;
  assign n9001 = ( n4353 & ~n8974 ) | ( n4353 & n9000 ) | ( ~n8974 & n9000 ) ;
  assign n9002 = n4053 &  n9001 ;
  assign n9248 = n8785 | n8839 ;
  assign n9249 = ( n8790 & ~n8785 ) | ( n8790 & n8798 ) | ( ~n8785 & n8798 ) ;
  assign n9251 = ( n8785 & n9248 ) | ( n8785 & n9249 ) | ( n9248 & n9249 ) ;
  assign n9250 = ( n8798 & ~n9249 ) | ( n8798 & n9248 ) | ( ~n9249 & n9248 ) ;
  assign n9252 = ( n8790 & ~n9251 ) | ( n8790 & n9250 ) | ( ~n9251 & n9250 ) ;
  assign n9182 = ~n8732 & n8839 ;
  assign n9183 = ( n8719 & n8724 ) | ( n8719 & n8839 ) | ( n8724 & n8839 ) ;
  assign n9185 = ( n9182 & ~n8719 ) | ( n9182 & n9183 ) | ( ~n8719 & n9183 ) ;
  assign n9184 = ( n8839 & ~n9183 ) | ( n8839 & n9182 ) | ( ~n9183 & n9182 ) ;
  assign n9186 = ( n8724 & ~n9185 ) | ( n8724 & n9184 ) | ( ~n9185 & n9184 ) ;
  assign n9116 = n8666 &  n8839 ;
  assign n9117 = ( n8653 & ~n9116 ) | ( n8653 & n8839 ) | ( ~n9116 & n8839 ) ;
  assign n9118 = ( n8658 & ~n8653 ) | ( n8658 & n9117 ) | ( ~n8653 & n9117 ) ;
  assign n9119 = ( n8653 & ~n9117 ) | ( n8653 & n8658 ) | ( ~n9117 & n8658 ) ;
  assign n9120 = ( n9118 & ~n8658 ) | ( n9118 & n9119 ) | ( ~n8658 & n9119 ) ;
  assign n9028 = ~n8578 & n8839 ;
  assign n9029 = ( n8565 & ~n9028 ) | ( n8565 & n8839 ) | ( ~n9028 & n8839 ) ;
  assign n9030 = ( n8570 & ~n8565 ) | ( n8570 & n9029 ) | ( ~n8565 & n9029 ) ;
  assign n9031 = ( n8565 & ~n9029 ) | ( n8565 & n8570 ) | ( ~n9029 & n8570 ) ;
  assign n9032 = ( n9030 & ~n8570 ) | ( n9030 & n9031 ) | ( ~n8570 & n9031 ) ;
  assign n9007 = ( n8544 & n8552 ) | ( n8544 & n8556 ) | ( n8552 & n8556 ) ;
  assign n9008 = ( n8839 & ~n8552 ) | ( n8839 & n9007 ) | ( ~n8552 & n9007 ) ;
  assign n9009 = ( n8544 & ~n9007 ) | ( n8544 & n8839 ) | ( ~n9007 & n8839 ) ;
  assign n9010 = ( n8556 & ~n9008 ) | ( n8556 & n9009 ) | ( ~n9008 & n9009 ) ;
  assign n8962 = n8947 | n8961 ;
  assign n8968 = ( n4668 & ~n8967 ) | ( n4668 & n8962 ) | ( ~n8967 & n8962 ) ;
  assign n8969 = n4353 &  n8968 ;
  assign n8981 = n4353 | n8980 ;
  assign n8982 = n8977 | n8981 ;
  assign n8983 = ~n8974 & n8982 ;
  assign n8984 = n8969 | n8983 ;
  assign n8990 = ( n4053 & n8984 ) | ( n4053 & n8989 ) | ( n8984 & n8989 ) ;
  assign n8991 = n3760 &  n8990 ;
  assign n8993 = ( n8546 & ~n8542 ) | ( n8546 & n8550 ) | ( ~n8542 & n8550 ) ;
  assign n8992 = n8550 | n8839 ;
  assign n8995 = ( n8550 & ~n8993 ) | ( n8550 & n8992 ) | ( ~n8993 & n8992 ) ;
  assign n8994 = ( n8992 & ~n8546 ) | ( n8992 & n8993 ) | ( ~n8546 & n8993 ) ;
  assign n8996 = ( n8542 & ~n8995 ) | ( n8542 & n8994 ) | ( ~n8995 & n8994 ) ;
  assign n8997 = n4053 | n8969 ;
  assign n8998 = n8983 | n8997 ;
  assign n8999 = n8989 &  n8998 ;
  assign n9003 = n3760 | n9002 ;
  assign n9004 = n8999 | n9003 ;
  assign n9005 = ~n8996 & n9004 ;
  assign n9006 = n8991 | n9005 ;
  assign n9011 = ( n3482 & ~n9010 ) | ( n3482 & n9006 ) | ( ~n9010 & n9006 ) ;
  assign n9012 = n3211 &  n9011 ;
  assign n9013 = n8576 | n8839 ;
  assign n9014 = ( n8563 & n8572 ) | ( n8563 & n8576 ) | ( n8572 & n8576 ) ;
  assign n9015 = ( n9013 & ~n8572 ) | ( n9013 & n9014 ) | ( ~n8572 & n9014 ) ;
  assign n9016 = ( n8576 & ~n9014 ) | ( n8576 & n9013 ) | ( ~n9014 & n9013 ) ;
  assign n9017 = ( n8563 & ~n9015 ) | ( n8563 & n9016 ) | ( ~n9015 & n9016 ) ;
  assign n9018 = n3482 | n8991 ;
  assign n9019 = n9005 | n9018 ;
  assign n9020 = ~n9010 & n9019 ;
  assign n9021 = n8999 | n9002 ;
  assign n9022 = ( n3760 & ~n8996 ) | ( n3760 & n9021 ) | ( ~n8996 & n9021 ) ;
  assign n9023 = n3482 &  n9022 ;
  assign n9024 = n3211 | n9023 ;
  assign n9025 = n9020 | n9024 ;
  assign n9026 = n9017 &  n9025 ;
  assign n9027 = n9012 | n9026 ;
  assign n9033 = ( n2955 & ~n9032 ) | ( n2955 & n9027 ) | ( ~n9032 & n9027 ) ;
  assign n9034 = n2706 &  n9033 ;
  assign n9035 = n8598 | n8839 ;
  assign n9036 = ( n8585 & n8594 ) | ( n8585 & n8598 ) | ( n8594 & n8598 ) ;
  assign n9037 = ( n9035 & ~n8594 ) | ( n9035 & n9036 ) | ( ~n8594 & n9036 ) ;
  assign n9038 = ( n8598 & ~n9036 ) | ( n8598 & n9035 ) | ( ~n9036 & n9035 ) ;
  assign n9039 = ( n8585 & ~n9037 ) | ( n8585 & n9038 ) | ( ~n9037 & n9038 ) ;
  assign n9040 = n2955 | n9012 ;
  assign n9041 = n9026 | n9040 ;
  assign n9042 = ~n9032 & n9041 ;
  assign n9043 = n9020 | n9023 ;
  assign n9044 = ( n3211 & n9017 ) | ( n3211 & n9043 ) | ( n9017 & n9043 ) ;
  assign n9045 = n2955 &  n9044 ;
  assign n9046 = n2706 | n9045 ;
  assign n9047 = n9042 | n9046 ;
  assign n9048 = n9039 &  n9047 ;
  assign n9049 = n9034 | n9048 ;
  assign n9051 = ( n8587 & ~n8592 ) | ( n8587 & n8839 ) | ( ~n8592 & n8839 ) ;
  assign n9050 = ~n8600 & n8839 ;
  assign n9052 = ( n8839 & ~n9051 ) | ( n8839 & n9050 ) | ( ~n9051 & n9050 ) ;
  assign n9053 = ( n9050 & ~n8587 ) | ( n9050 & n9051 ) | ( ~n8587 & n9051 ) ;
  assign n9054 = ( n8592 & ~n9052 ) | ( n8592 & n9053 ) | ( ~n9052 & n9053 ) ;
  assign n9055 = ( n2472 & n9049 ) | ( n2472 & n9054 ) | ( n9049 & n9054 ) ;
  assign n9056 = n2245 &  n9055 ;
  assign n9057 = n8620 | n8839 ;
  assign n9058 = ( n8607 & n8616 ) | ( n8607 & n8620 ) | ( n8616 & n8620 ) ;
  assign n9059 = ( n9057 & ~n8616 ) | ( n9057 & n9058 ) | ( ~n8616 & n9058 ) ;
  assign n9060 = ( n8620 & ~n9058 ) | ( n8620 & n9057 ) | ( ~n9058 & n9057 ) ;
  assign n9061 = ( n8607 & ~n9059 ) | ( n8607 & n9060 ) | ( ~n9059 & n9060 ) ;
  assign n9062 = n2472 | n9034 ;
  assign n9063 = n9048 | n9062 ;
  assign n9064 = n9054 &  n9063 ;
  assign n9065 = n9042 | n9045 ;
  assign n9066 = ( n2706 & n9039 ) | ( n2706 & n9065 ) | ( n9039 & n9065 ) ;
  assign n9067 = n2472 &  n9066 ;
  assign n9068 = n2245 | n9067 ;
  assign n9069 = n9064 | n9068 ;
  assign n9070 = n9061 &  n9069 ;
  assign n9071 = n9056 | n9070 ;
  assign n9073 = ( n8609 & ~n8614 ) | ( n8609 & n8839 ) | ( ~n8614 & n8839 ) ;
  assign n9072 = ~n8622 & n8839 ;
  assign n9074 = ( n8839 & ~n9073 ) | ( n8839 & n9072 ) | ( ~n9073 & n9072 ) ;
  assign n9075 = ( n9072 & ~n8609 ) | ( n9072 & n9073 ) | ( ~n8609 & n9073 ) ;
  assign n9076 = ( n8614 & ~n9074 ) | ( n8614 & n9075 ) | ( ~n9074 & n9075 ) ;
  assign n9077 = ( n9071 & ~n2033 ) | ( n9071 & n9076 ) | ( ~n2033 & n9076 ) ;
  assign n9078 = n1827 &  n9077 ;
  assign n9079 = n8642 | n8839 ;
  assign n9080 = ( n8629 & ~n8638 ) | ( n8629 & n8642 ) | ( ~n8638 & n8642 ) ;
  assign n9081 = ( n8638 & n9079 ) | ( n8638 & n9080 ) | ( n9079 & n9080 ) ;
  assign n9082 = ( n8642 & ~n9080 ) | ( n8642 & n9079 ) | ( ~n9080 & n9079 ) ;
  assign n9083 = ( n8629 & ~n9081 ) | ( n8629 & n9082 ) | ( ~n9081 & n9082 ) ;
  assign n9084 = ( n2033 & ~n9056 ) | ( n2033 & 1'b0 ) | ( ~n9056 & 1'b0 ) ;
  assign n9085 = ~n9070 & n9084 ;
  assign n9086 = ( n9076 & ~n9085 ) | ( n9076 & 1'b0 ) | ( ~n9085 & 1'b0 ) ;
  assign n9087 = n9064 | n9067 ;
  assign n9088 = ( n2245 & n9061 ) | ( n2245 & n9087 ) | ( n9061 & n9087 ) ;
  assign n9089 = ~n2033 & n9088 ;
  assign n9090 = n1827 | n9089 ;
  assign n9091 = n9086 | n9090 ;
  assign n9092 = n9083 &  n9091 ;
  assign n9093 = n9078 | n9092 ;
  assign n9094 = ~n8644 & n8839 ;
  assign n9095 = ( n8631 & n8636 ) | ( n8631 & n8839 ) | ( n8636 & n8839 ) ;
  assign n9097 = ( n9094 & ~n8631 ) | ( n9094 & n9095 ) | ( ~n8631 & n9095 ) ;
  assign n9096 = ( n8839 & ~n9095 ) | ( n8839 & n9094 ) | ( ~n9095 & n9094 ) ;
  assign n9098 = ( n8636 & ~n9097 ) | ( n8636 & n9096 ) | ( ~n9097 & n9096 ) ;
  assign n9099 = ( n9093 & ~n1636 ) | ( n9093 & n9098 ) | ( ~n1636 & n9098 ) ;
  assign n9100 = ~n1452 & n9099 ;
  assign n9101 = n8664 | n8839 ;
  assign n9102 = ( n8651 & ~n8660 ) | ( n8651 & n8664 ) | ( ~n8660 & n8664 ) ;
  assign n9103 = ( n8660 & n9101 ) | ( n8660 & n9102 ) | ( n9101 & n9102 ) ;
  assign n9104 = ( n8664 & ~n9102 ) | ( n8664 & n9101 ) | ( ~n9102 & n9101 ) ;
  assign n9105 = ( n8651 & ~n9103 ) | ( n8651 & n9104 ) | ( ~n9103 & n9104 ) ;
  assign n9106 = ( n1636 & ~n9078 ) | ( n1636 & 1'b0 ) | ( ~n9078 & 1'b0 ) ;
  assign n9107 = ~n9092 & n9106 ;
  assign n9108 = ( n9098 & ~n9107 ) | ( n9098 & 1'b0 ) | ( ~n9107 & 1'b0 ) ;
  assign n9109 = n9086 | n9089 ;
  assign n9110 = ( n1827 & n9083 ) | ( n1827 & n9109 ) | ( n9083 & n9109 ) ;
  assign n9111 = ~n1636 & n9110 ;
  assign n9112 = ( n1452 & ~n9111 ) | ( n1452 & 1'b0 ) | ( ~n9111 & 1'b0 ) ;
  assign n9113 = ~n9108 & n9112 ;
  assign n9114 = ( n9105 & ~n9113 ) | ( n9105 & 1'b0 ) | ( ~n9113 & 1'b0 ) ;
  assign n9115 = n9100 | n9114 ;
  assign n9121 = ( n1283 & ~n9120 ) | ( n1283 & n9115 ) | ( ~n9120 & n9115 ) ;
  assign n9122 = ~n1122 & n9121 ;
  assign n9123 = n8686 | n8839 ;
  assign n9124 = ( n8673 & ~n8686 ) | ( n8673 & n8682 ) | ( ~n8686 & n8682 ) ;
  assign n9126 = ( n8686 & n9123 ) | ( n8686 & n9124 ) | ( n9123 & n9124 ) ;
  assign n9125 = ( n8682 & ~n9124 ) | ( n8682 & n9123 ) | ( ~n9124 & n9123 ) ;
  assign n9127 = ( n8673 & ~n9126 ) | ( n8673 & n9125 ) | ( ~n9126 & n9125 ) ;
  assign n9128 = n1283 | n9100 ;
  assign n9129 = n9114 | n9128 ;
  assign n9130 = ~n9120 & n9129 ;
  assign n9131 = n9108 | n9111 ;
  assign n9132 = ( n9105 & ~n1452 ) | ( n9105 & n9131 ) | ( ~n1452 & n9131 ) ;
  assign n9133 = n1283 &  n9132 ;
  assign n9134 = ( n1122 & ~n9133 ) | ( n1122 & 1'b0 ) | ( ~n9133 & 1'b0 ) ;
  assign n9135 = ~n9130 & n9134 ;
  assign n9136 = n9127 | n9135 ;
  assign n9137 = ~n9122 & n9136 ;
  assign n9138 = n8688 &  n8839 ;
  assign n9139 = ( n8680 & ~n8675 ) | ( n8680 & n8839 ) | ( ~n8675 & n8839 ) ;
  assign n9141 = ( n8675 & n9138 ) | ( n8675 & n9139 ) | ( n9138 & n9139 ) ;
  assign n9140 = ( n8839 & ~n9139 ) | ( n8839 & n9138 ) | ( ~n9139 & n9138 ) ;
  assign n9142 = ( n8680 & ~n9141 ) | ( n8680 & n9140 ) | ( ~n9141 & n9140 ) ;
  assign n9143 = ( n976 & n9137 ) | ( n976 & n9142 ) | ( n9137 & n9142 ) ;
  assign n9144 = ( n837 & ~n9143 ) | ( n837 & 1'b0 ) | ( ~n9143 & 1'b0 ) ;
  assign n9145 = ( n8708 & ~n8839 ) | ( n8708 & 1'b0 ) | ( ~n8839 & 1'b0 ) ;
  assign n9146 = ( n8695 & n8704 ) | ( n8695 & n8708 ) | ( n8704 & n8708 ) ;
  assign n9147 = ( n9145 & ~n8704 ) | ( n9145 & n9146 ) | ( ~n8704 & n9146 ) ;
  assign n9148 = ( n8708 & ~n9146 ) | ( n8708 & n9145 ) | ( ~n9146 & n9145 ) ;
  assign n9149 = ( n8695 & ~n9147 ) | ( n8695 & n9148 ) | ( ~n9147 & n9148 ) ;
  assign n9150 = ( n976 & ~n9122 ) | ( n976 & 1'b0 ) | ( ~n9122 & 1'b0 ) ;
  assign n9151 = n9136 &  n9150 ;
  assign n9152 = n9142 | n9151 ;
  assign n9153 = n9130 | n9133 ;
  assign n9154 = ( n1122 & ~n9153 ) | ( n1122 & n9127 ) | ( ~n9153 & n9127 ) ;
  assign n9155 = n976 | n9154 ;
  assign n9156 = ~n837 & n9155 ;
  assign n9157 = n9152 &  n9156 ;
  assign n9158 = n9149 | n9157 ;
  assign n9159 = ~n9144 & n9158 ;
  assign n9161 = ( n8697 & ~n8702 ) | ( n8697 & n8839 ) | ( ~n8702 & n8839 ) ;
  assign n9160 = n8710 &  n8839 ;
  assign n9162 = ( n8839 & ~n9161 ) | ( n8839 & n9160 ) | ( ~n9161 & n9160 ) ;
  assign n9163 = ( n9160 & ~n8697 ) | ( n9160 & n9161 ) | ( ~n8697 & n9161 ) ;
  assign n9164 = ( n8702 & ~n9162 ) | ( n8702 & n9163 ) | ( ~n9162 & n9163 ) ;
  assign n9165 = ( n713 & ~n9159 ) | ( n713 & n9164 ) | ( ~n9159 & n9164 ) ;
  assign n9166 = n595 &  n9165 ;
  assign n9167 = n8730 | n8839 ;
  assign n9168 = ( n8717 & n8726 ) | ( n8717 & n8730 ) | ( n8726 & n8730 ) ;
  assign n9169 = ( n9167 & ~n8726 ) | ( n9167 & n9168 ) | ( ~n8726 & n9168 ) ;
  assign n9170 = ( n8730 & ~n9168 ) | ( n8730 & n9167 ) | ( ~n9168 & n9167 ) ;
  assign n9171 = ( n8717 & ~n9169 ) | ( n8717 & n9170 ) | ( ~n9169 & n9170 ) ;
  assign n9172 = n713 | n9144 ;
  assign n9173 = ( n9158 & ~n9172 ) | ( n9158 & 1'b0 ) | ( ~n9172 & 1'b0 ) ;
  assign n9174 = ( n9164 & ~n9173 ) | ( n9164 & 1'b0 ) | ( ~n9173 & 1'b0 ) ;
  assign n9175 = n9152 &  n9155 ;
  assign n9176 = ( n9149 & ~n837 ) | ( n9149 & n9175 ) | ( ~n837 & n9175 ) ;
  assign n9177 = ( n713 & ~n9176 ) | ( n713 & 1'b0 ) | ( ~n9176 & 1'b0 ) ;
  assign n9178 = n595 | n9177 ;
  assign n9179 = n9174 | n9178 ;
  assign n9180 = n9171 &  n9179 ;
  assign n9181 = n9166 | n9180 ;
  assign n9187 = ( n492 & ~n9186 ) | ( n492 & n9181 ) | ( ~n9186 & n9181 ) ;
  assign n9188 = n396 &  n9187 ;
  assign n9189 = n8752 | n8839 ;
  assign n9190 = ( n8739 & n8748 ) | ( n8739 & n8752 ) | ( n8748 & n8752 ) ;
  assign n9191 = ( n9189 & ~n8748 ) | ( n9189 & n9190 ) | ( ~n8748 & n9190 ) ;
  assign n9192 = ( n8752 & ~n9190 ) | ( n8752 & n9189 ) | ( ~n9190 & n9189 ) ;
  assign n9193 = ( n8739 & ~n9191 ) | ( n8739 & n9192 ) | ( ~n9191 & n9192 ) ;
  assign n9194 = n492 | n9166 ;
  assign n9195 = n9180 | n9194 ;
  assign n9196 = ~n9186 & n9195 ;
  assign n9197 = n9174 | n9177 ;
  assign n9198 = ( n595 & n9171 ) | ( n595 & n9197 ) | ( n9171 & n9197 ) ;
  assign n9199 = n492 &  n9198 ;
  assign n9200 = n396 | n9199 ;
  assign n9201 = n9196 | n9200 ;
  assign n9202 = n9193 &  n9201 ;
  assign n9203 = n9188 | n9202 ;
  assign n9205 = ( n8741 & ~n8746 ) | ( n8741 & n8839 ) | ( ~n8746 & n8839 ) ;
  assign n9204 = ~n8754 & n8839 ;
  assign n9206 = ( n8839 & ~n9205 ) | ( n8839 & n9204 ) | ( ~n9205 & n9204 ) ;
  assign n9207 = ( n9204 & ~n8741 ) | ( n9204 & n9205 ) | ( ~n8741 & n9205 ) ;
  assign n9208 = ( n8746 & ~n9206 ) | ( n8746 & n9207 ) | ( ~n9206 & n9207 ) ;
  assign n9209 = ( n315 & n9203 ) | ( n315 & n9208 ) | ( n9203 & n9208 ) ;
  assign n9210 = n240 &  n9209 ;
  assign n9212 = ( n8770 & ~n8761 ) | ( n8770 & n8774 ) | ( ~n8761 & n8774 ) ;
  assign n9211 = n8774 | n8839 ;
  assign n9214 = ( n8774 & ~n9212 ) | ( n8774 & n9211 ) | ( ~n9212 & n9211 ) ;
  assign n9213 = ( n9211 & ~n8770 ) | ( n9211 & n9212 ) | ( ~n8770 & n9212 ) ;
  assign n9215 = ( n8761 & ~n9214 ) | ( n8761 & n9213 ) | ( ~n9214 & n9213 ) ;
  assign n9216 = n315 | n9188 ;
  assign n9217 = n9202 | n9216 ;
  assign n9218 = n9208 &  n9217 ;
  assign n9219 = n9196 | n9199 ;
  assign n9220 = ( n396 & n9193 ) | ( n396 & n9219 ) | ( n9193 & n9219 ) ;
  assign n9221 = n315 &  n9220 ;
  assign n9222 = n240 | n9221 ;
  assign n9223 = n9218 | n9222 ;
  assign n9224 = ~n9215 & n9223 ;
  assign n9225 = n9210 | n9224 ;
  assign n9226 = ~n8776 & n8839 ;
  assign n9227 = ( n8763 & n8768 ) | ( n8763 & n8839 ) | ( n8768 & n8839 ) ;
  assign n9229 = ( n9226 & ~n8763 ) | ( n9226 & n9227 ) | ( ~n8763 & n9227 ) ;
  assign n9228 = ( n8839 & ~n9227 ) | ( n8839 & n9226 ) | ( ~n9227 & n9226 ) ;
  assign n9230 = ( n8768 & ~n9229 ) | ( n8768 & n9228 ) | ( ~n9229 & n9228 ) ;
  assign n9231 = ( n181 & n9225 ) | ( n181 & n9230 ) | ( n9225 & n9230 ) ;
  assign n9232 = ~n145 & n9231 ;
  assign n9234 = ( n8792 & ~n8783 ) | ( n8792 & n8796 ) | ( ~n8783 & n8796 ) ;
  assign n9233 = n8796 | n8839 ;
  assign n9236 = ( n8796 & ~n9234 ) | ( n8796 & n9233 ) | ( ~n9234 & n9233 ) ;
  assign n9235 = ( n9233 & ~n8792 ) | ( n9233 & n9234 ) | ( ~n8792 & n9234 ) ;
  assign n9237 = ( n8783 & ~n9236 ) | ( n8783 & n9235 ) | ( ~n9236 & n9235 ) ;
  assign n9238 = n181 | n9210 ;
  assign n9239 = n9224 | n9238 ;
  assign n9240 = n9230 &  n9239 ;
  assign n9241 = n9218 | n9221 ;
  assign n9242 = ( n240 & ~n9215 ) | ( n240 & n9241 ) | ( ~n9215 & n9241 ) ;
  assign n9243 = n181 &  n9242 ;
  assign n9244 = ( n145 & ~n9243 ) | ( n145 & 1'b0 ) | ( ~n9243 & 1'b0 ) ;
  assign n9245 = ~n9240 & n9244 ;
  assign n9246 = ( n9237 & ~n9245 ) | ( n9237 & 1'b0 ) | ( ~n9245 & 1'b0 ) ;
  assign n9247 = n9232 | n9246 ;
  assign n9253 = ( n150 & ~n9252 ) | ( n150 & n9247 ) | ( ~n9252 & n9247 ) ;
  assign n9254 = n8805 | n8821 ;
  assign n9255 = ( n8824 & ~n9254 ) | ( n8824 & n8839 ) | ( ~n9254 & n8839 ) ;
  assign n9256 = ~n8824 & n9255 ;
  assign n9257 = n8821 | n8824 ;
  assign n9258 = n8839 | n9257 ;
  assign n9259 = ( n8805 & ~n9258 ) | ( n8805 & n9257 ) | ( ~n9258 & n9257 ) ;
  assign n9260 = n9256 | n9259 ;
  assign n9261 = n8806 &  n8813 ;
  assign n9262 = ~n8839 & n9261 ;
  assign n9263 = ( n8827 & ~n9261 ) | ( n8827 & n9262 ) | ( ~n9261 & n9262 ) ;
  assign n9264 = n9260 &  n9263 ;
  assign n9265 = ~n9253 & n9264 ;
  assign n9266 = ( n133 & ~n9265 ) | ( n133 & n9264 ) | ( ~n9265 & n9264 ) ;
  assign n9269 = n9240 | n9243 ;
  assign n9270 = ( n9237 & ~n145 ) | ( n9237 & n9269 ) | ( ~n145 & n9269 ) ;
  assign n9271 = n150 &  n9270 ;
  assign n9272 = n9260 | n9271 ;
  assign n9267 = n150 | n9232 ;
  assign n9268 = n9246 | n9267 ;
  assign n9273 = n9252 | n9268 ;
  assign n9274 = ( n9272 & ~n9252 ) | ( n9272 & n9273 ) | ( ~n9252 & n9273 ) ;
  assign n9276 = ( n133 & n8806 ) | ( n133 & n8813 ) | ( n8806 & n8813 ) ;
  assign n9275 = ( n8806 & ~n8839 ) | ( n8806 & n8813 ) | ( ~n8839 & n8813 ) ;
  assign n9277 = ( n8813 & ~n9275 ) | ( n8813 & 1'b0 ) | ( ~n9275 & 1'b0 ) ;
  assign n9278 = ( n9276 & ~n8813 ) | ( n9276 & n9277 ) | ( ~n8813 & n9277 ) ;
  assign n9279 = n8809 | n8836 ;
  assign n9280 = ( n8831 & ~n8812 ) | ( n8831 & n9279 ) | ( ~n8812 & n9279 ) ;
  assign n9281 = n8812 | n9280 ;
  assign n9282 = ( n8819 & ~n8827 ) | ( n8819 & n9281 ) | ( ~n8827 & n9281 ) ;
  assign n9283 = ( n8819 & ~n9282 ) | ( n8819 & 1'b0 ) | ( ~n9282 & 1'b0 ) ;
  assign n9284 = n9278 | n9283 ;
  assign n9285 = ( n9274 & ~n9284 ) | ( n9274 & 1'b0 ) | ( ~n9284 & 1'b0 ) ;
  assign n9286 = ~n9266 | ~n9285 ;
  assign n9446 = n9002 | n9286 ;
  assign n9447 = ( n8989 & n8998 ) | ( n8989 & n9002 ) | ( n8998 & n9002 ) ;
  assign n9448 = ( n9446 & ~n8998 ) | ( n9446 & n9447 ) | ( ~n8998 & n9447 ) ;
  assign n9449 = ( n9002 & ~n9447 ) | ( n9002 & n9446 ) | ( ~n9447 & n9446 ) ;
  assign n9450 = ( n8989 & ~n9448 ) | ( n8989 & n9449 ) | ( ~n9448 & n9449 ) ;
  assign n9680 = ~n9223 & n9286 ;
  assign n9681 = ( n9210 & n9215 ) | ( n9210 & n9286 ) | ( n9215 & n9286 ) ;
  assign n9683 = ( n9680 & ~n9210 ) | ( n9680 & n9681 ) | ( ~n9210 & n9681 ) ;
  assign n9682 = ( n9286 & ~n9681 ) | ( n9286 & n9680 ) | ( ~n9681 & n9680 ) ;
  assign n9684 = ( n9215 & ~n9683 ) | ( n9215 & n9682 ) | ( ~n9683 & n9682 ) ;
  assign n9462 = ( n8991 & ~n8996 ) | ( n8991 & n9286 ) | ( ~n8996 & n9286 ) ;
  assign n9461 = ~n9004 & n9286 ;
  assign n9463 = ( n9286 & ~n9462 ) | ( n9286 & n9461 ) | ( ~n9462 & n9461 ) ;
  assign n9464 = ( n9461 & ~n8991 ) | ( n9461 & n9462 ) | ( ~n8991 & n9462 ) ;
  assign n9465 = ( n8996 & ~n9463 ) | ( n8996 & n9464 ) | ( ~n9463 & n9464 ) ;
  assign n9440 = ( n8969 & ~n8974 ) | ( n8969 & n9286 ) | ( ~n8974 & n9286 ) ;
  assign n9439 = ~n8982 & n9286 ;
  assign n9441 = ( n9286 & ~n9440 ) | ( n9286 & n9439 ) | ( ~n9440 & n9439 ) ;
  assign n9442 = ( n9439 & ~n8969 ) | ( n9439 & n9440 ) | ( ~n8969 & n9440 ) ;
  assign n9443 = ( n8974 & ~n9441 ) | ( n8974 & n9442 ) | ( ~n9441 & n9442 ) ;
  assign n9418 = ( n8947 & ~n8952 ) | ( n8947 & n8960 ) | ( ~n8952 & n8960 ) ;
  assign n9417 = n8947 | n9286 ;
  assign n9420 = ( n8947 & ~n9418 ) | ( n8947 & n9417 ) | ( ~n9418 & n9417 ) ;
  assign n9419 = ( n9417 & ~n8960 ) | ( n9417 & n9418 ) | ( ~n8960 & n9418 ) ;
  assign n9421 = ( n8952 & ~n9420 ) | ( n8952 & n9419 ) | ( ~n9420 & n9419 ) ;
  assign n8840 = x46 | x47 ;
  assign n8841 = x48 | n8840 ;
  assign n9287 = x48 &  n9286 ;
  assign n9288 = ( n8839 & ~n8841 ) | ( n8839 & n9287 ) | ( ~n8841 & n9287 ) ;
  assign n9289 = ( x48 & ~n9286 ) | ( x48 & x49 ) | ( ~n9286 & x49 ) ;
  assign n9295 = ( x48 & ~x49 ) | ( x48 & 1'b0 ) | ( ~x49 & 1'b0 ) ;
  assign n9290 = ~x48 & n8840 ;
  assign n9291 = ( x48 & ~n8837 ) | ( x48 & n9290 ) | ( ~n8837 & n9290 ) ;
  assign n9292 = ( n8827 & ~n8819 ) | ( n8827 & n9291 ) | ( ~n8819 & n9291 ) ;
  assign n9293 = n8819 &  n9292 ;
  assign n9294 = ( n9286 & ~x49 ) | ( n9286 & n9293 ) | ( ~x49 & n9293 ) ;
  assign n9296 = ( n9289 & ~n9295 ) | ( n9289 & n9294 ) | ( ~n9295 & n9294 ) ;
  assign n9297 = ~n9288 & n9296 ;
  assign n9299 = ( n8839 & ~n9283 ) | ( n8839 & 1'b0 ) | ( ~n9283 & 1'b0 ) ;
  assign n9300 = ( n9274 & ~n9299 ) | ( n9274 & n9278 ) | ( ~n9299 & n9278 ) ;
  assign n9301 = ( n9274 & ~n9300 ) | ( n9274 & 1'b0 ) | ( ~n9300 & 1'b0 ) ;
  assign n9302 = n9266 &  n9301 ;
  assign n9298 = ~n8842 & n9286 ;
  assign n9303 = ( n9298 & ~n9302 ) | ( n9298 & 1'b0 ) | ( ~n9302 & 1'b0 ) ;
  assign n9304 = ( x50 & n9302 ) | ( x50 & n9303 ) | ( n9302 & n9303 ) ;
  assign n9305 = x50 | n9302 ;
  assign n9306 = n9298 | n9305 ;
  assign n9307 = ~n9304 & n9306 ;
  assign n9308 = ( n9297 & ~n8407 ) | ( n9297 & n9307 ) | ( ~n8407 & n9307 ) ;
  assign n9309 = ( n7982 & ~n9308 ) | ( n7982 & 1'b0 ) | ( ~n9308 & 1'b0 ) ;
  assign n9313 = ~x50 & n8839 ;
  assign n9314 = ( x51 & ~n9313 ) | ( x51 & 1'b0 ) | ( ~n9313 & 1'b0 ) ;
  assign n9315 = n8858 | n9314 ;
  assign n9310 = ( n8839 & ~x50 ) | ( n8839 & n8850 ) | ( ~x50 & n8850 ) ;
  assign n9311 = x50 &  n9310 ;
  assign n9312 = ( n8845 & ~n9311 ) | ( n8845 & n8850 ) | ( ~n9311 & n8850 ) ;
  assign n9316 = ( n9286 & ~n9315 ) | ( n9286 & n9312 ) | ( ~n9315 & n9312 ) ;
  assign n9318 = ( n9286 & ~n9316 ) | ( n9286 & 1'b0 ) | ( ~n9316 & 1'b0 ) ;
  assign n9317 = ~n9312 & n9316 ;
  assign n9319 = ( n9315 & ~n9318 ) | ( n9315 & n9317 ) | ( ~n9318 & n9317 ) ;
  assign n9320 = n8407 | n9288 ;
  assign n9321 = ( n9296 & ~n9320 ) | ( n9296 & 1'b0 ) | ( ~n9320 & 1'b0 ) ;
  assign n9322 = n9307 | n9321 ;
  assign n9323 = n9288 &  n9296 ;
  assign n9324 = ( n8407 & ~n9296 ) | ( n8407 & n9323 ) | ( ~n9296 & n9323 ) ;
  assign n9325 = n7982 | n9324 ;
  assign n9326 = ( n9322 & ~n9325 ) | ( n9322 & 1'b0 ) | ( ~n9325 & 1'b0 ) ;
  assign n9327 = n9319 | n9326 ;
  assign n9328 = ~n9309 & n9327 ;
  assign n9329 = ( n8855 & ~n8857 ) | ( n8855 & 1'b0 ) | ( ~n8857 & 1'b0 ) ;
  assign n9330 = ( n8857 & ~n9329 ) | ( n8857 & n8867 ) | ( ~n9329 & n8867 ) ;
  assign n9332 = ( n9286 & n9329 ) | ( n9286 & n9330 ) | ( n9329 & n9330 ) ;
  assign n9331 = ( n8857 & ~n9330 ) | ( n8857 & n9286 ) | ( ~n9330 & n9286 ) ;
  assign n9333 = ( n8867 & ~n9332 ) | ( n8867 & n9331 ) | ( ~n9332 & n9331 ) ;
  assign n9334 = ( n7572 & n9328 ) | ( n7572 & n9333 ) | ( n9328 & n9333 ) ;
  assign n9335 = n7169 | n9334 ;
  assign n9336 = ( n8892 & ~n9286 ) | ( n8892 & 1'b0 ) | ( ~n9286 & 1'b0 ) ;
  assign n9337 = ( n8879 & n8888 ) | ( n8879 & n8892 ) | ( n8888 & n8892 ) ;
  assign n9338 = ( n9336 & ~n8888 ) | ( n9336 & n9337 ) | ( ~n8888 & n9337 ) ;
  assign n9339 = ( n8892 & ~n9337 ) | ( n8892 & n9336 ) | ( ~n9337 & n9336 ) ;
  assign n9340 = ( n8879 & ~n9338 ) | ( n8879 & n9339 ) | ( ~n9338 & n9339 ) ;
  assign n9341 = ( n7572 & ~n9309 ) | ( n7572 & 1'b0 ) | ( ~n9309 & 1'b0 ) ;
  assign n9342 = n9327 &  n9341 ;
  assign n9343 = n9333 | n9342 ;
  assign n9344 = ( n9322 & ~n9324 ) | ( n9322 & 1'b0 ) | ( ~n9324 & 1'b0 ) ;
  assign n9345 = ( n9319 & ~n7982 ) | ( n9319 & n9344 ) | ( ~n7982 & n9344 ) ;
  assign n9346 = n7572 | n9345 ;
  assign n9347 = n7169 &  n9346 ;
  assign n9348 = n9343 &  n9347 ;
  assign n9349 = n9340 | n9348 ;
  assign n9350 = n9335 &  n9349 ;
  assign n9351 = n8894 &  n9286 ;
  assign n9352 = ( n8881 & ~n9286 ) | ( n8881 & n8886 ) | ( ~n9286 & n8886 ) ;
  assign n9353 = ( n9286 & n9351 ) | ( n9286 & n9352 ) | ( n9351 & n9352 ) ;
  assign n9354 = ( n8881 & ~n9352 ) | ( n8881 & n9351 ) | ( ~n9352 & n9351 ) ;
  assign n9355 = ( n8886 & ~n9353 ) | ( n8886 & n9354 ) | ( ~n9353 & n9354 ) ;
  assign n9356 = ( n9350 & ~n6781 ) | ( n9350 & n9355 ) | ( ~n6781 & n9355 ) ;
  assign n9357 = n6399 | n9356 ;
  assign n9358 = n8914 | n9286 ;
  assign n9359 = ( n8901 & ~n8914 ) | ( n8901 & n8910 ) | ( ~n8914 & n8910 ) ;
  assign n9361 = ( n8914 & n9358 ) | ( n8914 & n9359 ) | ( n9358 & n9359 ) ;
  assign n9360 = ( n8910 & ~n9359 ) | ( n8910 & n9358 ) | ( ~n9359 & n9358 ) ;
  assign n9362 = ( n8901 & ~n9361 ) | ( n8901 & n9360 ) | ( ~n9361 & n9360 ) ;
  assign n9363 = ~n6781 & n9335 ;
  assign n9364 = n9349 &  n9363 ;
  assign n9365 = n9355 | n9364 ;
  assign n9366 = n9343 &  n9346 ;
  assign n9367 = ( n7169 & n9340 ) | ( n7169 & n9366 ) | ( n9340 & n9366 ) ;
  assign n9368 = ( n6781 & ~n9367 ) | ( n6781 & 1'b0 ) | ( ~n9367 & 1'b0 ) ;
  assign n9369 = ( n6399 & ~n9368 ) | ( n6399 & 1'b0 ) | ( ~n9368 & 1'b0 ) ;
  assign n9370 = n9365 &  n9369 ;
  assign n9371 = n9362 | n9370 ;
  assign n9372 = n9357 &  n9371 ;
  assign n9373 = n8916 &  n9286 ;
  assign n9374 = ( n8908 & ~n8903 ) | ( n8908 & n9286 ) | ( ~n8903 & n9286 ) ;
  assign n9376 = ( n8903 & n9373 ) | ( n8903 & n9374 ) | ( n9373 & n9374 ) ;
  assign n9375 = ( n9286 & ~n9374 ) | ( n9286 & n9373 ) | ( ~n9374 & n9373 ) ;
  assign n9377 = ( n8908 & ~n9376 ) | ( n8908 & n9375 ) | ( ~n9376 & n9375 ) ;
  assign n9378 = ( n9372 & ~n6032 ) | ( n9372 & n9377 ) | ( ~n6032 & n9377 ) ;
  assign n9379 = n5672 | n9378 ;
  assign n9380 = n8936 | n9286 ;
  assign n9381 = ( n8923 & ~n8936 ) | ( n8923 & n8932 ) | ( ~n8936 & n8932 ) ;
  assign n9383 = ( n8936 & n9380 ) | ( n8936 & n9381 ) | ( n9380 & n9381 ) ;
  assign n9382 = ( n8932 & ~n9381 ) | ( n8932 & n9380 ) | ( ~n9381 & n9380 ) ;
  assign n9384 = ( n8923 & ~n9383 ) | ( n8923 & n9382 ) | ( ~n9383 & n9382 ) ;
  assign n9385 = ~n6032 & n9357 ;
  assign n9386 = n9371 &  n9385 ;
  assign n9387 = n9377 | n9386 ;
  assign n9388 = ( n9365 & ~n9368 ) | ( n9365 & 1'b0 ) | ( ~n9368 & 1'b0 ) ;
  assign n9389 = ( n6399 & n9362 ) | ( n6399 & n9388 ) | ( n9362 & n9388 ) ;
  assign n9390 = ( n6032 & ~n9389 ) | ( n6032 & 1'b0 ) | ( ~n9389 & 1'b0 ) ;
  assign n9391 = ( n5672 & ~n9390 ) | ( n5672 & 1'b0 ) | ( ~n9390 & 1'b0 ) ;
  assign n9392 = n9387 &  n9391 ;
  assign n9393 = ( n9384 & ~n9392 ) | ( n9384 & 1'b0 ) | ( ~n9392 & 1'b0 ) ;
  assign n9394 = ( n9379 & ~n9393 ) | ( n9379 & 1'b0 ) | ( ~n9393 & 1'b0 ) ;
  assign n9395 = n8925 | n9286 ;
  assign n9396 = ( n8925 & ~n8938 ) | ( n8925 & n8930 ) | ( ~n8938 & n8930 ) ;
  assign n9397 = ( n8938 & n9395 ) | ( n8938 & n9396 ) | ( n9395 & n9396 ) ;
  assign n9398 = ( n8925 & ~n9396 ) | ( n8925 & n9395 ) | ( ~n9396 & n9395 ) ;
  assign n9399 = ( n8930 & ~n9397 ) | ( n8930 & n9398 ) | ( ~n9397 & n9398 ) ;
  assign n9400 = ( n5327 & ~n9394 ) | ( n5327 & n9399 ) | ( ~n9394 & n9399 ) ;
  assign n9401 = n4990 &  n9400 ;
  assign n9402 = n8958 | n9286 ;
  assign n9403 = ( n8945 & n8954 ) | ( n8945 & n8958 ) | ( n8954 & n8958 ) ;
  assign n9404 = ( n9402 & ~n8954 ) | ( n9402 & n9403 ) | ( ~n8954 & n9403 ) ;
  assign n9405 = ( n8958 & ~n9403 ) | ( n8958 & n9402 ) | ( ~n9403 & n9402 ) ;
  assign n9406 = ( n8945 & ~n9404 ) | ( n8945 & n9405 ) | ( ~n9404 & n9405 ) ;
  assign n9407 = ~n5327 & n9379 ;
  assign n9408 = ~n9393 & n9407 ;
  assign n9409 = ( n9399 & ~n9408 ) | ( n9399 & 1'b0 ) | ( ~n9408 & 1'b0 ) ;
  assign n9410 = ( n9387 & ~n9390 ) | ( n9387 & 1'b0 ) | ( ~n9390 & 1'b0 ) ;
  assign n9411 = ( n5672 & ~n9384 ) | ( n5672 & n9410 ) | ( ~n9384 & n9410 ) ;
  assign n9412 = ( n5327 & ~n9411 ) | ( n5327 & 1'b0 ) | ( ~n9411 & 1'b0 ) ;
  assign n9413 = n4990 | n9412 ;
  assign n9414 = n9409 | n9413 ;
  assign n9415 = ~n9406 & n9414 ;
  assign n9416 = n9401 | n9415 ;
  assign n9422 = ( n4668 & ~n9421 ) | ( n4668 & n9416 ) | ( ~n9421 & n9416 ) ;
  assign n9423 = n4353 &  n9422 ;
  assign n9425 = ( n8976 & ~n8967 ) | ( n8976 & n8980 ) | ( ~n8967 & n8980 ) ;
  assign n9424 = n8980 | n9286 ;
  assign n9427 = ( n8980 & ~n9425 ) | ( n8980 & n9424 ) | ( ~n9425 & n9424 ) ;
  assign n9426 = ( n9424 & ~n8976 ) | ( n9424 & n9425 ) | ( ~n8976 & n9425 ) ;
  assign n9428 = ( n8967 & ~n9427 ) | ( n8967 & n9426 ) | ( ~n9427 & n9426 ) ;
  assign n9429 = n4668 | n9401 ;
  assign n9430 = n9415 | n9429 ;
  assign n9431 = ~n9421 & n9430 ;
  assign n9432 = n9409 | n9412 ;
  assign n9433 = ( n4990 & ~n9406 ) | ( n4990 & n9432 ) | ( ~n9406 & n9432 ) ;
  assign n9434 = n4668 &  n9433 ;
  assign n9435 = n4353 | n9434 ;
  assign n9436 = n9431 | n9435 ;
  assign n9437 = ~n9428 & n9436 ;
  assign n9438 = n9423 | n9437 ;
  assign n9444 = ( n4053 & ~n9443 ) | ( n4053 & n9438 ) | ( ~n9443 & n9438 ) ;
  assign n9445 = n3760 &  n9444 ;
  assign n9451 = n4053 | n9423 ;
  assign n9452 = n9437 | n9451 ;
  assign n9453 = ~n9443 & n9452 ;
  assign n9454 = n9431 | n9434 ;
  assign n9455 = ( n4353 & ~n9428 ) | ( n4353 & n9454 ) | ( ~n9428 & n9454 ) ;
  assign n9456 = n4053 &  n9455 ;
  assign n9457 = n3760 | n9456 ;
  assign n9458 = n9453 | n9457 ;
  assign n9459 = n9450 &  n9458 ;
  assign n9460 = n9445 | n9459 ;
  assign n9466 = ( n3482 & ~n9465 ) | ( n3482 & n9460 ) | ( ~n9465 & n9460 ) ;
  assign n9467 = n3211 &  n9466 ;
  assign n9468 = n3482 | n9445 ;
  assign n9469 = n9459 | n9468 ;
  assign n9470 = ~n9465 & n9469 ;
  assign n9471 = n9453 | n9456 ;
  assign n9472 = ( n3760 & n9450 ) | ( n3760 & n9471 ) | ( n9450 & n9471 ) ;
  assign n9473 = n3482 &  n9472 ;
  assign n9474 = n3211 | n9473 ;
  assign n9475 = n9470 | n9474 ;
  assign n9476 = ( n9019 & ~n9286 ) | ( n9019 & n9023 ) | ( ~n9286 & n9023 ) ;
  assign n9477 = ( n9010 & ~n9476 ) | ( n9010 & n9019 ) | ( ~n9476 & n9019 ) ;
  assign n9478 = ( n9010 & ~n9019 ) | ( n9010 & n9476 ) | ( ~n9019 & n9476 ) ;
  assign n9479 = ( n9477 & ~n9010 ) | ( n9477 & n9478 ) | ( ~n9010 & n9478 ) ;
  assign n9480 = ( n9475 & ~n9479 ) | ( n9475 & 1'b0 ) | ( ~n9479 & 1'b0 ) ;
  assign n9481 = n9467 | n9480 ;
  assign n9482 = ~n9025 & n9286 ;
  assign n9483 = ( n9012 & n9017 ) | ( n9012 & n9286 ) | ( n9017 & n9286 ) ;
  assign n9485 = ( n9482 & ~n9012 ) | ( n9482 & n9483 ) | ( ~n9012 & n9483 ) ;
  assign n9484 = ( n9286 & ~n9483 ) | ( n9286 & n9482 ) | ( ~n9483 & n9482 ) ;
  assign n9486 = ( n9017 & ~n9485 ) | ( n9017 & n9484 ) | ( ~n9485 & n9484 ) ;
  assign n9487 = ( n2955 & n9481 ) | ( n2955 & n9486 ) | ( n9481 & n9486 ) ;
  assign n9488 = n2706 &  n9487 ;
  assign n9490 = ( n9041 & ~n9032 ) | ( n9041 & n9045 ) | ( ~n9032 & n9045 ) ;
  assign n9489 = n9045 | n9286 ;
  assign n9492 = ( n9045 & ~n9490 ) | ( n9045 & n9489 ) | ( ~n9490 & n9489 ) ;
  assign n9491 = ( n9489 & ~n9041 ) | ( n9489 & n9490 ) | ( ~n9041 & n9490 ) ;
  assign n9493 = ( n9032 & ~n9492 ) | ( n9032 & n9491 ) | ( ~n9492 & n9491 ) ;
  assign n9494 = n2955 | n9467 ;
  assign n9495 = n9480 | n9494 ;
  assign n9496 = n9486 &  n9495 ;
  assign n9497 = n9470 | n9473 ;
  assign n9498 = ( n3211 & ~n9479 ) | ( n3211 & n9497 ) | ( ~n9479 & n9497 ) ;
  assign n9499 = n2955 &  n9498 ;
  assign n9500 = n2706 | n9499 ;
  assign n9501 = n9496 | n9500 ;
  assign n9502 = ~n9493 & n9501 ;
  assign n9503 = n9488 | n9502 ;
  assign n9505 = ( n9034 & ~n9039 ) | ( n9034 & n9286 ) | ( ~n9039 & n9286 ) ;
  assign n9504 = ~n9047 & n9286 ;
  assign n9506 = ( n9286 & ~n9505 ) | ( n9286 & n9504 ) | ( ~n9505 & n9504 ) ;
  assign n9507 = ( n9504 & ~n9034 ) | ( n9504 & n9505 ) | ( ~n9034 & n9505 ) ;
  assign n9508 = ( n9039 & ~n9506 ) | ( n9039 & n9507 ) | ( ~n9506 & n9507 ) ;
  assign n9509 = ( n2472 & n9503 ) | ( n2472 & n9508 ) | ( n9503 & n9508 ) ;
  assign n9510 = n2245 &  n9509 ;
  assign n9511 = n9067 | n9286 ;
  assign n9512 = ( n9054 & n9063 ) | ( n9054 & n9067 ) | ( n9063 & n9067 ) ;
  assign n9513 = ( n9511 & ~n9063 ) | ( n9511 & n9512 ) | ( ~n9063 & n9512 ) ;
  assign n9514 = ( n9067 & ~n9512 ) | ( n9067 & n9511 ) | ( ~n9512 & n9511 ) ;
  assign n9515 = ( n9054 & ~n9513 ) | ( n9054 & n9514 ) | ( ~n9513 & n9514 ) ;
  assign n9516 = n2472 | n9488 ;
  assign n9517 = n9502 | n9516 ;
  assign n9518 = n9508 &  n9517 ;
  assign n9519 = n9496 | n9499 ;
  assign n9520 = ( n2706 & ~n9493 ) | ( n2706 & n9519 ) | ( ~n9493 & n9519 ) ;
  assign n9521 = n2472 &  n9520 ;
  assign n9522 = n2245 | n9521 ;
  assign n9523 = n9518 | n9522 ;
  assign n9524 = n9515 &  n9523 ;
  assign n9525 = n9510 | n9524 ;
  assign n9526 = ~n9069 & n9286 ;
  assign n9527 = ( n9056 & n9061 ) | ( n9056 & n9286 ) | ( n9061 & n9286 ) ;
  assign n9529 = ( n9526 & ~n9056 ) | ( n9526 & n9527 ) | ( ~n9056 & n9527 ) ;
  assign n9528 = ( n9286 & ~n9527 ) | ( n9286 & n9526 ) | ( ~n9527 & n9526 ) ;
  assign n9530 = ( n9061 & ~n9529 ) | ( n9061 & n9528 ) | ( ~n9529 & n9528 ) ;
  assign n9531 = ( n9525 & ~n2033 ) | ( n9525 & n9530 ) | ( ~n2033 & n9530 ) ;
  assign n9532 = n1827 &  n9531 ;
  assign n9533 = n9089 | n9286 ;
  assign n9534 = ( n9076 & ~n9085 ) | ( n9076 & n9089 ) | ( ~n9085 & n9089 ) ;
  assign n9535 = ( n9085 & n9533 ) | ( n9085 & n9534 ) | ( n9533 & n9534 ) ;
  assign n9536 = ( n9089 & ~n9534 ) | ( n9089 & n9533 ) | ( ~n9534 & n9533 ) ;
  assign n9537 = ( n9076 & ~n9535 ) | ( n9076 & n9536 ) | ( ~n9535 & n9536 ) ;
  assign n9538 = ( n2033 & ~n9510 ) | ( n2033 & 1'b0 ) | ( ~n9510 & 1'b0 ) ;
  assign n9539 = ~n9524 & n9538 ;
  assign n9540 = ( n9530 & ~n9539 ) | ( n9530 & 1'b0 ) | ( ~n9539 & 1'b0 ) ;
  assign n9541 = n9518 | n9521 ;
  assign n9542 = ( n2245 & n9515 ) | ( n2245 & n9541 ) | ( n9515 & n9541 ) ;
  assign n9543 = ~n2033 & n9542 ;
  assign n9544 = n1827 | n9543 ;
  assign n9545 = n9540 | n9544 ;
  assign n9546 = n9537 &  n9545 ;
  assign n9547 = n9532 | n9546 ;
  assign n9548 = ~n9091 & n9286 ;
  assign n9549 = ( n9078 & n9083 ) | ( n9078 & n9286 ) | ( n9083 & n9286 ) ;
  assign n9551 = ( n9548 & ~n9078 ) | ( n9548 & n9549 ) | ( ~n9078 & n9549 ) ;
  assign n9550 = ( n9286 & ~n9549 ) | ( n9286 & n9548 ) | ( ~n9549 & n9548 ) ;
  assign n9552 = ( n9083 & ~n9551 ) | ( n9083 & n9550 ) | ( ~n9551 & n9550 ) ;
  assign n9553 = ( n9547 & ~n1636 ) | ( n9547 & n9552 ) | ( ~n1636 & n9552 ) ;
  assign n9554 = ~n1452 & n9553 ;
  assign n9555 = n9111 | n9286 ;
  assign n9556 = ( n9098 & ~n9107 ) | ( n9098 & n9111 ) | ( ~n9107 & n9111 ) ;
  assign n9557 = ( n9107 & n9555 ) | ( n9107 & n9556 ) | ( n9555 & n9556 ) ;
  assign n9558 = ( n9111 & ~n9556 ) | ( n9111 & n9555 ) | ( ~n9556 & n9555 ) ;
  assign n9559 = ( n9098 & ~n9557 ) | ( n9098 & n9558 ) | ( ~n9557 & n9558 ) ;
  assign n9560 = ( n1636 & ~n9532 ) | ( n1636 & 1'b0 ) | ( ~n9532 & 1'b0 ) ;
  assign n9561 = ~n9546 & n9560 ;
  assign n9562 = ( n9552 & ~n9561 ) | ( n9552 & 1'b0 ) | ( ~n9561 & 1'b0 ) ;
  assign n9563 = n9540 | n9543 ;
  assign n9564 = ( n1827 & n9537 ) | ( n1827 & n9563 ) | ( n9537 & n9563 ) ;
  assign n9565 = ~n1636 & n9564 ;
  assign n9566 = ( n1452 & ~n9565 ) | ( n1452 & 1'b0 ) | ( ~n9565 & 1'b0 ) ;
  assign n9567 = ~n9562 & n9566 ;
  assign n9568 = ( n9559 & ~n9567 ) | ( n9559 & 1'b0 ) | ( ~n9567 & 1'b0 ) ;
  assign n9569 = n9554 | n9568 ;
  assign n9570 = n9113 &  n9286 ;
  assign n9571 = ( n9100 & n9105 ) | ( n9100 & n9286 ) | ( n9105 & n9286 ) ;
  assign n9573 = ( n9570 & ~n9100 ) | ( n9570 & n9571 ) | ( ~n9100 & n9571 ) ;
  assign n9572 = ( n9286 & ~n9571 ) | ( n9286 & n9570 ) | ( ~n9571 & n9570 ) ;
  assign n9574 = ( n9105 & ~n9573 ) | ( n9105 & n9572 ) | ( ~n9573 & n9572 ) ;
  assign n9575 = ( n1283 & n9569 ) | ( n1283 & n9574 ) | ( n9569 & n9574 ) ;
  assign n9576 = ~n1122 & n9575 ;
  assign n9578 = ( n9129 & ~n9120 ) | ( n9129 & n9133 ) | ( ~n9120 & n9133 ) ;
  assign n9577 = n9133 | n9286 ;
  assign n9580 = ( n9133 & ~n9578 ) | ( n9133 & n9577 ) | ( ~n9578 & n9577 ) ;
  assign n9579 = ( n9577 & ~n9129 ) | ( n9577 & n9578 ) | ( ~n9129 & n9578 ) ;
  assign n9581 = ( n9120 & ~n9580 ) | ( n9120 & n9579 ) | ( ~n9580 & n9579 ) ;
  assign n9582 = n1283 | n9554 ;
  assign n9583 = n9568 | n9582 ;
  assign n9584 = n9574 &  n9583 ;
  assign n9585 = n9562 | n9565 ;
  assign n9586 = ( n9559 & ~n1452 ) | ( n9559 & n9585 ) | ( ~n1452 & n9585 ) ;
  assign n9587 = n1283 &  n9586 ;
  assign n9588 = ( n1122 & ~n9587 ) | ( n1122 & 1'b0 ) | ( ~n9587 & 1'b0 ) ;
  assign n9589 = ~n9584 & n9588 ;
  assign n9590 = n9581 | n9589 ;
  assign n9591 = ~n9576 & n9590 ;
  assign n9593 = ( n9122 & ~n9127 ) | ( n9122 & n9286 ) | ( ~n9127 & n9286 ) ;
  assign n9592 = n9135 &  n9286 ;
  assign n9594 = ( n9286 & ~n9593 ) | ( n9286 & n9592 ) | ( ~n9593 & n9592 ) ;
  assign n9595 = ( n9592 & ~n9122 ) | ( n9592 & n9593 ) | ( ~n9122 & n9593 ) ;
  assign n9596 = ( n9127 & ~n9594 ) | ( n9127 & n9595 ) | ( ~n9594 & n9595 ) ;
  assign n9597 = ( n976 & n9591 ) | ( n976 & n9596 ) | ( n9591 & n9596 ) ;
  assign n9598 = ( n837 & ~n9597 ) | ( n837 & 1'b0 ) | ( ~n9597 & 1'b0 ) ;
  assign n9599 = ( n9155 & ~n9286 ) | ( n9155 & 1'b0 ) | ( ~n9286 & 1'b0 ) ;
  assign n9600 = ( n9142 & n9151 ) | ( n9142 & n9155 ) | ( n9151 & n9155 ) ;
  assign n9601 = ( n9599 & ~n9151 ) | ( n9599 & n9600 ) | ( ~n9151 & n9600 ) ;
  assign n9602 = ( n9155 & ~n9600 ) | ( n9155 & n9599 ) | ( ~n9600 & n9599 ) ;
  assign n9603 = ( n9142 & ~n9601 ) | ( n9142 & n9602 ) | ( ~n9601 & n9602 ) ;
  assign n9604 = ( n976 & ~n9576 ) | ( n976 & 1'b0 ) | ( ~n9576 & 1'b0 ) ;
  assign n9605 = n9590 &  n9604 ;
  assign n9606 = n9596 | n9605 ;
  assign n9607 = n9584 | n9587 ;
  assign n9608 = ( n1122 & ~n9607 ) | ( n1122 & n9581 ) | ( ~n9607 & n9581 ) ;
  assign n9609 = n976 | n9608 ;
  assign n9610 = ~n837 & n9609 ;
  assign n9611 = n9606 &  n9610 ;
  assign n9612 = n9603 | n9611 ;
  assign n9613 = ~n9598 & n9612 ;
  assign n9615 = ( n9144 & ~n9149 ) | ( n9144 & n9286 ) | ( ~n9149 & n9286 ) ;
  assign n9614 = n9157 &  n9286 ;
  assign n9616 = ( n9286 & ~n9615 ) | ( n9286 & n9614 ) | ( ~n9615 & n9614 ) ;
  assign n9617 = ( n9614 & ~n9144 ) | ( n9614 & n9615 ) | ( ~n9144 & n9615 ) ;
  assign n9618 = ( n9149 & ~n9616 ) | ( n9149 & n9617 ) | ( ~n9616 & n9617 ) ;
  assign n9619 = ( n9613 & ~n713 ) | ( n9613 & n9618 ) | ( ~n713 & n9618 ) ;
  assign n9620 = ( n595 & ~n9619 ) | ( n595 & 1'b0 ) | ( ~n9619 & 1'b0 ) ;
  assign n9621 = n9177 | n9286 ;
  assign n9622 = ( n9164 & ~n9173 ) | ( n9164 & n9177 ) | ( ~n9173 & n9177 ) ;
  assign n9623 = ( n9173 & n9621 ) | ( n9173 & n9622 ) | ( n9621 & n9622 ) ;
  assign n9624 = ( n9177 & ~n9622 ) | ( n9177 & n9621 ) | ( ~n9622 & n9621 ) ;
  assign n9625 = ( n9164 & ~n9623 ) | ( n9164 & n9624 ) | ( ~n9623 & n9624 ) ;
  assign n9626 = n713 | n9598 ;
  assign n9627 = ( n9612 & ~n9626 ) | ( n9612 & 1'b0 ) | ( ~n9626 & 1'b0 ) ;
  assign n9628 = n9618 | n9627 ;
  assign n9629 = n9606 &  n9609 ;
  assign n9630 = ( n9603 & ~n837 ) | ( n9603 & n9629 ) | ( ~n837 & n9629 ) ;
  assign n9631 = ( n713 & ~n9630 ) | ( n713 & 1'b0 ) | ( ~n9630 & 1'b0 ) ;
  assign n9632 = n595 | n9631 ;
  assign n9633 = ( n9628 & ~n9632 ) | ( n9628 & 1'b0 ) | ( ~n9632 & 1'b0 ) ;
  assign n9634 = ( n9625 & ~n9633 ) | ( n9625 & 1'b0 ) | ( ~n9633 & 1'b0 ) ;
  assign n9635 = n9620 | n9634 ;
  assign n9637 = ( n9166 & ~n9171 ) | ( n9166 & n9286 ) | ( ~n9171 & n9286 ) ;
  assign n9636 = ~n9179 & n9286 ;
  assign n9638 = ( n9286 & ~n9637 ) | ( n9286 & n9636 ) | ( ~n9637 & n9636 ) ;
  assign n9639 = ( n9636 & ~n9166 ) | ( n9636 & n9637 ) | ( ~n9166 & n9637 ) ;
  assign n9640 = ( n9171 & ~n9638 ) | ( n9171 & n9639 ) | ( ~n9638 & n9639 ) ;
  assign n9641 = ( n492 & n9635 ) | ( n492 & n9640 ) | ( n9635 & n9640 ) ;
  assign n9642 = n396 &  n9641 ;
  assign n9644 = ( n9195 & ~n9186 ) | ( n9195 & n9199 ) | ( ~n9186 & n9199 ) ;
  assign n9643 = n9199 | n9286 ;
  assign n9646 = ( n9199 & ~n9644 ) | ( n9199 & n9643 ) | ( ~n9644 & n9643 ) ;
  assign n9645 = ( n9643 & ~n9195 ) | ( n9643 & n9644 ) | ( ~n9195 & n9644 ) ;
  assign n9647 = ( n9186 & ~n9646 ) | ( n9186 & n9645 ) | ( ~n9646 & n9645 ) ;
  assign n9648 = n492 | n9620 ;
  assign n9649 = n9634 | n9648 ;
  assign n9650 = n9640 &  n9649 ;
  assign n9651 = ( n9628 & ~n9631 ) | ( n9628 & 1'b0 ) | ( ~n9631 & 1'b0 ) ;
  assign n9652 = ( n595 & ~n9651 ) | ( n595 & n9625 ) | ( ~n9651 & n9625 ) ;
  assign n9653 = n492 &  n9652 ;
  assign n9654 = n396 | n9653 ;
  assign n9655 = n9650 | n9654 ;
  assign n9656 = ~n9647 & n9655 ;
  assign n9657 = n9642 | n9656 ;
  assign n9658 = ~n9201 & n9286 ;
  assign n9659 = ( n9188 & ~n9658 ) | ( n9188 & n9286 ) | ( ~n9658 & n9286 ) ;
  assign n9660 = ( n9188 & ~n9659 ) | ( n9188 & n9193 ) | ( ~n9659 & n9193 ) ;
  assign n9661 = ( n9193 & ~n9188 ) | ( n9193 & n9659 ) | ( ~n9188 & n9659 ) ;
  assign n9662 = ( n9660 & ~n9193 ) | ( n9660 & n9661 ) | ( ~n9193 & n9661 ) ;
  assign n9663 = ( n315 & n9657 ) | ( n315 & n9662 ) | ( n9657 & n9662 ) ;
  assign n9664 = n240 &  n9663 ;
  assign n9665 = n9221 | n9286 ;
  assign n9666 = ( n9208 & n9217 ) | ( n9208 & n9221 ) | ( n9217 & n9221 ) ;
  assign n9667 = ( n9665 & ~n9217 ) | ( n9665 & n9666 ) | ( ~n9217 & n9666 ) ;
  assign n9668 = ( n9221 & ~n9666 ) | ( n9221 & n9665 ) | ( ~n9666 & n9665 ) ;
  assign n9669 = ( n9208 & ~n9667 ) | ( n9208 & n9668 ) | ( ~n9667 & n9668 ) ;
  assign n9670 = n315 | n9642 ;
  assign n9671 = n9656 | n9670 ;
  assign n9672 = n9662 &  n9671 ;
  assign n9673 = n9650 | n9653 ;
  assign n9674 = ( n396 & ~n9647 ) | ( n396 & n9673 ) | ( ~n9647 & n9673 ) ;
  assign n9675 = n315 &  n9674 ;
  assign n9676 = n240 | n9675 ;
  assign n9677 = n9672 | n9676 ;
  assign n9678 = n9669 &  n9677 ;
  assign n9679 = n9664 | n9678 ;
  assign n9685 = ( n181 & ~n9684 ) | ( n181 & n9679 ) | ( ~n9684 & n9679 ) ;
  assign n9686 = ~n145 & n9685 ;
  assign n9688 = ( n9239 & ~n9230 ) | ( n9239 & n9243 ) | ( ~n9230 & n9243 ) ;
  assign n9687 = n9243 | n9286 ;
  assign n9690 = ( n9243 & ~n9688 ) | ( n9243 & n9687 ) | ( ~n9688 & n9687 ) ;
  assign n9689 = ( n9687 & ~n9239 ) | ( n9687 & n9688 ) | ( ~n9239 & n9688 ) ;
  assign n9691 = ( n9230 & ~n9690 ) | ( n9230 & n9689 ) | ( ~n9690 & n9689 ) ;
  assign n9692 = n181 | n9664 ;
  assign n9693 = n9678 | n9692 ;
  assign n9694 = ~n9684 & n9693 ;
  assign n9695 = n9672 | n9675 ;
  assign n9696 = ( n240 & n9669 ) | ( n240 & n9695 ) | ( n9669 & n9695 ) ;
  assign n9697 = n181 &  n9696 ;
  assign n9698 = ( n145 & ~n9697 ) | ( n145 & 1'b0 ) | ( ~n9697 & 1'b0 ) ;
  assign n9699 = ~n9694 & n9698 ;
  assign n9700 = ( n9691 & ~n9699 ) | ( n9691 & 1'b0 ) | ( ~n9699 & 1'b0 ) ;
  assign n9701 = n9686 | n9700 ;
  assign n9702 = n9232 | n9286 ;
  assign n9703 = ( n9237 & ~n9232 ) | ( n9237 & n9245 ) | ( ~n9232 & n9245 ) ;
  assign n9705 = ( n9232 & n9702 ) | ( n9232 & n9703 ) | ( n9702 & n9703 ) ;
  assign n9704 = ( n9245 & ~n9703 ) | ( n9245 & n9702 ) | ( ~n9703 & n9702 ) ;
  assign n9706 = ( n9237 & ~n9705 ) | ( n9237 & n9704 ) | ( ~n9705 & n9704 ) ;
  assign n9707 = ( n150 & n9701 ) | ( n150 & n9706 ) | ( n9701 & n9706 ) ;
  assign n9708 = ( n9252 & ~n9271 ) | ( n9252 & 1'b0 ) | ( ~n9271 & 1'b0 ) ;
  assign n9709 = ( n9286 & ~n9268 ) | ( n9286 & n9708 ) | ( ~n9268 & n9708 ) ;
  assign n9710 = n9268 &  n9709 ;
  assign n9711 = ( n9268 & ~n9271 ) | ( n9268 & 1'b0 ) | ( ~n9271 & 1'b0 ) ;
  assign n9712 = ~n9286 & n9711 ;
  assign n9713 = ( n9252 & ~n9712 ) | ( n9252 & n9711 ) | ( ~n9712 & n9711 ) ;
  assign n9714 = ~n9710 & n9713 ;
  assign n9715 = n9253 &  n9260 ;
  assign n9716 = ~n9286 & n9715 ;
  assign n9717 = ( n9274 & ~n9715 ) | ( n9274 & n9716 ) | ( ~n9715 & n9716 ) ;
  assign n9718 = ~n9714 & n9717 ;
  assign n9719 = ~n9707 & n9718 ;
  assign n9720 = ( n133 & ~n9719 ) | ( n133 & n9718 ) | ( ~n9719 & n9718 ) ;
  assign n9723 = n9694 | n9697 ;
  assign n9724 = ( n9691 & ~n145 ) | ( n9691 & n9723 ) | ( ~n145 & n9723 ) ;
  assign n9725 = n150 &  n9724 ;
  assign n9726 = ( n9714 & ~n9725 ) | ( n9714 & 1'b0 ) | ( ~n9725 & 1'b0 ) ;
  assign n9721 = n150 | n9686 ;
  assign n9722 = n9700 | n9721 ;
  assign n9727 = ( n9706 & ~n9722 ) | ( n9706 & 1'b0 ) | ( ~n9722 & 1'b0 ) ;
  assign n9728 = ( n9726 & ~n9706 ) | ( n9726 & n9727 ) | ( ~n9706 & n9727 ) ;
  assign n9730 = ( n133 & n9253 ) | ( n133 & n9260 ) | ( n9253 & n9260 ) ;
  assign n9729 = ( n9253 & ~n9286 ) | ( n9253 & n9260 ) | ( ~n9286 & n9260 ) ;
  assign n9731 = ( n9260 & ~n9729 ) | ( n9260 & 1'b0 ) | ( ~n9729 & 1'b0 ) ;
  assign n9732 = ( n9730 & ~n9260 ) | ( n9730 & n9731 ) | ( ~n9260 & n9731 ) ;
  assign n9733 = n9256 | n9283 ;
  assign n9734 = ( n9278 & ~n9259 ) | ( n9278 & n9733 ) | ( ~n9259 & n9733 ) ;
  assign n9735 = n9259 | n9734 ;
  assign n9736 = ( n9266 & ~n9274 ) | ( n9266 & n9735 ) | ( ~n9274 & n9735 ) ;
  assign n9737 = ( n9266 & ~n9736 ) | ( n9266 & 1'b0 ) | ( ~n9736 & 1'b0 ) ;
  assign n9738 = n9732 | n9737 ;
  assign n9739 = n9728 | n9738 ;
  assign n9740 = ( n9720 & ~n9739 ) | ( n9720 & 1'b0 ) | ( ~n9739 & 1'b0 ) ;
  assign n9930 = n9458 | n9740 ;
  assign n9931 = ( n9445 & ~n9740 ) | ( n9445 & n9450 ) | ( ~n9740 & n9450 ) ;
  assign n9932 = ( n9740 & n9930 ) | ( n9740 & n9931 ) | ( n9930 & n9931 ) ;
  assign n9933 = ( n9445 & ~n9931 ) | ( n9445 & n9930 ) | ( ~n9931 & n9930 ) ;
  assign n9934 = ( n9450 & ~n9932 ) | ( n9450 & n9933 ) | ( ~n9932 & n9933 ) ;
  assign n9916 = ( n9452 & ~n9443 ) | ( n9452 & n9456 ) | ( ~n9443 & n9456 ) ;
  assign n9915 = ~n9456 & n9740 ;
  assign n9917 = ( n9452 & ~n9916 ) | ( n9452 & n9915 ) | ( ~n9916 & n9915 ) ;
  assign n9918 = ( n9915 & ~n9456 ) | ( n9915 & n9916 ) | ( ~n9456 & n9916 ) ;
  assign n9919 = ( n9443 & ~n9917 ) | ( n9443 & n9918 ) | ( ~n9917 & n9918 ) ;
  assign n9908 = n9436 | n9740 ;
  assign n9909 = ( n9428 & ~n9423 ) | ( n9428 & n9740 ) | ( ~n9423 & n9740 ) ;
  assign n9911 = ( n9423 & n9908 ) | ( n9423 & n9909 ) | ( n9908 & n9909 ) ;
  assign n9910 = ( n9740 & ~n9909 ) | ( n9740 & n9908 ) | ( ~n9909 & n9908 ) ;
  assign n9912 = ( n9428 & ~n9911 ) | ( n9428 & n9910 ) | ( ~n9911 & n9910 ) ;
  assign n9893 = ~n9434 & n9740 ;
  assign n9894 = ( n9421 & n9430 ) | ( n9421 & n9434 ) | ( n9430 & n9434 ) ;
  assign n9896 = ( n9893 & ~n9434 ) | ( n9893 & n9894 ) | ( ~n9434 & n9894 ) ;
  assign n9895 = ( n9430 & ~n9894 ) | ( n9430 & n9893 ) | ( ~n9894 & n9893 ) ;
  assign n9897 = ( n9421 & ~n9896 ) | ( n9421 & n9895 ) | ( ~n9896 & n9895 ) ;
  assign n9886 = n9414 | n9740 ;
  assign n9887 = ( n9401 & ~n9740 ) | ( n9401 & n9886 ) | ( ~n9740 & n9886 ) ;
  assign n9888 = ( n9406 & ~n9401 ) | ( n9406 & n9887 ) | ( ~n9401 & n9887 ) ;
  assign n9889 = ( n9401 & ~n9887 ) | ( n9401 & n9406 ) | ( ~n9887 & n9406 ) ;
  assign n9890 = ( n9888 & ~n9406 ) | ( n9888 & n9889 ) | ( ~n9406 & n9889 ) ;
  assign n9871 = ~n9412 & n9740 ;
  assign n9872 = ( n9399 & ~n9412 ) | ( n9399 & n9408 ) | ( ~n9412 & n9408 ) ;
  assign n9873 = ( n9871 & ~n9408 ) | ( n9871 & n9872 ) | ( ~n9408 & n9872 ) ;
  assign n9874 = ( n9412 & ~n9871 ) | ( n9412 & n9872 ) | ( ~n9871 & n9872 ) ;
  assign n9875 = ( n9873 & ~n9399 ) | ( n9873 & n9874 ) | ( ~n9399 & n9874 ) ;
  assign n9865 = ( n9379 & ~n9384 ) | ( n9379 & n9740 ) | ( ~n9384 & n9740 ) ;
  assign n9864 = ( n9392 & ~n9740 ) | ( n9392 & 1'b0 ) | ( ~n9740 & 1'b0 ) ;
  assign n9867 = ( n9379 & ~n9865 ) | ( n9379 & n9864 ) | ( ~n9865 & n9864 ) ;
  assign n9866 = ( n9864 & ~n9740 ) | ( n9864 & n9865 ) | ( ~n9740 & n9865 ) ;
  assign n9868 = ( n9384 & ~n9867 ) | ( n9384 & n9866 ) | ( ~n9867 & n9866 ) ;
  assign n9849 = ~n9390 & n9740 ;
  assign n9850 = ( n9377 & ~n9390 ) | ( n9377 & n9386 ) | ( ~n9390 & n9386 ) ;
  assign n9851 = ( n9849 & ~n9386 ) | ( n9849 & n9850 ) | ( ~n9386 & n9850 ) ;
  assign n9852 = ( n9390 & ~n9849 ) | ( n9390 & n9850 ) | ( ~n9849 & n9850 ) ;
  assign n9853 = ( n9851 & ~n9377 ) | ( n9851 & n9852 ) | ( ~n9377 & n9852 ) ;
  assign n9842 = ( n9370 & ~n9740 ) | ( n9370 & 1'b0 ) | ( ~n9740 & 1'b0 ) ;
  assign n9843 = ( n9357 & n9362 ) | ( n9357 & n9740 ) | ( n9362 & n9740 ) ;
  assign n9844 = ( n9842 & ~n9740 ) | ( n9842 & n9843 ) | ( ~n9740 & n9843 ) ;
  assign n9845 = ( n9357 & ~n9843 ) | ( n9357 & n9842 ) | ( ~n9843 & n9842 ) ;
  assign n9846 = ( n9362 & ~n9844 ) | ( n9362 & n9845 ) | ( ~n9844 & n9845 ) ;
  assign n9827 = ~n9368 & n9740 ;
  assign n9828 = ( n9355 & ~n9368 ) | ( n9355 & n9364 ) | ( ~n9368 & n9364 ) ;
  assign n9829 = ( n9827 & ~n9364 ) | ( n9827 & n9828 ) | ( ~n9364 & n9828 ) ;
  assign n9830 = ( n9368 & ~n9827 ) | ( n9368 & n9828 ) | ( ~n9827 & n9828 ) ;
  assign n9831 = ( n9829 & ~n9355 ) | ( n9829 & n9830 ) | ( ~n9355 & n9830 ) ;
  assign n9820 = ( n9348 & ~n9740 ) | ( n9348 & 1'b0 ) | ( ~n9740 & 1'b0 ) ;
  assign n9821 = ( n9335 & n9340 ) | ( n9335 & n9740 ) | ( n9340 & n9740 ) ;
  assign n9822 = ( n9820 & ~n9740 ) | ( n9820 & n9821 ) | ( ~n9740 & n9821 ) ;
  assign n9823 = ( n9335 & ~n9821 ) | ( n9335 & n9820 ) | ( ~n9821 & n9820 ) ;
  assign n9824 = ( n9340 & ~n9822 ) | ( n9340 & n9823 ) | ( ~n9822 & n9823 ) ;
  assign n9805 = n9346 &  n9740 ;
  assign n9806 = ( n9333 & n9342 ) | ( n9333 & n9346 ) | ( n9342 & n9346 ) ;
  assign n9807 = ( n9805 & ~n9342 ) | ( n9805 & n9806 ) | ( ~n9342 & n9806 ) ;
  assign n9808 = ( n9346 & ~n9806 ) | ( n9346 & n9805 ) | ( ~n9806 & n9805 ) ;
  assign n9809 = ( n9333 & ~n9807 ) | ( n9333 & n9808 ) | ( ~n9807 & n9808 ) ;
  assign n9798 = ~n9309 & n9740 ;
  assign n9799 = ( n9319 & ~n9309 ) | ( n9319 & n9326 ) | ( ~n9309 & n9326 ) ;
  assign n9800 = ( n9798 & ~n9326 ) | ( n9798 & n9799 ) | ( ~n9326 & n9799 ) ;
  assign n9801 = ( n9309 & ~n9798 ) | ( n9309 & n9799 ) | ( ~n9798 & n9799 ) ;
  assign n9802 = ( n9800 & ~n9319 ) | ( n9800 & n9801 ) | ( ~n9319 & n9801 ) ;
  assign n9783 = ~n9321 & n9324 ;
  assign n9784 = ( n9307 & ~n9321 ) | ( n9307 & n9783 ) | ( ~n9321 & n9783 ) ;
  assign n9785 = ( n9740 & ~n9783 ) | ( n9740 & n9784 ) | ( ~n9783 & n9784 ) ;
  assign n9786 = ( n9321 & ~n9740 ) | ( n9321 & n9784 ) | ( ~n9740 & n9784 ) ;
  assign n9787 = ( n9785 & ~n9307 ) | ( n9785 & n9786 ) | ( ~n9307 & n9786 ) ;
  assign n9771 = ( n9286 & ~x48 ) | ( n9286 & n9293 ) | ( ~x48 & n9293 ) ;
  assign n9772 = x48 &  n9771 ;
  assign n9773 = ( n9288 & ~n9772 ) | ( n9288 & n9293 ) | ( ~n9772 & n9293 ) ;
  assign n9774 = ~x48 & n9286 ;
  assign n9775 = ( x49 & ~n9774 ) | ( x49 & 1'b0 ) | ( ~n9774 & 1'b0 ) ;
  assign n9776 = n9298 | n9775 ;
  assign n9777 = ( n9740 & ~n9773 ) | ( n9740 & n9776 ) | ( ~n9773 & n9776 ) ;
  assign n9778 = n9773 | n9777 ;
  assign n9779 = ~n9740 & n9777 ;
  assign n9780 = ( n9778 & ~n9776 ) | ( n9778 & n9779 ) | ( ~n9776 & n9779 ) ;
  assign n9743 = x44 | x45 ;
  assign n9748 = ~x46 & n9743 ;
  assign n9749 = ( x46 & ~n9284 ) | ( x46 & n9748 ) | ( ~n9284 & n9748 ) ;
  assign n9750 = ( n9274 & ~n9266 ) | ( n9274 & n9749 ) | ( ~n9266 & n9749 ) ;
  assign n9751 = n9266 &  n9750 ;
  assign n9752 = ( x47 & ~n9751 ) | ( x47 & n9740 ) | ( ~n9751 & n9740 ) ;
  assign n9747 = ( x46 & x47 ) | ( x46 & n9740 ) | ( x47 & n9740 ) ;
  assign n9753 = ( x46 & ~x47 ) | ( x46 & 1'b0 ) | ( ~x47 & 1'b0 ) ;
  assign n9754 = ( n9752 & ~n9747 ) | ( n9752 & n9753 ) | ( ~n9747 & n9753 ) ;
  assign n9744 = x46 | n9743 ;
  assign n9745 = ( x46 & ~n9740 ) | ( x46 & 1'b0 ) | ( ~n9740 & 1'b0 ) ;
  assign n9746 = ( n9286 & ~n9744 ) | ( n9286 & n9745 ) | ( ~n9744 & n9745 ) ;
  assign n9757 = n8839 | n9746 ;
  assign n9758 = n9754 | n9757 ;
  assign n9759 = n8840 | n9740 ;
  assign n9760 = ( n9286 & ~n9737 ) | ( n9286 & 1'b0 ) | ( ~n9737 & 1'b0 ) ;
  assign n9761 = ( n9728 & ~n9732 ) | ( n9728 & n9760 ) | ( ~n9732 & n9760 ) ;
  assign n9762 = ~n9728 & n9761 ;
  assign n9763 = n9720 &  n9762 ;
  assign n9764 = n9759 | n9763 ;
  assign n9765 = ( x48 & ~n9764 ) | ( x48 & n9763 ) | ( ~n9764 & n9763 ) ;
  assign n9766 = x48 | n9763 ;
  assign n9767 = ( n9759 & ~n9766 ) | ( n9759 & 1'b0 ) | ( ~n9766 & 1'b0 ) ;
  assign n9768 = n9765 | n9767 ;
  assign n9769 = n9758 &  n9768 ;
  assign n9755 = ~n9754 & n9746 ;
  assign n9756 = ( n8839 & n9755 ) | ( n8839 & n9754 ) | ( n9755 & n9754 ) ;
  assign n9788 = n8407 | n9756 ;
  assign n9789 = n9769 | n9788 ;
  assign n9790 = n9780 &  n9789 ;
  assign n9791 = n9746 | n9754 ;
  assign n9792 = ( n8839 & n9768 ) | ( n8839 & n9791 ) | ( n9768 & n9791 ) ;
  assign n9793 = n8407 &  n9792 ;
  assign n9794 = n7982 | n9793 ;
  assign n9795 = n9790 | n9794 ;
  assign n9796 = n9787 &  n9795 ;
  assign n9770 = n9756 | n9769 ;
  assign n9781 = ( n8407 & n9770 ) | ( n8407 & n9780 ) | ( n9770 & n9780 ) ;
  assign n9782 = n7982 &  n9781 ;
  assign n9810 = ( n7572 & ~n9782 ) | ( n7572 & 1'b0 ) | ( ~n9782 & 1'b0 ) ;
  assign n9811 = ~n9796 & n9810 ;
  assign n9812 = ( n9802 & ~n9811 ) | ( n9802 & 1'b0 ) | ( ~n9811 & 1'b0 ) ;
  assign n9813 = n9790 | n9793 ;
  assign n9814 = ( n7982 & n9787 ) | ( n7982 & n9813 ) | ( n9787 & n9813 ) ;
  assign n9815 = ~n7572 & n9814 ;
  assign n9816 = ( n7169 & ~n9815 ) | ( n7169 & 1'b0 ) | ( ~n9815 & 1'b0 ) ;
  assign n9817 = ~n9812 & n9816 ;
  assign n9818 = n9809 | n9817 ;
  assign n9797 = n9782 | n9796 ;
  assign n9803 = ( n9797 & ~n7572 ) | ( n9797 & n9802 ) | ( ~n7572 & n9802 ) ;
  assign n9804 = ~n7169 & n9803 ;
  assign n9832 = n6781 | n9804 ;
  assign n9833 = ( n9818 & ~n9832 ) | ( n9818 & 1'b0 ) | ( ~n9832 & 1'b0 ) ;
  assign n9834 = n9824 | n9833 ;
  assign n9835 = n9812 | n9815 ;
  assign n9836 = ( n7169 & ~n9835 ) | ( n7169 & n9809 ) | ( ~n9835 & n9809 ) ;
  assign n9837 = ( n6781 & ~n9836 ) | ( n6781 & 1'b0 ) | ( ~n9836 & 1'b0 ) ;
  assign n9838 = ( n6399 & ~n9837 ) | ( n6399 & 1'b0 ) | ( ~n9837 & 1'b0 ) ;
  assign n9839 = n9834 &  n9838 ;
  assign n9840 = ( n9831 & ~n9839 ) | ( n9831 & 1'b0 ) | ( ~n9839 & 1'b0 ) ;
  assign n9819 = ~n9804 & n9818 ;
  assign n9825 = ( n9819 & ~n6781 ) | ( n9819 & n9824 ) | ( ~n6781 & n9824 ) ;
  assign n9826 = n6399 | n9825 ;
  assign n9854 = ~n6032 & n9826 ;
  assign n9855 = ~n9840 & n9854 ;
  assign n9856 = n9846 | n9855 ;
  assign n9857 = ( n9834 & ~n9837 ) | ( n9834 & 1'b0 ) | ( ~n9837 & 1'b0 ) ;
  assign n9858 = ( n6399 & ~n9831 ) | ( n6399 & n9857 ) | ( ~n9831 & n9857 ) ;
  assign n9859 = ( n6032 & ~n9858 ) | ( n6032 & 1'b0 ) | ( ~n9858 & 1'b0 ) ;
  assign n9860 = ( n5672 & ~n9859 ) | ( n5672 & 1'b0 ) | ( ~n9859 & 1'b0 ) ;
  assign n9861 = n9856 &  n9860 ;
  assign n9862 = ( n9853 & ~n9861 ) | ( n9853 & 1'b0 ) | ( ~n9861 & 1'b0 ) ;
  assign n9841 = ( n9826 & ~n9840 ) | ( n9826 & 1'b0 ) | ( ~n9840 & 1'b0 ) ;
  assign n9847 = ( n9841 & ~n6032 ) | ( n9841 & n9846 ) | ( ~n6032 & n9846 ) ;
  assign n9848 = n5672 | n9847 ;
  assign n9876 = ~n5327 & n9848 ;
  assign n9877 = ~n9862 & n9876 ;
  assign n9878 = ( n9868 & ~n9877 ) | ( n9868 & 1'b0 ) | ( ~n9877 & 1'b0 ) ;
  assign n9879 = ( n9856 & ~n9859 ) | ( n9856 & 1'b0 ) | ( ~n9859 & 1'b0 ) ;
  assign n9880 = ( n5672 & ~n9853 ) | ( n5672 & n9879 ) | ( ~n9853 & n9879 ) ;
  assign n9881 = ( n5327 & ~n9880 ) | ( n5327 & 1'b0 ) | ( ~n9880 & 1'b0 ) ;
  assign n9882 = n4990 | n9881 ;
  assign n9883 = n9878 | n9882 ;
  assign n9884 = ~n9875 & n9883 ;
  assign n9863 = ( n9848 & ~n9862 ) | ( n9848 & 1'b0 ) | ( ~n9862 & 1'b0 ) ;
  assign n9869 = ( n5327 & ~n9863 ) | ( n5327 & n9868 ) | ( ~n9863 & n9868 ) ;
  assign n9870 = n4990 &  n9869 ;
  assign n9898 = n4668 | n9870 ;
  assign n9899 = n9884 | n9898 ;
  assign n9900 = ~n9890 & n9899 ;
  assign n9901 = n9878 | n9881 ;
  assign n9902 = ( n4990 & ~n9875 ) | ( n4990 & n9901 ) | ( ~n9875 & n9901 ) ;
  assign n9903 = n4668 &  n9902 ;
  assign n9904 = n4353 | n9903 ;
  assign n9905 = n9900 | n9904 ;
  assign n9906 = ~n9897 & n9905 ;
  assign n9885 = n9870 | n9884 ;
  assign n9891 = ( n4668 & ~n9890 ) | ( n4668 & n9885 ) | ( ~n9890 & n9885 ) ;
  assign n9892 = n4353 &  n9891 ;
  assign n9920 = n4053 | n9892 ;
  assign n9921 = n9906 | n9920 ;
  assign n9922 = ~n9912 & n9921 ;
  assign n9923 = n9900 | n9903 ;
  assign n9924 = ( n4353 & ~n9897 ) | ( n4353 & n9923 ) | ( ~n9897 & n9923 ) ;
  assign n9925 = n4053 &  n9924 ;
  assign n9945 = n9922 | n9925 ;
  assign n9946 = ( n3760 & ~n9919 ) | ( n3760 & n9945 ) | ( ~n9919 & n9945 ) ;
  assign n9947 = n3482 &  n9946 ;
  assign n10127 = n9655 | n9740 ;
  assign n10128 = ( n9642 & ~n9740 ) | ( n9642 & n10127 ) | ( ~n9740 & n10127 ) ;
  assign n10129 = ( n9647 & ~n9642 ) | ( n9647 & n10128 ) | ( ~n9642 & n10128 ) ;
  assign n10130 = ( n9642 & ~n10128 ) | ( n9642 & n9647 ) | ( ~n10128 & n9647 ) ;
  assign n10131 = ( n10129 & ~n9647 ) | ( n10129 & n10130 ) | ( ~n9647 & n10130 ) ;
  assign n10105 = ( n9633 & ~n9740 ) | ( n9633 & 1'b0 ) | ( ~n9740 & 1'b0 ) ;
  assign n10106 = ( n9625 & ~n9620 ) | ( n9625 & n9740 ) | ( ~n9620 & n9740 ) ;
  assign n10107 = ( n10105 & ~n9740 ) | ( n10105 & n10106 ) | ( ~n9740 & n10106 ) ;
  assign n10108 = ( n9620 & ~n10105 ) | ( n9620 & n10106 ) | ( ~n10105 & n10106 ) ;
  assign n10109 = ( n10107 & ~n9625 ) | ( n10107 & n10108 ) | ( ~n9625 & n10108 ) ;
  assign n10061 = ( n9589 & ~n9740 ) | ( n9589 & 1'b0 ) | ( ~n9740 & 1'b0 ) ;
  assign n10062 = ( n9576 & ~n9740 ) | ( n9576 & n9581 ) | ( ~n9740 & n9581 ) ;
  assign n10063 = ( n9740 & ~n10061 ) | ( n9740 & n10062 ) | ( ~n10061 & n10062 ) ;
  assign n10064 = ( n10061 & ~n9576 ) | ( n10061 & n10062 ) | ( ~n9576 & n10062 ) ;
  assign n10065 = ( n10063 & ~n9581 ) | ( n10063 & n10064 ) | ( ~n9581 & n10064 ) ;
  assign n9973 = n9501 | n9740 ;
  assign n9974 = ( n9493 & ~n9488 ) | ( n9493 & n9740 ) | ( ~n9488 & n9740 ) ;
  assign n9976 = ( n9973 & n9488 ) | ( n9973 & n9974 ) | ( n9488 & n9974 ) ;
  assign n9975 = ( n9740 & ~n9974 ) | ( n9740 & n9973 ) | ( ~n9974 & n9973 ) ;
  assign n9977 = ( n9493 & ~n9976 ) | ( n9493 & n9975 ) | ( ~n9976 & n9975 ) ;
  assign n9952 = ( n9467 & n9475 ) | ( n9467 & n9479 ) | ( n9475 & n9479 ) ;
  assign n9954 = ( n9740 & ~n9467 ) | ( n9740 & n9952 ) | ( ~n9467 & n9952 ) ;
  assign n9953 = ( n9475 & ~n9952 ) | ( n9475 & n9740 ) | ( ~n9952 & n9740 ) ;
  assign n9955 = ( n9479 & ~n9954 ) | ( n9479 & n9953 ) | ( ~n9954 & n9953 ) ;
  assign n9907 = n9892 | n9906 ;
  assign n9913 = ( n4053 & ~n9912 ) | ( n4053 & n9907 ) | ( ~n9912 & n9907 ) ;
  assign n9914 = n3760 &  n9913 ;
  assign n9926 = n3760 | n9925 ;
  assign n9927 = n9922 | n9926 ;
  assign n9928 = ~n9919 & n9927 ;
  assign n9929 = n9914 | n9928 ;
  assign n9935 = ( n3482 & n9929 ) | ( n3482 & n9934 ) | ( n9929 & n9934 ) ;
  assign n9936 = n3211 &  n9935 ;
  assign n9938 = ( n9469 & ~n9465 ) | ( n9469 & n9473 ) | ( ~n9465 & n9473 ) ;
  assign n9937 = ~n9473 & n9740 ;
  assign n9939 = ( n9469 & ~n9938 ) | ( n9469 & n9937 ) | ( ~n9938 & n9937 ) ;
  assign n9940 = ( n9937 & ~n9473 ) | ( n9937 & n9938 ) | ( ~n9473 & n9938 ) ;
  assign n9941 = ( n9465 & ~n9939 ) | ( n9465 & n9940 ) | ( ~n9939 & n9940 ) ;
  assign n9942 = n3482 | n9914 ;
  assign n9943 = n9928 | n9942 ;
  assign n9944 = n9934 &  n9943 ;
  assign n9948 = n3211 | n9947 ;
  assign n9949 = n9944 | n9948 ;
  assign n9950 = ~n9941 & n9949 ;
  assign n9951 = n9936 | n9950 ;
  assign n9956 = ( n2955 & ~n9955 ) | ( n2955 & n9951 ) | ( ~n9955 & n9951 ) ;
  assign n9957 = n2706 &  n9956 ;
  assign n9958 = ~n9499 & n9740 ;
  assign n9959 = ( n9486 & n9495 ) | ( n9486 & n9499 ) | ( n9495 & n9499 ) ;
  assign n9961 = ( n9958 & ~n9499 ) | ( n9958 & n9959 ) | ( ~n9499 & n9959 ) ;
  assign n9960 = ( n9495 & ~n9959 ) | ( n9495 & n9958 ) | ( ~n9959 & n9958 ) ;
  assign n9962 = ( n9486 & ~n9961 ) | ( n9486 & n9960 ) | ( ~n9961 & n9960 ) ;
  assign n9963 = n2955 | n9936 ;
  assign n9964 = n9950 | n9963 ;
  assign n9965 = ~n9955 & n9964 ;
  assign n9966 = n9944 | n9947 ;
  assign n9967 = ( n3211 & ~n9941 ) | ( n3211 & n9966 ) | ( ~n9941 & n9966 ) ;
  assign n9968 = n2955 &  n9967 ;
  assign n9969 = n2706 | n9968 ;
  assign n9970 = n9965 | n9969 ;
  assign n9971 = n9962 &  n9970 ;
  assign n9972 = n9957 | n9971 ;
  assign n9978 = ( n2472 & ~n9977 ) | ( n2472 & n9972 ) | ( ~n9977 & n9972 ) ;
  assign n9979 = n2245 &  n9978 ;
  assign n9980 = ~n9521 & n9740 ;
  assign n9981 = ( n9508 & n9517 ) | ( n9508 & n9521 ) | ( n9517 & n9521 ) ;
  assign n9983 = ( n9980 & ~n9521 ) | ( n9980 & n9981 ) | ( ~n9521 & n9981 ) ;
  assign n9982 = ( n9517 & ~n9981 ) | ( n9517 & n9980 ) | ( ~n9981 & n9980 ) ;
  assign n9984 = ( n9508 & ~n9983 ) | ( n9508 & n9982 ) | ( ~n9983 & n9982 ) ;
  assign n9985 = n2472 | n9957 ;
  assign n9986 = n9971 | n9985 ;
  assign n9987 = ~n9977 & n9986 ;
  assign n9988 = n9965 | n9968 ;
  assign n9989 = ( n2706 & n9962 ) | ( n2706 & n9988 ) | ( n9962 & n9988 ) ;
  assign n9990 = n2472 &  n9989 ;
  assign n9991 = n2245 | n9990 ;
  assign n9992 = n9987 | n9991 ;
  assign n9993 = n9984 &  n9992 ;
  assign n9994 = n9979 | n9993 ;
  assign n9995 = n9523 | n9740 ;
  assign n9996 = ( n9510 & ~n9740 ) | ( n9510 & n9515 ) | ( ~n9740 & n9515 ) ;
  assign n9997 = ( n9740 & n9995 ) | ( n9740 & n9996 ) | ( n9995 & n9996 ) ;
  assign n9998 = ( n9510 & ~n9996 ) | ( n9510 & n9995 ) | ( ~n9996 & n9995 ) ;
  assign n9999 = ( n9515 & ~n9997 ) | ( n9515 & n9998 ) | ( ~n9997 & n9998 ) ;
  assign n10000 = ( n9994 & ~n2033 ) | ( n9994 & n9999 ) | ( ~n2033 & n9999 ) ;
  assign n10001 = n1827 &  n10000 ;
  assign n10002 = ~n9543 & n9740 ;
  assign n10003 = ( n9530 & ~n9539 ) | ( n9530 & n9543 ) | ( ~n9539 & n9543 ) ;
  assign n10004 = ( n9539 & ~n10002 ) | ( n9539 & n10003 ) | ( ~n10002 & n10003 ) ;
  assign n10005 = ( n10002 & ~n9543 ) | ( n10002 & n10003 ) | ( ~n9543 & n10003 ) ;
  assign n10006 = ( n10004 & ~n9530 ) | ( n10004 & n10005 ) | ( ~n9530 & n10005 ) ;
  assign n10007 = ( n2033 & ~n9979 ) | ( n2033 & 1'b0 ) | ( ~n9979 & 1'b0 ) ;
  assign n10008 = ~n9993 & n10007 ;
  assign n10009 = ( n9999 & ~n10008 ) | ( n9999 & 1'b0 ) | ( ~n10008 & 1'b0 ) ;
  assign n10010 = n9987 | n9990 ;
  assign n10011 = ( n2245 & n9984 ) | ( n2245 & n10010 ) | ( n9984 & n10010 ) ;
  assign n10012 = ~n2033 & n10011 ;
  assign n10013 = n1827 | n10012 ;
  assign n10014 = n10009 | n10013 ;
  assign n10015 = ~n10006 & n10014 ;
  assign n10016 = n10001 | n10015 ;
  assign n10017 = n9545 | n9740 ;
  assign n10018 = ( n9532 & ~n9740 ) | ( n9532 & n10017 ) | ( ~n9740 & n10017 ) ;
  assign n10019 = ( n9532 & ~n10018 ) | ( n9532 & n9537 ) | ( ~n10018 & n9537 ) ;
  assign n10020 = ( n9537 & ~n9532 ) | ( n9537 & n10018 ) | ( ~n9532 & n10018 ) ;
  assign n10021 = ( n10019 & ~n9537 ) | ( n10019 & n10020 ) | ( ~n9537 & n10020 ) ;
  assign n10022 = ( n10016 & ~n1636 ) | ( n10016 & n10021 ) | ( ~n1636 & n10021 ) ;
  assign n10023 = ~n1452 & n10022 ;
  assign n10024 = ~n9565 & n9740 ;
  assign n10025 = ( n9552 & ~n9561 ) | ( n9552 & n9565 ) | ( ~n9561 & n9565 ) ;
  assign n10026 = ( n9561 & ~n10024 ) | ( n9561 & n10025 ) | ( ~n10024 & n10025 ) ;
  assign n10027 = ( n10024 & ~n9565 ) | ( n10024 & n10025 ) | ( ~n9565 & n10025 ) ;
  assign n10028 = ( n10026 & ~n9552 ) | ( n10026 & n10027 ) | ( ~n9552 & n10027 ) ;
  assign n10029 = ( n1636 & ~n10001 ) | ( n1636 & 1'b0 ) | ( ~n10001 & 1'b0 ) ;
  assign n10030 = ~n10015 & n10029 ;
  assign n10031 = ( n10021 & ~n10030 ) | ( n10021 & 1'b0 ) | ( ~n10030 & 1'b0 ) ;
  assign n10032 = n10009 | n10012 ;
  assign n10033 = ( n1827 & ~n10006 ) | ( n1827 & n10032 ) | ( ~n10006 & n10032 ) ;
  assign n10034 = ~n1636 & n10033 ;
  assign n10035 = ( n1452 & ~n10034 ) | ( n1452 & 1'b0 ) | ( ~n10034 & 1'b0 ) ;
  assign n10036 = ~n10031 & n10035 ;
  assign n10037 = n10028 | n10036 ;
  assign n10038 = ~n10023 & n10037 ;
  assign n10039 = ( n9567 & ~n9740 ) | ( n9567 & 1'b0 ) | ( ~n9740 & 1'b0 ) ;
  assign n10040 = ( n9559 & ~n9554 ) | ( n9559 & n9740 ) | ( ~n9554 & n9740 ) ;
  assign n10041 = ( n10039 & ~n9740 ) | ( n10039 & n10040 ) | ( ~n9740 & n10040 ) ;
  assign n10042 = ( n9554 & ~n10039 ) | ( n9554 & n10040 ) | ( ~n10039 & n10040 ) ;
  assign n10043 = ( n10041 & ~n9559 ) | ( n10041 & n10042 ) | ( ~n9559 & n10042 ) ;
  assign n10044 = ( n10038 & ~n1283 ) | ( n10038 & n10043 ) | ( ~n1283 & n10043 ) ;
  assign n10045 = n1122 | n10044 ;
  assign n10046 = ~n9587 & n9740 ;
  assign n10047 = ( n9574 & n9583 ) | ( n9574 & n9587 ) | ( n9583 & n9587 ) ;
  assign n10049 = ( n10046 & ~n9587 ) | ( n10046 & n10047 ) | ( ~n9587 & n10047 ) ;
  assign n10048 = ( n9583 & ~n10047 ) | ( n9583 & n10046 ) | ( ~n10047 & n10046 ) ;
  assign n10050 = ( n9574 & ~n10049 ) | ( n9574 & n10048 ) | ( ~n10049 & n10048 ) ;
  assign n10051 = n1283 | n10023 ;
  assign n10052 = ( n10037 & ~n10051 ) | ( n10037 & 1'b0 ) | ( ~n10051 & 1'b0 ) ;
  assign n10053 = n10043 | n10052 ;
  assign n10054 = n10031 | n10034 ;
  assign n10055 = ( n1452 & ~n10054 ) | ( n1452 & n10028 ) | ( ~n10054 & n10028 ) ;
  assign n10056 = ( n1283 & ~n10055 ) | ( n1283 & 1'b0 ) | ( ~n10055 & 1'b0 ) ;
  assign n10057 = ( n1122 & ~n10056 ) | ( n1122 & 1'b0 ) | ( ~n10056 & 1'b0 ) ;
  assign n10058 = n10053 &  n10057 ;
  assign n10059 = ( n10050 & ~n10058 ) | ( n10050 & 1'b0 ) | ( ~n10058 & 1'b0 ) ;
  assign n10060 = ( n10045 & ~n10059 ) | ( n10045 & 1'b0 ) | ( ~n10059 & 1'b0 ) ;
  assign n10066 = ( n976 & ~n10065 ) | ( n976 & n10060 ) | ( ~n10065 & n10060 ) ;
  assign n10067 = ( n837 & ~n10066 ) | ( n837 & 1'b0 ) | ( ~n10066 & 1'b0 ) ;
  assign n10068 = n9609 &  n9740 ;
  assign n10069 = ( n9596 & n9605 ) | ( n9596 & n9609 ) | ( n9605 & n9609 ) ;
  assign n10070 = ( n10068 & ~n9605 ) | ( n10068 & n10069 ) | ( ~n9605 & n10069 ) ;
  assign n10071 = ( n9609 & ~n10069 ) | ( n9609 & n10068 ) | ( ~n10069 & n10068 ) ;
  assign n10072 = ( n9596 & ~n10070 ) | ( n9596 & n10071 ) | ( ~n10070 & n10071 ) ;
  assign n10073 = n976 &  n10045 ;
  assign n10074 = ~n10059 & n10073 ;
  assign n10075 = ( n10065 & ~n10074 ) | ( n10065 & 1'b0 ) | ( ~n10074 & 1'b0 ) ;
  assign n10076 = ( n10053 & ~n10056 ) | ( n10053 & 1'b0 ) | ( ~n10056 & 1'b0 ) ;
  assign n10077 = ( n1122 & ~n10050 ) | ( n1122 & n10076 ) | ( ~n10050 & n10076 ) ;
  assign n10078 = n976 | n10077 ;
  assign n10079 = ~n837 & n10078 ;
  assign n10080 = ~n10075 & n10079 ;
  assign n10081 = n10072 | n10080 ;
  assign n10082 = ~n10067 & n10081 ;
  assign n10084 = ( n9603 & ~n9598 ) | ( n9603 & n9740 ) | ( ~n9598 & n9740 ) ;
  assign n10083 = ( n9611 & ~n9740 ) | ( n9611 & 1'b0 ) | ( ~n9740 & 1'b0 ) ;
  assign n10085 = ( n10084 & ~n9740 ) | ( n10084 & n10083 ) | ( ~n9740 & n10083 ) ;
  assign n10086 = ( n9598 & ~n10083 ) | ( n9598 & n10084 ) | ( ~n10083 & n10084 ) ;
  assign n10087 = ( n10085 & ~n9603 ) | ( n10085 & n10086 ) | ( ~n9603 & n10086 ) ;
  assign n10088 = ( n713 & ~n10082 ) | ( n713 & n10087 ) | ( ~n10082 & n10087 ) ;
  assign n10089 = n595 &  n10088 ;
  assign n10090 = ~n9631 & n9740 ;
  assign n10091 = ( n9618 & ~n9631 ) | ( n9618 & n9627 ) | ( ~n9631 & n9627 ) ;
  assign n10092 = ( n10090 & ~n9627 ) | ( n10090 & n10091 ) | ( ~n9627 & n10091 ) ;
  assign n10093 = ( n9631 & ~n10090 ) | ( n9631 & n10091 ) | ( ~n10090 & n10091 ) ;
  assign n10094 = ( n10092 & ~n9618 ) | ( n10092 & n10093 ) | ( ~n9618 & n10093 ) ;
  assign n10095 = n713 | n10067 ;
  assign n10096 = ( n10081 & ~n10095 ) | ( n10081 & 1'b0 ) | ( ~n10095 & 1'b0 ) ;
  assign n10097 = ( n10087 & ~n10096 ) | ( n10087 & 1'b0 ) | ( ~n10096 & 1'b0 ) ;
  assign n10098 = ~n10075 & n10078 ;
  assign n10099 = ( n10072 & ~n837 ) | ( n10072 & n10098 ) | ( ~n837 & n10098 ) ;
  assign n10100 = ( n713 & ~n10099 ) | ( n713 & 1'b0 ) | ( ~n10099 & 1'b0 ) ;
  assign n10101 = n595 | n10100 ;
  assign n10102 = n10097 | n10101 ;
  assign n10103 = n10094 &  n10102 ;
  assign n10104 = n10089 | n10103 ;
  assign n10110 = ( n492 & ~n10109 ) | ( n492 & n10104 ) | ( ~n10109 & n10104 ) ;
  assign n10111 = n396 &  n10110 ;
  assign n10112 = ~n9653 & n9740 ;
  assign n10113 = ( n9640 & n9649 ) | ( n9640 & n9653 ) | ( n9649 & n9653 ) ;
  assign n10115 = ( n10112 & ~n9653 ) | ( n10112 & n10113 ) | ( ~n9653 & n10113 ) ;
  assign n10114 = ( n9649 & ~n10113 ) | ( n9649 & n10112 ) | ( ~n10113 & n10112 ) ;
  assign n10116 = ( n9640 & ~n10115 ) | ( n9640 & n10114 ) | ( ~n10115 & n10114 ) ;
  assign n10117 = n492 | n10089 ;
  assign n10118 = n10103 | n10117 ;
  assign n10119 = ~n10109 & n10118 ;
  assign n10120 = n10097 | n10100 ;
  assign n10121 = ( n595 & n10094 ) | ( n595 & n10120 ) | ( n10094 & n10120 ) ;
  assign n10122 = n492 &  n10121 ;
  assign n10123 = n396 | n10122 ;
  assign n10124 = n10119 | n10123 ;
  assign n10125 = n10116 &  n10124 ;
  assign n10126 = n10111 | n10125 ;
  assign n10132 = ( n315 & ~n10131 ) | ( n315 & n10126 ) | ( ~n10131 & n10126 ) ;
  assign n10133 = n240 &  n10132 ;
  assign n10134 = ~n9675 & n9740 ;
  assign n10135 = ( n9662 & n9671 ) | ( n9662 & n9675 ) | ( n9671 & n9675 ) ;
  assign n10137 = ( n10134 & ~n9675 ) | ( n10134 & n10135 ) | ( ~n9675 & n10135 ) ;
  assign n10136 = ( n9671 & ~n10135 ) | ( n9671 & n10134 ) | ( ~n10135 & n10134 ) ;
  assign n10138 = ( n9662 & ~n10137 ) | ( n9662 & n10136 ) | ( ~n10137 & n10136 ) ;
  assign n10139 = n315 | n10111 ;
  assign n10140 = n10125 | n10139 ;
  assign n10141 = ~n10131 & n10140 ;
  assign n10142 = n10119 | n10122 ;
  assign n10143 = ( n396 & n10116 ) | ( n396 & n10142 ) | ( n10116 & n10142 ) ;
  assign n10144 = n315 &  n10143 ;
  assign n10145 = n240 | n10144 ;
  assign n10146 = n10141 | n10145 ;
  assign n10147 = n10138 &  n10146 ;
  assign n10148 = n10133 | n10147 ;
  assign n10149 = n9677 | n9740 ;
  assign n10150 = ( n9669 & ~n9664 ) | ( n9669 & n9740 ) | ( ~n9664 & n9740 ) ;
  assign n10152 = ( n9664 & n10149 ) | ( n9664 & n10150 ) | ( n10149 & n10150 ) ;
  assign n10151 = ( n9740 & ~n10150 ) | ( n9740 & n10149 ) | ( ~n10150 & n10149 ) ;
  assign n10153 = ( n9669 & ~n10152 ) | ( n9669 & n10151 ) | ( ~n10152 & n10151 ) ;
  assign n10154 = ( n181 & n10148 ) | ( n181 & n10153 ) | ( n10148 & n10153 ) ;
  assign n10155 = ~n145 & n10154 ;
  assign n10156 = ~n9697 & n9740 ;
  assign n10157 = ( n9684 & n9693 ) | ( n9684 & n9697 ) | ( n9693 & n9697 ) ;
  assign n10159 = ( n10156 & ~n9697 ) | ( n10156 & n10157 ) | ( ~n9697 & n10157 ) ;
  assign n10158 = ( n9693 & ~n10157 ) | ( n9693 & n10156 ) | ( ~n10157 & n10156 ) ;
  assign n10160 = ( n9684 & ~n10159 ) | ( n9684 & n10158 ) | ( ~n10159 & n10158 ) ;
  assign n10161 = n181 | n10133 ;
  assign n10162 = n10147 | n10161 ;
  assign n10163 = n10153 &  n10162 ;
  assign n10164 = n10141 | n10144 ;
  assign n10165 = ( n240 & n10138 ) | ( n240 & n10164 ) | ( n10138 & n10164 ) ;
  assign n10166 = n181 &  n10165 ;
  assign n10167 = ( n145 & ~n10166 ) | ( n145 & 1'b0 ) | ( ~n10166 & 1'b0 ) ;
  assign n10168 = ~n10163 & n10167 ;
  assign n10169 = n10160 | n10168 ;
  assign n10170 = ~n10155 & n10169 ;
  assign n10171 = ~n9686 & n9740 ;
  assign n10172 = ( n9691 & ~n9686 ) | ( n9691 & n9699 ) | ( ~n9686 & n9699 ) ;
  assign n10173 = ( n10171 & ~n9699 ) | ( n10171 & n10172 ) | ( ~n9699 & n10172 ) ;
  assign n10174 = ( n9686 & ~n10171 ) | ( n9686 & n10172 ) | ( ~n10171 & n10172 ) ;
  assign n10175 = ( n10173 & ~n9691 ) | ( n10173 & n10174 ) | ( ~n9691 & n10174 ) ;
  assign n10176 = ( n10170 & ~n150 ) | ( n10170 & n10175 ) | ( ~n150 & n10175 ) ;
  assign n10177 = ~n9706 & n9722 ;
  assign n10178 = ( n9725 & ~n9740 ) | ( n9725 & n10177 ) | ( ~n9740 & n10177 ) ;
  assign n10179 = ~n9725 & n10178 ;
  assign n10180 = ( n9722 & ~n9725 ) | ( n9722 & 1'b0 ) | ( ~n9725 & 1'b0 ) ;
  assign n10181 = n9740 &  n10180 ;
  assign n10182 = ( n9706 & ~n10180 ) | ( n9706 & n10181 ) | ( ~n10180 & n10181 ) ;
  assign n10183 = n10179 | n10182 ;
  assign n10184 = ( n9707 & ~n9714 ) | ( n9707 & 1'b0 ) | ( ~n9714 & 1'b0 ) ;
  assign n10185 = n9740 &  n10184 ;
  assign n10186 = ( n9728 & ~n10185 ) | ( n9728 & n10184 ) | ( ~n10185 & n10184 ) ;
  assign n10187 = ( n10183 & ~n10186 ) | ( n10183 & 1'b0 ) | ( ~n10186 & 1'b0 ) ;
  assign n10188 = n10176 &  n10187 ;
  assign n10189 = ( n133 & ~n10188 ) | ( n133 & n10187 ) | ( ~n10188 & n10187 ) ;
  assign n10192 = n10163 | n10166 ;
  assign n10193 = ( n145 & ~n10192 ) | ( n145 & n10160 ) | ( ~n10192 & n10160 ) ;
  assign n10194 = ( n150 & ~n10193 ) | ( n150 & 1'b0 ) | ( ~n10193 & 1'b0 ) ;
  assign n10195 = n10183 | n10194 ;
  assign n10190 = n150 | n10155 ;
  assign n10191 = ( n10169 & ~n10190 ) | ( n10169 & 1'b0 ) | ( ~n10190 & 1'b0 ) ;
  assign n10196 = ~n10175 & n10191 ;
  assign n10197 = ( n10175 & ~n10195 ) | ( n10175 & n10196 ) | ( ~n10195 & n10196 ) ;
  assign n10198 = ( n9707 & ~n9714 ) | ( n9707 & n9740 ) | ( ~n9714 & n9740 ) ;
  assign n10200 = n9714 | n10198 ;
  assign n10199 = ( n133 & ~n9714 ) | ( n133 & n9707 ) | ( ~n9714 & n9707 ) ;
  assign n10201 = ( n9714 & ~n10200 ) | ( n9714 & n10199 ) | ( ~n10200 & n10199 ) ;
  assign n10202 = n9710 | n9737 ;
  assign n10203 = ( n9713 & n9732 ) | ( n9713 & n10202 ) | ( n9732 & n10202 ) ;
  assign n10204 = ( n9713 & ~n10203 ) | ( n9713 & 1'b0 ) | ( ~n10203 & 1'b0 ) ;
  assign n10205 = ( n9720 & ~n10204 ) | ( n9720 & n9728 ) | ( ~n10204 & n9728 ) ;
  assign n10206 = ( n9720 & ~n10205 ) | ( n9720 & 1'b0 ) | ( ~n10205 & 1'b0 ) ;
  assign n10207 = n10201 | n10206 ;
  assign n10208 = n10197 | n10207 ;
  assign n10209 = ~n10189 |  n10208 ;
  assign n10413 = n9947 | n10209 ;
  assign n10414 = ( n9934 & n9943 ) | ( n9934 & n9947 ) | ( n9943 & n9947 ) ;
  assign n10415 = ( n10413 & ~n9943 ) | ( n10413 & n10414 ) | ( ~n9943 & n10414 ) ;
  assign n10416 = ( n9947 & ~n10414 ) | ( n9947 & n10413 ) | ( ~n10414 & n10413 ) ;
  assign n10417 = ( n9934 & ~n10415 ) | ( n9934 & n10416 ) | ( ~n10415 & n10416 ) ;
  assign n10407 = ( n9914 & ~n9919 ) | ( n9914 & n10209 ) | ( ~n9919 & n10209 ) ;
  assign n10406 = ~n9927 & n10209 ;
  assign n10408 = ( n10209 & ~n10407 ) | ( n10209 & n10406 ) | ( ~n10407 & n10406 ) ;
  assign n10409 = ( n10406 & ~n9914 ) | ( n10406 & n10407 ) | ( ~n9914 & n10407 ) ;
  assign n10410 = ( n9919 & ~n10408 ) | ( n9919 & n10409 ) | ( ~n10408 & n10409 ) ;
  assign n10392 = ( n9921 & ~n9912 ) | ( n9921 & n9925 ) | ( ~n9912 & n9925 ) ;
  assign n10391 = n9925 | n10209 ;
  assign n10394 = ( n9925 & ~n10392 ) | ( n9925 & n10391 ) | ( ~n10392 & n10391 ) ;
  assign n10393 = ( n10391 & ~n9921 ) | ( n10391 & n10392 ) | ( ~n9921 & n10392 ) ;
  assign n10395 = ( n9912 & ~n10394 ) | ( n9912 & n10393 ) | ( ~n10394 & n10393 ) ;
  assign n10384 = ~n9905 & n10209 ;
  assign n10385 = ( n9892 & n9897 ) | ( n9892 & n10209 ) | ( n9897 & n10209 ) ;
  assign n10387 = ( n10384 & ~n9892 ) | ( n10384 & n10385 ) | ( ~n9892 & n10385 ) ;
  assign n10386 = ( n10209 & ~n10385 ) | ( n10209 & n10384 ) | ( ~n10385 & n10384 ) ;
  assign n10388 = ( n9897 & ~n10387 ) | ( n9897 & n10386 ) | ( ~n10387 & n10386 ) ;
  assign n10370 = ( n9899 & ~n9890 ) | ( n9899 & n9903 ) | ( ~n9890 & n9903 ) ;
  assign n10369 = n9903 | n10209 ;
  assign n10372 = ( n9903 & ~n10370 ) | ( n9903 & n10369 ) | ( ~n10370 & n10369 ) ;
  assign n10371 = ( n10369 & ~n9899 ) | ( n10369 & n10370 ) | ( ~n9899 & n10370 ) ;
  assign n10373 = ( n9890 & ~n10372 ) | ( n9890 & n10371 ) | ( ~n10372 & n10371 ) ;
  assign n10362 = ~n9883 & n10209 ;
  assign n10363 = ( n9870 & ~n10362 ) | ( n9870 & n10209 ) | ( ~n10362 & n10209 ) ;
  assign n10364 = ( n9875 & ~n9870 ) | ( n9875 & n10363 ) | ( ~n9870 & n10363 ) ;
  assign n10365 = ( n9870 & ~n10363 ) | ( n9870 & n9875 ) | ( ~n10363 & n9875 ) ;
  assign n10366 = ( n10364 & ~n9875 ) | ( n10364 & n10365 ) | ( ~n9875 & n10365 ) ;
  assign n10347 = n9881 | n10209 ;
  assign n10348 = ( n9868 & ~n9877 ) | ( n9868 & n9881 ) | ( ~n9877 & n9881 ) ;
  assign n10349 = ( n9877 & n10347 ) | ( n9877 & n10348 ) | ( n10347 & n10348 ) ;
  assign n10350 = ( n9881 & ~n10348 ) | ( n9881 & n10347 ) | ( ~n10348 & n10347 ) ;
  assign n10351 = ( n9868 & ~n10349 ) | ( n9868 & n10350 ) | ( ~n10349 & n10350 ) ;
  assign n10340 = n9861 &  n10209 ;
  assign n10341 = ( n9848 & ~n10209 ) | ( n9848 & n10340 ) | ( ~n10209 & n10340 ) ;
  assign n10342 = ( n9853 & ~n9848 ) | ( n9853 & n10341 ) | ( ~n9848 & n10341 ) ;
  assign n10343 = ( n9848 & ~n10341 ) | ( n9848 & n9853 ) | ( ~n10341 & n9853 ) ;
  assign n10344 = ( n10342 & ~n9853 ) | ( n10342 & n10343 ) | ( ~n9853 & n10343 ) ;
  assign n10325 = n9859 | n10209 ;
  assign n10326 = ( n9846 & ~n9859 ) | ( n9846 & n9855 ) | ( ~n9859 & n9855 ) ;
  assign n10328 = ( n9859 & n10325 ) | ( n9859 & n10326 ) | ( n10325 & n10326 ) ;
  assign n10327 = ( n9855 & ~n10326 ) | ( n9855 & n10325 ) | ( ~n10326 & n10325 ) ;
  assign n10329 = ( n9846 & ~n10328 ) | ( n9846 & n10327 ) | ( ~n10328 & n10327 ) ;
  assign n10318 = n9839 &  n10209 ;
  assign n10319 = ( n9826 & ~n10209 ) | ( n9826 & n10318 ) | ( ~n10209 & n10318 ) ;
  assign n10320 = ( n9831 & ~n9826 ) | ( n9831 & n10319 ) | ( ~n9826 & n10319 ) ;
  assign n10321 = ( n9826 & ~n10319 ) | ( n9826 & n9831 ) | ( ~n10319 & n9831 ) ;
  assign n10322 = ( n10320 & ~n9831 ) | ( n10320 & n10321 ) | ( ~n9831 & n10321 ) ;
  assign n10303 = n9837 | n10209 ;
  assign n10304 = ( n9824 & ~n9837 ) | ( n9824 & n9833 ) | ( ~n9837 & n9833 ) ;
  assign n10306 = ( n9837 & n10303 ) | ( n9837 & n10304 ) | ( n10303 & n10304 ) ;
  assign n10305 = ( n9833 & ~n10304 ) | ( n9833 & n10303 ) | ( ~n10304 & n10303 ) ;
  assign n10307 = ( n9824 & ~n10306 ) | ( n9824 & n10305 ) | ( ~n10306 & n10305 ) ;
  assign n10296 = n9804 | n10209 ;
  assign n10297 = ( n9809 & ~n9804 ) | ( n9809 & n9817 ) | ( ~n9804 & n9817 ) ;
  assign n10299 = ( n9804 & n10296 ) | ( n9804 & n10297 ) | ( n10296 & n10297 ) ;
  assign n10298 = ( n9817 & ~n10297 ) | ( n9817 & n10296 ) | ( ~n10297 & n10296 ) ;
  assign n10300 = ( n9809 & ~n10299 ) | ( n9809 & n10298 ) | ( ~n10299 & n10298 ) ;
  assign n10281 = n9815 | n10209 ;
  assign n10282 = ( n9802 & ~n9815 ) | ( n9802 & n9811 ) | ( ~n9815 & n9811 ) ;
  assign n10284 = ( n9815 & n10281 ) | ( n9815 & n10282 ) | ( n10281 & n10282 ) ;
  assign n10283 = ( n9811 & ~n10282 ) | ( n9811 & n10281 ) | ( ~n10282 & n10281 ) ;
  assign n10285 = ( n9802 & ~n10284 ) | ( n9802 & n10283 ) | ( ~n10284 & n10283 ) ;
  assign n10274 = n9782 | n10209 ;
  assign n10275 = ( n9782 & n9787 ) | ( n9782 & n9795 ) | ( n9787 & n9795 ) ;
  assign n10276 = ( n10274 & ~n9795 ) | ( n10274 & n10275 ) | ( ~n9795 & n10275 ) ;
  assign n10277 = ( n9782 & ~n10275 ) | ( n9782 & n10274 ) | ( ~n10275 & n10274 ) ;
  assign n10278 = ( n9787 & ~n10276 ) | ( n9787 & n10277 ) | ( ~n10276 & n10277 ) ;
  assign n10260 = ( n9789 & ~n9780 ) | ( n9789 & n9793 ) | ( ~n9780 & n9793 ) ;
  assign n10259 = n9793 | n10209 ;
  assign n10262 = ( n9793 & ~n10260 ) | ( n9793 & n10259 ) | ( ~n10260 & n10259 ) ;
  assign n10261 = ( n10259 & ~n9789 ) | ( n10259 & n10260 ) | ( ~n9789 & n10260 ) ;
  assign n10263 = ( n9780 & ~n10262 ) | ( n9780 & n10261 ) | ( ~n10262 & n10261 ) ;
  assign n10252 = n9756 &  n9758 ;
  assign n10253 = ( n9758 & n9768 ) | ( n9758 & n10252 ) | ( n9768 & n10252 ) ;
  assign n10254 = ( n10209 & ~n9758 ) | ( n10209 & n10253 ) | ( ~n9758 & n10253 ) ;
  assign n10255 = ( n10209 & ~n10253 ) | ( n10209 & n10252 ) | ( ~n10253 & n10252 ) ;
  assign n10256 = ( n9768 & ~n10254 ) | ( n9768 & n10255 ) | ( ~n10254 & n10255 ) ;
  assign n10236 = x46 | n9740 ;
  assign n10237 = x47 &  n10236 ;
  assign n10238 = ( n9759 & ~n10237 ) | ( n9759 & 1'b0 ) | ( ~n10237 & 1'b0 ) ;
  assign n10233 = ( x46 & ~n9751 ) | ( x46 & n9740 ) | ( ~n9751 & n9740 ) ;
  assign n10234 = ( x46 & ~n10233 ) | ( x46 & 1'b0 ) | ( ~n10233 & 1'b0 ) ;
  assign n10235 = ( n9746 & ~n10234 ) | ( n9746 & n9751 ) | ( ~n10234 & n9751 ) ;
  assign n10239 = ( n10209 & n10235 ) | ( n10209 & n10238 ) | ( n10235 & n10238 ) ;
  assign n10240 = ~n10235 & n10239 ;
  assign n10241 = ( n10209 & ~n10239 ) | ( n10209 & 1'b0 ) | ( ~n10239 & 1'b0 ) ;
  assign n10242 = ( n10238 & ~n10240 ) | ( n10238 & n10241 ) | ( ~n10240 & n10241 ) ;
  assign n10222 = n9740 | n10206 ;
  assign n10223 = ( n10201 & ~n10197 ) | ( n10201 & n10222 ) | ( ~n10197 & n10222 ) ;
  assign n10224 = n10197 | n10223 ;
  assign n10225 = ( n10189 & ~n10224 ) | ( n10189 & 1'b0 ) | ( ~n10224 & 1'b0 ) ;
  assign n10221 = ~n9743 & n10209 ;
  assign n10226 = ( n10221 & ~n10225 ) | ( n10221 & 1'b0 ) | ( ~n10225 & 1'b0 ) ;
  assign n10227 = ( x46 & n10225 ) | ( x46 & n10226 ) | ( n10225 & n10226 ) ;
  assign n10228 = x46 | n10225 ;
  assign n10229 = n10221 | n10228 ;
  assign n10230 = ~n10227 & n10229 ;
  assign n10212 = ( x44 & ~n10209 ) | ( x44 & x45 ) | ( ~n10209 & x45 ) ;
  assign n10218 = ( x44 & ~x45 ) | ( x44 & 1'b0 ) | ( ~x45 & 1'b0 ) ;
  assign n9741 = x42 | x43 ;
  assign n10213 = ~x44 & n9741 ;
  assign n10214 = ( x44 & ~n9738 ) | ( x44 & n10213 ) | ( ~n9738 & n10213 ) ;
  assign n10215 = ( n9720 & ~n10214 ) | ( n9720 & n9728 ) | ( ~n10214 & n9728 ) ;
  assign n10216 = ( n9720 & ~n10215 ) | ( n9720 & 1'b0 ) | ( ~n10215 & 1'b0 ) ;
  assign n10217 = ( n10209 & ~x45 ) | ( n10209 & n10216 ) | ( ~x45 & n10216 ) ;
  assign n10219 = ( n10212 & ~n10218 ) | ( n10212 & n10217 ) | ( ~n10218 & n10217 ) ;
  assign n10210 = x44 &  n10209 ;
  assign n9742 = x44 | n9741 ;
  assign n10211 = ( n9740 & ~n10210 ) | ( n9740 & n9742 ) | ( ~n10210 & n9742 ) ;
  assign n10243 = ~n9286 & n10211 ;
  assign n10244 = n10219 &  n10243 ;
  assign n10245 = n10230 | n10244 ;
  assign n10246 = ~n10211 & n10219 ;
  assign n10247 = ( n9286 & ~n10219 ) | ( n9286 & n10246 ) | ( ~n10219 & n10246 ) ;
  assign n10248 = n8839 | n10247 ;
  assign n10249 = ( n10245 & ~n10248 ) | ( n10245 & 1'b0 ) | ( ~n10248 & 1'b0 ) ;
  assign n10250 = ( n10242 & ~n10249 ) | ( n10242 & 1'b0 ) | ( ~n10249 & 1'b0 ) ;
  assign n10220 = n10211 &  n10219 ;
  assign n10231 = ( n10220 & ~n9286 ) | ( n10220 & n10230 ) | ( ~n9286 & n10230 ) ;
  assign n10232 = ( n8839 & ~n10231 ) | ( n8839 & 1'b0 ) | ( ~n10231 & 1'b0 ) ;
  assign n10264 = n8407 | n10232 ;
  assign n10265 = n10250 | n10264 ;
  assign n10266 = n10256 &  n10265 ;
  assign n10267 = ( n10245 & ~n10247 ) | ( n10245 & 1'b0 ) | ( ~n10247 & 1'b0 ) ;
  assign n10268 = ( n8839 & ~n10267 ) | ( n8839 & n10242 ) | ( ~n10267 & n10242 ) ;
  assign n10269 = n8407 &  n10268 ;
  assign n10270 = n7982 | n10269 ;
  assign n10271 = n10266 | n10270 ;
  assign n10272 = n10263 &  n10271 ;
  assign n10251 = n10232 | n10250 ;
  assign n10257 = ( n8407 & n10251 ) | ( n8407 & n10256 ) | ( n10251 & n10256 ) ;
  assign n10258 = n7982 &  n10257 ;
  assign n10286 = ( n7572 & ~n10258 ) | ( n7572 & 1'b0 ) | ( ~n10258 & 1'b0 ) ;
  assign n10287 = ~n10272 & n10286 ;
  assign n10288 = ( n10278 & ~n10287 ) | ( n10278 & 1'b0 ) | ( ~n10287 & 1'b0 ) ;
  assign n10289 = n10266 | n10269 ;
  assign n10290 = ( n7982 & n10263 ) | ( n7982 & n10289 ) | ( n10263 & n10289 ) ;
  assign n10291 = ~n7572 & n10290 ;
  assign n10292 = ( n7169 & ~n10291 ) | ( n7169 & 1'b0 ) | ( ~n10291 & 1'b0 ) ;
  assign n10293 = ~n10288 & n10292 ;
  assign n10294 = ( n10285 & ~n10293 ) | ( n10285 & 1'b0 ) | ( ~n10293 & 1'b0 ) ;
  assign n10273 = n10258 | n10272 ;
  assign n10279 = ( n10273 & ~n7572 ) | ( n10273 & n10278 ) | ( ~n7572 & n10278 ) ;
  assign n10280 = ~n7169 & n10279 ;
  assign n10308 = n6781 | n10280 ;
  assign n10309 = n10294 | n10308 ;
  assign n10310 = ~n10300 & n10309 ;
  assign n10311 = n10288 | n10291 ;
  assign n10312 = ( n10285 & ~n7169 ) | ( n10285 & n10311 ) | ( ~n7169 & n10311 ) ;
  assign n10313 = n6781 &  n10312 ;
  assign n10314 = ( n6399 & ~n10313 ) | ( n6399 & 1'b0 ) | ( ~n10313 & 1'b0 ) ;
  assign n10315 = ~n10310 & n10314 ;
  assign n10316 = n10307 | n10315 ;
  assign n10295 = n10280 | n10294 ;
  assign n10301 = ( n6781 & ~n10300 ) | ( n6781 & n10295 ) | ( ~n10300 & n10295 ) ;
  assign n10302 = ~n6399 & n10301 ;
  assign n10330 = n6032 | n10302 ;
  assign n10331 = ( n10316 & ~n10330 ) | ( n10316 & 1'b0 ) | ( ~n10330 & 1'b0 ) ;
  assign n10332 = ( n10322 & ~n10331 ) | ( n10322 & 1'b0 ) | ( ~n10331 & 1'b0 ) ;
  assign n10333 = n10310 | n10313 ;
  assign n10334 = ( n6399 & ~n10333 ) | ( n6399 & n10307 ) | ( ~n10333 & n10307 ) ;
  assign n10335 = ( n6032 & ~n10334 ) | ( n6032 & 1'b0 ) | ( ~n10334 & 1'b0 ) ;
  assign n10336 = ( n5672 & ~n10335 ) | ( n5672 & 1'b0 ) | ( ~n10335 & 1'b0 ) ;
  assign n10337 = ~n10332 & n10336 ;
  assign n10338 = n10329 | n10337 ;
  assign n10317 = ~n10302 & n10316 ;
  assign n10323 = ( n6032 & ~n10317 ) | ( n6032 & n10322 ) | ( ~n10317 & n10322 ) ;
  assign n10324 = ~n5672 & n10323 ;
  assign n10352 = n5327 | n10324 ;
  assign n10353 = ( n10338 & ~n10352 ) | ( n10338 & 1'b0 ) | ( ~n10352 & 1'b0 ) ;
  assign n10354 = ( n10344 & ~n10353 ) | ( n10344 & 1'b0 ) | ( ~n10353 & 1'b0 ) ;
  assign n10355 = n10332 | n10335 ;
  assign n10356 = ( n5672 & ~n10355 ) | ( n5672 & n10329 ) | ( ~n10355 & n10329 ) ;
  assign n10357 = ( n5327 & ~n10356 ) | ( n5327 & 1'b0 ) | ( ~n10356 & 1'b0 ) ;
  assign n10358 = n4990 | n10357 ;
  assign n10359 = n10354 | n10358 ;
  assign n10360 = n10351 &  n10359 ;
  assign n10339 = ~n10324 & n10338 ;
  assign n10345 = ( n5327 & ~n10339 ) | ( n5327 & n10344 ) | ( ~n10339 & n10344 ) ;
  assign n10346 = n4990 &  n10345 ;
  assign n10374 = n4668 | n10346 ;
  assign n10375 = n10360 | n10374 ;
  assign n10376 = ~n10366 & n10375 ;
  assign n10377 = n10354 | n10357 ;
  assign n10378 = ( n4990 & n10351 ) | ( n4990 & n10377 ) | ( n10351 & n10377 ) ;
  assign n10379 = n4668 &  n10378 ;
  assign n10380 = n4353 | n10379 ;
  assign n10381 = n10376 | n10380 ;
  assign n10382 = ~n10373 & n10381 ;
  assign n10361 = n10346 | n10360 ;
  assign n10367 = ( n4668 & ~n10366 ) | ( n4668 & n10361 ) | ( ~n10366 & n10361 ) ;
  assign n10368 = n4353 &  n10367 ;
  assign n10396 = n4053 | n10368 ;
  assign n10397 = n10382 | n10396 ;
  assign n10398 = ~n10388 & n10397 ;
  assign n10399 = n10376 | n10379 ;
  assign n10400 = ( n4353 & ~n10373 ) | ( n4353 & n10399 ) | ( ~n10373 & n10399 ) ;
  assign n10401 = n4053 &  n10400 ;
  assign n10402 = n3760 | n10401 ;
  assign n10403 = n10398 | n10402 ;
  assign n10404 = ~n10395 & n10403 ;
  assign n10383 = n10368 | n10382 ;
  assign n10389 = ( n4053 & ~n10388 ) | ( n4053 & n10383 ) | ( ~n10388 & n10383 ) ;
  assign n10390 = n3760 &  n10389 ;
  assign n10418 = n3482 | n10390 ;
  assign n10419 = n10404 | n10418 ;
  assign n10420 = ~n10410 & n10419 ;
  assign n10421 = n10398 | n10401 ;
  assign n10422 = ( n3760 & ~n10395 ) | ( n3760 & n10421 ) | ( ~n10395 & n10421 ) ;
  assign n10423 = n3482 &  n10422 ;
  assign n10424 = n3211 | n10423 ;
  assign n10425 = n10420 | n10424 ;
  assign n10653 = ( n10175 & ~n10194 ) | ( n10175 & 1'b0 ) | ( ~n10194 & 1'b0 ) ;
  assign n10654 = ( n10191 & n10209 ) | ( n10191 & n10653 ) | ( n10209 & n10653 ) ;
  assign n10655 = ~n10191 & n10654 ;
  assign n10656 = n10191 | n10194 ;
  assign n10657 = n10209 | n10656 ;
  assign n10658 = ( n10175 & ~n10656 ) | ( n10175 & n10657 ) | ( ~n10656 & n10657 ) ;
  assign n10659 = ~n10655 & n10658 ;
  assign n10660 = ~n10176 & n10183 ;
  assign n10661 = ~n10209 & n10660 ;
  assign n10662 = ( n10197 & ~n10661 ) | ( n10197 & n10660 ) | ( ~n10661 & n10660 ) ;
  assign n10663 = n10659 | n10662 ;
  assign n10647 = n10155 | n10209 ;
  assign n10648 = ( n10155 & ~n10168 ) | ( n10155 & n10160 ) | ( ~n10168 & n10160 ) ;
  assign n10649 = ( n10168 & n10647 ) | ( n10168 & n10648 ) | ( n10647 & n10648 ) ;
  assign n10650 = ( n10155 & ~n10648 ) | ( n10155 & n10647 ) | ( ~n10648 & n10647 ) ;
  assign n10651 = ( n10160 & ~n10649 ) | ( n10160 & n10650 ) | ( ~n10649 & n10650 ) ;
  assign n10560 = ( n10067 & ~n10072 ) | ( n10067 & n10209 ) | ( ~n10072 & n10209 ) ;
  assign n10559 = n10080 &  n10209 ;
  assign n10561 = ( n10209 & ~n10560 ) | ( n10209 & n10559 ) | ( ~n10560 & n10559 ) ;
  assign n10562 = ( n10559 & ~n10067 ) | ( n10559 & n10560 ) | ( ~n10067 & n10560 ) ;
  assign n10563 = ( n10072 & ~n10561 ) | ( n10072 & n10562 ) | ( ~n10561 & n10562 ) ;
  assign n10537 = n10058 &  n10209 ;
  assign n10538 = ( n10045 & ~n10209 ) | ( n10045 & n10537 ) | ( ~n10209 & n10537 ) ;
  assign n10539 = ( n10050 & ~n10045 ) | ( n10050 & n10538 ) | ( ~n10045 & n10538 ) ;
  assign n10540 = ( n10045 & ~n10538 ) | ( n10045 & n10050 ) | ( ~n10538 & n10050 ) ;
  assign n10541 = ( n10539 & ~n10050 ) | ( n10539 & n10540 ) | ( ~n10050 & n10540 ) ;
  assign n10429 = ( n9936 & ~n9941 ) | ( n9936 & n10209 ) | ( ~n9941 & n10209 ) ;
  assign n10428 = ~n9949 & n10209 ;
  assign n10430 = ( n10209 & ~n10429 ) | ( n10209 & n10428 ) | ( ~n10429 & n10428 ) ;
  assign n10431 = ( n10428 & ~n9936 ) | ( n10428 & n10429 ) | ( ~n9936 & n10429 ) ;
  assign n10432 = ( n9941 & ~n10430 ) | ( n9941 & n10431 ) | ( ~n10430 & n10431 ) ;
  assign n10405 = n10390 | n10404 ;
  assign n10411 = ( n3482 & ~n10410 ) | ( n3482 & n10405 ) | ( ~n10410 & n10405 ) ;
  assign n10412 = n3211 &  n10411 ;
  assign n10426 = n10417 &  n10425 ;
  assign n10427 = n10412 | n10426 ;
  assign n10433 = ( n2955 & ~n10432 ) | ( n2955 & n10427 ) | ( ~n10432 & n10427 ) ;
  assign n10434 = n2706 &  n10433 ;
  assign n10435 = n2955 | n10412 ;
  assign n10436 = n10426 | n10435 ;
  assign n10437 = ~n10432 & n10436 ;
  assign n10438 = n10420 | n10423 ;
  assign n10439 = ( n3211 & n10417 ) | ( n3211 & n10438 ) | ( n10417 & n10438 ) ;
  assign n10440 = n2955 &  n10439 ;
  assign n10441 = n2706 | n10440 ;
  assign n10442 = n10437 | n10441 ;
  assign n10443 = ( n9955 & n9964 ) | ( n9955 & n9968 ) | ( n9964 & n9968 ) ;
  assign n10444 = ( n10209 & ~n9964 ) | ( n10209 & n10443 ) | ( ~n9964 & n10443 ) ;
  assign n10445 = ( n9968 & ~n10443 ) | ( n9968 & n10209 ) | ( ~n10443 & n10209 ) ;
  assign n10446 = ( n9955 & ~n10444 ) | ( n9955 & n10445 ) | ( ~n10444 & n10445 ) ;
  assign n10447 = ( n10442 & ~n10446 ) | ( n10442 & 1'b0 ) | ( ~n10446 & 1'b0 ) ;
  assign n10448 = n10434 | n10447 ;
  assign n10450 = ( n9957 & ~n9962 ) | ( n9957 & n10209 ) | ( ~n9962 & n10209 ) ;
  assign n10449 = ~n9970 & n10209 ;
  assign n10451 = ( n10209 & ~n10450 ) | ( n10209 & n10449 ) | ( ~n10450 & n10449 ) ;
  assign n10452 = ( n10449 & ~n9957 ) | ( n10449 & n10450 ) | ( ~n9957 & n10450 ) ;
  assign n10453 = ( n9962 & ~n10451 ) | ( n9962 & n10452 ) | ( ~n10451 & n10452 ) ;
  assign n10454 = ( n2472 & n10448 ) | ( n2472 & n10453 ) | ( n10448 & n10453 ) ;
  assign n10455 = n2245 &  n10454 ;
  assign n10457 = ( n9986 & ~n9977 ) | ( n9986 & n9990 ) | ( ~n9977 & n9990 ) ;
  assign n10456 = n9990 | n10209 ;
  assign n10459 = ( n9990 & ~n10457 ) | ( n9990 & n10456 ) | ( ~n10457 & n10456 ) ;
  assign n10458 = ( n10456 & ~n9986 ) | ( n10456 & n10457 ) | ( ~n9986 & n10457 ) ;
  assign n10460 = ( n9977 & ~n10459 ) | ( n9977 & n10458 ) | ( ~n10459 & n10458 ) ;
  assign n10461 = n2472 | n10434 ;
  assign n10462 = n10447 | n10461 ;
  assign n10463 = n10453 &  n10462 ;
  assign n10464 = n10437 | n10440 ;
  assign n10465 = ( n2706 & ~n10446 ) | ( n2706 & n10464 ) | ( ~n10446 & n10464 ) ;
  assign n10466 = n2472 &  n10465 ;
  assign n10467 = n2245 | n10466 ;
  assign n10468 = n10463 | n10467 ;
  assign n10469 = ~n10460 & n10468 ;
  assign n10470 = n10455 | n10469 ;
  assign n10471 = ~n9992 & n10209 ;
  assign n10472 = ( n9979 & ~n10471 ) | ( n9979 & n10209 ) | ( ~n10471 & n10209 ) ;
  assign n10473 = ( n9979 & ~n10472 ) | ( n9979 & n9984 ) | ( ~n10472 & n9984 ) ;
  assign n10474 = ( n9984 & ~n9979 ) | ( n9984 & n10472 ) | ( ~n9979 & n10472 ) ;
  assign n10475 = ( n10473 & ~n9984 ) | ( n10473 & n10474 ) | ( ~n9984 & n10474 ) ;
  assign n10476 = ( n10470 & ~n2033 ) | ( n10470 & n10475 ) | ( ~n2033 & n10475 ) ;
  assign n10477 = n1827 &  n10476 ;
  assign n10478 = n10012 | n10209 ;
  assign n10479 = ( n9999 & ~n10008 ) | ( n9999 & n10012 ) | ( ~n10008 & n10012 ) ;
  assign n10480 = ( n10008 & n10478 ) | ( n10008 & n10479 ) | ( n10478 & n10479 ) ;
  assign n10481 = ( n10012 & ~n10479 ) | ( n10012 & n10478 ) | ( ~n10479 & n10478 ) ;
  assign n10482 = ( n9999 & ~n10480 ) | ( n9999 & n10481 ) | ( ~n10480 & n10481 ) ;
  assign n10483 = ( n2033 & ~n10455 ) | ( n2033 & 1'b0 ) | ( ~n10455 & 1'b0 ) ;
  assign n10484 = ~n10469 & n10483 ;
  assign n10485 = ( n10475 & ~n10484 ) | ( n10475 & 1'b0 ) | ( ~n10484 & 1'b0 ) ;
  assign n10486 = n10463 | n10466 ;
  assign n10487 = ( n2245 & ~n10460 ) | ( n2245 & n10486 ) | ( ~n10460 & n10486 ) ;
  assign n10488 = ~n2033 & n10487 ;
  assign n10489 = n1827 | n10488 ;
  assign n10490 = n10485 | n10489 ;
  assign n10491 = n10482 &  n10490 ;
  assign n10492 = n10477 | n10491 ;
  assign n10493 = ~n10014 & n10209 ;
  assign n10494 = ( n10001 & n10006 ) | ( n10001 & n10209 ) | ( n10006 & n10209 ) ;
  assign n10496 = ( n10493 & ~n10001 ) | ( n10493 & n10494 ) | ( ~n10001 & n10494 ) ;
  assign n10495 = ( n10209 & ~n10494 ) | ( n10209 & n10493 ) | ( ~n10494 & n10493 ) ;
  assign n10497 = ( n10006 & ~n10496 ) | ( n10006 & n10495 ) | ( ~n10496 & n10495 ) ;
  assign n10498 = ( n1636 & ~n10492 ) | ( n1636 & n10497 ) | ( ~n10492 & n10497 ) ;
  assign n10499 = n1452 | n10498 ;
  assign n10500 = n10034 | n10209 ;
  assign n10501 = ( n10021 & ~n10030 ) | ( n10021 & n10034 ) | ( ~n10030 & n10034 ) ;
  assign n10502 = ( n10030 & n10500 ) | ( n10030 & n10501 ) | ( n10500 & n10501 ) ;
  assign n10503 = ( n10034 & ~n10501 ) | ( n10034 & n10500 ) | ( ~n10501 & n10500 ) ;
  assign n10504 = ( n10021 & ~n10502 ) | ( n10021 & n10503 ) | ( ~n10502 & n10503 ) ;
  assign n10505 = ( n1636 & ~n10477 ) | ( n1636 & 1'b0 ) | ( ~n10477 & 1'b0 ) ;
  assign n10506 = ~n10491 & n10505 ;
  assign n10507 = n10497 | n10506 ;
  assign n10508 = n10485 | n10488 ;
  assign n10509 = ( n1827 & n10482 ) | ( n1827 & n10508 ) | ( n10482 & n10508 ) ;
  assign n10510 = ~n1636 & n10509 ;
  assign n10511 = ( n1452 & ~n10510 ) | ( n1452 & 1'b0 ) | ( ~n10510 & 1'b0 ) ;
  assign n10512 = n10507 &  n10511 ;
  assign n10513 = ( n10504 & ~n10512 ) | ( n10504 & 1'b0 ) | ( ~n10512 & 1'b0 ) ;
  assign n10514 = ( n10499 & ~n10513 ) | ( n10499 & 1'b0 ) | ( ~n10513 & 1'b0 ) ;
  assign n10515 = n10036 &  n10209 ;
  assign n10516 = ( n10023 & ~n10515 ) | ( n10023 & n10209 ) | ( ~n10515 & n10209 ) ;
  assign n10517 = ( n10028 & ~n10023 ) | ( n10028 & n10516 ) | ( ~n10023 & n10516 ) ;
  assign n10518 = ( n10023 & ~n10516 ) | ( n10023 & n10028 ) | ( ~n10516 & n10028 ) ;
  assign n10519 = ( n10517 & ~n10028 ) | ( n10517 & n10518 ) | ( ~n10028 & n10518 ) ;
  assign n10520 = ( n10514 & ~n1283 ) | ( n10514 & n10519 ) | ( ~n1283 & n10519 ) ;
  assign n10521 = n1122 | n10520 ;
  assign n10522 = n10056 | n10209 ;
  assign n10523 = ( n10043 & ~n10056 ) | ( n10043 & n10052 ) | ( ~n10056 & n10052 ) ;
  assign n10525 = ( n10056 & n10522 ) | ( n10056 & n10523 ) | ( n10522 & n10523 ) ;
  assign n10524 = ( n10052 & ~n10523 ) | ( n10052 & n10522 ) | ( ~n10523 & n10522 ) ;
  assign n10526 = ( n10043 & ~n10525 ) | ( n10043 & n10524 ) | ( ~n10525 & n10524 ) ;
  assign n10527 = ~n1283 & n10499 ;
  assign n10528 = ~n10513 & n10527 ;
  assign n10529 = n10519 | n10528 ;
  assign n10530 = ( n10507 & ~n10510 ) | ( n10507 & 1'b0 ) | ( ~n10510 & 1'b0 ) ;
  assign n10531 = ( n1452 & ~n10504 ) | ( n1452 & n10530 ) | ( ~n10504 & n10530 ) ;
  assign n10532 = ( n1283 & ~n10531 ) | ( n1283 & 1'b0 ) | ( ~n10531 & 1'b0 ) ;
  assign n10533 = ( n1122 & ~n10532 ) | ( n1122 & 1'b0 ) | ( ~n10532 & 1'b0 ) ;
  assign n10534 = n10529 &  n10533 ;
  assign n10535 = n10526 | n10534 ;
  assign n10536 = n10521 &  n10535 ;
  assign n10542 = ( n976 & ~n10541 ) | ( n976 & n10536 ) | ( ~n10541 & n10536 ) ;
  assign n10543 = ( n837 & ~n10542 ) | ( n837 & 1'b0 ) | ( ~n10542 & 1'b0 ) ;
  assign n10545 = ( n10074 & ~n10065 ) | ( n10074 & n10078 ) | ( ~n10065 & n10078 ) ;
  assign n10544 = ( n10078 & ~n10209 ) | ( n10078 & 1'b0 ) | ( ~n10209 & 1'b0 ) ;
  assign n10547 = ( n10078 & ~n10545 ) | ( n10078 & n10544 ) | ( ~n10545 & n10544 ) ;
  assign n10546 = ( n10544 & ~n10074 ) | ( n10544 & n10545 ) | ( ~n10074 & n10545 ) ;
  assign n10548 = ( n10065 & ~n10547 ) | ( n10065 & n10546 ) | ( ~n10547 & n10546 ) ;
  assign n10549 = n976 &  n10521 ;
  assign n10550 = n10535 &  n10549 ;
  assign n10551 = ( n10541 & ~n10550 ) | ( n10541 & 1'b0 ) | ( ~n10550 & 1'b0 ) ;
  assign n10552 = ( n10529 & ~n10532 ) | ( n10529 & 1'b0 ) | ( ~n10532 & 1'b0 ) ;
  assign n10553 = ( n1122 & n10526 ) | ( n1122 & n10552 ) | ( n10526 & n10552 ) ;
  assign n10554 = n976 | n10553 ;
  assign n10555 = ~n837 & n10554 ;
  assign n10556 = ~n10551 & n10555 ;
  assign n10557 = ( n10548 & ~n10556 ) | ( n10548 & 1'b0 ) | ( ~n10556 & 1'b0 ) ;
  assign n10558 = n10543 | n10557 ;
  assign n10564 = ( n713 & ~n10563 ) | ( n713 & n10558 ) | ( ~n10563 & n10558 ) ;
  assign n10565 = n595 &  n10564 ;
  assign n10566 = n10100 | n10209 ;
  assign n10567 = ( n10087 & ~n10096 ) | ( n10087 & n10100 ) | ( ~n10096 & n10100 ) ;
  assign n10568 = ( n10096 & n10566 ) | ( n10096 & n10567 ) | ( n10566 & n10567 ) ;
  assign n10569 = ( n10100 & ~n10567 ) | ( n10100 & n10566 ) | ( ~n10567 & n10566 ) ;
  assign n10570 = ( n10087 & ~n10568 ) | ( n10087 & n10569 ) | ( ~n10568 & n10569 ) ;
  assign n10571 = n713 | n10543 ;
  assign n10572 = n10557 | n10571 ;
  assign n10573 = ~n10563 & n10572 ;
  assign n10574 = ~n10551 & n10554 ;
  assign n10575 = ( n837 & ~n10574 ) | ( n837 & n10548 ) | ( ~n10574 & n10548 ) ;
  assign n10576 = n713 &  n10575 ;
  assign n10577 = n595 | n10576 ;
  assign n10578 = n10573 | n10577 ;
  assign n10579 = n10570 &  n10578 ;
  assign n10580 = n10565 | n10579 ;
  assign n10581 = ~n10102 & n10209 ;
  assign n10582 = ( n10089 & ~n10581 ) | ( n10089 & n10209 ) | ( ~n10581 & n10209 ) ;
  assign n10583 = ( n10089 & ~n10582 ) | ( n10089 & n10094 ) | ( ~n10582 & n10094 ) ;
  assign n10584 = ( n10094 & ~n10089 ) | ( n10094 & n10582 ) | ( ~n10089 & n10582 ) ;
  assign n10585 = ( n10583 & ~n10094 ) | ( n10583 & n10584 ) | ( ~n10094 & n10584 ) ;
  assign n10586 = ( n492 & n10580 ) | ( n492 & n10585 ) | ( n10580 & n10585 ) ;
  assign n10587 = n396 &  n10586 ;
  assign n10589 = ( n10118 & ~n10109 ) | ( n10118 & n10122 ) | ( ~n10109 & n10122 ) ;
  assign n10588 = n10122 | n10209 ;
  assign n10591 = ( n10122 & ~n10589 ) | ( n10122 & n10588 ) | ( ~n10589 & n10588 ) ;
  assign n10590 = ( n10588 & ~n10118 ) | ( n10588 & n10589 ) | ( ~n10118 & n10589 ) ;
  assign n10592 = ( n10109 & ~n10591 ) | ( n10109 & n10590 ) | ( ~n10591 & n10590 ) ;
  assign n10593 = n492 | n10565 ;
  assign n10594 = n10579 | n10593 ;
  assign n10595 = n10585 &  n10594 ;
  assign n10596 = n10573 | n10576 ;
  assign n10597 = ( n595 & n10570 ) | ( n595 & n10596 ) | ( n10570 & n10596 ) ;
  assign n10598 = n492 &  n10597 ;
  assign n10599 = n396 | n10598 ;
  assign n10600 = n10595 | n10599 ;
  assign n10601 = ~n10592 & n10600 ;
  assign n10602 = n10587 | n10601 ;
  assign n10604 = ( n10111 & ~n10116 ) | ( n10111 & n10209 ) | ( ~n10116 & n10209 ) ;
  assign n10603 = ~n10124 & n10209 ;
  assign n10605 = ( n10209 & ~n10604 ) | ( n10209 & n10603 ) | ( ~n10604 & n10603 ) ;
  assign n10606 = ( n10603 & ~n10111 ) | ( n10603 & n10604 ) | ( ~n10111 & n10604 ) ;
  assign n10607 = ( n10116 & ~n10605 ) | ( n10116 & n10606 ) | ( ~n10605 & n10606 ) ;
  assign n10608 = ( n315 & n10602 ) | ( n315 & n10607 ) | ( n10602 & n10607 ) ;
  assign n10609 = n240 &  n10608 ;
  assign n10611 = ( n10140 & ~n10131 ) | ( n10140 & n10144 ) | ( ~n10131 & n10144 ) ;
  assign n10610 = n10144 | n10209 ;
  assign n10613 = ( n10144 & ~n10611 ) | ( n10144 & n10610 ) | ( ~n10611 & n10610 ) ;
  assign n10612 = ( n10610 & ~n10140 ) | ( n10610 & n10611 ) | ( ~n10140 & n10611 ) ;
  assign n10614 = ( n10131 & ~n10613 ) | ( n10131 & n10612 ) | ( ~n10613 & n10612 ) ;
  assign n10615 = n315 | n10587 ;
  assign n10616 = n10601 | n10615 ;
  assign n10617 = n10607 &  n10616 ;
  assign n10618 = n10595 | n10598 ;
  assign n10619 = ( n396 & ~n10592 ) | ( n396 & n10618 ) | ( ~n10592 & n10618 ) ;
  assign n10620 = n315 &  n10619 ;
  assign n10621 = n240 | n10620 ;
  assign n10622 = n10617 | n10621 ;
  assign n10623 = ~n10614 & n10622 ;
  assign n10624 = n10609 | n10623 ;
  assign n10625 = ~n10146 & n10209 ;
  assign n10626 = ( n10133 & ~n10625 ) | ( n10133 & n10209 ) | ( ~n10625 & n10209 ) ;
  assign n10627 = ( n10133 & ~n10626 ) | ( n10133 & n10138 ) | ( ~n10626 & n10138 ) ;
  assign n10628 = ( n10138 & ~n10133 ) | ( n10138 & n10626 ) | ( ~n10133 & n10626 ) ;
  assign n10629 = ( n10627 & ~n10138 ) | ( n10627 & n10628 ) | ( ~n10138 & n10628 ) ;
  assign n10630 = ( n181 & n10624 ) | ( n181 & n10629 ) | ( n10624 & n10629 ) ;
  assign n10631 = ~n145 & n10630 ;
  assign n10633 = ( n10162 & ~n10153 ) | ( n10162 & n10166 ) | ( ~n10153 & n10166 ) ;
  assign n10632 = n10166 | n10209 ;
  assign n10635 = ( n10166 & ~n10633 ) | ( n10166 & n10632 ) | ( ~n10633 & n10632 ) ;
  assign n10634 = ( n10632 & ~n10162 ) | ( n10632 & n10633 ) | ( ~n10162 & n10633 ) ;
  assign n10636 = ( n10153 & ~n10635 ) | ( n10153 & n10634 ) | ( ~n10635 & n10634 ) ;
  assign n10637 = n181 | n10609 ;
  assign n10638 = n10623 | n10637 ;
  assign n10639 = n10629 &  n10638 ;
  assign n10640 = n10617 | n10620 ;
  assign n10641 = ( n240 & ~n10614 ) | ( n240 & n10640 ) | ( ~n10614 & n10640 ) ;
  assign n10642 = n181 &  n10641 ;
  assign n10643 = ( n145 & ~n10642 ) | ( n145 & 1'b0 ) | ( ~n10642 & 1'b0 ) ;
  assign n10644 = ~n10639 & n10643 ;
  assign n10645 = ( n10636 & ~n10644 ) | ( n10636 & 1'b0 ) | ( ~n10644 & 1'b0 ) ;
  assign n10646 = n10631 | n10645 ;
  assign n10652 = ( n150 & ~n10651 ) | ( n150 & n10646 ) | ( ~n10651 & n10646 ) ;
  assign n10664 = n10652 | n10663 ;
  assign n10665 = ( n133 & ~n10663 ) | ( n133 & n10664 ) | ( ~n10663 & n10664 ) ;
  assign n10666 = n150 | n10631 ;
  assign n10667 = n10645 | n10666 ;
  assign n10672 = n10651 | n10667 ;
  assign n10668 = n10639 | n10642 ;
  assign n10669 = ( n10636 & ~n145 ) | ( n10636 & n10668 ) | ( ~n145 & n10668 ) ;
  assign n10670 = n150 &  n10669 ;
  assign n10671 = ( n10659 & ~n10670 ) | ( n10659 & 1'b0 ) | ( ~n10670 & 1'b0 ) ;
  assign n10673 = ( n10651 & ~n10672 ) | ( n10651 & n10671 ) | ( ~n10672 & n10671 ) ;
  assign n10675 = ( n133 & ~n10176 ) | ( n133 & n10183 ) | ( ~n10176 & n10183 ) ;
  assign n10674 = ( n10176 & ~n10183 ) | ( n10176 & n10209 ) | ( ~n10183 & n10209 ) ;
  assign n10676 = n10183 &  n10674 ;
  assign n10677 = ( n10675 & ~n10183 ) | ( n10675 & n10676 ) | ( ~n10183 & n10676 ) ;
  assign n10678 = n10179 | n10206 ;
  assign n10679 = ( n10201 & ~n10182 ) | ( n10201 & n10678 ) | ( ~n10182 & n10678 ) ;
  assign n10680 = n10182 | n10679 ;
  assign n10681 = ( n10189 & n10197 ) | ( n10189 & n10680 ) | ( n10197 & n10680 ) ;
  assign n10682 = ( n10189 & ~n10681 ) | ( n10189 & 1'b0 ) | ( ~n10681 & 1'b0 ) ;
  assign n10683 = n10677 | n10682 ;
  assign n10684 = n10673 | n10683 ;
  assign n10685 = ~n10665 |  n10684 ;
  assign n10919 = ~n10425 & n10685 ;
  assign n10920 = ( n10412 & n10417 ) | ( n10412 & n10685 ) | ( n10417 & n10685 ) ;
  assign n10922 = ( n10919 & ~n10412 ) | ( n10919 & n10920 ) | ( ~n10412 & n10920 ) ;
  assign n10921 = ( n10685 & ~n10920 ) | ( n10685 & n10919 ) | ( ~n10920 & n10919 ) ;
  assign n10923 = ( n10417 & ~n10922 ) | ( n10417 & n10921 ) | ( ~n10922 & n10921 ) ;
  assign n10905 = ( n10419 & ~n10410 ) | ( n10419 & n10423 ) | ( ~n10410 & n10423 ) ;
  assign n10904 = n10423 | n10685 ;
  assign n10907 = ( n10423 & ~n10905 ) | ( n10423 & n10904 ) | ( ~n10905 & n10904 ) ;
  assign n10906 = ( n10904 & ~n10419 ) | ( n10904 & n10905 ) | ( ~n10419 & n10905 ) ;
  assign n10908 = ( n10410 & ~n10907 ) | ( n10410 & n10906 ) | ( ~n10907 & n10906 ) ;
  assign n10898 = ( n10390 & ~n10395 ) | ( n10390 & n10685 ) | ( ~n10395 & n10685 ) ;
  assign n10897 = ~n10403 & n10685 ;
  assign n10899 = ( n10685 & ~n10898 ) | ( n10685 & n10897 ) | ( ~n10898 & n10897 ) ;
  assign n10900 = ( n10897 & ~n10390 ) | ( n10897 & n10898 ) | ( ~n10390 & n10898 ) ;
  assign n10901 = ( n10395 & ~n10899 ) | ( n10395 & n10900 ) | ( ~n10899 & n10900 ) ;
  assign n10883 = ( n10397 & ~n10388 ) | ( n10397 & n10401 ) | ( ~n10388 & n10401 ) ;
  assign n10882 = n10401 | n10685 ;
  assign n10885 = ( n10401 & ~n10883 ) | ( n10401 & n10882 ) | ( ~n10883 & n10882 ) ;
  assign n10884 = ( n10882 & ~n10397 ) | ( n10882 & n10883 ) | ( ~n10397 & n10883 ) ;
  assign n10886 = ( n10388 & ~n10885 ) | ( n10388 & n10884 ) | ( ~n10885 & n10884 ) ;
  assign n10875 = ~n10381 & n10685 ;
  assign n10876 = ( n10368 & n10373 ) | ( n10368 & n10685 ) | ( n10373 & n10685 ) ;
  assign n10878 = ( n10875 & ~n10368 ) | ( n10875 & n10876 ) | ( ~n10368 & n10876 ) ;
  assign n10877 = ( n10685 & ~n10876 ) | ( n10685 & n10875 ) | ( ~n10876 & n10875 ) ;
  assign n10879 = ( n10373 & ~n10878 ) | ( n10373 & n10877 ) | ( ~n10878 & n10877 ) ;
  assign n10861 = ( n10375 & ~n10366 ) | ( n10375 & n10379 ) | ( ~n10366 & n10379 ) ;
  assign n10860 = n10379 | n10685 ;
  assign n10863 = ( n10379 & ~n10861 ) | ( n10379 & n10860 ) | ( ~n10861 & n10860 ) ;
  assign n10862 = ( n10860 & ~n10375 ) | ( n10860 & n10861 ) | ( ~n10375 & n10861 ) ;
  assign n10864 = ( n10366 & ~n10863 ) | ( n10366 & n10862 ) | ( ~n10863 & n10862 ) ;
  assign n10853 = ~n10359 & n10685 ;
  assign n10854 = ( n10346 & ~n10853 ) | ( n10346 & n10685 ) | ( ~n10853 & n10685 ) ;
  assign n10855 = ( n10346 & ~n10854 ) | ( n10346 & n10351 ) | ( ~n10854 & n10351 ) ;
  assign n10856 = ( n10351 & ~n10346 ) | ( n10351 & n10854 ) | ( ~n10346 & n10854 ) ;
  assign n10857 = ( n10855 & ~n10351 ) | ( n10855 & n10856 ) | ( ~n10351 & n10856 ) ;
  assign n10838 = n10357 | n10685 ;
  assign n10839 = ( n10344 & ~n10353 ) | ( n10344 & n10357 ) | ( ~n10353 & n10357 ) ;
  assign n10840 = ( n10353 & n10838 ) | ( n10353 & n10839 ) | ( n10838 & n10839 ) ;
  assign n10841 = ( n10357 & ~n10839 ) | ( n10357 & n10838 ) | ( ~n10839 & n10838 ) ;
  assign n10842 = ( n10344 & ~n10840 ) | ( n10344 & n10841 ) | ( ~n10840 & n10841 ) ;
  assign n10831 = n10337 &  n10685 ;
  assign n10832 = ( n10324 & n10329 ) | ( n10324 & n10685 ) | ( n10329 & n10685 ) ;
  assign n10834 = ( n10831 & ~n10324 ) | ( n10831 & n10832 ) | ( ~n10324 & n10832 ) ;
  assign n10833 = ( n10685 & ~n10832 ) | ( n10685 & n10831 ) | ( ~n10832 & n10831 ) ;
  assign n10835 = ( n10329 & ~n10834 ) | ( n10329 & n10833 ) | ( ~n10834 & n10833 ) ;
  assign n10816 = n10335 | n10685 ;
  assign n10817 = ( n10322 & ~n10331 ) | ( n10322 & n10335 ) | ( ~n10331 & n10335 ) ;
  assign n10818 = ( n10331 & n10816 ) | ( n10331 & n10817 ) | ( n10816 & n10817 ) ;
  assign n10819 = ( n10335 & ~n10817 ) | ( n10335 & n10816 ) | ( ~n10817 & n10816 ) ;
  assign n10820 = ( n10322 & ~n10818 ) | ( n10322 & n10819 ) | ( ~n10818 & n10819 ) ;
  assign n10809 = n10302 | n10685 ;
  assign n10810 = ( n10307 & ~n10302 ) | ( n10307 & n10315 ) | ( ~n10302 & n10315 ) ;
  assign n10812 = ( n10302 & n10809 ) | ( n10302 & n10810 ) | ( n10809 & n10810 ) ;
  assign n10811 = ( n10315 & ~n10810 ) | ( n10315 & n10809 ) | ( ~n10810 & n10809 ) ;
  assign n10813 = ( n10307 & ~n10812 ) | ( n10307 & n10811 ) | ( ~n10812 & n10811 ) ;
  assign n10794 = n10313 | n10685 ;
  assign n10795 = ( n10300 & n10309 ) | ( n10300 & n10313 ) | ( n10309 & n10313 ) ;
  assign n10796 = ( n10794 & ~n10309 ) | ( n10794 & n10795 ) | ( ~n10309 & n10795 ) ;
  assign n10797 = ( n10313 & ~n10795 ) | ( n10313 & n10794 ) | ( ~n10795 & n10794 ) ;
  assign n10798 = ( n10300 & ~n10796 ) | ( n10300 & n10797 ) | ( ~n10796 & n10797 ) ;
  assign n10787 = n10280 | n10685 ;
  assign n10788 = ( n10280 & ~n10293 ) | ( n10280 & n10285 ) | ( ~n10293 & n10285 ) ;
  assign n10789 = ( n10293 & n10787 ) | ( n10293 & n10788 ) | ( n10787 & n10788 ) ;
  assign n10790 = ( n10280 & ~n10788 ) | ( n10280 & n10787 ) | ( ~n10788 & n10787 ) ;
  assign n10791 = ( n10285 & ~n10789 ) | ( n10285 & n10790 ) | ( ~n10789 & n10790 ) ;
  assign n10772 = n10291 | n10685 ;
  assign n10773 = ( n10278 & ~n10291 ) | ( n10278 & n10287 ) | ( ~n10291 & n10287 ) ;
  assign n10775 = ( n10291 & n10772 ) | ( n10291 & n10773 ) | ( n10772 & n10773 ) ;
  assign n10774 = ( n10287 & ~n10773 ) | ( n10287 & n10772 ) | ( ~n10773 & n10772 ) ;
  assign n10776 = ( n10278 & ~n10775 ) | ( n10278 & n10774 ) | ( ~n10775 & n10774 ) ;
  assign n10765 = n10258 | n10685 ;
  assign n10766 = ( n10258 & n10263 ) | ( n10258 & n10271 ) | ( n10263 & n10271 ) ;
  assign n10767 = ( n10765 & ~n10271 ) | ( n10765 & n10766 ) | ( ~n10271 & n10766 ) ;
  assign n10768 = ( n10258 & ~n10766 ) | ( n10258 & n10765 ) | ( ~n10766 & n10765 ) ;
  assign n10769 = ( n10263 & ~n10767 ) | ( n10263 & n10768 ) | ( ~n10767 & n10768 ) ;
  assign n10750 = n10269 | n10685 ;
  assign n10751 = ( n10256 & n10265 ) | ( n10256 & n10269 ) | ( n10265 & n10269 ) ;
  assign n10752 = ( n10750 & ~n10265 ) | ( n10750 & n10751 ) | ( ~n10265 & n10751 ) ;
  assign n10753 = ( n10269 & ~n10751 ) | ( n10269 & n10750 ) | ( ~n10751 & n10750 ) ;
  assign n10754 = ( n10256 & ~n10752 ) | ( n10256 & n10753 ) | ( ~n10752 & n10753 ) ;
  assign n10743 = n10232 | n10685 ;
  assign n10744 = ( n10242 & ~n10232 ) | ( n10242 & n10249 ) | ( ~n10232 & n10249 ) ;
  assign n10746 = ( n10232 & n10743 ) | ( n10232 & n10744 ) | ( n10743 & n10744 ) ;
  assign n10745 = ( n10249 & ~n10744 ) | ( n10249 & n10743 ) | ( ~n10744 & n10743 ) ;
  assign n10747 = ( n10242 & ~n10746 ) | ( n10242 & n10745 ) | ( ~n10746 & n10745 ) ;
  assign n10728 = ~n10244 & n10247 ;
  assign n10729 = ( n10230 & ~n10728 ) | ( n10230 & n10244 ) | ( ~n10728 & n10244 ) ;
  assign n10730 = ( n10685 & n10728 ) | ( n10685 & n10729 ) | ( n10728 & n10729 ) ;
  assign n10731 = ( n10244 & ~n10729 ) | ( n10244 & n10685 ) | ( ~n10729 & n10685 ) ;
  assign n10732 = ( n10230 & ~n10730 ) | ( n10230 & n10731 ) | ( ~n10730 & n10731 ) ;
  assign n10719 = ~x44 & n10209 ;
  assign n10720 = ( x45 & ~n10719 ) | ( x45 & 1'b0 ) | ( ~n10719 & 1'b0 ) ;
  assign n10721 = n10221 | n10720 ;
  assign n10716 = ( n10209 & ~x44 ) | ( n10209 & n10216 ) | ( ~x44 & n10216 ) ;
  assign n10717 = x44 &  n10716 ;
  assign n10718 = ( n10211 & ~n10216 ) | ( n10211 & n10717 ) | ( ~n10216 & n10717 ) ;
  assign n10722 = ( n10718 & ~n10685 ) | ( n10718 & n10721 ) | ( ~n10685 & n10721 ) ;
  assign n10724 = n10685 &  n10722 ;
  assign n10723 = ( n10718 & ~n10722 ) | ( n10718 & 1'b0 ) | ( ~n10722 & 1'b0 ) ;
  assign n10725 = ( n10721 & ~n10724 ) | ( n10721 & n10723 ) | ( ~n10724 & n10723 ) ;
  assign n10692 = ( x42 & ~n10685 ) | ( x42 & x43 ) | ( ~n10685 & x43 ) ;
  assign n10698 = ( x42 & ~x43 ) | ( x42 & 1'b0 ) | ( ~x43 & 1'b0 ) ;
  assign n10688 = x40 | x41 ;
  assign n10693 = ~x42 & n10688 ;
  assign n10694 = ( x42 & ~n10207 ) | ( x42 & n10693 ) | ( ~n10207 & n10693 ) ;
  assign n10695 = ( n10189 & ~n10694 ) | ( n10189 & n10197 ) | ( ~n10694 & n10197 ) ;
  assign n10696 = ( n10189 & ~n10695 ) | ( n10189 & 1'b0 ) | ( ~n10695 & 1'b0 ) ;
  assign n10697 = ( n10685 & ~x43 ) | ( n10685 & n10696 ) | ( ~x43 & n10696 ) ;
  assign n10699 = ( n10692 & ~n10698 ) | ( n10692 & n10697 ) | ( ~n10698 & n10697 ) ;
  assign n10689 = x42 | n10688 ;
  assign n10690 = x42 &  n10685 ;
  assign n10691 = ( n10209 & ~n10689 ) | ( n10209 & n10690 ) | ( ~n10689 & n10690 ) ;
  assign n10702 = ( n9740 & ~n10691 ) | ( n9740 & 1'b0 ) | ( ~n10691 & 1'b0 ) ;
  assign n10703 = n10699 &  n10702 ;
  assign n10705 = ( n10209 & ~n10682 ) | ( n10209 & 1'b0 ) | ( ~n10682 & 1'b0 ) ;
  assign n10706 = ( n10673 & ~n10677 ) | ( n10673 & n10705 ) | ( ~n10677 & n10705 ) ;
  assign n10707 = ~n10673 & n10706 ;
  assign n10708 = n10665 &  n10707 ;
  assign n10704 = ~n9741 & n10685 ;
  assign n10709 = ( n10704 & ~n10708 ) | ( n10704 & 1'b0 ) | ( ~n10708 & 1'b0 ) ;
  assign n10710 = ( x44 & n10708 ) | ( x44 & n10709 ) | ( n10708 & n10709 ) ;
  assign n10711 = x44 | n10708 ;
  assign n10712 = n10704 | n10711 ;
  assign n10713 = ~n10710 & n10712 ;
  assign n10714 = n10703 | n10713 ;
  assign n10700 = n10691 &  n10699 ;
  assign n10701 = ( n9740 & ~n10700 ) | ( n9740 & n10699 ) | ( ~n10700 & n10699 ) ;
  assign n10733 = ~n9286 & n10701 ;
  assign n10734 = n10714 &  n10733 ;
  assign n10735 = n10725 | n10734 ;
  assign n10736 = ~n10691 & n10699 ;
  assign n10737 = ( n9740 & n10713 ) | ( n9740 & n10736 ) | ( n10713 & n10736 ) ;
  assign n10738 = ( n9286 & ~n10737 ) | ( n9286 & 1'b0 ) | ( ~n10737 & 1'b0 ) ;
  assign n10739 = n8839 | n10738 ;
  assign n10740 = ( n10735 & ~n10739 ) | ( n10735 & 1'b0 ) | ( ~n10739 & 1'b0 ) ;
  assign n10741 = n10732 | n10740 ;
  assign n10715 = n10701 &  n10714 ;
  assign n10726 = ( n10715 & ~n9286 ) | ( n10715 & n10725 ) | ( ~n9286 & n10725 ) ;
  assign n10727 = ( n8839 & ~n10726 ) | ( n8839 & 1'b0 ) | ( ~n10726 & 1'b0 ) ;
  assign n10755 = n8407 | n10727 ;
  assign n10756 = ( n10741 & ~n10755 ) | ( n10741 & 1'b0 ) | ( ~n10755 & 1'b0 ) ;
  assign n10757 = ( n10747 & ~n10756 ) | ( n10747 & 1'b0 ) | ( ~n10756 & 1'b0 ) ;
  assign n10758 = ( n10735 & ~n10738 ) | ( n10735 & 1'b0 ) | ( ~n10738 & 1'b0 ) ;
  assign n10759 = ( n10732 & ~n8839 ) | ( n10732 & n10758 ) | ( ~n8839 & n10758 ) ;
  assign n10760 = ( n8407 & ~n10759 ) | ( n8407 & 1'b0 ) | ( ~n10759 & 1'b0 ) ;
  assign n10761 = n7982 | n10760 ;
  assign n10762 = n10757 | n10761 ;
  assign n10763 = n10754 &  n10762 ;
  assign n10742 = ~n10727 & n10741 ;
  assign n10748 = ( n8407 & ~n10742 ) | ( n8407 & n10747 ) | ( ~n10742 & n10747 ) ;
  assign n10749 = n7982 &  n10748 ;
  assign n10777 = ( n7572 & ~n10749 ) | ( n7572 & 1'b0 ) | ( ~n10749 & 1'b0 ) ;
  assign n10778 = ~n10763 & n10777 ;
  assign n10779 = ( n10769 & ~n10778 ) | ( n10769 & 1'b0 ) | ( ~n10778 & 1'b0 ) ;
  assign n10780 = n10757 | n10760 ;
  assign n10781 = ( n7982 & n10754 ) | ( n7982 & n10780 ) | ( n10754 & n10780 ) ;
  assign n10782 = ~n7572 & n10781 ;
  assign n10783 = ( n7169 & ~n10782 ) | ( n7169 & 1'b0 ) | ( ~n10782 & 1'b0 ) ;
  assign n10784 = ~n10779 & n10783 ;
  assign n10785 = ( n10776 & ~n10784 ) | ( n10776 & 1'b0 ) | ( ~n10784 & 1'b0 ) ;
  assign n10764 = n10749 | n10763 ;
  assign n10770 = ( n10764 & ~n7572 ) | ( n10764 & n10769 ) | ( ~n7572 & n10769 ) ;
  assign n10771 = ~n7169 & n10770 ;
  assign n10799 = n6781 | n10771 ;
  assign n10800 = n10785 | n10799 ;
  assign n10801 = n10791 &  n10800 ;
  assign n10802 = n10779 | n10782 ;
  assign n10803 = ( n10776 & ~n7169 ) | ( n10776 & n10802 ) | ( ~n7169 & n10802 ) ;
  assign n10804 = n6781 &  n10803 ;
  assign n10805 = ( n6399 & ~n10804 ) | ( n6399 & 1'b0 ) | ( ~n10804 & 1'b0 ) ;
  assign n10806 = ~n10801 & n10805 ;
  assign n10807 = n10798 | n10806 ;
  assign n10786 = n10771 | n10785 ;
  assign n10792 = ( n6781 & n10786 ) | ( n6781 & n10791 ) | ( n10786 & n10791 ) ;
  assign n10793 = ~n6399 & n10792 ;
  assign n10821 = n6032 | n10793 ;
  assign n10822 = ( n10807 & ~n10821 ) | ( n10807 & 1'b0 ) | ( ~n10821 & 1'b0 ) ;
  assign n10823 = n10813 | n10822 ;
  assign n10824 = n10801 | n10804 ;
  assign n10825 = ( n6399 & ~n10824 ) | ( n6399 & n10798 ) | ( ~n10824 & n10798 ) ;
  assign n10826 = ( n6032 & ~n10825 ) | ( n6032 & 1'b0 ) | ( ~n10825 & 1'b0 ) ;
  assign n10827 = ( n5672 & ~n10826 ) | ( n5672 & 1'b0 ) | ( ~n10826 & 1'b0 ) ;
  assign n10828 = n10823 &  n10827 ;
  assign n10829 = ( n10820 & ~n10828 ) | ( n10820 & 1'b0 ) | ( ~n10828 & 1'b0 ) ;
  assign n10808 = ~n10793 & n10807 ;
  assign n10814 = ( n10808 & ~n6032 ) | ( n10808 & n10813 ) | ( ~n6032 & n10813 ) ;
  assign n10815 = n5672 | n10814 ;
  assign n10843 = ~n5327 & n10815 ;
  assign n10844 = ~n10829 & n10843 ;
  assign n10845 = n10835 | n10844 ;
  assign n10846 = ( n10823 & ~n10826 ) | ( n10823 & 1'b0 ) | ( ~n10826 & 1'b0 ) ;
  assign n10847 = ( n5672 & ~n10820 ) | ( n5672 & n10846 ) | ( ~n10820 & n10846 ) ;
  assign n10848 = ( n5327 & ~n10847 ) | ( n5327 & 1'b0 ) | ( ~n10847 & 1'b0 ) ;
  assign n10849 = n4990 | n10848 ;
  assign n10850 = ( n10845 & ~n10849 ) | ( n10845 & 1'b0 ) | ( ~n10849 & 1'b0 ) ;
  assign n10851 = ( n10842 & ~n10850 ) | ( n10842 & 1'b0 ) | ( ~n10850 & 1'b0 ) ;
  assign n10830 = ( n10815 & ~n10829 ) | ( n10815 & 1'b0 ) | ( ~n10829 & 1'b0 ) ;
  assign n10836 = ( n10830 & ~n5327 ) | ( n10830 & n10835 ) | ( ~n5327 & n10835 ) ;
  assign n10837 = ( n4990 & ~n10836 ) | ( n4990 & 1'b0 ) | ( ~n10836 & 1'b0 ) ;
  assign n10865 = n4668 | n10837 ;
  assign n10866 = n10851 | n10865 ;
  assign n10867 = n10857 &  n10866 ;
  assign n10868 = ( n10845 & ~n10848 ) | ( n10845 & 1'b0 ) | ( ~n10848 & 1'b0 ) ;
  assign n10869 = ( n4990 & ~n10868 ) | ( n4990 & n10842 ) | ( ~n10868 & n10842 ) ;
  assign n10870 = n4668 &  n10869 ;
  assign n10871 = n4353 | n10870 ;
  assign n10872 = n10867 | n10871 ;
  assign n10873 = ~n10864 & n10872 ;
  assign n10852 = n10837 | n10851 ;
  assign n10858 = ( n4668 & n10852 ) | ( n4668 & n10857 ) | ( n10852 & n10857 ) ;
  assign n10859 = n4353 &  n10858 ;
  assign n10887 = n4053 | n10859 ;
  assign n10888 = n10873 | n10887 ;
  assign n10889 = ~n10879 & n10888 ;
  assign n10890 = n10867 | n10870 ;
  assign n10891 = ( n4353 & ~n10864 ) | ( n4353 & n10890 ) | ( ~n10864 & n10890 ) ;
  assign n10892 = n4053 &  n10891 ;
  assign n10893 = n3760 | n10892 ;
  assign n10894 = n10889 | n10893 ;
  assign n10895 = ~n10886 & n10894 ;
  assign n10874 = n10859 | n10873 ;
  assign n10880 = ( n4053 & ~n10879 ) | ( n4053 & n10874 ) | ( ~n10879 & n10874 ) ;
  assign n10881 = n3760 &  n10880 ;
  assign n10909 = n3482 | n10881 ;
  assign n10910 = n10895 | n10909 ;
  assign n10911 = ~n10901 & n10910 ;
  assign n10912 = n10889 | n10892 ;
  assign n10913 = ( n3760 & ~n10886 ) | ( n3760 & n10912 ) | ( ~n10886 & n10912 ) ;
  assign n10914 = n3482 &  n10913 ;
  assign n10934 = n10911 | n10914 ;
  assign n10935 = ( n3211 & ~n10908 ) | ( n3211 & n10934 ) | ( ~n10908 & n10934 ) ;
  assign n10936 = n2955 &  n10935 ;
  assign n11144 = n10651 &  n10667 ;
  assign n11145 = ( n10670 & n10685 ) | ( n10670 & n11144 ) | ( n10685 & n11144 ) ;
  assign n11146 = ~n10670 & n11145 ;
  assign n11147 = ( n10667 & ~n10670 ) | ( n10667 & 1'b0 ) | ( ~n10670 & 1'b0 ) ;
  assign n11148 = ~n10685 & n11147 ;
  assign n11149 = ( n10651 & ~n11148 ) | ( n10651 & n11147 ) | ( ~n11148 & n11147 ) ;
  assign n11150 = ~n11146 & n11149 ;
  assign n11151 = ( n10652 & ~n10659 ) | ( n10652 & 1'b0 ) | ( ~n10659 & 1'b0 ) ;
  assign n11152 = ~n10685 & n11151 ;
  assign n11153 = ( n10673 & ~n11152 ) | ( n10673 & n11151 ) | ( ~n11152 & n11151 ) ;
  assign n11154 = n11150 | n11153 ;
  assign n11116 = ~n10622 & n10685 ;
  assign n11117 = ( n10609 & ~n11116 ) | ( n10609 & n10685 ) | ( ~n11116 & n10685 ) ;
  assign n11118 = ( n10614 & ~n10609 ) | ( n10614 & n11117 ) | ( ~n10609 & n11117 ) ;
  assign n11119 = ( n10609 & ~n11117 ) | ( n10609 & n10614 ) | ( ~n11117 & n10614 ) ;
  assign n11120 = ( n11118 & ~n10614 ) | ( n11118 & n11119 ) | ( ~n10614 & n11119 ) ;
  assign n11094 = ~n10600 & n10685 ;
  assign n11095 = ( n10587 & ~n11094 ) | ( n10587 & n10685 ) | ( ~n11094 & n10685 ) ;
  assign n11096 = ( n10592 & ~n10587 ) | ( n10592 & n11095 ) | ( ~n10587 & n11095 ) ;
  assign n11097 = ( n10587 & ~n11095 ) | ( n10587 & n10592 ) | ( ~n11095 & n10592 ) ;
  assign n11098 = ( n11096 & ~n10592 ) | ( n11096 & n11097 ) | ( ~n10592 & n11097 ) ;
  assign n10941 = ( n10434 & n10442 ) | ( n10434 & n10446 ) | ( n10442 & n10446 ) ;
  assign n10942 = ( n10685 & ~n10442 ) | ( n10685 & n10941 ) | ( ~n10442 & n10941 ) ;
  assign n10943 = ( n10434 & ~n10941 ) | ( n10434 & n10685 ) | ( ~n10941 & n10685 ) ;
  assign n10944 = ( n10446 & ~n10942 ) | ( n10446 & n10943 ) | ( ~n10942 & n10943 ) ;
  assign n10896 = n10881 | n10895 ;
  assign n10902 = ( n3482 & ~n10901 ) | ( n3482 & n10896 ) | ( ~n10901 & n10896 ) ;
  assign n10903 = n3211 &  n10902 ;
  assign n10915 = n3211 | n10914 ;
  assign n10916 = n10911 | n10915 ;
  assign n10917 = ~n10908 & n10916 ;
  assign n10918 = n10903 | n10917 ;
  assign n10924 = ( n2955 & n10918 ) | ( n2955 & n10923 ) | ( n10918 & n10923 ) ;
  assign n10925 = n2706 &  n10924 ;
  assign n10927 = ( n10436 & ~n10432 ) | ( n10436 & n10440 ) | ( ~n10432 & n10440 ) ;
  assign n10926 = n10440 | n10685 ;
  assign n10929 = ( n10440 & ~n10927 ) | ( n10440 & n10926 ) | ( ~n10927 & n10926 ) ;
  assign n10928 = ( n10926 & ~n10436 ) | ( n10926 & n10927 ) | ( ~n10436 & n10927 ) ;
  assign n10930 = ( n10432 & ~n10929 ) | ( n10432 & n10928 ) | ( ~n10929 & n10928 ) ;
  assign n10931 = n2955 | n10903 ;
  assign n10932 = n10917 | n10931 ;
  assign n10933 = n10923 &  n10932 ;
  assign n10937 = n2706 | n10936 ;
  assign n10938 = n10933 | n10937 ;
  assign n10939 = ~n10930 & n10938 ;
  assign n10940 = n10925 | n10939 ;
  assign n10945 = ( n2472 & ~n10944 ) | ( n2472 & n10940 ) | ( ~n10944 & n10940 ) ;
  assign n10946 = n2245 &  n10945 ;
  assign n10947 = n10466 | n10685 ;
  assign n10948 = ( n10453 & n10462 ) | ( n10453 & n10466 ) | ( n10462 & n10466 ) ;
  assign n10949 = ( n10947 & ~n10462 ) | ( n10947 & n10948 ) | ( ~n10462 & n10948 ) ;
  assign n10950 = ( n10466 & ~n10948 ) | ( n10466 & n10947 ) | ( ~n10948 & n10947 ) ;
  assign n10951 = ( n10453 & ~n10949 ) | ( n10453 & n10950 ) | ( ~n10949 & n10950 ) ;
  assign n10952 = n2472 | n10925 ;
  assign n10953 = n10939 | n10952 ;
  assign n10954 = ~n10944 & n10953 ;
  assign n10955 = n10933 | n10936 ;
  assign n10956 = ( n2706 & ~n10930 ) | ( n2706 & n10955 ) | ( ~n10930 & n10955 ) ;
  assign n10957 = n2472 &  n10956 ;
  assign n10958 = n2245 | n10957 ;
  assign n10959 = n10954 | n10958 ;
  assign n10960 = n10951 &  n10959 ;
  assign n10961 = n10946 | n10960 ;
  assign n10962 = ~n10468 & n10685 ;
  assign n10963 = ( n10455 & ~n10962 ) | ( n10455 & n10685 ) | ( ~n10962 & n10685 ) ;
  assign n10964 = ( n10460 & ~n10455 ) | ( n10460 & n10963 ) | ( ~n10455 & n10963 ) ;
  assign n10965 = ( n10455 & ~n10963 ) | ( n10455 & n10460 ) | ( ~n10963 & n10460 ) ;
  assign n10966 = ( n10964 & ~n10460 ) | ( n10964 & n10965 ) | ( ~n10460 & n10965 ) ;
  assign n10967 = ( n2033 & ~n10961 ) | ( n2033 & n10966 ) | ( ~n10961 & n10966 ) ;
  assign n10968 = ( n1827 & ~n10967 ) | ( n1827 & 1'b0 ) | ( ~n10967 & 1'b0 ) ;
  assign n10969 = n10488 | n10685 ;
  assign n10970 = ( n10475 & ~n10484 ) | ( n10475 & n10488 ) | ( ~n10484 & n10488 ) ;
  assign n10971 = ( n10484 & n10969 ) | ( n10484 & n10970 ) | ( n10969 & n10970 ) ;
  assign n10972 = ( n10488 & ~n10970 ) | ( n10488 & n10969 ) | ( ~n10970 & n10969 ) ;
  assign n10973 = ( n10475 & ~n10971 ) | ( n10475 & n10972 ) | ( ~n10971 & n10972 ) ;
  assign n10974 = ( n2033 & ~n10946 ) | ( n2033 & 1'b0 ) | ( ~n10946 & 1'b0 ) ;
  assign n10975 = ~n10960 & n10974 ;
  assign n10976 = n10966 | n10975 ;
  assign n10977 = n10954 | n10957 ;
  assign n10978 = ( n2245 & n10951 ) | ( n2245 & n10977 ) | ( n10951 & n10977 ) ;
  assign n10979 = ~n2033 & n10978 ;
  assign n10980 = n1827 | n10979 ;
  assign n10981 = ( n10976 & ~n10980 ) | ( n10976 & 1'b0 ) | ( ~n10980 & 1'b0 ) ;
  assign n10982 = ( n10973 & ~n10981 ) | ( n10973 & 1'b0 ) | ( ~n10981 & 1'b0 ) ;
  assign n10983 = n10968 | n10982 ;
  assign n10984 = ~n10490 & n10685 ;
  assign n10985 = ( n10477 & n10482 ) | ( n10477 & n10685 ) | ( n10482 & n10685 ) ;
  assign n10987 = ( n10984 & ~n10477 ) | ( n10984 & n10985 ) | ( ~n10477 & n10985 ) ;
  assign n10986 = ( n10685 & ~n10985 ) | ( n10685 & n10984 ) | ( ~n10985 & n10984 ) ;
  assign n10988 = ( n10482 & ~n10987 ) | ( n10482 & n10986 ) | ( ~n10987 & n10986 ) ;
  assign n10989 = ( n10983 & ~n1636 ) | ( n10983 & n10988 ) | ( ~n1636 & n10988 ) ;
  assign n10990 = ~n1452 & n10989 ;
  assign n10991 = n10510 | n10685 ;
  assign n10992 = ( n10497 & ~n10510 ) | ( n10497 & n10506 ) | ( ~n10510 & n10506 ) ;
  assign n10994 = ( n10510 & n10991 ) | ( n10510 & n10992 ) | ( n10991 & n10992 ) ;
  assign n10993 = ( n10506 & ~n10992 ) | ( n10506 & n10991 ) | ( ~n10992 & n10991 ) ;
  assign n10995 = ( n10497 & ~n10994 ) | ( n10497 & n10993 ) | ( ~n10994 & n10993 ) ;
  assign n10996 = ( n1636 & ~n10968 ) | ( n1636 & 1'b0 ) | ( ~n10968 & 1'b0 ) ;
  assign n10997 = ~n10982 & n10996 ;
  assign n10998 = ( n10988 & ~n10997 ) | ( n10988 & 1'b0 ) | ( ~n10997 & 1'b0 ) ;
  assign n10999 = ( n10976 & ~n10979 ) | ( n10976 & 1'b0 ) | ( ~n10979 & 1'b0 ) ;
  assign n11000 = ( n1827 & ~n10999 ) | ( n1827 & n10973 ) | ( ~n10999 & n10973 ) ;
  assign n11001 = ~n1636 & n11000 ;
  assign n11002 = ( n1452 & ~n11001 ) | ( n1452 & 1'b0 ) | ( ~n11001 & 1'b0 ) ;
  assign n11003 = ~n10998 & n11002 ;
  assign n11004 = n10995 | n11003 ;
  assign n11005 = ~n10990 & n11004 ;
  assign n11006 = n10512 &  n10685 ;
  assign n11007 = ( n10499 & ~n10685 ) | ( n10499 & n11006 ) | ( ~n10685 & n11006 ) ;
  assign n11008 = ( n10504 & ~n10499 ) | ( n10504 & n11007 ) | ( ~n10499 & n11007 ) ;
  assign n11009 = ( n10499 & ~n11007 ) | ( n10499 & n10504 ) | ( ~n11007 & n10504 ) ;
  assign n11010 = ( n11008 & ~n10504 ) | ( n11008 & n11009 ) | ( ~n10504 & n11009 ) ;
  assign n11011 = ( n1283 & ~n11005 ) | ( n1283 & n11010 ) | ( ~n11005 & n11010 ) ;
  assign n11012 = ~n1122 & n11011 ;
  assign n11013 = n10532 | n10685 ;
  assign n11014 = ( n10519 & ~n10532 ) | ( n10519 & n10528 ) | ( ~n10532 & n10528 ) ;
  assign n11016 = ( n10532 & n11013 ) | ( n10532 & n11014 ) | ( n11013 & n11014 ) ;
  assign n11015 = ( n10528 & ~n11014 ) | ( n10528 & n11013 ) | ( ~n11014 & n11013 ) ;
  assign n11017 = ( n10519 & ~n11016 ) | ( n10519 & n11015 ) | ( ~n11016 & n11015 ) ;
  assign n11018 = n1283 | n10990 ;
  assign n11019 = ( n11004 & ~n11018 ) | ( n11004 & 1'b0 ) | ( ~n11018 & 1'b0 ) ;
  assign n11020 = ( n11010 & ~n11019 ) | ( n11010 & 1'b0 ) | ( ~n11019 & 1'b0 ) ;
  assign n11021 = n10998 | n11001 ;
  assign n11022 = ( n1452 & ~n11021 ) | ( n1452 & n10995 ) | ( ~n11021 & n10995 ) ;
  assign n11023 = ( n1283 & ~n11022 ) | ( n1283 & 1'b0 ) | ( ~n11022 & 1'b0 ) ;
  assign n11024 = ( n1122 & ~n11023 ) | ( n1122 & 1'b0 ) | ( ~n11023 & 1'b0 ) ;
  assign n11025 = ~n11020 & n11024 ;
  assign n11026 = n11017 | n11025 ;
  assign n11027 = ~n11012 & n11026 ;
  assign n11028 = n10534 &  n10685 ;
  assign n11029 = ( n10521 & ~n10685 ) | ( n10521 & n11028 ) | ( ~n10685 & n11028 ) ;
  assign n11030 = ( n10521 & ~n11029 ) | ( n10521 & n10526 ) | ( ~n11029 & n10526 ) ;
  assign n11031 = ( n10526 & ~n10521 ) | ( n10526 & n11029 ) | ( ~n10521 & n11029 ) ;
  assign n11032 = ( n11030 & ~n10526 ) | ( n11030 & n11031 ) | ( ~n10526 & n11031 ) ;
  assign n11033 = ( n976 & n11027 ) | ( n976 & n11032 ) | ( n11027 & n11032 ) ;
  assign n11034 = ( n837 & ~n11033 ) | ( n837 & 1'b0 ) | ( ~n11033 & 1'b0 ) ;
  assign n11036 = ( n10550 & ~n10541 ) | ( n10550 & n10554 ) | ( ~n10541 & n10554 ) ;
  assign n11035 = ( n10554 & ~n10685 ) | ( n10554 & 1'b0 ) | ( ~n10685 & 1'b0 ) ;
  assign n11038 = ( n10554 & ~n11036 ) | ( n10554 & n11035 ) | ( ~n11036 & n11035 ) ;
  assign n11037 = ( n11035 & ~n10550 ) | ( n11035 & n11036 ) | ( ~n10550 & n11036 ) ;
  assign n11039 = ( n10541 & ~n11038 ) | ( n10541 & n11037 ) | ( ~n11038 & n11037 ) ;
  assign n11040 = ( n976 & ~n11012 ) | ( n976 & 1'b0 ) | ( ~n11012 & 1'b0 ) ;
  assign n11041 = n11026 &  n11040 ;
  assign n11042 = n11032 | n11041 ;
  assign n11043 = n11020 | n11023 ;
  assign n11044 = ( n1122 & ~n11043 ) | ( n1122 & n11017 ) | ( ~n11043 & n11017 ) ;
  assign n11045 = n976 | n11044 ;
  assign n11046 = ~n837 & n11045 ;
  assign n11047 = n11042 &  n11046 ;
  assign n11048 = ( n11039 & ~n11047 ) | ( n11039 & 1'b0 ) | ( ~n11047 & 1'b0 ) ;
  assign n11049 = n11034 | n11048 ;
  assign n11050 = n10556 &  n10685 ;
  assign n11051 = ( n10543 & ~n11050 ) | ( n10543 & n10685 ) | ( ~n11050 & n10685 ) ;
  assign n11052 = ( n10543 & ~n11051 ) | ( n10543 & n10548 ) | ( ~n11051 & n10548 ) ;
  assign n11053 = ( n10548 & ~n10543 ) | ( n10548 & n11051 ) | ( ~n10543 & n11051 ) ;
  assign n11054 = ( n11052 & ~n10548 ) | ( n11052 & n11053 ) | ( ~n10548 & n11053 ) ;
  assign n11055 = ( n713 & n11049 ) | ( n713 & n11054 ) | ( n11049 & n11054 ) ;
  assign n11056 = n595 &  n11055 ;
  assign n11058 = ( n10572 & ~n10563 ) | ( n10572 & n10576 ) | ( ~n10563 & n10576 ) ;
  assign n11057 = n10576 | n10685 ;
  assign n11060 = ( n10576 & ~n11058 ) | ( n10576 & n11057 ) | ( ~n11058 & n11057 ) ;
  assign n11059 = ( n11057 & ~n10572 ) | ( n11057 & n11058 ) | ( ~n10572 & n11058 ) ;
  assign n11061 = ( n10563 & ~n11060 ) | ( n10563 & n11059 ) | ( ~n11060 & n11059 ) ;
  assign n11062 = n713 | n11034 ;
  assign n11063 = n11048 | n11062 ;
  assign n11064 = n11054 &  n11063 ;
  assign n11065 = n11042 &  n11045 ;
  assign n11066 = ( n837 & ~n11065 ) | ( n837 & n11039 ) | ( ~n11065 & n11039 ) ;
  assign n11067 = n713 &  n11066 ;
  assign n11068 = n595 | n11067 ;
  assign n11069 = n11064 | n11068 ;
  assign n11070 = ~n11061 & n11069 ;
  assign n11071 = n11056 | n11070 ;
  assign n11072 = ~n10578 & n10685 ;
  assign n11073 = ( n10565 & ~n11072 ) | ( n10565 & n10685 ) | ( ~n11072 & n10685 ) ;
  assign n11074 = ( n10565 & ~n11073 ) | ( n10565 & n10570 ) | ( ~n11073 & n10570 ) ;
  assign n11075 = ( n10570 & ~n10565 ) | ( n10570 & n11073 ) | ( ~n10565 & n11073 ) ;
  assign n11076 = ( n11074 & ~n10570 ) | ( n11074 & n11075 ) | ( ~n10570 & n11075 ) ;
  assign n11077 = ( n492 & n11071 ) | ( n492 & n11076 ) | ( n11071 & n11076 ) ;
  assign n11078 = n396 &  n11077 ;
  assign n11079 = n10598 | n10685 ;
  assign n11080 = ( n10585 & n10594 ) | ( n10585 & n10598 ) | ( n10594 & n10598 ) ;
  assign n11081 = ( n11079 & ~n10594 ) | ( n11079 & n11080 ) | ( ~n10594 & n11080 ) ;
  assign n11082 = ( n10598 & ~n11080 ) | ( n10598 & n11079 ) | ( ~n11080 & n11079 ) ;
  assign n11083 = ( n10585 & ~n11081 ) | ( n10585 & n11082 ) | ( ~n11081 & n11082 ) ;
  assign n11084 = n492 | n11056 ;
  assign n11085 = n11070 | n11084 ;
  assign n11086 = n11076 &  n11085 ;
  assign n11087 = n11064 | n11067 ;
  assign n11088 = ( n595 & ~n11061 ) | ( n595 & n11087 ) | ( ~n11061 & n11087 ) ;
  assign n11089 = n492 &  n11088 ;
  assign n11090 = n396 | n11089 ;
  assign n11091 = n11086 | n11090 ;
  assign n11092 = n11083 &  n11091 ;
  assign n11093 = n11078 | n11092 ;
  assign n11099 = ( n315 & ~n11098 ) | ( n315 & n11093 ) | ( ~n11098 & n11093 ) ;
  assign n11100 = n240 &  n11099 ;
  assign n11101 = n10620 | n10685 ;
  assign n11102 = ( n10607 & n10616 ) | ( n10607 & n10620 ) | ( n10616 & n10620 ) ;
  assign n11103 = ( n11101 & ~n10616 ) | ( n11101 & n11102 ) | ( ~n10616 & n11102 ) ;
  assign n11104 = ( n10620 & ~n11102 ) | ( n10620 & n11101 ) | ( ~n11102 & n11101 ) ;
  assign n11105 = ( n10607 & ~n11103 ) | ( n10607 & n11104 ) | ( ~n11103 & n11104 ) ;
  assign n11106 = n315 | n11078 ;
  assign n11107 = n11092 | n11106 ;
  assign n11108 = ~n11098 & n11107 ;
  assign n11109 = n11086 | n11089 ;
  assign n11110 = ( n396 & n11083 ) | ( n396 & n11109 ) | ( n11083 & n11109 ) ;
  assign n11111 = n315 &  n11110 ;
  assign n11112 = n240 | n11111 ;
  assign n11113 = n11108 | n11112 ;
  assign n11114 = n11105 &  n11113 ;
  assign n11115 = n11100 | n11114 ;
  assign n11121 = ( n181 & ~n11120 ) | ( n181 & n11115 ) | ( ~n11120 & n11115 ) ;
  assign n11122 = ~n145 & n11121 ;
  assign n11124 = ( n10638 & ~n10629 ) | ( n10638 & n10642 ) | ( ~n10629 & n10642 ) ;
  assign n11123 = n10642 | n10685 ;
  assign n11126 = ( n10642 & ~n11124 ) | ( n10642 & n11123 ) | ( ~n11124 & n11123 ) ;
  assign n11125 = ( n11123 & ~n10638 ) | ( n11123 & n11124 ) | ( ~n10638 & n11124 ) ;
  assign n11127 = ( n10629 & ~n11126 ) | ( n10629 & n11125 ) | ( ~n11126 & n11125 ) ;
  assign n11128 = n181 | n11100 ;
  assign n11129 = n11114 | n11128 ;
  assign n11130 = ~n11120 & n11129 ;
  assign n11131 = n11108 | n11111 ;
  assign n11132 = ( n240 & n11105 ) | ( n240 & n11131 ) | ( n11105 & n11131 ) ;
  assign n11133 = n181 &  n11132 ;
  assign n11134 = ( n145 & ~n11133 ) | ( n145 & 1'b0 ) | ( ~n11133 & 1'b0 ) ;
  assign n11135 = ~n11130 & n11134 ;
  assign n11136 = ( n11127 & ~n11135 ) | ( n11127 & 1'b0 ) | ( ~n11135 & 1'b0 ) ;
  assign n11137 = n11122 | n11136 ;
  assign n11138 = n10631 | n10685 ;
  assign n11139 = ( n10636 & ~n10631 ) | ( n10636 & n10644 ) | ( ~n10631 & n10644 ) ;
  assign n11141 = ( n10631 & n11138 ) | ( n10631 & n11139 ) | ( n11138 & n11139 ) ;
  assign n11140 = ( n10644 & ~n11139 ) | ( n10644 & n11138 ) | ( ~n11139 & n11138 ) ;
  assign n11142 = ( n10636 & ~n11141 ) | ( n10636 & n11140 ) | ( ~n11141 & n11140 ) ;
  assign n11143 = ( n150 & n11137 ) | ( n150 & n11142 ) | ( n11137 & n11142 ) ;
  assign n11155 = n11143 | n11154 ;
  assign n11156 = ( n133 & ~n11154 ) | ( n133 & n11155 ) | ( ~n11154 & n11155 ) ;
  assign n11159 = n11130 | n11133 ;
  assign n11160 = ( n11127 & ~n145 ) | ( n11127 & n11159 ) | ( ~n145 & n11159 ) ;
  assign n11161 = n150 &  n11160 ;
  assign n11162 = ( n11150 & ~n11161 ) | ( n11150 & 1'b0 ) | ( ~n11161 & 1'b0 ) ;
  assign n11157 = n150 | n11122 ;
  assign n11158 = n11136 | n11157 ;
  assign n11163 = ( n11142 & ~n11158 ) | ( n11142 & 1'b0 ) | ( ~n11158 & 1'b0 ) ;
  assign n11164 = ( n11162 & ~n11142 ) | ( n11162 & n11163 ) | ( ~n11142 & n11163 ) ;
  assign n11166 = ( n133 & ~n10659 ) | ( n133 & n10652 ) | ( ~n10659 & n10652 ) ;
  assign n11165 = ( n10659 & ~n10652 ) | ( n10659 & n10685 ) | ( ~n10652 & n10685 ) ;
  assign n11167 = ~n10659 & n11165 ;
  assign n11168 = ( n10659 & n11166 ) | ( n10659 & n11167 ) | ( n11166 & n11167 ) ;
  assign n11169 = n10655 | n10682 ;
  assign n11170 = ( n10658 & n10677 ) | ( n10658 & n11169 ) | ( n10677 & n11169 ) ;
  assign n11171 = ( n10658 & ~n11170 ) | ( n10658 & 1'b0 ) | ( ~n11170 & 1'b0 ) ;
  assign n11172 = ( n10665 & ~n11171 ) | ( n10665 & n10673 ) | ( ~n11171 & n10673 ) ;
  assign n11173 = ( n10665 & ~n11172 ) | ( n10665 & 1'b0 ) | ( ~n11172 & 1'b0 ) ;
  assign n11174 = n11168 | n11173 ;
  assign n11175 = n11164 | n11174 ;
  assign n11176 = ~n11156 |  n11175 ;
  assign n11424 = n10936 | n11176 ;
  assign n11425 = ( n10923 & n10932 ) | ( n10923 & n10936 ) | ( n10932 & n10936 ) ;
  assign n11426 = ( n11424 & ~n10932 ) | ( n11424 & n11425 ) | ( ~n10932 & n11425 ) ;
  assign n11427 = ( n10936 & ~n11425 ) | ( n10936 & n11424 ) | ( ~n11425 & n11424 ) ;
  assign n11428 = ( n10923 & ~n11426 ) | ( n10923 & n11427 ) | ( ~n11426 & n11427 ) ;
  assign n11418 = ( n10903 & ~n10908 ) | ( n10903 & n11176 ) | ( ~n10908 & n11176 ) ;
  assign n11417 = ~n10916 & n11176 ;
  assign n11419 = ( n11176 & ~n11418 ) | ( n11176 & n11417 ) | ( ~n11418 & n11417 ) ;
  assign n11420 = ( n11417 & ~n10903 ) | ( n11417 & n11418 ) | ( ~n10903 & n11418 ) ;
  assign n11421 = ( n10908 & ~n11419 ) | ( n10908 & n11420 ) | ( ~n11419 & n11420 ) ;
  assign n11403 = ( n10910 & ~n10901 ) | ( n10910 & n10914 ) | ( ~n10901 & n10914 ) ;
  assign n11402 = n10914 | n11176 ;
  assign n11405 = ( n10914 & ~n11403 ) | ( n10914 & n11402 ) | ( ~n11403 & n11402 ) ;
  assign n11404 = ( n11402 & ~n10910 ) | ( n11402 & n11403 ) | ( ~n10910 & n11403 ) ;
  assign n11406 = ( n10901 & ~n11405 ) | ( n10901 & n11404 ) | ( ~n11405 & n11404 ) ;
  assign n11396 = ( n10881 & ~n10886 ) | ( n10881 & n11176 ) | ( ~n10886 & n11176 ) ;
  assign n11395 = ~n10894 & n11176 ;
  assign n11397 = ( n11176 & ~n11396 ) | ( n11176 & n11395 ) | ( ~n11396 & n11395 ) ;
  assign n11398 = ( n11395 & ~n10881 ) | ( n11395 & n11396 ) | ( ~n10881 & n11396 ) ;
  assign n11399 = ( n10886 & ~n11397 ) | ( n10886 & n11398 ) | ( ~n11397 & n11398 ) ;
  assign n11381 = ( n10888 & ~n10879 ) | ( n10888 & n10892 ) | ( ~n10879 & n10892 ) ;
  assign n11380 = n10892 | n11176 ;
  assign n11383 = ( n10892 & ~n11381 ) | ( n10892 & n11380 ) | ( ~n11381 & n11380 ) ;
  assign n11382 = ( n11380 & ~n10888 ) | ( n11380 & n11381 ) | ( ~n10888 & n11381 ) ;
  assign n11384 = ( n10879 & ~n11383 ) | ( n10879 & n11382 ) | ( ~n11383 & n11382 ) ;
  assign n11374 = ( n10859 & ~n10864 ) | ( n10859 & n11176 ) | ( ~n10864 & n11176 ) ;
  assign n11373 = ~n10872 & n11176 ;
  assign n11375 = ( n11176 & ~n11374 ) | ( n11176 & n11373 ) | ( ~n11374 & n11373 ) ;
  assign n11376 = ( n11373 & ~n10859 ) | ( n11373 & n11374 ) | ( ~n10859 & n11374 ) ;
  assign n11377 = ( n10864 & ~n11375 ) | ( n10864 & n11376 ) | ( ~n11375 & n11376 ) ;
  assign n11358 = n10870 | n11176 ;
  assign n11359 = ( n10857 & n10866 ) | ( n10857 & n10870 ) | ( n10866 & n10870 ) ;
  assign n11360 = ( n11358 & ~n10866 ) | ( n11358 & n11359 ) | ( ~n10866 & n11359 ) ;
  assign n11361 = ( n10870 & ~n11359 ) | ( n10870 & n11358 ) | ( ~n11359 & n11358 ) ;
  assign n11362 = ( n10857 & ~n11360 ) | ( n10857 & n11361 ) | ( ~n11360 & n11361 ) ;
  assign n11351 = n10850 &  n11176 ;
  assign n11352 = ( n10837 & n10842 ) | ( n10837 & n11176 ) | ( n10842 & n11176 ) ;
  assign n11354 = ( n11351 & ~n10837 ) | ( n11351 & n11352 ) | ( ~n10837 & n11352 ) ;
  assign n11353 = ( n11176 & ~n11352 ) | ( n11176 & n11351 ) | ( ~n11352 & n11351 ) ;
  assign n11355 = ( n10842 & ~n11354 ) | ( n10842 & n11353 ) | ( ~n11354 & n11353 ) ;
  assign n11336 = n10848 | n11176 ;
  assign n11337 = ( n10835 & ~n10848 ) | ( n10835 & n10844 ) | ( ~n10848 & n10844 ) ;
  assign n11339 = ( n10848 & n11336 ) | ( n10848 & n11337 ) | ( n11336 & n11337 ) ;
  assign n11338 = ( n10844 & ~n11337 ) | ( n10844 & n11336 ) | ( ~n11337 & n11336 ) ;
  assign n11340 = ( n10835 & ~n11339 ) | ( n10835 & n11338 ) | ( ~n11339 & n11338 ) ;
  assign n11330 = ( n10815 & ~n10820 ) | ( n10815 & n10828 ) | ( ~n10820 & n10828 ) ;
  assign n11329 = ( n10815 & ~n11176 ) | ( n10815 & 1'b0 ) | ( ~n11176 & 1'b0 ) ;
  assign n11332 = ( n10815 & ~n11330 ) | ( n10815 & n11329 ) | ( ~n11330 & n11329 ) ;
  assign n11331 = ( n11329 & ~n10828 ) | ( n11329 & n11330 ) | ( ~n10828 & n11330 ) ;
  assign n11333 = ( n10820 & ~n11332 ) | ( n10820 & n11331 ) | ( ~n11332 & n11331 ) ;
  assign n11314 = n10826 | n11176 ;
  assign n11315 = ( n10813 & ~n10822 ) | ( n10813 & n10826 ) | ( ~n10822 & n10826 ) ;
  assign n11316 = ( n10822 & n11314 ) | ( n10822 & n11315 ) | ( n11314 & n11315 ) ;
  assign n11317 = ( n10826 & ~n11315 ) | ( n10826 & n11314 ) | ( ~n11315 & n11314 ) ;
  assign n11318 = ( n10813 & ~n11316 ) | ( n10813 & n11317 ) | ( ~n11316 & n11317 ) ;
  assign n11307 = n10793 | n11176 ;
  assign n11308 = ( n10798 & ~n10793 ) | ( n10798 & n10806 ) | ( ~n10793 & n10806 ) ;
  assign n11310 = ( n10793 & n11307 ) | ( n10793 & n11308 ) | ( n11307 & n11308 ) ;
  assign n11309 = ( n10806 & ~n11308 ) | ( n10806 & n11307 ) | ( ~n11308 & n11307 ) ;
  assign n11311 = ( n10798 & ~n11310 ) | ( n10798 & n11309 ) | ( ~n11310 & n11309 ) ;
  assign n11293 = ( n10800 & ~n10791 ) | ( n10800 & n10804 ) | ( ~n10791 & n10804 ) ;
  assign n11292 = n10804 | n11176 ;
  assign n11295 = ( n10804 & ~n11293 ) | ( n10804 & n11292 ) | ( ~n11293 & n11292 ) ;
  assign n11294 = ( n11292 & ~n10800 ) | ( n11292 & n11293 ) | ( ~n10800 & n11293 ) ;
  assign n11296 = ( n10791 & ~n11295 ) | ( n10791 & n11294 ) | ( ~n11295 & n11294 ) ;
  assign n11285 = n10771 | n11176 ;
  assign n11286 = ( n10771 & ~n10784 ) | ( n10771 & n10776 ) | ( ~n10784 & n10776 ) ;
  assign n11287 = ( n10784 & n11285 ) | ( n10784 & n11286 ) | ( n11285 & n11286 ) ;
  assign n11288 = ( n10771 & ~n11286 ) | ( n10771 & n11285 ) | ( ~n11286 & n11285 ) ;
  assign n11289 = ( n10776 & ~n11287 ) | ( n10776 & n11288 ) | ( ~n11287 & n11288 ) ;
  assign n11270 = n10782 | n11176 ;
  assign n11271 = ( n10769 & ~n10782 ) | ( n10769 & n10778 ) | ( ~n10782 & n10778 ) ;
  assign n11273 = ( n10782 & n11270 ) | ( n10782 & n11271 ) | ( n11270 & n11271 ) ;
  assign n11272 = ( n10778 & ~n11271 ) | ( n10778 & n11270 ) | ( ~n11271 & n11270 ) ;
  assign n11274 = ( n10769 & ~n11273 ) | ( n10769 & n11272 ) | ( ~n11273 & n11272 ) ;
  assign n11263 = n10749 | n11176 ;
  assign n11264 = ( n10749 & n10754 ) | ( n10749 & n10762 ) | ( n10754 & n10762 ) ;
  assign n11265 = ( n11263 & ~n10762 ) | ( n11263 & n11264 ) | ( ~n10762 & n11264 ) ;
  assign n11266 = ( n10749 & ~n11264 ) | ( n10749 & n11263 ) | ( ~n11264 & n11263 ) ;
  assign n11267 = ( n10754 & ~n11265 ) | ( n10754 & n11266 ) | ( ~n11265 & n11266 ) ;
  assign n11248 = n10760 | n11176 ;
  assign n11249 = ( n10747 & ~n10760 ) | ( n10747 & n10756 ) | ( ~n10760 & n10756 ) ;
  assign n11251 = ( n10760 & n11248 ) | ( n10760 & n11249 ) | ( n11248 & n11249 ) ;
  assign n11250 = ( n10756 & ~n11249 ) | ( n10756 & n11248 ) | ( ~n11249 & n11248 ) ;
  assign n11252 = ( n10747 & ~n11251 ) | ( n10747 & n11250 ) | ( ~n11251 & n11250 ) ;
  assign n11241 = n10727 | n11176 ;
  assign n11242 = ( n10732 & ~n10727 ) | ( n10732 & n10740 ) | ( ~n10727 & n10740 ) ;
  assign n11244 = ( n10727 & n11241 ) | ( n10727 & n11242 ) | ( n11241 & n11242 ) ;
  assign n11243 = ( n10740 & ~n11242 ) | ( n10740 & n11241 ) | ( ~n11242 & n11241 ) ;
  assign n11245 = ( n10732 & ~n11244 ) | ( n10732 & n11243 ) | ( ~n11244 & n11243 ) ;
  assign n11226 = n10738 | n11176 ;
  assign n11227 = ( n10725 & ~n10734 ) | ( n10725 & n10738 ) | ( ~n10734 & n10738 ) ;
  assign n11228 = ( n10734 & n11226 ) | ( n10734 & n11227 ) | ( n11226 & n11227 ) ;
  assign n11229 = ( n10738 & ~n11227 ) | ( n10738 & n11226 ) | ( ~n11227 & n11226 ) ;
  assign n11230 = ( n10725 & ~n11228 ) | ( n10725 & n11229 ) | ( ~n11228 & n11229 ) ;
  assign n11219 = n10701 | n10703 ;
  assign n11220 = ( n10703 & n10713 ) | ( n10703 & n11219 ) | ( n10713 & n11219 ) ;
  assign n11222 = ( n11176 & ~n11219 ) | ( n11176 & n11220 ) | ( ~n11219 & n11220 ) ;
  assign n11221 = ( n10703 & ~n11220 ) | ( n10703 & n11176 ) | ( ~n11220 & n11176 ) ;
  assign n11223 = ( n10713 & ~n11222 ) | ( n10713 & n11221 ) | ( ~n11222 & n11221 ) ;
  assign n11203 = ~x42 & n10685 ;
  assign n11204 = ( x43 & ~n11203 ) | ( x43 & 1'b0 ) | ( ~n11203 & 1'b0 ) ;
  assign n11205 = n10704 | n11204 ;
  assign n11200 = ( n10685 & ~x42 ) | ( n10685 & n10696 ) | ( ~x42 & n10696 ) ;
  assign n11201 = x42 &  n11200 ;
  assign n11202 = ( n10691 & ~n11201 ) | ( n10691 & n10696 ) | ( ~n11201 & n10696 ) ;
  assign n11206 = ( n11176 & ~n11205 ) | ( n11176 & n11202 ) | ( ~n11205 & n11202 ) ;
  assign n11208 = ( n11176 & ~n11206 ) | ( n11176 & 1'b0 ) | ( ~n11206 & 1'b0 ) ;
  assign n11207 = ~n11202 & n11206 ;
  assign n11209 = ( n11205 & ~n11208 ) | ( n11205 & n11207 ) | ( ~n11208 & n11207 ) ;
  assign n11189 = ( n10685 & ~n11173 ) | ( n10685 & 1'b0 ) | ( ~n11173 & 1'b0 ) ;
  assign n11190 = ( n11164 & ~n11168 ) | ( n11164 & n11189 ) | ( ~n11168 & n11189 ) ;
  assign n11191 = ~n11164 & n11190 ;
  assign n11192 = n11156 &  n11191 ;
  assign n11188 = ~n10688 & n11176 ;
  assign n11193 = ( n11188 & ~n11192 ) | ( n11188 & 1'b0 ) | ( ~n11192 & 1'b0 ) ;
  assign n11194 = ( x42 & n11192 ) | ( x42 & n11193 ) | ( n11192 & n11193 ) ;
  assign n11195 = x42 | n11192 ;
  assign n11196 = n11188 | n11195 ;
  assign n11197 = ~n11194 & n11196 ;
  assign n11179 = ( x40 & ~n11176 ) | ( x40 & x41 ) | ( ~n11176 & x41 ) ;
  assign n11185 = ( x40 & ~x41 ) | ( x40 & 1'b0 ) | ( ~x41 & 1'b0 ) ;
  assign n10686 = x38 | x39 ;
  assign n11180 = ~x40 & n10686 ;
  assign n11181 = ( x40 & ~n10683 ) | ( x40 & n11180 ) | ( ~n10683 & n11180 ) ;
  assign n11182 = ( n10665 & ~n11181 ) | ( n10665 & n10673 ) | ( ~n11181 & n10673 ) ;
  assign n11183 = ( n10665 & ~n11182 ) | ( n10665 & 1'b0 ) | ( ~n11182 & 1'b0 ) ;
  assign n11184 = ( n11176 & ~x41 ) | ( n11176 & n11183 ) | ( ~x41 & n11183 ) ;
  assign n11186 = ( n11179 & ~n11185 ) | ( n11179 & n11184 ) | ( ~n11185 & n11184 ) ;
  assign n10687 = x40 | n10686 ;
  assign n11177 = x40 &  n11176 ;
  assign n11178 = ( n10685 & ~n10687 ) | ( n10685 & n11177 ) | ( ~n10687 & n11177 ) ;
  assign n11210 = n10209 | n11178 ;
  assign n11211 = ( n11186 & ~n11210 ) | ( n11186 & 1'b0 ) | ( ~n11210 & 1'b0 ) ;
  assign n11212 = n11197 | n11211 ;
  assign n11213 = n11178 &  n11186 ;
  assign n11214 = ( n10209 & ~n11186 ) | ( n10209 & n11213 ) | ( ~n11186 & n11213 ) ;
  assign n11215 = ( n9740 & ~n11214 ) | ( n9740 & 1'b0 ) | ( ~n11214 & 1'b0 ) ;
  assign n11216 = n11212 &  n11215 ;
  assign n11217 = n11209 | n11216 ;
  assign n11187 = ~n11178 & n11186 ;
  assign n11198 = ( n11187 & ~n10209 ) | ( n11187 & n11197 ) | ( ~n10209 & n11197 ) ;
  assign n11199 = n9740 | n11198 ;
  assign n11231 = ~n9286 & n11199 ;
  assign n11232 = n11217 &  n11231 ;
  assign n11233 = n11223 | n11232 ;
  assign n11234 = ( n11212 & ~n11214 ) | ( n11212 & 1'b0 ) | ( ~n11214 & 1'b0 ) ;
  assign n11235 = ( n9740 & n11209 ) | ( n9740 & n11234 ) | ( n11209 & n11234 ) ;
  assign n11236 = ( n9286 & ~n11235 ) | ( n9286 & 1'b0 ) | ( ~n11235 & 1'b0 ) ;
  assign n11237 = n8839 | n11236 ;
  assign n11238 = ( n11233 & ~n11237 ) | ( n11233 & 1'b0 ) | ( ~n11237 & 1'b0 ) ;
  assign n11239 = n11230 | n11238 ;
  assign n11218 = n11199 &  n11217 ;
  assign n11224 = ( n11218 & ~n9286 ) | ( n11218 & n11223 ) | ( ~n9286 & n11223 ) ;
  assign n11225 = ( n8839 & ~n11224 ) | ( n8839 & 1'b0 ) | ( ~n11224 & 1'b0 ) ;
  assign n11253 = n8407 | n11225 ;
  assign n11254 = ( n11239 & ~n11253 ) | ( n11239 & 1'b0 ) | ( ~n11253 & 1'b0 ) ;
  assign n11255 = n11245 | n11254 ;
  assign n11256 = ( n11233 & ~n11236 ) | ( n11233 & 1'b0 ) | ( ~n11236 & 1'b0 ) ;
  assign n11257 = ( n11230 & ~n8839 ) | ( n11230 & n11256 ) | ( ~n8839 & n11256 ) ;
  assign n11258 = ( n8407 & ~n11257 ) | ( n8407 & 1'b0 ) | ( ~n11257 & 1'b0 ) ;
  assign n11259 = n7982 | n11258 ;
  assign n11260 = ( n11255 & ~n11259 ) | ( n11255 & 1'b0 ) | ( ~n11259 & 1'b0 ) ;
  assign n11261 = ( n11252 & ~n11260 ) | ( n11252 & 1'b0 ) | ( ~n11260 & 1'b0 ) ;
  assign n11240 = ~n11225 & n11239 ;
  assign n11246 = ( n11240 & ~n8407 ) | ( n11240 & n11245 ) | ( ~n8407 & n11245 ) ;
  assign n11247 = ( n7982 & ~n11246 ) | ( n7982 & 1'b0 ) | ( ~n11246 & 1'b0 ) ;
  assign n11275 = ( n7572 & ~n11247 ) | ( n7572 & 1'b0 ) | ( ~n11247 & 1'b0 ) ;
  assign n11276 = ~n11261 & n11275 ;
  assign n11277 = ( n11267 & ~n11276 ) | ( n11267 & 1'b0 ) | ( ~n11276 & 1'b0 ) ;
  assign n11278 = ( n11255 & ~n11258 ) | ( n11255 & 1'b0 ) | ( ~n11258 & 1'b0 ) ;
  assign n11279 = ( n7982 & ~n11278 ) | ( n7982 & n11252 ) | ( ~n11278 & n11252 ) ;
  assign n11280 = ~n7572 & n11279 ;
  assign n11281 = ( n7169 & ~n11280 ) | ( n7169 & 1'b0 ) | ( ~n11280 & 1'b0 ) ;
  assign n11282 = ~n11277 & n11281 ;
  assign n11283 = ( n11274 & ~n11282 ) | ( n11274 & 1'b0 ) | ( ~n11282 & 1'b0 ) ;
  assign n11262 = n11247 | n11261 ;
  assign n11268 = ( n11262 & ~n7572 ) | ( n11262 & n11267 ) | ( ~n7572 & n11267 ) ;
  assign n11269 = ~n7169 & n11268 ;
  assign n11297 = n6781 | n11269 ;
  assign n11298 = n11283 | n11297 ;
  assign n11299 = n11289 &  n11298 ;
  assign n11300 = n11277 | n11280 ;
  assign n11301 = ( n11274 & ~n7169 ) | ( n11274 & n11300 ) | ( ~n7169 & n11300 ) ;
  assign n11302 = n6781 &  n11301 ;
  assign n11303 = ( n6399 & ~n11302 ) | ( n6399 & 1'b0 ) | ( ~n11302 & 1'b0 ) ;
  assign n11304 = ~n11299 & n11303 ;
  assign n11305 = ( n11296 & ~n11304 ) | ( n11296 & 1'b0 ) | ( ~n11304 & 1'b0 ) ;
  assign n11284 = n11269 | n11283 ;
  assign n11290 = ( n6781 & n11284 ) | ( n6781 & n11289 ) | ( n11284 & n11289 ) ;
  assign n11291 = ~n6399 & n11290 ;
  assign n11319 = n6032 | n11291 ;
  assign n11320 = n11305 | n11319 ;
  assign n11321 = ~n11311 & n11320 ;
  assign n11322 = n11299 | n11302 ;
  assign n11323 = ( n11296 & ~n6399 ) | ( n11296 & n11322 ) | ( ~n6399 & n11322 ) ;
  assign n11324 = n6032 &  n11323 ;
  assign n11325 = ( n5672 & ~n11324 ) | ( n5672 & 1'b0 ) | ( ~n11324 & 1'b0 ) ;
  assign n11326 = ~n11321 & n11325 ;
  assign n11327 = n11318 | n11326 ;
  assign n11306 = n11291 | n11305 ;
  assign n11312 = ( n6032 & ~n11311 ) | ( n6032 & n11306 ) | ( ~n11311 & n11306 ) ;
  assign n11313 = ~n5672 & n11312 ;
  assign n11341 = n5327 | n11313 ;
  assign n11342 = ( n11327 & ~n11341 ) | ( n11327 & 1'b0 ) | ( ~n11341 & 1'b0 ) ;
  assign n11343 = ( n11333 & ~n11342 ) | ( n11333 & 1'b0 ) | ( ~n11342 & 1'b0 ) ;
  assign n11344 = n11321 | n11324 ;
  assign n11345 = ( n5672 & ~n11344 ) | ( n5672 & n11318 ) | ( ~n11344 & n11318 ) ;
  assign n11346 = ( n5327 & ~n11345 ) | ( n5327 & 1'b0 ) | ( ~n11345 & 1'b0 ) ;
  assign n11347 = n4990 | n11346 ;
  assign n11348 = n11343 | n11347 ;
  assign n11349 = ~n11340 & n11348 ;
  assign n11328 = ~n11313 & n11327 ;
  assign n11334 = ( n5327 & ~n11328 ) | ( n5327 & n11333 ) | ( ~n11328 & n11333 ) ;
  assign n11335 = n4990 &  n11334 ;
  assign n11363 = n4668 | n11335 ;
  assign n11364 = n11349 | n11363 ;
  assign n11365 = n11355 &  n11364 ;
  assign n11366 = n11343 | n11346 ;
  assign n11367 = ( n4990 & ~n11340 ) | ( n4990 & n11366 ) | ( ~n11340 & n11366 ) ;
  assign n11368 = n4668 &  n11367 ;
  assign n11369 = n4353 | n11368 ;
  assign n11370 = n11365 | n11369 ;
  assign n11371 = n11362 &  n11370 ;
  assign n11350 = n11335 | n11349 ;
  assign n11356 = ( n4668 & n11350 ) | ( n4668 & n11355 ) | ( n11350 & n11355 ) ;
  assign n11357 = n4353 &  n11356 ;
  assign n11385 = n4053 | n11357 ;
  assign n11386 = n11371 | n11385 ;
  assign n11387 = ~n11377 & n11386 ;
  assign n11388 = n11365 | n11368 ;
  assign n11389 = ( n4353 & n11362 ) | ( n4353 & n11388 ) | ( n11362 & n11388 ) ;
  assign n11390 = n4053 &  n11389 ;
  assign n11391 = n3760 | n11390 ;
  assign n11392 = n11387 | n11391 ;
  assign n11393 = ~n11384 & n11392 ;
  assign n11372 = n11357 | n11371 ;
  assign n11378 = ( n4053 & ~n11377 ) | ( n4053 & n11372 ) | ( ~n11377 & n11372 ) ;
  assign n11379 = n3760 &  n11378 ;
  assign n11407 = n3482 | n11379 ;
  assign n11408 = n11393 | n11407 ;
  assign n11409 = ~n11399 & n11408 ;
  assign n11410 = n11387 | n11390 ;
  assign n11411 = ( n3760 & ~n11384 ) | ( n3760 & n11410 ) | ( ~n11384 & n11410 ) ;
  assign n11412 = n3482 &  n11411 ;
  assign n11413 = n3211 | n11412 ;
  assign n11414 = n11409 | n11413 ;
  assign n11415 = ~n11406 & n11414 ;
  assign n11394 = n11379 | n11393 ;
  assign n11400 = ( n3482 & ~n11399 ) | ( n3482 & n11394 ) | ( ~n11399 & n11394 ) ;
  assign n11401 = n3211 &  n11400 ;
  assign n11429 = n2955 | n11401 ;
  assign n11430 = n11415 | n11429 ;
  assign n11431 = ~n11421 & n11430 ;
  assign n11432 = n11409 | n11412 ;
  assign n11433 = ( n3211 & ~n11406 ) | ( n3211 & n11432 ) | ( ~n11406 & n11432 ) ;
  assign n11434 = n2955 &  n11433 ;
  assign n11435 = n2706 | n11434 ;
  assign n11436 = n11431 | n11435 ;
  assign n11571 = ( n11056 & ~n11061 ) | ( n11056 & n11176 ) | ( ~n11061 & n11176 ) ;
  assign n11570 = ~n11069 & n11176 ;
  assign n11572 = ( n11176 & ~n11571 ) | ( n11176 & n11570 ) | ( ~n11571 & n11570 ) ;
  assign n11573 = ( n11570 & ~n11056 ) | ( n11570 & n11571 ) | ( ~n11056 & n11571 ) ;
  assign n11574 = ( n11061 & ~n11572 ) | ( n11061 & n11573 ) | ( ~n11572 & n11573 ) ;
  assign n11504 = n11003 &  n11176 ;
  assign n11505 = ( n10990 & ~n11504 ) | ( n10990 & n11176 ) | ( ~n11504 & n11176 ) ;
  assign n11506 = ( n10995 & ~n10990 ) | ( n10995 & n11505 ) | ( ~n10990 & n11505 ) ;
  assign n11507 = ( n10990 & ~n11505 ) | ( n10990 & n10995 ) | ( ~n11505 & n10995 ) ;
  assign n11508 = ( n11506 & ~n10995 ) | ( n11506 & n11507 ) | ( ~n10995 & n11507 ) ;
  assign n11439 = ~n10938 & n11176 ;
  assign n11440 = ( n10925 & n10930 ) | ( n10925 & n11176 ) | ( n10930 & n11176 ) ;
  assign n11442 = ( n11439 & ~n10925 ) | ( n11439 & n11440 ) | ( ~n10925 & n11440 ) ;
  assign n11441 = ( n11176 & ~n11440 ) | ( n11176 & n11439 ) | ( ~n11440 & n11439 ) ;
  assign n11443 = ( n10930 & ~n11442 ) | ( n10930 & n11441 ) | ( ~n11442 & n11441 ) ;
  assign n11416 = n11401 | n11415 ;
  assign n11422 = ( n2955 & ~n11421 ) | ( n2955 & n11416 ) | ( ~n11421 & n11416 ) ;
  assign n11423 = n2706 &  n11422 ;
  assign n11437 = n11428 &  n11436 ;
  assign n11438 = n11423 | n11437 ;
  assign n11444 = ( n2472 & ~n11443 ) | ( n2472 & n11438 ) | ( ~n11443 & n11438 ) ;
  assign n11445 = n2245 &  n11444 ;
  assign n11446 = n2472 | n11423 ;
  assign n11447 = n11437 | n11446 ;
  assign n11448 = ~n11443 & n11447 ;
  assign n11449 = n11431 | n11434 ;
  assign n11450 = ( n2706 & n11428 ) | ( n2706 & n11449 ) | ( n11428 & n11449 ) ;
  assign n11451 = n2472 &  n11450 ;
  assign n11452 = n2245 | n11451 ;
  assign n11453 = n11448 | n11452 ;
  assign n11454 = ( n10953 & ~n11176 ) | ( n10953 & n10957 ) | ( ~n11176 & n10957 ) ;
  assign n11455 = ( n10944 & ~n11454 ) | ( n10944 & n10953 ) | ( ~n11454 & n10953 ) ;
  assign n11456 = ( n10944 & ~n10953 ) | ( n10944 & n11454 ) | ( ~n10953 & n11454 ) ;
  assign n11457 = ( n11455 & ~n10944 ) | ( n11455 & n11456 ) | ( ~n10944 & n11456 ) ;
  assign n11458 = ( n11453 & ~n11457 ) | ( n11453 & 1'b0 ) | ( ~n11457 & 1'b0 ) ;
  assign n11459 = n11445 | n11458 ;
  assign n11460 = ~n10959 & n11176 ;
  assign n11461 = ( n10946 & n10951 ) | ( n10946 & n11176 ) | ( n10951 & n11176 ) ;
  assign n11463 = ( n11460 & ~n10946 ) | ( n11460 & n11461 ) | ( ~n10946 & n11461 ) ;
  assign n11462 = ( n11176 & ~n11461 ) | ( n11176 & n11460 ) | ( ~n11461 & n11460 ) ;
  assign n11464 = ( n10951 & ~n11463 ) | ( n10951 & n11462 ) | ( ~n11463 & n11462 ) ;
  assign n11465 = ( n11459 & ~n2033 ) | ( n11459 & n11464 ) | ( ~n2033 & n11464 ) ;
  assign n11466 = n1827 &  n11465 ;
  assign n11467 = n10979 | n11176 ;
  assign n11468 = ( n10966 & ~n10979 ) | ( n10966 & n10975 ) | ( ~n10979 & n10975 ) ;
  assign n11470 = ( n10979 & n11467 ) | ( n10979 & n11468 ) | ( n11467 & n11468 ) ;
  assign n11469 = ( n10975 & ~n11468 ) | ( n10975 & n11467 ) | ( ~n11468 & n11467 ) ;
  assign n11471 = ( n10966 & ~n11470 ) | ( n10966 & n11469 ) | ( ~n11470 & n11469 ) ;
  assign n11472 = ( n2033 & ~n11445 ) | ( n2033 & 1'b0 ) | ( ~n11445 & 1'b0 ) ;
  assign n11473 = ~n11458 & n11472 ;
  assign n11474 = ( n11464 & ~n11473 ) | ( n11464 & 1'b0 ) | ( ~n11473 & 1'b0 ) ;
  assign n11475 = n11448 | n11451 ;
  assign n11476 = ( n2245 & ~n11457 ) | ( n2245 & n11475 ) | ( ~n11457 & n11475 ) ;
  assign n11477 = ~n2033 & n11476 ;
  assign n11478 = n1827 | n11477 ;
  assign n11479 = n11474 | n11478 ;
  assign n11480 = ~n11471 & n11479 ;
  assign n11481 = n11466 | n11480 ;
  assign n11483 = ( n10968 & ~n10973 ) | ( n10968 & n11176 ) | ( ~n10973 & n11176 ) ;
  assign n11482 = n10981 &  n11176 ;
  assign n11484 = ( n11176 & ~n11483 ) | ( n11176 & n11482 ) | ( ~n11483 & n11482 ) ;
  assign n11485 = ( n11482 & ~n10968 ) | ( n11482 & n11483 ) | ( ~n10968 & n11483 ) ;
  assign n11486 = ( n10973 & ~n11484 ) | ( n10973 & n11485 ) | ( ~n11484 & n11485 ) ;
  assign n11487 = ( n11481 & ~n1636 ) | ( n11481 & n11486 ) | ( ~n1636 & n11486 ) ;
  assign n11488 = ~n1452 & n11487 ;
  assign n11489 = n11001 | n11176 ;
  assign n11490 = ( n10988 & ~n10997 ) | ( n10988 & n11001 ) | ( ~n10997 & n11001 ) ;
  assign n11491 = ( n10997 & n11489 ) | ( n10997 & n11490 ) | ( n11489 & n11490 ) ;
  assign n11492 = ( n11001 & ~n11490 ) | ( n11001 & n11489 ) | ( ~n11490 & n11489 ) ;
  assign n11493 = ( n10988 & ~n11491 ) | ( n10988 & n11492 ) | ( ~n11491 & n11492 ) ;
  assign n11494 = ( n1636 & ~n11466 ) | ( n1636 & 1'b0 ) | ( ~n11466 & 1'b0 ) ;
  assign n11495 = ~n11480 & n11494 ;
  assign n11496 = ( n11486 & ~n11495 ) | ( n11486 & 1'b0 ) | ( ~n11495 & 1'b0 ) ;
  assign n11497 = n11474 | n11477 ;
  assign n11498 = ( n1827 & ~n11471 ) | ( n1827 & n11497 ) | ( ~n11471 & n11497 ) ;
  assign n11499 = ~n1636 & n11498 ;
  assign n11500 = ( n1452 & ~n11499 ) | ( n1452 & 1'b0 ) | ( ~n11499 & 1'b0 ) ;
  assign n11501 = ~n11496 & n11500 ;
  assign n11502 = ( n11493 & ~n11501 ) | ( n11493 & 1'b0 ) | ( ~n11501 & 1'b0 ) ;
  assign n11503 = n11488 | n11502 ;
  assign n11509 = ( n1283 & ~n11508 ) | ( n1283 & n11503 ) | ( ~n11508 & n11503 ) ;
  assign n11510 = ~n1122 & n11509 ;
  assign n11511 = n11023 | n11176 ;
  assign n11512 = ( n11010 & ~n11019 ) | ( n11010 & n11023 ) | ( ~n11019 & n11023 ) ;
  assign n11513 = ( n11019 & n11511 ) | ( n11019 & n11512 ) | ( n11511 & n11512 ) ;
  assign n11514 = ( n11023 & ~n11512 ) | ( n11023 & n11511 ) | ( ~n11512 & n11511 ) ;
  assign n11515 = ( n11010 & ~n11513 ) | ( n11010 & n11514 ) | ( ~n11513 & n11514 ) ;
  assign n11516 = n1283 | n11488 ;
  assign n11517 = n11502 | n11516 ;
  assign n11518 = ~n11508 & n11517 ;
  assign n11519 = n11496 | n11499 ;
  assign n11520 = ( n11493 & ~n1452 ) | ( n11493 & n11519 ) | ( ~n1452 & n11519 ) ;
  assign n11521 = n1283 &  n11520 ;
  assign n11522 = ( n1122 & ~n11521 ) | ( n1122 & 1'b0 ) | ( ~n11521 & 1'b0 ) ;
  assign n11523 = ~n11518 & n11522 ;
  assign n11524 = ( n11515 & ~n11523 ) | ( n11515 & 1'b0 ) | ( ~n11523 & 1'b0 ) ;
  assign n11525 = n11510 | n11524 ;
  assign n11527 = ( n11012 & ~n11017 ) | ( n11012 & n11176 ) | ( ~n11017 & n11176 ) ;
  assign n11526 = n11025 &  n11176 ;
  assign n11528 = ( n11176 & ~n11527 ) | ( n11176 & n11526 ) | ( ~n11527 & n11526 ) ;
  assign n11529 = ( n11526 & ~n11012 ) | ( n11526 & n11527 ) | ( ~n11012 & n11527 ) ;
  assign n11530 = ( n11017 & ~n11528 ) | ( n11017 & n11529 ) | ( ~n11528 & n11529 ) ;
  assign n11531 = ( n976 & ~n11525 ) | ( n976 & n11530 ) | ( ~n11525 & n11530 ) ;
  assign n11532 = ( n837 & ~n11531 ) | ( n837 & 1'b0 ) | ( ~n11531 & 1'b0 ) ;
  assign n11533 = ( n11045 & ~n11176 ) | ( n11045 & 1'b0 ) | ( ~n11176 & 1'b0 ) ;
  assign n11534 = ( n11032 & n11041 ) | ( n11032 & n11045 ) | ( n11041 & n11045 ) ;
  assign n11535 = ( n11533 & ~n11041 ) | ( n11533 & n11534 ) | ( ~n11041 & n11534 ) ;
  assign n11536 = ( n11045 & ~n11534 ) | ( n11045 & n11533 ) | ( ~n11534 & n11533 ) ;
  assign n11537 = ( n11032 & ~n11535 ) | ( n11032 & n11536 ) | ( ~n11535 & n11536 ) ;
  assign n11538 = ( n976 & ~n11510 ) | ( n976 & 1'b0 ) | ( ~n11510 & 1'b0 ) ;
  assign n11539 = ~n11524 & n11538 ;
  assign n11540 = n11530 | n11539 ;
  assign n11541 = n11518 | n11521 ;
  assign n11542 = ( n11515 & ~n1122 ) | ( n11515 & n11541 ) | ( ~n1122 & n11541 ) ;
  assign n11543 = ~n976 & n11542 ;
  assign n11544 = n837 | n11543 ;
  assign n11545 = ( n11540 & ~n11544 ) | ( n11540 & 1'b0 ) | ( ~n11544 & 1'b0 ) ;
  assign n11546 = n11537 | n11545 ;
  assign n11547 = ~n11532 & n11546 ;
  assign n11548 = n11047 &  n11176 ;
  assign n11549 = ( n11034 & n11039 ) | ( n11034 & n11176 ) | ( n11039 & n11176 ) ;
  assign n11551 = ( n11548 & ~n11034 ) | ( n11548 & n11549 ) | ( ~n11034 & n11549 ) ;
  assign n11550 = ( n11176 & ~n11549 ) | ( n11176 & n11548 ) | ( ~n11549 & n11548 ) ;
  assign n11552 = ( n11039 & ~n11551 ) | ( n11039 & n11550 ) | ( ~n11551 & n11550 ) ;
  assign n11553 = ( n713 & ~n11547 ) | ( n713 & n11552 ) | ( ~n11547 & n11552 ) ;
  assign n11554 = n595 &  n11553 ;
  assign n11555 = n11067 | n11176 ;
  assign n11556 = ( n11054 & n11063 ) | ( n11054 & n11067 ) | ( n11063 & n11067 ) ;
  assign n11557 = ( n11555 & ~n11063 ) | ( n11555 & n11556 ) | ( ~n11063 & n11556 ) ;
  assign n11558 = ( n11067 & ~n11556 ) | ( n11067 & n11555 ) | ( ~n11556 & n11555 ) ;
  assign n11559 = ( n11054 & ~n11557 ) | ( n11054 & n11558 ) | ( ~n11557 & n11558 ) ;
  assign n11560 = n713 | n11532 ;
  assign n11561 = ( n11546 & ~n11560 ) | ( n11546 & 1'b0 ) | ( ~n11560 & 1'b0 ) ;
  assign n11562 = ( n11552 & ~n11561 ) | ( n11552 & 1'b0 ) | ( ~n11561 & 1'b0 ) ;
  assign n11563 = ( n11540 & ~n11543 ) | ( n11540 & 1'b0 ) | ( ~n11543 & 1'b0 ) ;
  assign n11564 = ( n11537 & ~n837 ) | ( n11537 & n11563 ) | ( ~n837 & n11563 ) ;
  assign n11565 = ( n713 & ~n11564 ) | ( n713 & 1'b0 ) | ( ~n11564 & 1'b0 ) ;
  assign n11566 = n595 | n11565 ;
  assign n11567 = n11562 | n11566 ;
  assign n11568 = n11559 &  n11567 ;
  assign n11569 = n11554 | n11568 ;
  assign n11575 = ( n492 & ~n11574 ) | ( n492 & n11569 ) | ( ~n11574 & n11569 ) ;
  assign n11576 = n396 &  n11575 ;
  assign n11577 = n11089 | n11176 ;
  assign n11578 = ( n11076 & n11085 ) | ( n11076 & n11089 ) | ( n11085 & n11089 ) ;
  assign n11579 = ( n11577 & ~n11085 ) | ( n11577 & n11578 ) | ( ~n11085 & n11578 ) ;
  assign n11580 = ( n11089 & ~n11578 ) | ( n11089 & n11577 ) | ( ~n11578 & n11577 ) ;
  assign n11581 = ( n11076 & ~n11579 ) | ( n11076 & n11580 ) | ( ~n11579 & n11580 ) ;
  assign n11582 = n492 | n11554 ;
  assign n11583 = n11568 | n11582 ;
  assign n11584 = ~n11574 & n11583 ;
  assign n11585 = n11562 | n11565 ;
  assign n11586 = ( n595 & n11559 ) | ( n595 & n11585 ) | ( n11559 & n11585 ) ;
  assign n11587 = n492 &  n11586 ;
  assign n11588 = n396 | n11587 ;
  assign n11589 = n11584 | n11588 ;
  assign n11590 = n11581 &  n11589 ;
  assign n11591 = n11576 | n11590 ;
  assign n11592 = ~n11091 & n11176 ;
  assign n11593 = ( n11078 & n11083 ) | ( n11078 & n11176 ) | ( n11083 & n11176 ) ;
  assign n11595 = ( n11592 & ~n11078 ) | ( n11592 & n11593 ) | ( ~n11078 & n11593 ) ;
  assign n11594 = ( n11176 & ~n11593 ) | ( n11176 & n11592 ) | ( ~n11593 & n11592 ) ;
  assign n11596 = ( n11083 & ~n11595 ) | ( n11083 & n11594 ) | ( ~n11595 & n11594 ) ;
  assign n11597 = ( n315 & n11591 ) | ( n315 & n11596 ) | ( n11591 & n11596 ) ;
  assign n11598 = n240 &  n11597 ;
  assign n11600 = ( n11107 & ~n11098 ) | ( n11107 & n11111 ) | ( ~n11098 & n11111 ) ;
  assign n11599 = n11111 | n11176 ;
  assign n11602 = ( n11111 & ~n11600 ) | ( n11111 & n11599 ) | ( ~n11600 & n11599 ) ;
  assign n11601 = ( n11599 & ~n11107 ) | ( n11599 & n11600 ) | ( ~n11107 & n11600 ) ;
  assign n11603 = ( n11098 & ~n11602 ) | ( n11098 & n11601 ) | ( ~n11602 & n11601 ) ;
  assign n11604 = n315 | n11576 ;
  assign n11605 = n11590 | n11604 ;
  assign n11606 = n11596 &  n11605 ;
  assign n11607 = n11584 | n11587 ;
  assign n11608 = ( n396 & n11581 ) | ( n396 & n11607 ) | ( n11581 & n11607 ) ;
  assign n11609 = n315 &  n11608 ;
  assign n11610 = n240 | n11609 ;
  assign n11611 = n11606 | n11610 ;
  assign n11612 = ~n11603 & n11611 ;
  assign n11613 = n11598 | n11612 ;
  assign n11614 = ~n11113 & n11176 ;
  assign n11615 = ( n11100 & n11105 ) | ( n11100 & n11176 ) | ( n11105 & n11176 ) ;
  assign n11617 = ( n11614 & ~n11100 ) | ( n11614 & n11615 ) | ( ~n11100 & n11615 ) ;
  assign n11616 = ( n11176 & ~n11615 ) | ( n11176 & n11614 ) | ( ~n11615 & n11614 ) ;
  assign n11618 = ( n11105 & ~n11617 ) | ( n11105 & n11616 ) | ( ~n11617 & n11616 ) ;
  assign n11619 = ( n181 & n11613 ) | ( n181 & n11618 ) | ( n11613 & n11618 ) ;
  assign n11620 = ~n145 & n11619 ;
  assign n11621 = n11133 | n11176 ;
  assign n11622 = ( n11120 & n11129 ) | ( n11120 & n11133 ) | ( n11129 & n11133 ) ;
  assign n11623 = ( n11621 & ~n11129 ) | ( n11621 & n11622 ) | ( ~n11129 & n11622 ) ;
  assign n11624 = ( n11133 & ~n11622 ) | ( n11133 & n11621 ) | ( ~n11622 & n11621 ) ;
  assign n11625 = ( n11120 & ~n11623 ) | ( n11120 & n11624 ) | ( ~n11623 & n11624 ) ;
  assign n11626 = n181 | n11598 ;
  assign n11627 = n11612 | n11626 ;
  assign n11628 = n11618 &  n11627 ;
  assign n11629 = n11606 | n11609 ;
  assign n11630 = ( n240 & ~n11603 ) | ( n240 & n11629 ) | ( ~n11603 & n11629 ) ;
  assign n11631 = n181 &  n11630 ;
  assign n11632 = ( n145 & ~n11631 ) | ( n145 & 1'b0 ) | ( ~n11631 & 1'b0 ) ;
  assign n11633 = ~n11628 & n11632 ;
  assign n11634 = n11625 | n11633 ;
  assign n11635 = ~n11620 & n11634 ;
  assign n11636 = n11122 | n11176 ;
  assign n11637 = ( n11127 & ~n11122 ) | ( n11127 & n11135 ) | ( ~n11122 & n11135 ) ;
  assign n11639 = ( n11122 & n11636 ) | ( n11122 & n11637 ) | ( n11636 & n11637 ) ;
  assign n11638 = ( n11135 & ~n11637 ) | ( n11135 & n11636 ) | ( ~n11637 & n11636 ) ;
  assign n11640 = ( n11127 & ~n11639 ) | ( n11127 & n11638 ) | ( ~n11639 & n11638 ) ;
  assign n11641 = ( n150 & ~n11635 ) | ( n150 & n11640 ) | ( ~n11635 & n11640 ) ;
  assign n11642 = n11142 | n11161 ;
  assign n11643 = ( n11158 & ~n11176 ) | ( n11158 & n11642 ) | ( ~n11176 & n11642 ) ;
  assign n11644 = ( n11158 & ~n11643 ) | ( n11158 & 1'b0 ) | ( ~n11643 & 1'b0 ) ;
  assign n11645 = ( n11158 & ~n11161 ) | ( n11158 & 1'b0 ) | ( ~n11161 & 1'b0 ) ;
  assign n11646 = ~n11176 & n11645 ;
  assign n11647 = ( n11142 & ~n11645 ) | ( n11142 & n11646 ) | ( ~n11645 & n11646 ) ;
  assign n11648 = n11644 | n11647 ;
  assign n11649 = ( n11143 & ~n11150 ) | ( n11143 & 1'b0 ) | ( ~n11150 & 1'b0 ) ;
  assign n11650 = ~n11176 & n11649 ;
  assign n11651 = ( n11164 & ~n11650 ) | ( n11164 & n11649 ) | ( ~n11650 & n11649 ) ;
  assign n11652 = ( n11648 & ~n11651 ) | ( n11648 & 1'b0 ) | ( ~n11651 & 1'b0 ) ;
  assign n11653 = ~n11641 & n11652 ;
  assign n11654 = ( n133 & ~n11653 ) | ( n133 & n11652 ) | ( ~n11653 & n11652 ) ;
  assign n11655 = n150 | n11620 ;
  assign n11656 = ( n11634 & ~n11655 ) | ( n11634 & 1'b0 ) | ( ~n11655 & 1'b0 ) ;
  assign n11661 = n11640 &  n11656 ;
  assign n11657 = n11628 | n11631 ;
  assign n11658 = ( n145 & ~n11657 ) | ( n145 & n11625 ) | ( ~n11657 & n11625 ) ;
  assign n11659 = ( n150 & ~n11658 ) | ( n150 & 1'b0 ) | ( ~n11658 & 1'b0 ) ;
  assign n11660 = n11648 | n11659 ;
  assign n11662 = ( n11640 & ~n11661 ) | ( n11640 & n11660 ) | ( ~n11661 & n11660 ) ;
  assign n11664 = ( n133 & ~n11150 ) | ( n133 & n11143 ) | ( ~n11150 & n11143 ) ;
  assign n11663 = ( n11150 & ~n11143 ) | ( n11150 & n11176 ) | ( ~n11143 & n11176 ) ;
  assign n11665 = ~n11150 & n11663 ;
  assign n11666 = ( n11150 & n11664 ) | ( n11150 & n11665 ) | ( n11664 & n11665 ) ;
  assign n11667 = n11146 | n11173 ;
  assign n11668 = ( n11149 & n11168 ) | ( n11149 & n11667 ) | ( n11168 & n11667 ) ;
  assign n11669 = ( n11149 & ~n11668 ) | ( n11149 & 1'b0 ) | ( ~n11668 & 1'b0 ) ;
  assign n11670 = ( n11156 & ~n11669 ) | ( n11156 & n11164 ) | ( ~n11669 & n11164 ) ;
  assign n11671 = ( n11156 & ~n11670 ) | ( n11156 & 1'b0 ) | ( ~n11670 & 1'b0 ) ;
  assign n11672 = n11666 | n11671 ;
  assign n11673 = ( n11662 & ~n11672 ) | ( n11662 & 1'b0 ) | ( ~n11672 & 1'b0 ) ;
  assign n11674 = ~n11654 | ~n11673 ;
  assign n11952 = ~n11436 & n11674 ;
  assign n11953 = ( n11423 & n11428 ) | ( n11423 & n11674 ) | ( n11428 & n11674 ) ;
  assign n11955 = ( n11952 & ~n11423 ) | ( n11952 & n11953 ) | ( ~n11423 & n11953 ) ;
  assign n11954 = ( n11674 & ~n11953 ) | ( n11674 & n11952 ) | ( ~n11953 & n11952 ) ;
  assign n11956 = ( n11428 & ~n11955 ) | ( n11428 & n11954 ) | ( ~n11955 & n11954 ) ;
  assign n11938 = ( n11430 & ~n11421 ) | ( n11430 & n11434 ) | ( ~n11421 & n11434 ) ;
  assign n11937 = n11434 | n11674 ;
  assign n11940 = ( n11434 & ~n11938 ) | ( n11434 & n11937 ) | ( ~n11938 & n11937 ) ;
  assign n11939 = ( n11937 & ~n11430 ) | ( n11937 & n11938 ) | ( ~n11430 & n11938 ) ;
  assign n11941 = ( n11421 & ~n11940 ) | ( n11421 & n11939 ) | ( ~n11940 & n11939 ) ;
  assign n11931 = ( n11401 & ~n11406 ) | ( n11401 & n11674 ) | ( ~n11406 & n11674 ) ;
  assign n11930 = ~n11414 & n11674 ;
  assign n11932 = ( n11674 & ~n11931 ) | ( n11674 & n11930 ) | ( ~n11931 & n11930 ) ;
  assign n11933 = ( n11930 & ~n11401 ) | ( n11930 & n11931 ) | ( ~n11401 & n11931 ) ;
  assign n11934 = ( n11406 & ~n11932 ) | ( n11406 & n11933 ) | ( ~n11932 & n11933 ) ;
  assign n11916 = ( n11408 & ~n11399 ) | ( n11408 & n11412 ) | ( ~n11399 & n11412 ) ;
  assign n11915 = n11412 | n11674 ;
  assign n11918 = ( n11412 & ~n11916 ) | ( n11412 & n11915 ) | ( ~n11916 & n11915 ) ;
  assign n11917 = ( n11915 & ~n11408 ) | ( n11915 & n11916 ) | ( ~n11408 & n11916 ) ;
  assign n11919 = ( n11399 & ~n11918 ) | ( n11399 & n11917 ) | ( ~n11918 & n11917 ) ;
  assign n11909 = ( n11379 & ~n11384 ) | ( n11379 & n11674 ) | ( ~n11384 & n11674 ) ;
  assign n11908 = ~n11392 & n11674 ;
  assign n11910 = ( n11674 & ~n11909 ) | ( n11674 & n11908 ) | ( ~n11909 & n11908 ) ;
  assign n11911 = ( n11908 & ~n11379 ) | ( n11908 & n11909 ) | ( ~n11379 & n11909 ) ;
  assign n11912 = ( n11384 & ~n11910 ) | ( n11384 & n11911 ) | ( ~n11910 & n11911 ) ;
  assign n11894 = ( n11386 & ~n11377 ) | ( n11386 & n11390 ) | ( ~n11377 & n11390 ) ;
  assign n11893 = n11390 | n11674 ;
  assign n11896 = ( n11390 & ~n11894 ) | ( n11390 & n11893 ) | ( ~n11894 & n11893 ) ;
  assign n11895 = ( n11893 & ~n11386 ) | ( n11893 & n11894 ) | ( ~n11386 & n11894 ) ;
  assign n11897 = ( n11377 & ~n11896 ) | ( n11377 & n11895 ) | ( ~n11896 & n11895 ) ;
  assign n11886 = ~n11370 & n11674 ;
  assign n11887 = ( n11357 & n11362 ) | ( n11357 & n11674 ) | ( n11362 & n11674 ) ;
  assign n11889 = ( n11886 & ~n11357 ) | ( n11886 & n11887 ) | ( ~n11357 & n11887 ) ;
  assign n11888 = ( n11674 & ~n11887 ) | ( n11674 & n11886 ) | ( ~n11887 & n11886 ) ;
  assign n11890 = ( n11362 & ~n11889 ) | ( n11362 & n11888 ) | ( ~n11889 & n11888 ) ;
  assign n11871 = n11368 | n11674 ;
  assign n11872 = ( n11355 & n11364 ) | ( n11355 & n11368 ) | ( n11364 & n11368 ) ;
  assign n11873 = ( n11871 & ~n11364 ) | ( n11871 & n11872 ) | ( ~n11364 & n11872 ) ;
  assign n11874 = ( n11368 & ~n11872 ) | ( n11368 & n11871 ) | ( ~n11872 & n11871 ) ;
  assign n11875 = ( n11355 & ~n11873 ) | ( n11355 & n11874 ) | ( ~n11873 & n11874 ) ;
  assign n11865 = ( n11335 & ~n11340 ) | ( n11335 & n11348 ) | ( ~n11340 & n11348 ) ;
  assign n11864 = n11335 | n11674 ;
  assign n11867 = ( n11335 & ~n11865 ) | ( n11335 & n11864 ) | ( ~n11865 & n11864 ) ;
  assign n11866 = ( n11864 & ~n11348 ) | ( n11864 & n11865 ) | ( ~n11348 & n11865 ) ;
  assign n11868 = ( n11340 & ~n11867 ) | ( n11340 & n11866 ) | ( ~n11867 & n11866 ) ;
  assign n11849 = n11346 | n11674 ;
  assign n11850 = ( n11333 & ~n11346 ) | ( n11333 & n11342 ) | ( ~n11346 & n11342 ) ;
  assign n11852 = ( n11346 & n11849 ) | ( n11346 & n11850 ) | ( n11849 & n11850 ) ;
  assign n11851 = ( n11342 & ~n11850 ) | ( n11342 & n11849 ) | ( ~n11850 & n11849 ) ;
  assign n11853 = ( n11333 & ~n11852 ) | ( n11333 & n11851 ) | ( ~n11852 & n11851 ) ;
  assign n11842 = n11313 | n11674 ;
  assign n11843 = ( n11318 & ~n11313 ) | ( n11318 & n11326 ) | ( ~n11313 & n11326 ) ;
  assign n11845 = ( n11313 & n11842 ) | ( n11313 & n11843 ) | ( n11842 & n11843 ) ;
  assign n11844 = ( n11326 & ~n11843 ) | ( n11326 & n11842 ) | ( ~n11843 & n11842 ) ;
  assign n11846 = ( n11318 & ~n11845 ) | ( n11318 & n11844 ) | ( ~n11845 & n11844 ) ;
  assign n11827 = n11324 | n11674 ;
  assign n11828 = ( n11311 & n11320 ) | ( n11311 & n11324 ) | ( n11320 & n11324 ) ;
  assign n11829 = ( n11827 & ~n11320 ) | ( n11827 & n11828 ) | ( ~n11320 & n11828 ) ;
  assign n11830 = ( n11324 & ~n11828 ) | ( n11324 & n11827 ) | ( ~n11828 & n11827 ) ;
  assign n11831 = ( n11311 & ~n11829 ) | ( n11311 & n11830 ) | ( ~n11829 & n11830 ) ;
  assign n11820 = n11291 | n11674 ;
  assign n11821 = ( n11291 & ~n11304 ) | ( n11291 & n11296 ) | ( ~n11304 & n11296 ) ;
  assign n11822 = ( n11304 & n11820 ) | ( n11304 & n11821 ) | ( n11820 & n11821 ) ;
  assign n11823 = ( n11291 & ~n11821 ) | ( n11291 & n11820 ) | ( ~n11821 & n11820 ) ;
  assign n11824 = ( n11296 & ~n11822 ) | ( n11296 & n11823 ) | ( ~n11822 & n11823 ) ;
  assign n11806 = ( n11298 & ~n11289 ) | ( n11298 & n11302 ) | ( ~n11289 & n11302 ) ;
  assign n11805 = n11302 | n11674 ;
  assign n11808 = ( n11302 & ~n11806 ) | ( n11302 & n11805 ) | ( ~n11806 & n11805 ) ;
  assign n11807 = ( n11805 & ~n11298 ) | ( n11805 & n11806 ) | ( ~n11298 & n11806 ) ;
  assign n11809 = ( n11289 & ~n11808 ) | ( n11289 & n11807 ) | ( ~n11808 & n11807 ) ;
  assign n11798 = n11269 | n11674 ;
  assign n11799 = ( n11269 & ~n11282 ) | ( n11269 & n11274 ) | ( ~n11282 & n11274 ) ;
  assign n11800 = ( n11282 & n11798 ) | ( n11282 & n11799 ) | ( n11798 & n11799 ) ;
  assign n11801 = ( n11269 & ~n11799 ) | ( n11269 & n11798 ) | ( ~n11799 & n11798 ) ;
  assign n11802 = ( n11274 & ~n11800 ) | ( n11274 & n11801 ) | ( ~n11800 & n11801 ) ;
  assign n11783 = n11280 | n11674 ;
  assign n11784 = ( n11267 & ~n11280 ) | ( n11267 & n11276 ) | ( ~n11280 & n11276 ) ;
  assign n11786 = ( n11280 & n11783 ) | ( n11280 & n11784 ) | ( n11783 & n11784 ) ;
  assign n11785 = ( n11276 & ~n11784 ) | ( n11276 & n11783 ) | ( ~n11784 & n11783 ) ;
  assign n11787 = ( n11267 & ~n11786 ) | ( n11267 & n11785 ) | ( ~n11786 & n11785 ) ;
  assign n11776 = n11247 | n11674 ;
  assign n11777 = ( n11247 & ~n11260 ) | ( n11247 & n11252 ) | ( ~n11260 & n11252 ) ;
  assign n11778 = ( n11260 & n11776 ) | ( n11260 & n11777 ) | ( n11776 & n11777 ) ;
  assign n11779 = ( n11247 & ~n11777 ) | ( n11247 & n11776 ) | ( ~n11777 & n11776 ) ;
  assign n11780 = ( n11252 & ~n11778 ) | ( n11252 & n11779 ) | ( ~n11778 & n11779 ) ;
  assign n11761 = n11258 | n11674 ;
  assign n11762 = ( n11245 & ~n11254 ) | ( n11245 & n11258 ) | ( ~n11254 & n11258 ) ;
  assign n11763 = ( n11254 & n11761 ) | ( n11254 & n11762 ) | ( n11761 & n11762 ) ;
  assign n11764 = ( n11258 & ~n11762 ) | ( n11258 & n11761 ) | ( ~n11762 & n11761 ) ;
  assign n11765 = ( n11245 & ~n11763 ) | ( n11245 & n11764 ) | ( ~n11763 & n11764 ) ;
  assign n11754 = n11238 &  n11674 ;
  assign n11755 = ( n11225 & n11230 ) | ( n11225 & n11674 ) | ( n11230 & n11674 ) ;
  assign n11757 = ( n11754 & ~n11225 ) | ( n11754 & n11755 ) | ( ~n11225 & n11755 ) ;
  assign n11756 = ( n11674 & ~n11755 ) | ( n11674 & n11754 ) | ( ~n11755 & n11754 ) ;
  assign n11758 = ( n11230 & ~n11757 ) | ( n11230 & n11756 ) | ( ~n11757 & n11756 ) ;
  assign n11739 = n11236 | n11674 ;
  assign n11740 = ( n11223 & ~n11236 ) | ( n11223 & n11232 ) | ( ~n11236 & n11232 ) ;
  assign n11742 = ( n11236 & n11739 ) | ( n11236 & n11740 ) | ( n11739 & n11740 ) ;
  assign n11741 = ( n11232 & ~n11740 ) | ( n11232 & n11739 ) | ( ~n11740 & n11739 ) ;
  assign n11743 = ( n11223 & ~n11742 ) | ( n11223 & n11741 ) | ( ~n11742 & n11741 ) ;
  assign n11733 = ( n11199 & ~n11209 ) | ( n11199 & n11216 ) | ( ~n11209 & n11216 ) ;
  assign n11732 = ( n11199 & ~n11674 ) | ( n11199 & 1'b0 ) | ( ~n11674 & 1'b0 ) ;
  assign n11735 = ( n11199 & ~n11733 ) | ( n11199 & n11732 ) | ( ~n11733 & n11732 ) ;
  assign n11734 = ( n11732 & ~n11216 ) | ( n11732 & n11733 ) | ( ~n11216 & n11733 ) ;
  assign n11736 = ( n11209 & ~n11735 ) | ( n11209 & n11734 ) | ( ~n11735 & n11734 ) ;
  assign n11717 = ~n11211 & n11214 ;
  assign n11718 = ( n11197 & ~n11211 ) | ( n11197 & n11717 ) | ( ~n11211 & n11717 ) ;
  assign n11720 = ( n11674 & n11211 ) | ( n11674 & n11718 ) | ( n11211 & n11718 ) ;
  assign n11719 = ( n11674 & ~n11718 ) | ( n11674 & n11717 ) | ( ~n11718 & n11717 ) ;
  assign n11721 = ( n11197 & ~n11720 ) | ( n11197 & n11719 ) | ( ~n11720 & n11719 ) ;
  assign n11708 = ~x40 & n11176 ;
  assign n11709 = ( x41 & ~n11708 ) | ( x41 & 1'b0 ) | ( ~n11708 & 1'b0 ) ;
  assign n11710 = n11188 | n11709 ;
  assign n11705 = ( n11176 & ~x40 ) | ( n11176 & n11183 ) | ( ~x40 & n11183 ) ;
  assign n11706 = x40 &  n11705 ;
  assign n11707 = ( n11178 & ~n11706 ) | ( n11178 & n11183 ) | ( ~n11706 & n11183 ) ;
  assign n11711 = ( n11674 & ~n11710 ) | ( n11674 & n11707 ) | ( ~n11710 & n11707 ) ;
  assign n11713 = ( n11674 & ~n11711 ) | ( n11674 & 1'b0 ) | ( ~n11711 & 1'b0 ) ;
  assign n11712 = ~n11707 & n11711 ;
  assign n11714 = ( n11710 & ~n11713 ) | ( n11710 & n11712 ) | ( ~n11713 & n11712 ) ;
  assign n11681 = ( x38 & ~n11674 ) | ( x38 & x39 ) | ( ~n11674 & x39 ) ;
  assign n11687 = ( x38 & ~x39 ) | ( x38 & 1'b0 ) | ( ~x39 & 1'b0 ) ;
  assign n11677 = x36 | x37 ;
  assign n11682 = ~x38 & n11677 ;
  assign n11683 = ( x38 & ~n11174 ) | ( x38 & n11682 ) | ( ~n11174 & n11682 ) ;
  assign n11684 = ( n11156 & ~n11683 ) | ( n11156 & n11164 ) | ( ~n11683 & n11164 ) ;
  assign n11685 = ( n11156 & ~n11684 ) | ( n11156 & 1'b0 ) | ( ~n11684 & 1'b0 ) ;
  assign n11686 = ( n11674 & ~x39 ) | ( n11674 & n11685 ) | ( ~x39 & n11685 ) ;
  assign n11688 = ( n11681 & ~n11687 ) | ( n11681 & n11686 ) | ( ~n11687 & n11686 ) ;
  assign n11678 = x38 | n11677 ;
  assign n11679 = x38 &  n11674 ;
  assign n11680 = ( n11176 & ~n11678 ) | ( n11176 & n11679 ) | ( ~n11678 & n11679 ) ;
  assign n11691 = n10685 | n11680 ;
  assign n11692 = ( n11688 & ~n11691 ) | ( n11688 & 1'b0 ) | ( ~n11691 & 1'b0 ) ;
  assign n11694 = ( n11176 & ~n11671 ) | ( n11176 & 1'b0 ) | ( ~n11671 & 1'b0 ) ;
  assign n11695 = ( n11662 & ~n11694 ) | ( n11662 & n11666 ) | ( ~n11694 & n11666 ) ;
  assign n11696 = ( n11662 & ~n11695 ) | ( n11662 & 1'b0 ) | ( ~n11695 & 1'b0 ) ;
  assign n11697 = n11654 &  n11696 ;
  assign n11693 = ~n10686 & n11674 ;
  assign n11698 = ( n11693 & ~n11697 ) | ( n11693 & 1'b0 ) | ( ~n11697 & 1'b0 ) ;
  assign n11699 = ( x40 & n11697 ) | ( x40 & n11698 ) | ( n11697 & n11698 ) ;
  assign n11700 = x40 | n11697 ;
  assign n11701 = n11693 | n11700 ;
  assign n11702 = ~n11699 & n11701 ;
  assign n11703 = n11692 | n11702 ;
  assign n11689 = n11680 &  n11688 ;
  assign n11690 = ( n10685 & ~n11688 ) | ( n10685 & n11689 ) | ( ~n11688 & n11689 ) ;
  assign n11722 = n10209 | n11690 ;
  assign n11723 = ( n11703 & ~n11722 ) | ( n11703 & 1'b0 ) | ( ~n11722 & 1'b0 ) ;
  assign n11724 = n11714 | n11723 ;
  assign n11725 = ~n11680 & n11688 ;
  assign n11726 = ( n11702 & ~n10685 ) | ( n11702 & n11725 ) | ( ~n10685 & n11725 ) ;
  assign n11727 = ( n10209 & ~n11726 ) | ( n10209 & 1'b0 ) | ( ~n11726 & 1'b0 ) ;
  assign n11728 = ( n9740 & ~n11727 ) | ( n9740 & 1'b0 ) | ( ~n11727 & 1'b0 ) ;
  assign n11729 = n11724 &  n11728 ;
  assign n11730 = n11721 | n11729 ;
  assign n11704 = ~n11690 & n11703 ;
  assign n11715 = ( n11704 & ~n10209 ) | ( n11704 & n11714 ) | ( ~n10209 & n11714 ) ;
  assign n11716 = n9740 | n11715 ;
  assign n11744 = ~n9286 & n11716 ;
  assign n11745 = n11730 &  n11744 ;
  assign n11746 = n11736 | n11745 ;
  assign n11747 = ( n11724 & ~n11727 ) | ( n11724 & 1'b0 ) | ( ~n11727 & 1'b0 ) ;
  assign n11748 = ( n9740 & n11721 ) | ( n9740 & n11747 ) | ( n11721 & n11747 ) ;
  assign n11749 = ( n9286 & ~n11748 ) | ( n9286 & 1'b0 ) | ( ~n11748 & 1'b0 ) ;
  assign n11750 = n8839 | n11749 ;
  assign n11751 = ( n11746 & ~n11750 ) | ( n11746 & 1'b0 ) | ( ~n11750 & 1'b0 ) ;
  assign n11752 = n11743 | n11751 ;
  assign n11731 = n11716 &  n11730 ;
  assign n11737 = ( n11731 & ~n9286 ) | ( n11731 & n11736 ) | ( ~n9286 & n11736 ) ;
  assign n11738 = ( n8839 & ~n11737 ) | ( n8839 & 1'b0 ) | ( ~n11737 & 1'b0 ) ;
  assign n11766 = n8407 | n11738 ;
  assign n11767 = ( n11752 & ~n11766 ) | ( n11752 & 1'b0 ) | ( ~n11766 & 1'b0 ) ;
  assign n11768 = n11758 | n11767 ;
  assign n11769 = ( n11746 & ~n11749 ) | ( n11746 & 1'b0 ) | ( ~n11749 & 1'b0 ) ;
  assign n11770 = ( n11743 & ~n8839 ) | ( n11743 & n11769 ) | ( ~n8839 & n11769 ) ;
  assign n11771 = ( n8407 & ~n11770 ) | ( n8407 & 1'b0 ) | ( ~n11770 & 1'b0 ) ;
  assign n11772 = n7982 | n11771 ;
  assign n11773 = ( n11768 & ~n11772 ) | ( n11768 & 1'b0 ) | ( ~n11772 & 1'b0 ) ;
  assign n11774 = n11765 | n11773 ;
  assign n11753 = ~n11738 & n11752 ;
  assign n11759 = ( n11753 & ~n8407 ) | ( n11753 & n11758 ) | ( ~n8407 & n11758 ) ;
  assign n11760 = ( n7982 & ~n11759 ) | ( n7982 & 1'b0 ) | ( ~n11759 & 1'b0 ) ;
  assign n11788 = ( n7572 & ~n11760 ) | ( n7572 & 1'b0 ) | ( ~n11760 & 1'b0 ) ;
  assign n11789 = n11774 &  n11788 ;
  assign n11790 = ( n11780 & ~n11789 ) | ( n11780 & 1'b0 ) | ( ~n11789 & 1'b0 ) ;
  assign n11791 = ( n11768 & ~n11771 ) | ( n11768 & 1'b0 ) | ( ~n11771 & 1'b0 ) ;
  assign n11792 = ( n11765 & ~n7982 ) | ( n11765 & n11791 ) | ( ~n7982 & n11791 ) ;
  assign n11793 = n7572 | n11792 ;
  assign n11794 = n7169 &  n11793 ;
  assign n11795 = ~n11790 & n11794 ;
  assign n11796 = ( n11787 & ~n11795 ) | ( n11787 & 1'b0 ) | ( ~n11795 & 1'b0 ) ;
  assign n11775 = ~n11760 & n11774 ;
  assign n11781 = ( n7572 & ~n11780 ) | ( n7572 & n11775 ) | ( ~n11780 & n11775 ) ;
  assign n11782 = n7169 | n11781 ;
  assign n11810 = ~n6781 & n11782 ;
  assign n11811 = ~n11796 & n11810 ;
  assign n11812 = ( n11802 & ~n11811 ) | ( n11802 & 1'b0 ) | ( ~n11811 & 1'b0 ) ;
  assign n11813 = ~n11790 & n11793 ;
  assign n11814 = ( n7169 & ~n11787 ) | ( n7169 & n11813 ) | ( ~n11787 & n11813 ) ;
  assign n11815 = ( n6781 & ~n11814 ) | ( n6781 & 1'b0 ) | ( ~n11814 & 1'b0 ) ;
  assign n11816 = ( n6399 & ~n11815 ) | ( n6399 & 1'b0 ) | ( ~n11815 & 1'b0 ) ;
  assign n11817 = ~n11812 & n11816 ;
  assign n11818 = ( n11809 & ~n11817 ) | ( n11809 & 1'b0 ) | ( ~n11817 & 1'b0 ) ;
  assign n11797 = ( n11782 & ~n11796 ) | ( n11782 & 1'b0 ) | ( ~n11796 & 1'b0 ) ;
  assign n11803 = ( n6781 & ~n11797 ) | ( n6781 & n11802 ) | ( ~n11797 & n11802 ) ;
  assign n11804 = ~n6399 & n11803 ;
  assign n11832 = n6032 | n11804 ;
  assign n11833 = n11818 | n11832 ;
  assign n11834 = n11824 &  n11833 ;
  assign n11835 = n11812 | n11815 ;
  assign n11836 = ( n11809 & ~n6399 ) | ( n11809 & n11835 ) | ( ~n6399 & n11835 ) ;
  assign n11837 = n6032 &  n11836 ;
  assign n11838 = ( n5672 & ~n11837 ) | ( n5672 & 1'b0 ) | ( ~n11837 & 1'b0 ) ;
  assign n11839 = ~n11834 & n11838 ;
  assign n11840 = n11831 | n11839 ;
  assign n11819 = n11804 | n11818 ;
  assign n11825 = ( n6032 & n11819 ) | ( n6032 & n11824 ) | ( n11819 & n11824 ) ;
  assign n11826 = ~n5672 & n11825 ;
  assign n11854 = n5327 | n11826 ;
  assign n11855 = ( n11840 & ~n11854 ) | ( n11840 & 1'b0 ) | ( ~n11854 & 1'b0 ) ;
  assign n11856 = n11846 | n11855 ;
  assign n11857 = n11834 | n11837 ;
  assign n11858 = ( n5672 & ~n11857 ) | ( n5672 & n11831 ) | ( ~n11857 & n11831 ) ;
  assign n11859 = ( n5327 & ~n11858 ) | ( n5327 & 1'b0 ) | ( ~n11858 & 1'b0 ) ;
  assign n11860 = n4990 | n11859 ;
  assign n11861 = ( n11856 & ~n11860 ) | ( n11856 & 1'b0 ) | ( ~n11860 & 1'b0 ) ;
  assign n11862 = ( n11853 & ~n11861 ) | ( n11853 & 1'b0 ) | ( ~n11861 & 1'b0 ) ;
  assign n11841 = ~n11826 & n11840 ;
  assign n11847 = ( n11841 & ~n5327 ) | ( n11841 & n11846 ) | ( ~n5327 & n11846 ) ;
  assign n11848 = ( n4990 & ~n11847 ) | ( n4990 & 1'b0 ) | ( ~n11847 & 1'b0 ) ;
  assign n11876 = n4668 | n11848 ;
  assign n11877 = n11862 | n11876 ;
  assign n11878 = ~n11868 & n11877 ;
  assign n11879 = ( n11856 & ~n11859 ) | ( n11856 & 1'b0 ) | ( ~n11859 & 1'b0 ) ;
  assign n11880 = ( n4990 & ~n11879 ) | ( n4990 & n11853 ) | ( ~n11879 & n11853 ) ;
  assign n11881 = n4668 &  n11880 ;
  assign n11882 = n4353 | n11881 ;
  assign n11883 = n11878 | n11882 ;
  assign n11884 = n11875 &  n11883 ;
  assign n11863 = n11848 | n11862 ;
  assign n11869 = ( n4668 & ~n11868 ) | ( n4668 & n11863 ) | ( ~n11868 & n11863 ) ;
  assign n11870 = n4353 &  n11869 ;
  assign n11898 = n4053 | n11870 ;
  assign n11899 = n11884 | n11898 ;
  assign n11900 = n11890 &  n11899 ;
  assign n11901 = n11878 | n11881 ;
  assign n11902 = ( n4353 & n11875 ) | ( n4353 & n11901 ) | ( n11875 & n11901 ) ;
  assign n11903 = n4053 &  n11902 ;
  assign n11904 = n3760 | n11903 ;
  assign n11905 = n11900 | n11904 ;
  assign n11906 = ~n11897 & n11905 ;
  assign n11885 = n11870 | n11884 ;
  assign n11891 = ( n4053 & n11885 ) | ( n4053 & n11890 ) | ( n11885 & n11890 ) ;
  assign n11892 = n3760 &  n11891 ;
  assign n11920 = n3482 | n11892 ;
  assign n11921 = n11906 | n11920 ;
  assign n11922 = ~n11912 & n11921 ;
  assign n11923 = n11900 | n11903 ;
  assign n11924 = ( n3760 & ~n11897 ) | ( n3760 & n11923 ) | ( ~n11897 & n11923 ) ;
  assign n11925 = n3482 &  n11924 ;
  assign n11926 = n3211 | n11925 ;
  assign n11927 = n11922 | n11926 ;
  assign n11928 = ~n11919 & n11927 ;
  assign n11907 = n11892 | n11906 ;
  assign n11913 = ( n3482 & ~n11912 ) | ( n3482 & n11907 ) | ( ~n11912 & n11907 ) ;
  assign n11914 = n3211 &  n11913 ;
  assign n11942 = n2955 | n11914 ;
  assign n11943 = n11928 | n11942 ;
  assign n11944 = ~n11934 & n11943 ;
  assign n11945 = n11922 | n11925 ;
  assign n11946 = ( n3211 & ~n11919 ) | ( n3211 & n11945 ) | ( ~n11919 & n11945 ) ;
  assign n11947 = n2955 &  n11946 ;
  assign n11967 = n11944 | n11947 ;
  assign n11968 = ( n2706 & ~n11941 ) | ( n2706 & n11967 ) | ( ~n11941 & n11967 ) ;
  assign n11969 = n2472 &  n11968 ;
  assign n12149 = n11620 | n11674 ;
  assign n12150 = ( n11620 & ~n11633 ) | ( n11620 & n11625 ) | ( ~n11633 & n11625 ) ;
  assign n12151 = ( n11633 & n12149 ) | ( n11633 & n12150 ) | ( n12149 & n12150 ) ;
  assign n12152 = ( n11620 & ~n12150 ) | ( n11620 & n12149 ) | ( ~n12150 & n12149 ) ;
  assign n12153 = ( n11625 & ~n12151 ) | ( n11625 & n12152 ) | ( ~n12151 & n12152 ) ;
  assign n12128 = ( n11598 & ~n11603 ) | ( n11598 & n11674 ) | ( ~n11603 & n11674 ) ;
  assign n12127 = ~n11611 & n11674 ;
  assign n12129 = ( n11674 & ~n12128 ) | ( n11674 & n12127 ) | ( ~n12128 & n12127 ) ;
  assign n12130 = ( n12127 & ~n11598 ) | ( n12127 & n12128 ) | ( ~n11598 & n12128 ) ;
  assign n12131 = ( n11603 & ~n12129 ) | ( n11603 & n12130 ) | ( ~n12129 & n12130 ) ;
  assign n12039 = n11523 &  n11674 ;
  assign n12040 = ( n11510 & n11515 ) | ( n11510 & n11674 ) | ( n11515 & n11674 ) ;
  assign n12042 = ( n12039 & ~n11510 ) | ( n12039 & n12040 ) | ( ~n11510 & n12040 ) ;
  assign n12041 = ( n11674 & ~n12040 ) | ( n11674 & n12039 ) | ( ~n12040 & n12039 ) ;
  assign n12043 = ( n11515 & ~n12042 ) | ( n11515 & n12041 ) | ( ~n12042 & n12041 ) ;
  assign n11929 = n11914 | n11928 ;
  assign n11935 = ( n2955 & ~n11934 ) | ( n2955 & n11929 ) | ( ~n11934 & n11929 ) ;
  assign n11936 = n2706 &  n11935 ;
  assign n11948 = n2706 | n11947 ;
  assign n11949 = n11944 | n11948 ;
  assign n11950 = ~n11941 & n11949 ;
  assign n11951 = n11936 | n11950 ;
  assign n11957 = ( n2472 & n11951 ) | ( n2472 & n11956 ) | ( n11951 & n11956 ) ;
  assign n11958 = n2245 &  n11957 ;
  assign n11960 = ( n11447 & ~n11443 ) | ( n11447 & n11451 ) | ( ~n11443 & n11451 ) ;
  assign n11959 = n11451 | n11674 ;
  assign n11962 = ( n11451 & ~n11960 ) | ( n11451 & n11959 ) | ( ~n11960 & n11959 ) ;
  assign n11961 = ( n11959 & ~n11447 ) | ( n11959 & n11960 ) | ( ~n11447 & n11960 ) ;
  assign n11963 = ( n11443 & ~n11962 ) | ( n11443 & n11961 ) | ( ~n11962 & n11961 ) ;
  assign n11964 = n2472 | n11936 ;
  assign n11965 = n11950 | n11964 ;
  assign n11966 = n11956 &  n11965 ;
  assign n11970 = n2245 | n11969 ;
  assign n11971 = n11966 | n11970 ;
  assign n11972 = ~n11963 & n11971 ;
  assign n11973 = n11958 | n11972 ;
  assign n11974 = ( n11445 & n11453 ) | ( n11445 & n11457 ) | ( n11453 & n11457 ) ;
  assign n11975 = ( n11674 & ~n11453 ) | ( n11674 & n11974 ) | ( ~n11453 & n11974 ) ;
  assign n11976 = ( n11445 & ~n11974 ) | ( n11445 & n11674 ) | ( ~n11974 & n11674 ) ;
  assign n11977 = ( n11457 & ~n11975 ) | ( n11457 & n11976 ) | ( ~n11975 & n11976 ) ;
  assign n11978 = ( n2033 & ~n11973 ) | ( n2033 & n11977 ) | ( ~n11973 & n11977 ) ;
  assign n11979 = ( n1827 & ~n11978 ) | ( n1827 & 1'b0 ) | ( ~n11978 & 1'b0 ) ;
  assign n11980 = n11477 | n11674 ;
  assign n11981 = ( n11464 & ~n11473 ) | ( n11464 & n11477 ) | ( ~n11473 & n11477 ) ;
  assign n11982 = ( n11473 & n11980 ) | ( n11473 & n11981 ) | ( n11980 & n11981 ) ;
  assign n11983 = ( n11477 & ~n11981 ) | ( n11477 & n11980 ) | ( ~n11981 & n11980 ) ;
  assign n11984 = ( n11464 & ~n11982 ) | ( n11464 & n11983 ) | ( ~n11982 & n11983 ) ;
  assign n11985 = ( n2033 & ~n11958 ) | ( n2033 & 1'b0 ) | ( ~n11958 & 1'b0 ) ;
  assign n11986 = ~n11972 & n11985 ;
  assign n11987 = n11977 | n11986 ;
  assign n11988 = n11966 | n11969 ;
  assign n11989 = ( n2245 & ~n11963 ) | ( n2245 & n11988 ) | ( ~n11963 & n11988 ) ;
  assign n11990 = ~n2033 & n11989 ;
  assign n11991 = n1827 | n11990 ;
  assign n11992 = ( n11987 & ~n11991 ) | ( n11987 & 1'b0 ) | ( ~n11991 & 1'b0 ) ;
  assign n11993 = ( n11984 & ~n11992 ) | ( n11984 & 1'b0 ) | ( ~n11992 & 1'b0 ) ;
  assign n11994 = n11979 | n11993 ;
  assign n11995 = ~n11479 & n11674 ;
  assign n11996 = ( n11466 & n11471 ) | ( n11466 & n11674 ) | ( n11471 & n11674 ) ;
  assign n11998 = ( n11995 & ~n11466 ) | ( n11995 & n11996 ) | ( ~n11466 & n11996 ) ;
  assign n11997 = ( n11674 & ~n11996 ) | ( n11674 & n11995 ) | ( ~n11996 & n11995 ) ;
  assign n11999 = ( n11471 & ~n11998 ) | ( n11471 & n11997 ) | ( ~n11998 & n11997 ) ;
  assign n12000 = ( n1636 & ~n11994 ) | ( n1636 & n11999 ) | ( ~n11994 & n11999 ) ;
  assign n12001 = n1452 | n12000 ;
  assign n12002 = n11499 | n11674 ;
  assign n12003 = ( n11486 & ~n11495 ) | ( n11486 & n11499 ) | ( ~n11495 & n11499 ) ;
  assign n12004 = ( n11495 & n12002 ) | ( n11495 & n12003 ) | ( n12002 & n12003 ) ;
  assign n12005 = ( n11499 & ~n12003 ) | ( n11499 & n12002 ) | ( ~n12003 & n12002 ) ;
  assign n12006 = ( n11486 & ~n12004 ) | ( n11486 & n12005 ) | ( ~n12004 & n12005 ) ;
  assign n12007 = ( n1636 & ~n11979 ) | ( n1636 & 1'b0 ) | ( ~n11979 & 1'b0 ) ;
  assign n12008 = ~n11993 & n12007 ;
  assign n12009 = n11999 | n12008 ;
  assign n12010 = ( n11987 & ~n11990 ) | ( n11987 & 1'b0 ) | ( ~n11990 & 1'b0 ) ;
  assign n12011 = ( n1827 & ~n12010 ) | ( n1827 & n11984 ) | ( ~n12010 & n11984 ) ;
  assign n12012 = ~n1636 & n12011 ;
  assign n12013 = ( n1452 & ~n12012 ) | ( n1452 & 1'b0 ) | ( ~n12012 & 1'b0 ) ;
  assign n12014 = n12009 &  n12013 ;
  assign n12015 = ( n12006 & ~n12014 ) | ( n12006 & 1'b0 ) | ( ~n12014 & 1'b0 ) ;
  assign n12016 = ( n12001 & ~n12015 ) | ( n12001 & 1'b0 ) | ( ~n12015 & 1'b0 ) ;
  assign n12017 = n11501 &  n11674 ;
  assign n12018 = ( n11488 & n11493 ) | ( n11488 & n11674 ) | ( n11493 & n11674 ) ;
  assign n12020 = ( n12017 & ~n11488 ) | ( n12017 & n12018 ) | ( ~n11488 & n12018 ) ;
  assign n12019 = ( n11674 & ~n12018 ) | ( n11674 & n12017 ) | ( ~n12018 & n12017 ) ;
  assign n12021 = ( n11493 & ~n12020 ) | ( n11493 & n12019 ) | ( ~n12020 & n12019 ) ;
  assign n12022 = ( n1283 & ~n12016 ) | ( n1283 & n12021 ) | ( ~n12016 & n12021 ) ;
  assign n12023 = ~n1122 & n12022 ;
  assign n12025 = ( n11517 & ~n11508 ) | ( n11517 & n11521 ) | ( ~n11508 & n11521 ) ;
  assign n12024 = n11521 | n11674 ;
  assign n12027 = ( n11521 & ~n12025 ) | ( n11521 & n12024 ) | ( ~n12025 & n12024 ) ;
  assign n12026 = ( n12024 & ~n11517 ) | ( n12024 & n12025 ) | ( ~n11517 & n12025 ) ;
  assign n12028 = ( n11508 & ~n12027 ) | ( n11508 & n12026 ) | ( ~n12027 & n12026 ) ;
  assign n12029 = ~n1283 & n12001 ;
  assign n12030 = ~n12015 & n12029 ;
  assign n12031 = ( n12021 & ~n12030 ) | ( n12021 & 1'b0 ) | ( ~n12030 & 1'b0 ) ;
  assign n12032 = ( n12009 & ~n12012 ) | ( n12009 & 1'b0 ) | ( ~n12012 & 1'b0 ) ;
  assign n12033 = ( n1452 & ~n12006 ) | ( n1452 & n12032 ) | ( ~n12006 & n12032 ) ;
  assign n12034 = ( n1283 & ~n12033 ) | ( n1283 & 1'b0 ) | ( ~n12033 & 1'b0 ) ;
  assign n12035 = ( n1122 & ~n12034 ) | ( n1122 & 1'b0 ) | ( ~n12034 & 1'b0 ) ;
  assign n12036 = ~n12031 & n12035 ;
  assign n12037 = n12028 | n12036 ;
  assign n12038 = ~n12023 & n12037 ;
  assign n12044 = ( n976 & ~n12043 ) | ( n976 & n12038 ) | ( ~n12043 & n12038 ) ;
  assign n12045 = ( n837 & ~n12044 ) | ( n837 & 1'b0 ) | ( ~n12044 & 1'b0 ) ;
  assign n12046 = n11543 | n11674 ;
  assign n12047 = ( n11530 & ~n11543 ) | ( n11530 & n11539 ) | ( ~n11543 & n11539 ) ;
  assign n12049 = ( n11543 & n12046 ) | ( n11543 & n12047 ) | ( n12046 & n12047 ) ;
  assign n12048 = ( n11539 & ~n12047 ) | ( n11539 & n12046 ) | ( ~n12047 & n12046 ) ;
  assign n12050 = ( n11530 & ~n12049 ) | ( n11530 & n12048 ) | ( ~n12049 & n12048 ) ;
  assign n12051 = ( n976 & ~n12023 ) | ( n976 & 1'b0 ) | ( ~n12023 & 1'b0 ) ;
  assign n12052 = n12037 &  n12051 ;
  assign n12053 = ( n12043 & ~n12052 ) | ( n12043 & 1'b0 ) | ( ~n12052 & 1'b0 ) ;
  assign n12054 = n12031 | n12034 ;
  assign n12055 = ( n1122 & ~n12054 ) | ( n1122 & n12028 ) | ( ~n12054 & n12028 ) ;
  assign n12056 = n976 | n12055 ;
  assign n12057 = ~n837 & n12056 ;
  assign n12058 = ~n12053 & n12057 ;
  assign n12059 = n12050 | n12058 ;
  assign n12060 = ~n12045 & n12059 ;
  assign n12062 = ( n11532 & ~n11537 ) | ( n11532 & n11674 ) | ( ~n11537 & n11674 ) ;
  assign n12061 = n11545 &  n11674 ;
  assign n12063 = ( n11674 & ~n12062 ) | ( n11674 & n12061 ) | ( ~n12062 & n12061 ) ;
  assign n12064 = ( n12061 & ~n11532 ) | ( n12061 & n12062 ) | ( ~n11532 & n12062 ) ;
  assign n12065 = ( n11537 & ~n12063 ) | ( n11537 & n12064 ) | ( ~n12063 & n12064 ) ;
  assign n12066 = ( n12060 & ~n713 ) | ( n12060 & n12065 ) | ( ~n713 & n12065 ) ;
  assign n12067 = ( n595 & ~n12066 ) | ( n595 & 1'b0 ) | ( ~n12066 & 1'b0 ) ;
  assign n12068 = n11565 | n11674 ;
  assign n12069 = ( n11552 & ~n11561 ) | ( n11552 & n11565 ) | ( ~n11561 & n11565 ) ;
  assign n12070 = ( n11561 & n12068 ) | ( n11561 & n12069 ) | ( n12068 & n12069 ) ;
  assign n12071 = ( n11565 & ~n12069 ) | ( n11565 & n12068 ) | ( ~n12069 & n12068 ) ;
  assign n12072 = ( n11552 & ~n12070 ) | ( n11552 & n12071 ) | ( ~n12070 & n12071 ) ;
  assign n12073 = n713 | n12045 ;
  assign n12074 = ( n12059 & ~n12073 ) | ( n12059 & 1'b0 ) | ( ~n12073 & 1'b0 ) ;
  assign n12075 = n12065 | n12074 ;
  assign n12076 = ~n12053 & n12056 ;
  assign n12077 = ( n12050 & ~n837 ) | ( n12050 & n12076 ) | ( ~n837 & n12076 ) ;
  assign n12078 = ( n713 & ~n12077 ) | ( n713 & 1'b0 ) | ( ~n12077 & 1'b0 ) ;
  assign n12079 = n595 | n12078 ;
  assign n12080 = ( n12075 & ~n12079 ) | ( n12075 & 1'b0 ) | ( ~n12079 & 1'b0 ) ;
  assign n12081 = ( n12072 & ~n12080 ) | ( n12072 & 1'b0 ) | ( ~n12080 & 1'b0 ) ;
  assign n12082 = n12067 | n12081 ;
  assign n12083 = ~n11567 & n11674 ;
  assign n12084 = ( n11554 & n11559 ) | ( n11554 & n11674 ) | ( n11559 & n11674 ) ;
  assign n12086 = ( n12083 & ~n11554 ) | ( n12083 & n12084 ) | ( ~n11554 & n12084 ) ;
  assign n12085 = ( n11674 & ~n12084 ) | ( n11674 & n12083 ) | ( ~n12084 & n12083 ) ;
  assign n12087 = ( n11559 & ~n12086 ) | ( n11559 & n12085 ) | ( ~n12086 & n12085 ) ;
  assign n12088 = ( n492 & n12082 ) | ( n492 & n12087 ) | ( n12082 & n12087 ) ;
  assign n12089 = n396 &  n12088 ;
  assign n12091 = ( n11583 & ~n11574 ) | ( n11583 & n11587 ) | ( ~n11574 & n11587 ) ;
  assign n12090 = n11587 | n11674 ;
  assign n12093 = ( n11587 & ~n12091 ) | ( n11587 & n12090 ) | ( ~n12091 & n12090 ) ;
  assign n12092 = ( n12090 & ~n11583 ) | ( n12090 & n12091 ) | ( ~n11583 & n12091 ) ;
  assign n12094 = ( n11574 & ~n12093 ) | ( n11574 & n12092 ) | ( ~n12093 & n12092 ) ;
  assign n12095 = n492 | n12067 ;
  assign n12096 = n12081 | n12095 ;
  assign n12097 = n12087 &  n12096 ;
  assign n12098 = ( n12075 & ~n12078 ) | ( n12075 & 1'b0 ) | ( ~n12078 & 1'b0 ) ;
  assign n12099 = ( n595 & ~n12098 ) | ( n595 & n12072 ) | ( ~n12098 & n12072 ) ;
  assign n12100 = n492 &  n12099 ;
  assign n12101 = n396 | n12100 ;
  assign n12102 = n12097 | n12101 ;
  assign n12103 = ~n12094 & n12102 ;
  assign n12104 = n12089 | n12103 ;
  assign n12105 = ~n11589 & n11674 ;
  assign n12106 = ( n11576 & n11581 ) | ( n11576 & n11674 ) | ( n11581 & n11674 ) ;
  assign n12108 = ( n12105 & ~n11576 ) | ( n12105 & n12106 ) | ( ~n11576 & n12106 ) ;
  assign n12107 = ( n11674 & ~n12106 ) | ( n11674 & n12105 ) | ( ~n12106 & n12105 ) ;
  assign n12109 = ( n11581 & ~n12108 ) | ( n11581 & n12107 ) | ( ~n12108 & n12107 ) ;
  assign n12110 = ( n315 & n12104 ) | ( n315 & n12109 ) | ( n12104 & n12109 ) ;
  assign n12111 = n240 &  n12110 ;
  assign n12112 = n11609 | n11674 ;
  assign n12113 = ( n11596 & n11605 ) | ( n11596 & n11609 ) | ( n11605 & n11609 ) ;
  assign n12114 = ( n12112 & ~n11605 ) | ( n12112 & n12113 ) | ( ~n11605 & n12113 ) ;
  assign n12115 = ( n11609 & ~n12113 ) | ( n11609 & n12112 ) | ( ~n12113 & n12112 ) ;
  assign n12116 = ( n11596 & ~n12114 ) | ( n11596 & n12115 ) | ( ~n12114 & n12115 ) ;
  assign n12117 = n315 | n12089 ;
  assign n12118 = n12103 | n12117 ;
  assign n12119 = n12109 &  n12118 ;
  assign n12120 = n12097 | n12100 ;
  assign n12121 = ( n396 & ~n12094 ) | ( n396 & n12120 ) | ( ~n12094 & n12120 ) ;
  assign n12122 = n315 &  n12121 ;
  assign n12123 = n240 | n12122 ;
  assign n12124 = n12119 | n12123 ;
  assign n12125 = n12116 &  n12124 ;
  assign n12126 = n12111 | n12125 ;
  assign n12132 = ( n181 & ~n12131 ) | ( n181 & n12126 ) | ( ~n12131 & n12126 ) ;
  assign n12133 = ~n145 & n12132 ;
  assign n12135 = ( n11627 & ~n11618 ) | ( n11627 & n11631 ) | ( ~n11618 & n11631 ) ;
  assign n12134 = n11631 | n11674 ;
  assign n12137 = ( n11631 & ~n12135 ) | ( n11631 & n12134 ) | ( ~n12135 & n12134 ) ;
  assign n12136 = ( n12134 & ~n11627 ) | ( n12134 & n12135 ) | ( ~n11627 & n12135 ) ;
  assign n12138 = ( n11618 & ~n12137 ) | ( n11618 & n12136 ) | ( ~n12137 & n12136 ) ;
  assign n12139 = n181 | n12111 ;
  assign n12140 = n12125 | n12139 ;
  assign n12141 = ~n12131 & n12140 ;
  assign n12142 = n12119 | n12122 ;
  assign n12143 = ( n240 & n12116 ) | ( n240 & n12142 ) | ( n12116 & n12142 ) ;
  assign n12144 = n181 &  n12143 ;
  assign n12145 = ( n145 & ~n12144 ) | ( n145 & 1'b0 ) | ( ~n12144 & 1'b0 ) ;
  assign n12146 = ~n12141 & n12145 ;
  assign n12147 = ( n12138 & ~n12146 ) | ( n12138 & 1'b0 ) | ( ~n12146 & 1'b0 ) ;
  assign n12148 = n12133 | n12147 ;
  assign n12154 = ( n150 & ~n12153 ) | ( n150 & n12148 ) | ( ~n12153 & n12148 ) ;
  assign n12155 = n11640 | n11656 ;
  assign n12156 = ( n11659 & ~n12155 ) | ( n11659 & n11674 ) | ( ~n12155 & n11674 ) ;
  assign n12157 = ~n11659 & n12156 ;
  assign n12158 = n11656 | n11659 ;
  assign n12159 = n11674 | n12158 ;
  assign n12160 = ( n11640 & ~n12159 ) | ( n11640 & n12158 ) | ( ~n12159 & n12158 ) ;
  assign n12161 = n12157 | n12160 ;
  assign n12162 = n11641 &  n11648 ;
  assign n12163 = ~n11674 & n12162 ;
  assign n12164 = ( n11662 & ~n12162 ) | ( n11662 & n12163 ) | ( ~n12162 & n12163 ) ;
  assign n12165 = n12161 &  n12164 ;
  assign n12166 = ~n12154 & n12165 ;
  assign n12167 = ( n133 & ~n12166 ) | ( n133 & n12165 ) | ( ~n12166 & n12165 ) ;
  assign n12170 = n12141 | n12144 ;
  assign n12171 = ( n12138 & ~n145 ) | ( n12138 & n12170 ) | ( ~n145 & n12170 ) ;
  assign n12172 = n150 &  n12171 ;
  assign n12173 = n12161 | n12172 ;
  assign n12168 = n150 | n12133 ;
  assign n12169 = n12147 | n12168 ;
  assign n12174 = n12153 | n12169 ;
  assign n12175 = ( n12173 & ~n12153 ) | ( n12173 & n12174 ) | ( ~n12153 & n12174 ) ;
  assign n12177 = ( n133 & n11641 ) | ( n133 & n11648 ) | ( n11641 & n11648 ) ;
  assign n12176 = ( n11641 & ~n11674 ) | ( n11641 & n11648 ) | ( ~n11674 & n11648 ) ;
  assign n12178 = ( n11648 & ~n12176 ) | ( n11648 & 1'b0 ) | ( ~n12176 & 1'b0 ) ;
  assign n12179 = ( n12177 & ~n11648 ) | ( n12177 & n12178 ) | ( ~n11648 & n12178 ) ;
  assign n12180 = n11644 | n11671 ;
  assign n12181 = ( n11666 & ~n11647 ) | ( n11666 & n12180 ) | ( ~n11647 & n12180 ) ;
  assign n12182 = n11647 | n12181 ;
  assign n12183 = ( n11654 & ~n11662 ) | ( n11654 & n12182 ) | ( ~n11662 & n12182 ) ;
  assign n12184 = ( n11654 & ~n12183 ) | ( n11654 & 1'b0 ) | ( ~n12183 & 1'b0 ) ;
  assign n12185 = n12179 | n12184 ;
  assign n12186 = ( n12175 & ~n12185 ) | ( n12175 & 1'b0 ) | ( ~n12185 & 1'b0 ) ;
  assign n12187 = ~n12167 | ~n12186 ;
  assign n12479 = n11969 | n12187 ;
  assign n12480 = ( n11956 & n11965 ) | ( n11956 & n11969 ) | ( n11965 & n11969 ) ;
  assign n12481 = ( n12479 & ~n11965 ) | ( n12479 & n12480 ) | ( ~n11965 & n12480 ) ;
  assign n12482 = ( n11969 & ~n12480 ) | ( n11969 & n12479 ) | ( ~n12480 & n12479 ) ;
  assign n12483 = ( n11956 & ~n12481 ) | ( n11956 & n12482 ) | ( ~n12481 & n12482 ) ;
  assign n12473 = ( n11936 & ~n11941 ) | ( n11936 & n12187 ) | ( ~n11941 & n12187 ) ;
  assign n12472 = ~n11949 & n12187 ;
  assign n12474 = ( n12187 & ~n12473 ) | ( n12187 & n12472 ) | ( ~n12473 & n12472 ) ;
  assign n12475 = ( n12472 & ~n11936 ) | ( n12472 & n12473 ) | ( ~n11936 & n12473 ) ;
  assign n12476 = ( n11941 & ~n12474 ) | ( n11941 & n12475 ) | ( ~n12474 & n12475 ) ;
  assign n12458 = ( n11943 & ~n11934 ) | ( n11943 & n11947 ) | ( ~n11934 & n11947 ) ;
  assign n12457 = n11947 | n12187 ;
  assign n12460 = ( n11947 & ~n12458 ) | ( n11947 & n12457 ) | ( ~n12458 & n12457 ) ;
  assign n12459 = ( n12457 & ~n11943 ) | ( n12457 & n12458 ) | ( ~n11943 & n12458 ) ;
  assign n12461 = ( n11934 & ~n12460 ) | ( n11934 & n12459 ) | ( ~n12460 & n12459 ) ;
  assign n12451 = ( n11914 & ~n11919 ) | ( n11914 & n12187 ) | ( ~n11919 & n12187 ) ;
  assign n12450 = ~n11927 & n12187 ;
  assign n12452 = ( n12187 & ~n12451 ) | ( n12187 & n12450 ) | ( ~n12451 & n12450 ) ;
  assign n12453 = ( n12450 & ~n11914 ) | ( n12450 & n12451 ) | ( ~n11914 & n12451 ) ;
  assign n12454 = ( n11919 & ~n12452 ) | ( n11919 & n12453 ) | ( ~n12452 & n12453 ) ;
  assign n12436 = ( n11921 & ~n11912 ) | ( n11921 & n11925 ) | ( ~n11912 & n11925 ) ;
  assign n12435 = n11925 | n12187 ;
  assign n12438 = ( n11925 & ~n12436 ) | ( n11925 & n12435 ) | ( ~n12436 & n12435 ) ;
  assign n12437 = ( n12435 & ~n11921 ) | ( n12435 & n12436 ) | ( ~n11921 & n12436 ) ;
  assign n12439 = ( n11912 & ~n12438 ) | ( n11912 & n12437 ) | ( ~n12438 & n12437 ) ;
  assign n12429 = ( n11892 & ~n11897 ) | ( n11892 & n12187 ) | ( ~n11897 & n12187 ) ;
  assign n12428 = ~n11905 & n12187 ;
  assign n12430 = ( n12187 & ~n12429 ) | ( n12187 & n12428 ) | ( ~n12429 & n12428 ) ;
  assign n12431 = ( n12428 & ~n11892 ) | ( n12428 & n12429 ) | ( ~n11892 & n12429 ) ;
  assign n12432 = ( n11897 & ~n12430 ) | ( n11897 & n12431 ) | ( ~n12430 & n12431 ) ;
  assign n12413 = n11903 | n12187 ;
  assign n12414 = ( n11890 & n11899 ) | ( n11890 & n11903 ) | ( n11899 & n11903 ) ;
  assign n12415 = ( n12413 & ~n11899 ) | ( n12413 & n12414 ) | ( ~n11899 & n12414 ) ;
  assign n12416 = ( n11903 & ~n12414 ) | ( n11903 & n12413 ) | ( ~n12414 & n12413 ) ;
  assign n12417 = ( n11890 & ~n12415 ) | ( n11890 & n12416 ) | ( ~n12415 & n12416 ) ;
  assign n12406 = n11870 | n12187 ;
  assign n12407 = ( n11870 & n11875 ) | ( n11870 & n11883 ) | ( n11875 & n11883 ) ;
  assign n12408 = ( n12406 & ~n11883 ) | ( n12406 & n12407 ) | ( ~n11883 & n12407 ) ;
  assign n12409 = ( n11870 & ~n12407 ) | ( n11870 & n12406 ) | ( ~n12407 & n12406 ) ;
  assign n12410 = ( n11875 & ~n12408 ) | ( n11875 & n12409 ) | ( ~n12408 & n12409 ) ;
  assign n12391 = n11881 | n12187 ;
  assign n12392 = ( n11868 & n11877 ) | ( n11868 & n11881 ) | ( n11877 & n11881 ) ;
  assign n12393 = ( n12391 & ~n11877 ) | ( n12391 & n12392 ) | ( ~n11877 & n12392 ) ;
  assign n12394 = ( n11881 & ~n12392 ) | ( n11881 & n12391 ) | ( ~n12392 & n12391 ) ;
  assign n12395 = ( n11868 & ~n12393 ) | ( n11868 & n12394 ) | ( ~n12393 & n12394 ) ;
  assign n12384 = n11848 | n12187 ;
  assign n12385 = ( n11848 & ~n11861 ) | ( n11848 & n11853 ) | ( ~n11861 & n11853 ) ;
  assign n12386 = ( n11861 & n12384 ) | ( n11861 & n12385 ) | ( n12384 & n12385 ) ;
  assign n12387 = ( n11848 & ~n12385 ) | ( n11848 & n12384 ) | ( ~n12385 & n12384 ) ;
  assign n12388 = ( n11853 & ~n12386 ) | ( n11853 & n12387 ) | ( ~n12386 & n12387 ) ;
  assign n12369 = n11859 | n12187 ;
  assign n12370 = ( n11846 & ~n11855 ) | ( n11846 & n11859 ) | ( ~n11855 & n11859 ) ;
  assign n12371 = ( n11855 & n12369 ) | ( n11855 & n12370 ) | ( n12369 & n12370 ) ;
  assign n12372 = ( n11859 & ~n12370 ) | ( n11859 & n12369 ) | ( ~n12370 & n12369 ) ;
  assign n12373 = ( n11846 & ~n12371 ) | ( n11846 & n12372 ) | ( ~n12371 & n12372 ) ;
  assign n12362 = n11826 | n12187 ;
  assign n12363 = ( n11831 & ~n11826 ) | ( n11831 & n11839 ) | ( ~n11826 & n11839 ) ;
  assign n12365 = ( n11826 & n12362 ) | ( n11826 & n12363 ) | ( n12362 & n12363 ) ;
  assign n12364 = ( n11839 & ~n12363 ) | ( n11839 & n12362 ) | ( ~n12363 & n12362 ) ;
  assign n12366 = ( n11831 & ~n12365 ) | ( n11831 & n12364 ) | ( ~n12365 & n12364 ) ;
  assign n12348 = ( n11833 & ~n11824 ) | ( n11833 & n11837 ) | ( ~n11824 & n11837 ) ;
  assign n12347 = n11837 | n12187 ;
  assign n12350 = ( n11837 & ~n12348 ) | ( n11837 & n12347 ) | ( ~n12348 & n12347 ) ;
  assign n12349 = ( n12347 & ~n11833 ) | ( n12347 & n12348 ) | ( ~n11833 & n12348 ) ;
  assign n12351 = ( n11824 & ~n12350 ) | ( n11824 & n12349 ) | ( ~n12350 & n12349 ) ;
  assign n12340 = n11804 | n12187 ;
  assign n12341 = ( n11804 & ~n11817 ) | ( n11804 & n11809 ) | ( ~n11817 & n11809 ) ;
  assign n12342 = ( n11817 & n12340 ) | ( n11817 & n12341 ) | ( n12340 & n12341 ) ;
  assign n12343 = ( n11804 & ~n12341 ) | ( n11804 & n12340 ) | ( ~n12341 & n12340 ) ;
  assign n12344 = ( n11809 & ~n12342 ) | ( n11809 & n12343 ) | ( ~n12342 & n12343 ) ;
  assign n12325 = n11815 | n12187 ;
  assign n12326 = ( n11802 & ~n11815 ) | ( n11802 & n11811 ) | ( ~n11815 & n11811 ) ;
  assign n12328 = ( n11815 & n12325 ) | ( n11815 & n12326 ) | ( n12325 & n12326 ) ;
  assign n12327 = ( n11811 & ~n12326 ) | ( n11811 & n12325 ) | ( ~n12326 & n12325 ) ;
  assign n12329 = ( n11802 & ~n12328 ) | ( n11802 & n12327 ) | ( ~n12328 & n12327 ) ;
  assign n12319 = ( n11782 & ~n11787 ) | ( n11782 & n11795 ) | ( ~n11787 & n11795 ) ;
  assign n12318 = ( n11782 & ~n12187 ) | ( n11782 & 1'b0 ) | ( ~n12187 & 1'b0 ) ;
  assign n12321 = ( n11782 & ~n12319 ) | ( n11782 & n12318 ) | ( ~n12319 & n12318 ) ;
  assign n12320 = ( n12318 & ~n11795 ) | ( n12318 & n12319 ) | ( ~n11795 & n12319 ) ;
  assign n12322 = ( n11787 & ~n12321 ) | ( n11787 & n12320 ) | ( ~n12321 & n12320 ) ;
  assign n12303 = ( n11793 & ~n12187 ) | ( n11793 & 1'b0 ) | ( ~n12187 & 1'b0 ) ;
  assign n12304 = ( n11780 & n11789 ) | ( n11780 & n11793 ) | ( n11789 & n11793 ) ;
  assign n12305 = ( n12303 & ~n11789 ) | ( n12303 & n12304 ) | ( ~n11789 & n12304 ) ;
  assign n12306 = ( n11793 & ~n12304 ) | ( n11793 & n12303 ) | ( ~n12304 & n12303 ) ;
  assign n12307 = ( n11780 & ~n12305 ) | ( n11780 & n12306 ) | ( ~n12305 & n12306 ) ;
  assign n12296 = n11760 | n12187 ;
  assign n12297 = ( n11765 & ~n11760 ) | ( n11765 & n11773 ) | ( ~n11760 & n11773 ) ;
  assign n12299 = ( n11760 & n12296 ) | ( n11760 & n12297 ) | ( n12296 & n12297 ) ;
  assign n12298 = ( n11773 & ~n12297 ) | ( n11773 & n12296 ) | ( ~n12297 & n12296 ) ;
  assign n12300 = ( n11765 & ~n12299 ) | ( n11765 & n12298 ) | ( ~n12299 & n12298 ) ;
  assign n12281 = n11771 | n12187 ;
  assign n12282 = ( n11758 & ~n11771 ) | ( n11758 & n11767 ) | ( ~n11771 & n11767 ) ;
  assign n12284 = ( n11771 & n12281 ) | ( n11771 & n12282 ) | ( n12281 & n12282 ) ;
  assign n12283 = ( n11767 & ~n12282 ) | ( n11767 & n12281 ) | ( ~n12282 & n12281 ) ;
  assign n12285 = ( n11758 & ~n12284 ) | ( n11758 & n12283 ) | ( ~n12284 & n12283 ) ;
  assign n12274 = n11738 | n12187 ;
  assign n12275 = ( n11738 & ~n11751 ) | ( n11738 & n11743 ) | ( ~n11751 & n11743 ) ;
  assign n12276 = ( n11751 & n12274 ) | ( n11751 & n12275 ) | ( n12274 & n12275 ) ;
  assign n12277 = ( n11738 & ~n12275 ) | ( n11738 & n12274 ) | ( ~n12275 & n12274 ) ;
  assign n12278 = ( n11743 & ~n12276 ) | ( n11743 & n12277 ) | ( ~n12276 & n12277 ) ;
  assign n12259 = n11749 | n12187 ;
  assign n12260 = ( n11736 & ~n11745 ) | ( n11736 & n11749 ) | ( ~n11745 & n11749 ) ;
  assign n12261 = ( n11745 & n12259 ) | ( n11745 & n12260 ) | ( n12259 & n12260 ) ;
  assign n12262 = ( n11749 & ~n12260 ) | ( n11749 & n12259 ) | ( ~n12260 & n12259 ) ;
  assign n12263 = ( n11736 & ~n12261 ) | ( n11736 & n12262 ) | ( ~n12261 & n12262 ) ;
  assign n12252 = ( n11716 & ~n12187 ) | ( n11716 & 1'b0 ) | ( ~n12187 & 1'b0 ) ;
  assign n12253 = ( n11716 & n11721 ) | ( n11716 & n11729 ) | ( n11721 & n11729 ) ;
  assign n12254 = ( n12252 & ~n11729 ) | ( n12252 & n12253 ) | ( ~n11729 & n12253 ) ;
  assign n12255 = ( n11716 & ~n12253 ) | ( n11716 & n12252 ) | ( ~n12253 & n12252 ) ;
  assign n12256 = ( n11721 & ~n12254 ) | ( n11721 & n12255 ) | ( ~n12254 & n12255 ) ;
  assign n12237 = n11727 | n12187 ;
  assign n12238 = ( n11714 & ~n11723 ) | ( n11714 & n11727 ) | ( ~n11723 & n11727 ) ;
  assign n12239 = ( n11723 & n12237 ) | ( n11723 & n12238 ) | ( n12237 & n12238 ) ;
  assign n12240 = ( n11727 & ~n12238 ) | ( n11727 & n12237 ) | ( ~n12238 & n12237 ) ;
  assign n12241 = ( n11714 & ~n12239 ) | ( n11714 & n12240 ) | ( ~n12239 & n12240 ) ;
  assign n12230 = ( n11690 & ~n11692 ) | ( n11690 & 1'b0 ) | ( ~n11692 & 1'b0 ) ;
  assign n12231 = ( n11692 & ~n12230 ) | ( n11692 & n11702 ) | ( ~n12230 & n11702 ) ;
  assign n12233 = ( n12187 & n12230 ) | ( n12187 & n12231 ) | ( n12230 & n12231 ) ;
  assign n12232 = ( n11692 & ~n12231 ) | ( n11692 & n12187 ) | ( ~n12231 & n12187 ) ;
  assign n12234 = ( n11702 & ~n12233 ) | ( n11702 & n12232 ) | ( ~n12233 & n12232 ) ;
  assign n12214 = ~x38 & n11674 ;
  assign n12215 = ( x39 & ~n12214 ) | ( x39 & 1'b0 ) | ( ~n12214 & 1'b0 ) ;
  assign n12216 = n11693 | n12215 ;
  assign n12211 = ( n11674 & ~x38 ) | ( n11674 & n11685 ) | ( ~x38 & n11685 ) ;
  assign n12212 = x38 &  n12211 ;
  assign n12213 = ( n11680 & ~n12212 ) | ( n11680 & n11685 ) | ( ~n12212 & n11685 ) ;
  assign n12217 = ( n12187 & ~n12216 ) | ( n12187 & n12213 ) | ( ~n12216 & n12213 ) ;
  assign n12219 = ( n12187 & ~n12217 ) | ( n12187 & 1'b0 ) | ( ~n12217 & 1'b0 ) ;
  assign n12218 = ~n12213 & n12217 ;
  assign n12220 = ( n12216 & ~n12219 ) | ( n12216 & n12218 ) | ( ~n12219 & n12218 ) ;
  assign n12200 = ( n11674 & ~n12184 ) | ( n11674 & 1'b0 ) | ( ~n12184 & 1'b0 ) ;
  assign n12201 = ( n12175 & ~n12200 ) | ( n12175 & n12179 ) | ( ~n12200 & n12179 ) ;
  assign n12202 = ( n12175 & ~n12201 ) | ( n12175 & 1'b0 ) | ( ~n12201 & 1'b0 ) ;
  assign n12203 = n12167 &  n12202 ;
  assign n12199 = ~n11677 & n12187 ;
  assign n12204 = ( n12199 & ~n12203 ) | ( n12199 & 1'b0 ) | ( ~n12203 & 1'b0 ) ;
  assign n12205 = ( x38 & n12203 ) | ( x38 & n12204 ) | ( n12203 & n12204 ) ;
  assign n12206 = x38 | n12203 ;
  assign n12207 = n12199 | n12206 ;
  assign n12208 = ~n12205 & n12207 ;
  assign n12190 = ( x36 & ~n12187 ) | ( x36 & x37 ) | ( ~n12187 & x37 ) ;
  assign n12196 = ( x36 & ~x37 ) | ( x36 & 1'b0 ) | ( ~x37 & 1'b0 ) ;
  assign n11675 = x34 | x35 ;
  assign n12191 = ~x36 & n11675 ;
  assign n12192 = ( x36 & ~n11672 ) | ( x36 & n12191 ) | ( ~n11672 & n12191 ) ;
  assign n12193 = ( n11662 & ~n11654 ) | ( n11662 & n12192 ) | ( ~n11654 & n12192 ) ;
  assign n12194 = n11654 &  n12193 ;
  assign n12195 = ( n12187 & ~x37 ) | ( n12187 & n12194 ) | ( ~x37 & n12194 ) ;
  assign n12197 = ( n12190 & ~n12196 ) | ( n12190 & n12195 ) | ( ~n12196 & n12195 ) ;
  assign n11676 = x36 | n11675 ;
  assign n12188 = x36 &  n12187 ;
  assign n12189 = ( n11674 & ~n11676 ) | ( n11674 & n12188 ) | ( ~n11676 & n12188 ) ;
  assign n12221 = n11176 | n12189 ;
  assign n12222 = ( n12197 & ~n12221 ) | ( n12197 & 1'b0 ) | ( ~n12221 & 1'b0 ) ;
  assign n12223 = n12208 | n12222 ;
  assign n12224 = n12189 &  n12197 ;
  assign n12225 = ( n11176 & ~n12197 ) | ( n11176 & n12224 ) | ( ~n12197 & n12224 ) ;
  assign n12226 = n10685 | n12225 ;
  assign n12227 = ( n12223 & ~n12226 ) | ( n12223 & 1'b0 ) | ( ~n12226 & 1'b0 ) ;
  assign n12228 = n12220 | n12227 ;
  assign n12198 = ~n12189 & n12197 ;
  assign n12209 = ( n12198 & ~n11176 ) | ( n12198 & n12208 ) | ( ~n11176 & n12208 ) ;
  assign n12210 = ( n10685 & ~n12209 ) | ( n10685 & 1'b0 ) | ( ~n12209 & 1'b0 ) ;
  assign n12242 = n10209 | n12210 ;
  assign n12243 = ( n12228 & ~n12242 ) | ( n12228 & 1'b0 ) | ( ~n12242 & 1'b0 ) ;
  assign n12244 = n12234 | n12243 ;
  assign n12245 = ( n12223 & ~n12225 ) | ( n12223 & 1'b0 ) | ( ~n12225 & 1'b0 ) ;
  assign n12246 = ( n12220 & ~n10685 ) | ( n12220 & n12245 ) | ( ~n10685 & n12245 ) ;
  assign n12247 = ( n10209 & ~n12246 ) | ( n10209 & 1'b0 ) | ( ~n12246 & 1'b0 ) ;
  assign n12248 = ( n9740 & ~n12247 ) | ( n9740 & 1'b0 ) | ( ~n12247 & 1'b0 ) ;
  assign n12249 = n12244 &  n12248 ;
  assign n12250 = n12241 | n12249 ;
  assign n12229 = ~n12210 & n12228 ;
  assign n12235 = ( n12229 & ~n10209 ) | ( n12229 & n12234 ) | ( ~n10209 & n12234 ) ;
  assign n12236 = n9740 | n12235 ;
  assign n12264 = ~n9286 & n12236 ;
  assign n12265 = n12250 &  n12264 ;
  assign n12266 = n12256 | n12265 ;
  assign n12267 = ( n12244 & ~n12247 ) | ( n12244 & 1'b0 ) | ( ~n12247 & 1'b0 ) ;
  assign n12268 = ( n9740 & n12241 ) | ( n9740 & n12267 ) | ( n12241 & n12267 ) ;
  assign n12269 = ( n9286 & ~n12268 ) | ( n9286 & 1'b0 ) | ( ~n12268 & 1'b0 ) ;
  assign n12270 = n8839 | n12269 ;
  assign n12271 = ( n12266 & ~n12270 ) | ( n12266 & 1'b0 ) | ( ~n12270 & 1'b0 ) ;
  assign n12272 = n12263 | n12271 ;
  assign n12251 = n12236 &  n12250 ;
  assign n12257 = ( n12251 & ~n9286 ) | ( n12251 & n12256 ) | ( ~n9286 & n12256 ) ;
  assign n12258 = ( n8839 & ~n12257 ) | ( n8839 & 1'b0 ) | ( ~n12257 & 1'b0 ) ;
  assign n12286 = n8407 | n12258 ;
  assign n12287 = ( n12272 & ~n12286 ) | ( n12272 & 1'b0 ) | ( ~n12286 & 1'b0 ) ;
  assign n12288 = n12278 | n12287 ;
  assign n12289 = ( n12266 & ~n12269 ) | ( n12266 & 1'b0 ) | ( ~n12269 & 1'b0 ) ;
  assign n12290 = ( n12263 & ~n8839 ) | ( n12263 & n12289 ) | ( ~n8839 & n12289 ) ;
  assign n12291 = ( n8407 & ~n12290 ) | ( n8407 & 1'b0 ) | ( ~n12290 & 1'b0 ) ;
  assign n12292 = n7982 | n12291 ;
  assign n12293 = ( n12288 & ~n12292 ) | ( n12288 & 1'b0 ) | ( ~n12292 & 1'b0 ) ;
  assign n12294 = n12285 | n12293 ;
  assign n12273 = ~n12258 & n12272 ;
  assign n12279 = ( n12273 & ~n8407 ) | ( n12273 & n12278 ) | ( ~n8407 & n12278 ) ;
  assign n12280 = ( n7982 & ~n12279 ) | ( n7982 & 1'b0 ) | ( ~n12279 & 1'b0 ) ;
  assign n12308 = ( n7572 & ~n12280 ) | ( n7572 & 1'b0 ) | ( ~n12280 & 1'b0 ) ;
  assign n12309 = n12294 &  n12308 ;
  assign n12310 = n12300 | n12309 ;
  assign n12311 = ( n12288 & ~n12291 ) | ( n12288 & 1'b0 ) | ( ~n12291 & 1'b0 ) ;
  assign n12312 = ( n12285 & ~n7982 ) | ( n12285 & n12311 ) | ( ~n7982 & n12311 ) ;
  assign n12313 = n7572 | n12312 ;
  assign n12314 = n7169 &  n12313 ;
  assign n12315 = n12310 &  n12314 ;
  assign n12316 = ( n12307 & ~n12315 ) | ( n12307 & 1'b0 ) | ( ~n12315 & 1'b0 ) ;
  assign n12295 = ~n12280 & n12294 ;
  assign n12301 = ( n7572 & n12295 ) | ( n7572 & n12300 ) | ( n12295 & n12300 ) ;
  assign n12302 = n7169 | n12301 ;
  assign n12330 = ~n6781 & n12302 ;
  assign n12331 = ~n12316 & n12330 ;
  assign n12332 = ( n12322 & ~n12331 ) | ( n12322 & 1'b0 ) | ( ~n12331 & 1'b0 ) ;
  assign n12333 = n12310 &  n12313 ;
  assign n12334 = ( n7169 & ~n12307 ) | ( n7169 & n12333 ) | ( ~n12307 & n12333 ) ;
  assign n12335 = ( n6781 & ~n12334 ) | ( n6781 & 1'b0 ) | ( ~n12334 & 1'b0 ) ;
  assign n12336 = ( n6399 & ~n12335 ) | ( n6399 & 1'b0 ) | ( ~n12335 & 1'b0 ) ;
  assign n12337 = ~n12332 & n12336 ;
  assign n12338 = ( n12329 & ~n12337 ) | ( n12329 & 1'b0 ) | ( ~n12337 & 1'b0 ) ;
  assign n12317 = ( n12302 & ~n12316 ) | ( n12302 & 1'b0 ) | ( ~n12316 & 1'b0 ) ;
  assign n12323 = ( n6781 & ~n12317 ) | ( n6781 & n12322 ) | ( ~n12317 & n12322 ) ;
  assign n12324 = ~n6399 & n12323 ;
  assign n12352 = n6032 | n12324 ;
  assign n12353 = n12338 | n12352 ;
  assign n12354 = n12344 &  n12353 ;
  assign n12355 = n12332 | n12335 ;
  assign n12356 = ( n12329 & ~n6399 ) | ( n12329 & n12355 ) | ( ~n6399 & n12355 ) ;
  assign n12357 = n6032 &  n12356 ;
  assign n12358 = ( n5672 & ~n12357 ) | ( n5672 & 1'b0 ) | ( ~n12357 & 1'b0 ) ;
  assign n12359 = ~n12354 & n12358 ;
  assign n12360 = ( n12351 & ~n12359 ) | ( n12351 & 1'b0 ) | ( ~n12359 & 1'b0 ) ;
  assign n12339 = n12324 | n12338 ;
  assign n12345 = ( n6032 & n12339 ) | ( n6032 & n12344 ) | ( n12339 & n12344 ) ;
  assign n12346 = ~n5672 & n12345 ;
  assign n12374 = n5327 | n12346 ;
  assign n12375 = n12360 | n12374 ;
  assign n12376 = ~n12366 & n12375 ;
  assign n12377 = n12354 | n12357 ;
  assign n12378 = ( n12351 & ~n5672 ) | ( n12351 & n12377 ) | ( ~n5672 & n12377 ) ;
  assign n12379 = n5327 &  n12378 ;
  assign n12380 = n4990 | n12379 ;
  assign n12381 = n12376 | n12380 ;
  assign n12382 = ~n12373 & n12381 ;
  assign n12361 = n12346 | n12360 ;
  assign n12367 = ( n5327 & ~n12366 ) | ( n5327 & n12361 ) | ( ~n12366 & n12361 ) ;
  assign n12368 = n4990 &  n12367 ;
  assign n12396 = n4668 | n12368 ;
  assign n12397 = n12382 | n12396 ;
  assign n12398 = n12388 &  n12397 ;
  assign n12399 = n12376 | n12379 ;
  assign n12400 = ( n4990 & ~n12373 ) | ( n4990 & n12399 ) | ( ~n12373 & n12399 ) ;
  assign n12401 = n4668 &  n12400 ;
  assign n12402 = n4353 | n12401 ;
  assign n12403 = n12398 | n12402 ;
  assign n12404 = ~n12395 & n12403 ;
  assign n12383 = n12368 | n12382 ;
  assign n12389 = ( n4668 & n12383 ) | ( n4668 & n12388 ) | ( n12383 & n12388 ) ;
  assign n12390 = n4353 &  n12389 ;
  assign n12418 = n4053 | n12390 ;
  assign n12419 = n12404 | n12418 ;
  assign n12420 = n12410 &  n12419 ;
  assign n12421 = n12398 | n12401 ;
  assign n12422 = ( n4353 & ~n12395 ) | ( n4353 & n12421 ) | ( ~n12395 & n12421 ) ;
  assign n12423 = n4053 &  n12422 ;
  assign n12424 = n3760 | n12423 ;
  assign n12425 = n12420 | n12424 ;
  assign n12426 = n12417 &  n12425 ;
  assign n12405 = n12390 | n12404 ;
  assign n12411 = ( n4053 & n12405 ) | ( n4053 & n12410 ) | ( n12405 & n12410 ) ;
  assign n12412 = n3760 &  n12411 ;
  assign n12440 = n3482 | n12412 ;
  assign n12441 = n12426 | n12440 ;
  assign n12442 = ~n12432 & n12441 ;
  assign n12443 = n12420 | n12423 ;
  assign n12444 = ( n3760 & n12417 ) | ( n3760 & n12443 ) | ( n12417 & n12443 ) ;
  assign n12445 = n3482 &  n12444 ;
  assign n12446 = n3211 | n12445 ;
  assign n12447 = n12442 | n12446 ;
  assign n12448 = ~n12439 & n12447 ;
  assign n12427 = n12412 | n12426 ;
  assign n12433 = ( n3482 & ~n12432 ) | ( n3482 & n12427 ) | ( ~n12432 & n12427 ) ;
  assign n12434 = n3211 &  n12433 ;
  assign n12462 = n2955 | n12434 ;
  assign n12463 = n12448 | n12462 ;
  assign n12464 = ~n12454 & n12463 ;
  assign n12465 = n12442 | n12445 ;
  assign n12466 = ( n3211 & ~n12439 ) | ( n3211 & n12465 ) | ( ~n12439 & n12465 ) ;
  assign n12467 = n2955 &  n12466 ;
  assign n12468 = n2706 | n12467 ;
  assign n12469 = n12464 | n12468 ;
  assign n12470 = ~n12461 & n12469 ;
  assign n12449 = n12434 | n12448 ;
  assign n12455 = ( n2955 & ~n12454 ) | ( n2955 & n12449 ) | ( ~n12454 & n12449 ) ;
  assign n12456 = n2706 &  n12455 ;
  assign n12484 = n2472 | n12456 ;
  assign n12485 = n12470 | n12484 ;
  assign n12486 = ~n12476 & n12485 ;
  assign n12487 = n12464 | n12467 ;
  assign n12488 = ( n2706 & ~n12461 ) | ( n2706 & n12487 ) | ( ~n12461 & n12487 ) ;
  assign n12489 = n2472 &  n12488 ;
  assign n12490 = n2245 | n12489 ;
  assign n12491 = n12486 | n12490 ;
  assign n12625 = ~n12102 & n12187 ;
  assign n12626 = ( n12089 & n12094 ) | ( n12089 & n12187 ) | ( n12094 & n12187 ) ;
  assign n12628 = ( n12625 & ~n12089 ) | ( n12625 & n12626 ) | ( ~n12089 & n12626 ) ;
  assign n12627 = ( n12187 & ~n12626 ) | ( n12187 & n12625 ) | ( ~n12626 & n12625 ) ;
  assign n12629 = ( n12094 & ~n12628 ) | ( n12094 & n12627 ) | ( ~n12628 & n12627 ) ;
  assign n12582 = ( n12045 & ~n12050 ) | ( n12045 & n12187 ) | ( ~n12050 & n12187 ) ;
  assign n12581 = n12058 &  n12187 ;
  assign n12583 = ( n12187 & ~n12582 ) | ( n12187 & n12581 ) | ( ~n12582 & n12581 ) ;
  assign n12584 = ( n12581 & ~n12045 ) | ( n12581 & n12582 ) | ( ~n12045 & n12582 ) ;
  assign n12585 = ( n12050 & ~n12583 ) | ( n12050 & n12584 ) | ( ~n12583 & n12584 ) ;
  assign n12516 = ( n11979 & ~n11984 ) | ( n11979 & n12187 ) | ( ~n11984 & n12187 ) ;
  assign n12515 = n11992 &  n12187 ;
  assign n12517 = ( n12187 & ~n12516 ) | ( n12187 & n12515 ) | ( ~n12516 & n12515 ) ;
  assign n12518 = ( n12515 & ~n11979 ) | ( n12515 & n12516 ) | ( ~n11979 & n12516 ) ;
  assign n12519 = ( n11984 & ~n12517 ) | ( n11984 & n12518 ) | ( ~n12517 & n12518 ) ;
  assign n12471 = n12456 | n12470 ;
  assign n12477 = ( n2472 & ~n12476 ) | ( n2472 & n12471 ) | ( ~n12476 & n12471 ) ;
  assign n12478 = n2245 &  n12477 ;
  assign n12492 = n12483 &  n12491 ;
  assign n12493 = n12478 | n12492 ;
  assign n12494 = ~n11971 & n12187 ;
  assign n12495 = ( n11958 & n11963 ) | ( n11958 & n12187 ) | ( n11963 & n12187 ) ;
  assign n12497 = ( n12494 & ~n11958 ) | ( n12494 & n12495 ) | ( ~n11958 & n12495 ) ;
  assign n12496 = ( n12187 & ~n12495 ) | ( n12187 & n12494 ) | ( ~n12495 & n12494 ) ;
  assign n12498 = ( n11963 & ~n12497 ) | ( n11963 & n12496 ) | ( ~n12497 & n12496 ) ;
  assign n12499 = ( n2033 & ~n12493 ) | ( n2033 & n12498 ) | ( ~n12493 & n12498 ) ;
  assign n12500 = ( n1827 & ~n12499 ) | ( n1827 & 1'b0 ) | ( ~n12499 & 1'b0 ) ;
  assign n12501 = ( n2033 & ~n12478 ) | ( n2033 & 1'b0 ) | ( ~n12478 & 1'b0 ) ;
  assign n12502 = ~n12492 & n12501 ;
  assign n12503 = n12498 | n12502 ;
  assign n12504 = n12486 | n12489 ;
  assign n12505 = ( n2245 & n12483 ) | ( n2245 & n12504 ) | ( n12483 & n12504 ) ;
  assign n12506 = ~n2033 & n12505 ;
  assign n12507 = n1827 | n12506 ;
  assign n12508 = ( n12503 & ~n12507 ) | ( n12503 & 1'b0 ) | ( ~n12507 & 1'b0 ) ;
  assign n12509 = ( n11977 & ~n11986 ) | ( n11977 & n11990 ) | ( ~n11986 & n11990 ) ;
  assign n12510 = ( n11986 & n12187 ) | ( n11986 & n12509 ) | ( n12187 & n12509 ) ;
  assign n12511 = ( n11990 & ~n12509 ) | ( n11990 & n12187 ) | ( ~n12509 & n12187 ) ;
  assign n12512 = ( n11977 & ~n12510 ) | ( n11977 & n12511 ) | ( ~n12510 & n12511 ) ;
  assign n12513 = n12508 | n12512 ;
  assign n12514 = ~n12500 & n12513 ;
  assign n12520 = ( n1636 & ~n12519 ) | ( n1636 & n12514 ) | ( ~n12519 & n12514 ) ;
  assign n12521 = n1452 | n12520 ;
  assign n12522 = n12012 | n12187 ;
  assign n12523 = ( n11999 & ~n12012 ) | ( n11999 & n12008 ) | ( ~n12012 & n12008 ) ;
  assign n12525 = ( n12012 & n12522 ) | ( n12012 & n12523 ) | ( n12522 & n12523 ) ;
  assign n12524 = ( n12008 & ~n12523 ) | ( n12008 & n12522 ) | ( ~n12523 & n12522 ) ;
  assign n12526 = ( n11999 & ~n12525 ) | ( n11999 & n12524 ) | ( ~n12525 & n12524 ) ;
  assign n12527 = ( n1636 & ~n12500 ) | ( n1636 & 1'b0 ) | ( ~n12500 & 1'b0 ) ;
  assign n12528 = n12513 &  n12527 ;
  assign n12529 = ( n12519 & ~n12528 ) | ( n12519 & 1'b0 ) | ( ~n12528 & 1'b0 ) ;
  assign n12530 = ( n12503 & ~n12506 ) | ( n12503 & 1'b0 ) | ( ~n12506 & 1'b0 ) ;
  assign n12531 = ( n12512 & ~n1827 ) | ( n12512 & n12530 ) | ( ~n1827 & n12530 ) ;
  assign n12532 = n1636 | n12531 ;
  assign n12533 = n1452 &  n12532 ;
  assign n12534 = ~n12529 & n12533 ;
  assign n12535 = n12526 | n12534 ;
  assign n12536 = n12521 &  n12535 ;
  assign n12537 = n12014 &  n12187 ;
  assign n12538 = ( n12001 & ~n12187 ) | ( n12001 & n12006 ) | ( ~n12187 & n12006 ) ;
  assign n12539 = ( n12187 & n12537 ) | ( n12187 & n12538 ) | ( n12537 & n12538 ) ;
  assign n12540 = ( n12001 & ~n12538 ) | ( n12001 & n12537 ) | ( ~n12538 & n12537 ) ;
  assign n12541 = ( n12006 & ~n12539 ) | ( n12006 & n12540 ) | ( ~n12539 & n12540 ) ;
  assign n12542 = ( n1283 & ~n12536 ) | ( n1283 & n12541 ) | ( ~n12536 & n12541 ) ;
  assign n12543 = ~n1122 & n12542 ;
  assign n12544 = n12034 | n12187 ;
  assign n12545 = ( n12021 & ~n12030 ) | ( n12021 & n12034 ) | ( ~n12030 & n12034 ) ;
  assign n12546 = ( n12030 & n12544 ) | ( n12030 & n12545 ) | ( n12544 & n12545 ) ;
  assign n12547 = ( n12034 & ~n12545 ) | ( n12034 & n12544 ) | ( ~n12545 & n12544 ) ;
  assign n12548 = ( n12021 & ~n12546 ) | ( n12021 & n12547 ) | ( ~n12546 & n12547 ) ;
  assign n12549 = ~n1283 & n12521 ;
  assign n12550 = n12535 &  n12549 ;
  assign n12551 = ( n12541 & ~n12550 ) | ( n12541 & 1'b0 ) | ( ~n12550 & 1'b0 ) ;
  assign n12552 = ~n12529 & n12532 ;
  assign n12553 = ( n1452 & n12526 ) | ( n1452 & n12552 ) | ( n12526 & n12552 ) ;
  assign n12554 = ( n1283 & ~n12553 ) | ( n1283 & 1'b0 ) | ( ~n12553 & 1'b0 ) ;
  assign n12555 = ( n1122 & ~n12554 ) | ( n1122 & 1'b0 ) | ( ~n12554 & 1'b0 ) ;
  assign n12556 = ~n12551 & n12555 ;
  assign n12557 = ( n12548 & ~n12556 ) | ( n12548 & 1'b0 ) | ( ~n12556 & 1'b0 ) ;
  assign n12558 = n12543 | n12557 ;
  assign n12560 = ( n12023 & ~n12028 ) | ( n12023 & n12187 ) | ( ~n12028 & n12187 ) ;
  assign n12559 = n12036 &  n12187 ;
  assign n12561 = ( n12187 & ~n12560 ) | ( n12187 & n12559 ) | ( ~n12560 & n12559 ) ;
  assign n12562 = ( n12559 & ~n12023 ) | ( n12559 & n12560 ) | ( ~n12023 & n12560 ) ;
  assign n12563 = ( n12028 & ~n12561 ) | ( n12028 & n12562 ) | ( ~n12561 & n12562 ) ;
  assign n12564 = ( n976 & ~n12558 ) | ( n976 & n12563 ) | ( ~n12558 & n12563 ) ;
  assign n12565 = ( n837 & ~n12564 ) | ( n837 & 1'b0 ) | ( ~n12564 & 1'b0 ) ;
  assign n12567 = ( n12052 & ~n12043 ) | ( n12052 & n12056 ) | ( ~n12043 & n12056 ) ;
  assign n12566 = ( n12056 & ~n12187 ) | ( n12056 & 1'b0 ) | ( ~n12187 & 1'b0 ) ;
  assign n12569 = ( n12056 & ~n12567 ) | ( n12056 & n12566 ) | ( ~n12567 & n12566 ) ;
  assign n12568 = ( n12566 & ~n12052 ) | ( n12566 & n12567 ) | ( ~n12052 & n12567 ) ;
  assign n12570 = ( n12043 & ~n12569 ) | ( n12043 & n12568 ) | ( ~n12569 & n12568 ) ;
  assign n12571 = ( n976 & ~n12543 ) | ( n976 & 1'b0 ) | ( ~n12543 & 1'b0 ) ;
  assign n12572 = ~n12557 & n12571 ;
  assign n12573 = n12563 | n12572 ;
  assign n12574 = n12551 | n12554 ;
  assign n12575 = ( n12548 & ~n1122 ) | ( n12548 & n12574 ) | ( ~n1122 & n12574 ) ;
  assign n12576 = ~n976 & n12575 ;
  assign n12577 = n837 | n12576 ;
  assign n12578 = ( n12573 & ~n12577 ) | ( n12573 & 1'b0 ) | ( ~n12577 & 1'b0 ) ;
  assign n12579 = ( n12570 & ~n12578 ) | ( n12570 & 1'b0 ) | ( ~n12578 & 1'b0 ) ;
  assign n12580 = n12565 | n12579 ;
  assign n12586 = ( n713 & ~n12585 ) | ( n713 & n12580 ) | ( ~n12585 & n12580 ) ;
  assign n12587 = n595 &  n12586 ;
  assign n12588 = n12078 | n12187 ;
  assign n12589 = ( n12065 & ~n12078 ) | ( n12065 & n12074 ) | ( ~n12078 & n12074 ) ;
  assign n12591 = ( n12078 & n12588 ) | ( n12078 & n12589 ) | ( n12588 & n12589 ) ;
  assign n12590 = ( n12074 & ~n12589 ) | ( n12074 & n12588 ) | ( ~n12589 & n12588 ) ;
  assign n12592 = ( n12065 & ~n12591 ) | ( n12065 & n12590 ) | ( ~n12591 & n12590 ) ;
  assign n12593 = n713 | n12565 ;
  assign n12594 = n12579 | n12593 ;
  assign n12595 = ~n12585 & n12594 ;
  assign n12596 = ( n12573 & ~n12576 ) | ( n12573 & 1'b0 ) | ( ~n12576 & 1'b0 ) ;
  assign n12597 = ( n837 & ~n12596 ) | ( n837 & n12570 ) | ( ~n12596 & n12570 ) ;
  assign n12598 = n713 &  n12597 ;
  assign n12599 = n595 | n12598 ;
  assign n12600 = n12595 | n12599 ;
  assign n12601 = ~n12592 & n12600 ;
  assign n12602 = n12587 | n12601 ;
  assign n12603 = n12080 &  n12187 ;
  assign n12604 = ( n12067 & n12072 ) | ( n12067 & n12187 ) | ( n12072 & n12187 ) ;
  assign n12606 = ( n12603 & ~n12067 ) | ( n12603 & n12604 ) | ( ~n12067 & n12604 ) ;
  assign n12605 = ( n12187 & ~n12604 ) | ( n12187 & n12603 ) | ( ~n12604 & n12603 ) ;
  assign n12607 = ( n12072 & ~n12606 ) | ( n12072 & n12605 ) | ( ~n12606 & n12605 ) ;
  assign n12608 = ( n492 & n12602 ) | ( n492 & n12607 ) | ( n12602 & n12607 ) ;
  assign n12609 = n396 &  n12608 ;
  assign n12610 = n12100 | n12187 ;
  assign n12611 = ( n12087 & n12096 ) | ( n12087 & n12100 ) | ( n12096 & n12100 ) ;
  assign n12612 = ( n12610 & ~n12096 ) | ( n12610 & n12611 ) | ( ~n12096 & n12611 ) ;
  assign n12613 = ( n12100 & ~n12611 ) | ( n12100 & n12610 ) | ( ~n12611 & n12610 ) ;
  assign n12614 = ( n12087 & ~n12612 ) | ( n12087 & n12613 ) | ( ~n12612 & n12613 ) ;
  assign n12615 = n492 | n12587 ;
  assign n12616 = n12601 | n12615 ;
  assign n12617 = n12607 &  n12616 ;
  assign n12618 = n12595 | n12598 ;
  assign n12619 = ( n595 & ~n12592 ) | ( n595 & n12618 ) | ( ~n12592 & n12618 ) ;
  assign n12620 = n492 &  n12619 ;
  assign n12621 = n396 | n12620 ;
  assign n12622 = n12617 | n12621 ;
  assign n12623 = n12614 &  n12622 ;
  assign n12624 = n12609 | n12623 ;
  assign n12630 = ( n315 & ~n12629 ) | ( n315 & n12624 ) | ( ~n12629 & n12624 ) ;
  assign n12631 = n240 &  n12630 ;
  assign n12632 = n12122 | n12187 ;
  assign n12633 = ( n12109 & n12118 ) | ( n12109 & n12122 ) | ( n12118 & n12122 ) ;
  assign n12634 = ( n12632 & ~n12118 ) | ( n12632 & n12633 ) | ( ~n12118 & n12633 ) ;
  assign n12635 = ( n12122 & ~n12633 ) | ( n12122 & n12632 ) | ( ~n12633 & n12632 ) ;
  assign n12636 = ( n12109 & ~n12634 ) | ( n12109 & n12635 ) | ( ~n12634 & n12635 ) ;
  assign n12637 = n315 | n12609 ;
  assign n12638 = n12623 | n12637 ;
  assign n12639 = ~n12629 & n12638 ;
  assign n12640 = n12617 | n12620 ;
  assign n12641 = ( n396 & n12614 ) | ( n396 & n12640 ) | ( n12614 & n12640 ) ;
  assign n12642 = n315 &  n12641 ;
  assign n12643 = n240 | n12642 ;
  assign n12644 = n12639 | n12643 ;
  assign n12645 = n12636 &  n12644 ;
  assign n12646 = n12631 | n12645 ;
  assign n12648 = ( n12111 & ~n12116 ) | ( n12111 & n12187 ) | ( ~n12116 & n12187 ) ;
  assign n12647 = ~n12124 & n12187 ;
  assign n12649 = ( n12187 & ~n12648 ) | ( n12187 & n12647 ) | ( ~n12648 & n12647 ) ;
  assign n12650 = ( n12647 & ~n12111 ) | ( n12647 & n12648 ) | ( ~n12111 & n12648 ) ;
  assign n12651 = ( n12116 & ~n12649 ) | ( n12116 & n12650 ) | ( ~n12649 & n12650 ) ;
  assign n12652 = ( n181 & n12646 ) | ( n181 & n12651 ) | ( n12646 & n12651 ) ;
  assign n12653 = ~n145 & n12652 ;
  assign n12654 = n12144 | n12187 ;
  assign n12655 = ( n12131 & n12140 ) | ( n12131 & n12144 ) | ( n12140 & n12144 ) ;
  assign n12656 = ( n12654 & ~n12140 ) | ( n12654 & n12655 ) | ( ~n12140 & n12655 ) ;
  assign n12657 = ( n12144 & ~n12655 ) | ( n12144 & n12654 ) | ( ~n12655 & n12654 ) ;
  assign n12658 = ( n12131 & ~n12656 ) | ( n12131 & n12657 ) | ( ~n12656 & n12657 ) ;
  assign n12659 = n181 | n12631 ;
  assign n12660 = n12645 | n12659 ;
  assign n12661 = n12651 &  n12660 ;
  assign n12662 = n12639 | n12642 ;
  assign n12663 = ( n240 & n12636 ) | ( n240 & n12662 ) | ( n12636 & n12662 ) ;
  assign n12664 = n181 &  n12663 ;
  assign n12665 = ( n145 & ~n12664 ) | ( n145 & 1'b0 ) | ( ~n12664 & 1'b0 ) ;
  assign n12666 = ~n12661 & n12665 ;
  assign n12667 = n12658 | n12666 ;
  assign n12668 = ~n12653 & n12667 ;
  assign n12669 = n12133 | n12187 ;
  assign n12670 = ( n12138 & ~n12133 ) | ( n12138 & n12146 ) | ( ~n12133 & n12146 ) ;
  assign n12672 = ( n12133 & n12669 ) | ( n12133 & n12670 ) | ( n12669 & n12670 ) ;
  assign n12671 = ( n12146 & ~n12670 ) | ( n12146 & n12669 ) | ( ~n12670 & n12669 ) ;
  assign n12673 = ( n12138 & ~n12672 ) | ( n12138 & n12671 ) | ( ~n12672 & n12671 ) ;
  assign n12674 = ( n150 & ~n12668 ) | ( n150 & n12673 ) | ( ~n12668 & n12673 ) ;
  assign n12675 = ( n12153 & ~n12172 ) | ( n12153 & 1'b0 ) | ( ~n12172 & 1'b0 ) ;
  assign n12676 = ( n12187 & ~n12169 ) | ( n12187 & n12675 ) | ( ~n12169 & n12675 ) ;
  assign n12677 = n12169 &  n12676 ;
  assign n12678 = ( n12169 & ~n12172 ) | ( n12169 & 1'b0 ) | ( ~n12172 & 1'b0 ) ;
  assign n12679 = ~n12187 & n12678 ;
  assign n12680 = ( n12153 & ~n12679 ) | ( n12153 & n12678 ) | ( ~n12679 & n12678 ) ;
  assign n12681 = ~n12677 & n12680 ;
  assign n12682 = n12154 &  n12161 ;
  assign n12683 = ~n12187 & n12682 ;
  assign n12684 = ( n12175 & ~n12682 ) | ( n12175 & n12683 ) | ( ~n12682 & n12683 ) ;
  assign n12685 = ~n12681 & n12684 ;
  assign n12686 = ~n12674 & n12685 ;
  assign n12687 = ( n133 & ~n12686 ) | ( n133 & n12685 ) | ( ~n12686 & n12685 ) ;
  assign n12690 = n12661 | n12664 ;
  assign n12691 = ( n145 & ~n12690 ) | ( n145 & n12658 ) | ( ~n12690 & n12658 ) ;
  assign n12692 = ( n150 & ~n12691 ) | ( n150 & 1'b0 ) | ( ~n12691 & 1'b0 ) ;
  assign n12693 = ( n12681 & ~n12692 ) | ( n12681 & 1'b0 ) | ( ~n12692 & 1'b0 ) ;
  assign n12688 = n150 | n12653 ;
  assign n12689 = ( n12667 & ~n12688 ) | ( n12667 & 1'b0 ) | ( ~n12688 & 1'b0 ) ;
  assign n12694 = n12673 &  n12689 ;
  assign n12695 = ( n12693 & ~n12673 ) | ( n12693 & n12694 ) | ( ~n12673 & n12694 ) ;
  assign n12697 = ( n133 & n12154 ) | ( n133 & n12161 ) | ( n12154 & n12161 ) ;
  assign n12696 = ( n12154 & ~n12187 ) | ( n12154 & n12161 ) | ( ~n12187 & n12161 ) ;
  assign n12698 = ( n12161 & ~n12696 ) | ( n12161 & 1'b0 ) | ( ~n12696 & 1'b0 ) ;
  assign n12699 = ( n12697 & ~n12161 ) | ( n12697 & n12698 ) | ( ~n12161 & n12698 ) ;
  assign n12700 = n12157 | n12184 ;
  assign n12701 = ( n12179 & ~n12160 ) | ( n12179 & n12700 ) | ( ~n12160 & n12700 ) ;
  assign n12702 = n12160 | n12701 ;
  assign n12703 = ( n12167 & ~n12175 ) | ( n12167 & n12702 ) | ( ~n12175 & n12702 ) ;
  assign n12704 = ( n12167 & ~n12703 ) | ( n12167 & 1'b0 ) | ( ~n12703 & 1'b0 ) ;
  assign n12705 = n12699 | n12704 ;
  assign n12706 = n12695 | n12705 ;
  assign n12707 = ~n12687 |  n12706 ;
  assign n13029 = ~n12491 & n12707 ;
  assign n13030 = ( n12478 & n12483 ) | ( n12478 & n12707 ) | ( n12483 & n12707 ) ;
  assign n13032 = ( n13029 & ~n12478 ) | ( n13029 & n13030 ) | ( ~n12478 & n13030 ) ;
  assign n13031 = ( n12707 & ~n13030 ) | ( n12707 & n13029 ) | ( ~n13030 & n13029 ) ;
  assign n13033 = ( n12483 & ~n13032 ) | ( n12483 & n13031 ) | ( ~n13032 & n13031 ) ;
  assign n13015 = ( n12485 & ~n12476 ) | ( n12485 & n12489 ) | ( ~n12476 & n12489 ) ;
  assign n13014 = n12489 | n12707 ;
  assign n13017 = ( n12489 & ~n13015 ) | ( n12489 & n13014 ) | ( ~n13015 & n13014 ) ;
  assign n13016 = ( n13014 & ~n12485 ) | ( n13014 & n13015 ) | ( ~n12485 & n13015 ) ;
  assign n13018 = ( n12476 & ~n13017 ) | ( n12476 & n13016 ) | ( ~n13017 & n13016 ) ;
  assign n13008 = ( n12456 & ~n12461 ) | ( n12456 & n12707 ) | ( ~n12461 & n12707 ) ;
  assign n13007 = ~n12469 & n12707 ;
  assign n13009 = ( n12707 & ~n13008 ) | ( n12707 & n13007 ) | ( ~n13008 & n13007 ) ;
  assign n13010 = ( n13007 & ~n12456 ) | ( n13007 & n13008 ) | ( ~n12456 & n13008 ) ;
  assign n13011 = ( n12461 & ~n13009 ) | ( n12461 & n13010 ) | ( ~n13009 & n13010 ) ;
  assign n12993 = ( n12463 & ~n12454 ) | ( n12463 & n12467 ) | ( ~n12454 & n12467 ) ;
  assign n12992 = n12467 | n12707 ;
  assign n12995 = ( n12467 & ~n12993 ) | ( n12467 & n12992 ) | ( ~n12993 & n12992 ) ;
  assign n12994 = ( n12992 & ~n12463 ) | ( n12992 & n12993 ) | ( ~n12463 & n12993 ) ;
  assign n12996 = ( n12454 & ~n12995 ) | ( n12454 & n12994 ) | ( ~n12995 & n12994 ) ;
  assign n12986 = ( n12434 & ~n12439 ) | ( n12434 & n12707 ) | ( ~n12439 & n12707 ) ;
  assign n12985 = ~n12447 & n12707 ;
  assign n12987 = ( n12707 & ~n12986 ) | ( n12707 & n12985 ) | ( ~n12986 & n12985 ) ;
  assign n12988 = ( n12985 & ~n12434 ) | ( n12985 & n12986 ) | ( ~n12434 & n12986 ) ;
  assign n12989 = ( n12439 & ~n12987 ) | ( n12439 & n12988 ) | ( ~n12987 & n12988 ) ;
  assign n12971 = ( n12441 & ~n12432 ) | ( n12441 & n12445 ) | ( ~n12432 & n12445 ) ;
  assign n12970 = n12445 | n12707 ;
  assign n12973 = ( n12445 & ~n12971 ) | ( n12445 & n12970 ) | ( ~n12971 & n12970 ) ;
  assign n12972 = ( n12970 & ~n12441 ) | ( n12970 & n12971 ) | ( ~n12441 & n12971 ) ;
  assign n12974 = ( n12432 & ~n12973 ) | ( n12432 & n12972 ) | ( ~n12973 & n12972 ) ;
  assign n12963 = n12412 | n12707 ;
  assign n12964 = ( n12412 & n12417 ) | ( n12412 & n12425 ) | ( n12417 & n12425 ) ;
  assign n12965 = ( n12963 & ~n12425 ) | ( n12963 & n12964 ) | ( ~n12425 & n12964 ) ;
  assign n12966 = ( n12412 & ~n12964 ) | ( n12412 & n12963 ) | ( ~n12964 & n12963 ) ;
  assign n12967 = ( n12417 & ~n12965 ) | ( n12417 & n12966 ) | ( ~n12965 & n12966 ) ;
  assign n12949 = ( n12419 & ~n12410 ) | ( n12419 & n12423 ) | ( ~n12410 & n12423 ) ;
  assign n12948 = n12423 | n12707 ;
  assign n12951 = ( n12423 & ~n12949 ) | ( n12423 & n12948 ) | ( ~n12949 & n12948 ) ;
  assign n12950 = ( n12948 & ~n12419 ) | ( n12948 & n12949 ) | ( ~n12419 & n12949 ) ;
  assign n12952 = ( n12410 & ~n12951 ) | ( n12410 & n12950 ) | ( ~n12951 & n12950 ) ;
  assign n12942 = ( n12390 & ~n12395 ) | ( n12390 & n12403 ) | ( ~n12395 & n12403 ) ;
  assign n12941 = n12390 | n12707 ;
  assign n12944 = ( n12390 & ~n12942 ) | ( n12390 & n12941 ) | ( ~n12942 & n12941 ) ;
  assign n12943 = ( n12941 & ~n12403 ) | ( n12941 & n12942 ) | ( ~n12403 & n12942 ) ;
  assign n12945 = ( n12395 & ~n12944 ) | ( n12395 & n12943 ) | ( ~n12944 & n12943 ) ;
  assign n12927 = ( n12397 & ~n12388 ) | ( n12397 & n12401 ) | ( ~n12388 & n12401 ) ;
  assign n12926 = n12401 | n12707 ;
  assign n12929 = ( n12401 & ~n12927 ) | ( n12401 & n12926 ) | ( ~n12927 & n12926 ) ;
  assign n12928 = ( n12926 & ~n12397 ) | ( n12926 & n12927 ) | ( ~n12397 & n12927 ) ;
  assign n12930 = ( n12388 & ~n12929 ) | ( n12388 & n12928 ) | ( ~n12929 & n12928 ) ;
  assign n12920 = ( n12368 & ~n12373 ) | ( n12368 & n12381 ) | ( ~n12373 & n12381 ) ;
  assign n12919 = n12368 | n12707 ;
  assign n12922 = ( n12368 & ~n12920 ) | ( n12368 & n12919 ) | ( ~n12920 & n12919 ) ;
  assign n12921 = ( n12919 & ~n12381 ) | ( n12919 & n12920 ) | ( ~n12381 & n12920 ) ;
  assign n12923 = ( n12373 & ~n12922 ) | ( n12373 & n12921 ) | ( ~n12922 & n12921 ) ;
  assign n12904 = n12379 | n12707 ;
  assign n12905 = ( n12366 & n12375 ) | ( n12366 & n12379 ) | ( n12375 & n12379 ) ;
  assign n12906 = ( n12904 & ~n12375 ) | ( n12904 & n12905 ) | ( ~n12375 & n12905 ) ;
  assign n12907 = ( n12379 & ~n12905 ) | ( n12379 & n12904 ) | ( ~n12905 & n12904 ) ;
  assign n12908 = ( n12366 & ~n12906 ) | ( n12366 & n12907 ) | ( ~n12906 & n12907 ) ;
  assign n12897 = n12346 | n12707 ;
  assign n12898 = ( n12346 & ~n12359 ) | ( n12346 & n12351 ) | ( ~n12359 & n12351 ) ;
  assign n12899 = ( n12359 & n12897 ) | ( n12359 & n12898 ) | ( n12897 & n12898 ) ;
  assign n12900 = ( n12346 & ~n12898 ) | ( n12346 & n12897 ) | ( ~n12898 & n12897 ) ;
  assign n12901 = ( n12351 & ~n12899 ) | ( n12351 & n12900 ) | ( ~n12899 & n12900 ) ;
  assign n12883 = ( n12353 & ~n12344 ) | ( n12353 & n12357 ) | ( ~n12344 & n12357 ) ;
  assign n12882 = n12357 | n12707 ;
  assign n12885 = ( n12357 & ~n12883 ) | ( n12357 & n12882 ) | ( ~n12883 & n12882 ) ;
  assign n12884 = ( n12882 & ~n12353 ) | ( n12882 & n12883 ) | ( ~n12353 & n12883 ) ;
  assign n12886 = ( n12344 & ~n12885 ) | ( n12344 & n12884 ) | ( ~n12885 & n12884 ) ;
  assign n12875 = n12324 | n12707 ;
  assign n12876 = ( n12324 & ~n12337 ) | ( n12324 & n12329 ) | ( ~n12337 & n12329 ) ;
  assign n12877 = ( n12337 & n12875 ) | ( n12337 & n12876 ) | ( n12875 & n12876 ) ;
  assign n12878 = ( n12324 & ~n12876 ) | ( n12324 & n12875 ) | ( ~n12876 & n12875 ) ;
  assign n12879 = ( n12329 & ~n12877 ) | ( n12329 & n12878 ) | ( ~n12877 & n12878 ) ;
  assign n12860 = n12335 | n12707 ;
  assign n12861 = ( n12322 & ~n12335 ) | ( n12322 & n12331 ) | ( ~n12335 & n12331 ) ;
  assign n12863 = ( n12335 & n12860 ) | ( n12335 & n12861 ) | ( n12860 & n12861 ) ;
  assign n12862 = ( n12331 & ~n12861 ) | ( n12331 & n12860 ) | ( ~n12861 & n12860 ) ;
  assign n12864 = ( n12322 & ~n12863 ) | ( n12322 & n12862 ) | ( ~n12863 & n12862 ) ;
  assign n12854 = ( n12302 & ~n12307 ) | ( n12302 & n12315 ) | ( ~n12307 & n12315 ) ;
  assign n12853 = ( n12302 & ~n12707 ) | ( n12302 & 1'b0 ) | ( ~n12707 & 1'b0 ) ;
  assign n12856 = ( n12302 & ~n12854 ) | ( n12302 & n12853 ) | ( ~n12854 & n12853 ) ;
  assign n12855 = ( n12853 & ~n12315 ) | ( n12853 & n12854 ) | ( ~n12315 & n12854 ) ;
  assign n12857 = ( n12307 & ~n12856 ) | ( n12307 & n12855 ) | ( ~n12856 & n12855 ) ;
  assign n12839 = ( n12309 & ~n12300 ) | ( n12309 & n12313 ) | ( ~n12300 & n12313 ) ;
  assign n12838 = ( n12313 & ~n12707 ) | ( n12313 & 1'b0 ) | ( ~n12707 & 1'b0 ) ;
  assign n12841 = ( n12313 & ~n12839 ) | ( n12313 & n12838 ) | ( ~n12839 & n12838 ) ;
  assign n12840 = ( n12838 & ~n12309 ) | ( n12838 & n12839 ) | ( ~n12309 & n12839 ) ;
  assign n12842 = ( n12300 & ~n12841 ) | ( n12300 & n12840 ) | ( ~n12841 & n12840 ) ;
  assign n12831 = n12280 | n12707 ;
  assign n12832 = ( n12285 & ~n12280 ) | ( n12285 & n12293 ) | ( ~n12280 & n12293 ) ;
  assign n12834 = ( n12280 & n12831 ) | ( n12280 & n12832 ) | ( n12831 & n12832 ) ;
  assign n12833 = ( n12293 & ~n12832 ) | ( n12293 & n12831 ) | ( ~n12832 & n12831 ) ;
  assign n12835 = ( n12285 & ~n12834 ) | ( n12285 & n12833 ) | ( ~n12834 & n12833 ) ;
  assign n12816 = n12291 | n12707 ;
  assign n12817 = ( n12278 & ~n12287 ) | ( n12278 & n12291 ) | ( ~n12287 & n12291 ) ;
  assign n12818 = ( n12287 & n12816 ) | ( n12287 & n12817 ) | ( n12816 & n12817 ) ;
  assign n12819 = ( n12291 & ~n12817 ) | ( n12291 & n12816 ) | ( ~n12817 & n12816 ) ;
  assign n12820 = ( n12278 & ~n12818 ) | ( n12278 & n12819 ) | ( ~n12818 & n12819 ) ;
  assign n12809 = n12258 | n12707 ;
  assign n12810 = ( n12263 & ~n12258 ) | ( n12263 & n12271 ) | ( ~n12258 & n12271 ) ;
  assign n12812 = ( n12258 & n12809 ) | ( n12258 & n12810 ) | ( n12809 & n12810 ) ;
  assign n12811 = ( n12271 & ~n12810 ) | ( n12271 & n12809 ) | ( ~n12810 & n12809 ) ;
  assign n12813 = ( n12263 & ~n12812 ) | ( n12263 & n12811 ) | ( ~n12812 & n12811 ) ;
  assign n12794 = n12269 | n12707 ;
  assign n12795 = ( n12256 & ~n12265 ) | ( n12256 & n12269 ) | ( ~n12265 & n12269 ) ;
  assign n12796 = ( n12265 & n12794 ) | ( n12265 & n12795 ) | ( n12794 & n12795 ) ;
  assign n12797 = ( n12269 & ~n12795 ) | ( n12269 & n12794 ) | ( ~n12795 & n12794 ) ;
  assign n12798 = ( n12256 & ~n12796 ) | ( n12256 & n12797 ) | ( ~n12796 & n12797 ) ;
  assign n12787 = n12249 &  n12707 ;
  assign n12788 = ( n12241 & ~n12236 ) | ( n12241 & n12707 ) | ( ~n12236 & n12707 ) ;
  assign n12790 = ( n12787 & n12236 ) | ( n12787 & n12788 ) | ( n12236 & n12788 ) ;
  assign n12789 = ( n12707 & ~n12788 ) | ( n12707 & n12787 ) | ( ~n12788 & n12787 ) ;
  assign n12791 = ( n12241 & ~n12790 ) | ( n12241 & n12789 ) | ( ~n12790 & n12789 ) ;
  assign n12772 = n12247 | n12707 ;
  assign n12773 = ( n12234 & ~n12247 ) | ( n12234 & n12243 ) | ( ~n12247 & n12243 ) ;
  assign n12775 = ( n12247 & n12772 ) | ( n12247 & n12773 ) | ( n12772 & n12773 ) ;
  assign n12774 = ( n12243 & ~n12773 ) | ( n12243 & n12772 ) | ( ~n12773 & n12772 ) ;
  assign n12776 = ( n12234 & ~n12775 ) | ( n12234 & n12774 ) | ( ~n12775 & n12774 ) ;
  assign n12765 = n12210 | n12707 ;
  assign n12766 = ( n12210 & ~n12227 ) | ( n12210 & n12220 ) | ( ~n12227 & n12220 ) ;
  assign n12767 = ( n12227 & n12765 ) | ( n12227 & n12766 ) | ( n12765 & n12766 ) ;
  assign n12768 = ( n12210 & ~n12766 ) | ( n12210 & n12765 ) | ( ~n12766 & n12765 ) ;
  assign n12769 = ( n12220 & ~n12767 ) | ( n12220 & n12768 ) | ( ~n12767 & n12768 ) ;
  assign n12750 = ~n12222 & n12225 ;
  assign n12751 = ( n12208 & ~n12222 ) | ( n12208 & n12750 ) | ( ~n12222 & n12750 ) ;
  assign n12753 = ( n12222 & n12707 ) | ( n12222 & n12751 ) | ( n12707 & n12751 ) ;
  assign n12752 = ( n12707 & ~n12751 ) | ( n12707 & n12750 ) | ( ~n12751 & n12750 ) ;
  assign n12754 = ( n12208 & ~n12753 ) | ( n12208 & n12752 ) | ( ~n12753 & n12752 ) ;
  assign n12741 = ~x36 & n12187 ;
  assign n12742 = ( x37 & ~n12741 ) | ( x37 & 1'b0 ) | ( ~n12741 & 1'b0 ) ;
  assign n12743 = n12199 | n12742 ;
  assign n12738 = ( n12187 & ~x36 ) | ( n12187 & n12194 ) | ( ~x36 & n12194 ) ;
  assign n12739 = x36 &  n12738 ;
  assign n12740 = ( n12189 & ~n12739 ) | ( n12189 & n12194 ) | ( ~n12739 & n12194 ) ;
  assign n12744 = ( n12707 & ~n12743 ) | ( n12707 & n12740 ) | ( ~n12743 & n12740 ) ;
  assign n12746 = ( n12707 & ~n12744 ) | ( n12707 & 1'b0 ) | ( ~n12744 & 1'b0 ) ;
  assign n12745 = ~n12740 & n12744 ;
  assign n12747 = ( n12743 & ~n12746 ) | ( n12743 & n12745 ) | ( ~n12746 & n12745 ) ;
  assign n12714 = ( x34 & ~n12707 ) | ( x34 & x35 ) | ( ~n12707 & x35 ) ;
  assign n12720 = ( x34 & ~x35 ) | ( x34 & 1'b0 ) | ( ~x35 & 1'b0 ) ;
  assign n12710 = x32 | x33 ;
  assign n12715 = ~x34 & n12710 ;
  assign n12716 = ( x34 & ~n12185 ) | ( x34 & n12715 ) | ( ~n12185 & n12715 ) ;
  assign n12717 = ( n12175 & ~n12167 ) | ( n12175 & n12716 ) | ( ~n12167 & n12716 ) ;
  assign n12718 = n12167 &  n12717 ;
  assign n12719 = ( n12707 & ~x35 ) | ( n12707 & n12718 ) | ( ~x35 & n12718 ) ;
  assign n12721 = ( n12714 & ~n12720 ) | ( n12714 & n12719 ) | ( ~n12720 & n12719 ) ;
  assign n12711 = x34 | n12710 ;
  assign n12712 = x34 &  n12707 ;
  assign n12713 = ( n12187 & ~n12711 ) | ( n12187 & n12712 ) | ( ~n12711 & n12712 ) ;
  assign n12724 = n11674 | n12713 ;
  assign n12725 = ( n12721 & ~n12724 ) | ( n12721 & 1'b0 ) | ( ~n12724 & 1'b0 ) ;
  assign n12727 = ( n12187 & ~n12704 ) | ( n12187 & 1'b0 ) | ( ~n12704 & 1'b0 ) ;
  assign n12728 = ( n12695 & ~n12699 ) | ( n12695 & n12727 ) | ( ~n12699 & n12727 ) ;
  assign n12729 = ~n12695 & n12728 ;
  assign n12730 = n12687 &  n12729 ;
  assign n12726 = ~n11675 & n12707 ;
  assign n12731 = ( n12726 & ~n12730 ) | ( n12726 & 1'b0 ) | ( ~n12730 & 1'b0 ) ;
  assign n12732 = ( x36 & n12730 ) | ( x36 & n12731 ) | ( n12730 & n12731 ) ;
  assign n12733 = x36 | n12730 ;
  assign n12734 = n12726 | n12733 ;
  assign n12735 = ~n12732 & n12734 ;
  assign n12736 = n12725 | n12735 ;
  assign n12722 = n12713 &  n12721 ;
  assign n12723 = ( n11674 & ~n12721 ) | ( n11674 & n12722 ) | ( ~n12721 & n12722 ) ;
  assign n12755 = n11176 | n12723 ;
  assign n12756 = ( n12736 & ~n12755 ) | ( n12736 & 1'b0 ) | ( ~n12755 & 1'b0 ) ;
  assign n12757 = n12747 | n12756 ;
  assign n12758 = ~n12713 & n12721 ;
  assign n12759 = ( n12735 & ~n11674 ) | ( n12735 & n12758 ) | ( ~n11674 & n12758 ) ;
  assign n12760 = ( n11176 & ~n12759 ) | ( n11176 & 1'b0 ) | ( ~n12759 & 1'b0 ) ;
  assign n12761 = n10685 | n12760 ;
  assign n12762 = ( n12757 & ~n12761 ) | ( n12757 & 1'b0 ) | ( ~n12761 & 1'b0 ) ;
  assign n12763 = n12754 | n12762 ;
  assign n12737 = ~n12723 & n12736 ;
  assign n12748 = ( n12737 & ~n11176 ) | ( n12737 & n12747 ) | ( ~n11176 & n12747 ) ;
  assign n12749 = ( n10685 & ~n12748 ) | ( n10685 & 1'b0 ) | ( ~n12748 & 1'b0 ) ;
  assign n12777 = n10209 | n12749 ;
  assign n12778 = ( n12763 & ~n12777 ) | ( n12763 & 1'b0 ) | ( ~n12777 & 1'b0 ) ;
  assign n12779 = n12769 | n12778 ;
  assign n12780 = ( n12757 & ~n12760 ) | ( n12757 & 1'b0 ) | ( ~n12760 & 1'b0 ) ;
  assign n12781 = ( n12754 & ~n10685 ) | ( n12754 & n12780 ) | ( ~n10685 & n12780 ) ;
  assign n12782 = ( n10209 & ~n12781 ) | ( n10209 & 1'b0 ) | ( ~n12781 & 1'b0 ) ;
  assign n12783 = ( n9740 & ~n12782 ) | ( n9740 & 1'b0 ) | ( ~n12782 & 1'b0 ) ;
  assign n12784 = n12779 &  n12783 ;
  assign n12785 = n12776 | n12784 ;
  assign n12764 = ~n12749 & n12763 ;
  assign n12770 = ( n12764 & ~n10209 ) | ( n12764 & n12769 ) | ( ~n10209 & n12769 ) ;
  assign n12771 = n9740 | n12770 ;
  assign n12799 = ~n9286 & n12771 ;
  assign n12800 = n12785 &  n12799 ;
  assign n12801 = n12791 | n12800 ;
  assign n12802 = ( n12779 & ~n12782 ) | ( n12779 & 1'b0 ) | ( ~n12782 & 1'b0 ) ;
  assign n12803 = ( n9740 & n12776 ) | ( n9740 & n12802 ) | ( n12776 & n12802 ) ;
  assign n12804 = ( n9286 & ~n12803 ) | ( n9286 & 1'b0 ) | ( ~n12803 & 1'b0 ) ;
  assign n12805 = n8839 | n12804 ;
  assign n12806 = ( n12801 & ~n12805 ) | ( n12801 & 1'b0 ) | ( ~n12805 & 1'b0 ) ;
  assign n12807 = n12798 | n12806 ;
  assign n12786 = n12771 &  n12785 ;
  assign n12792 = ( n12786 & ~n9286 ) | ( n12786 & n12791 ) | ( ~n9286 & n12791 ) ;
  assign n12793 = ( n8839 & ~n12792 ) | ( n8839 & 1'b0 ) | ( ~n12792 & 1'b0 ) ;
  assign n12821 = n8407 | n12793 ;
  assign n12822 = ( n12807 & ~n12821 ) | ( n12807 & 1'b0 ) | ( ~n12821 & 1'b0 ) ;
  assign n12823 = n12813 | n12822 ;
  assign n12824 = ( n12801 & ~n12804 ) | ( n12801 & 1'b0 ) | ( ~n12804 & 1'b0 ) ;
  assign n12825 = ( n12798 & ~n8839 ) | ( n12798 & n12824 ) | ( ~n8839 & n12824 ) ;
  assign n12826 = ( n8407 & ~n12825 ) | ( n8407 & 1'b0 ) | ( ~n12825 & 1'b0 ) ;
  assign n12827 = n7982 | n12826 ;
  assign n12828 = ( n12823 & ~n12827 ) | ( n12823 & 1'b0 ) | ( ~n12827 & 1'b0 ) ;
  assign n12829 = n12820 | n12828 ;
  assign n12808 = ~n12793 & n12807 ;
  assign n12814 = ( n12808 & ~n8407 ) | ( n12808 & n12813 ) | ( ~n8407 & n12813 ) ;
  assign n12815 = ( n7982 & ~n12814 ) | ( n7982 & 1'b0 ) | ( ~n12814 & 1'b0 ) ;
  assign n12843 = ( n7572 & ~n12815 ) | ( n7572 & 1'b0 ) | ( ~n12815 & 1'b0 ) ;
  assign n12844 = n12829 &  n12843 ;
  assign n12845 = n12835 | n12844 ;
  assign n12846 = ( n12823 & ~n12826 ) | ( n12823 & 1'b0 ) | ( ~n12826 & 1'b0 ) ;
  assign n12847 = ( n12820 & ~n7982 ) | ( n12820 & n12846 ) | ( ~n7982 & n12846 ) ;
  assign n12848 = n7572 | n12847 ;
  assign n12849 = n7169 &  n12848 ;
  assign n12850 = n12845 &  n12849 ;
  assign n12851 = n12842 | n12850 ;
  assign n12830 = ~n12815 & n12829 ;
  assign n12836 = ( n7572 & n12830 ) | ( n7572 & n12835 ) | ( n12830 & n12835 ) ;
  assign n12837 = n7169 | n12836 ;
  assign n12865 = ~n6781 & n12837 ;
  assign n12866 = n12851 &  n12865 ;
  assign n12867 = ( n12857 & ~n12866 ) | ( n12857 & 1'b0 ) | ( ~n12866 & 1'b0 ) ;
  assign n12868 = n12845 &  n12848 ;
  assign n12869 = ( n7169 & n12842 ) | ( n7169 & n12868 ) | ( n12842 & n12868 ) ;
  assign n12870 = ( n6781 & ~n12869 ) | ( n6781 & 1'b0 ) | ( ~n12869 & 1'b0 ) ;
  assign n12871 = ( n6399 & ~n12870 ) | ( n6399 & 1'b0 ) | ( ~n12870 & 1'b0 ) ;
  assign n12872 = ~n12867 & n12871 ;
  assign n12873 = ( n12864 & ~n12872 ) | ( n12864 & 1'b0 ) | ( ~n12872 & 1'b0 ) ;
  assign n12852 = n12837 &  n12851 ;
  assign n12858 = ( n6781 & ~n12852 ) | ( n6781 & n12857 ) | ( ~n12852 & n12857 ) ;
  assign n12859 = ~n6399 & n12858 ;
  assign n12887 = n6032 | n12859 ;
  assign n12888 = n12873 | n12887 ;
  assign n12889 = n12879 &  n12888 ;
  assign n12890 = n12867 | n12870 ;
  assign n12891 = ( n12864 & ~n6399 ) | ( n12864 & n12890 ) | ( ~n6399 & n12890 ) ;
  assign n12892 = n6032 &  n12891 ;
  assign n12893 = ( n5672 & ~n12892 ) | ( n5672 & 1'b0 ) | ( ~n12892 & 1'b0 ) ;
  assign n12894 = ~n12889 & n12893 ;
  assign n12895 = ( n12886 & ~n12894 ) | ( n12886 & 1'b0 ) | ( ~n12894 & 1'b0 ) ;
  assign n12874 = n12859 | n12873 ;
  assign n12880 = ( n6032 & n12874 ) | ( n6032 & n12879 ) | ( n12874 & n12879 ) ;
  assign n12881 = ~n5672 & n12880 ;
  assign n12909 = n5327 | n12881 ;
  assign n12910 = n12895 | n12909 ;
  assign n12911 = n12901 &  n12910 ;
  assign n12912 = n12889 | n12892 ;
  assign n12913 = ( n12886 & ~n5672 ) | ( n12886 & n12912 ) | ( ~n5672 & n12912 ) ;
  assign n12914 = n5327 &  n12913 ;
  assign n12915 = n4990 | n12914 ;
  assign n12916 = n12911 | n12915 ;
  assign n12917 = ~n12908 & n12916 ;
  assign n12896 = n12881 | n12895 ;
  assign n12902 = ( n5327 & n12896 ) | ( n5327 & n12901 ) | ( n12896 & n12901 ) ;
  assign n12903 = n4990 &  n12902 ;
  assign n12931 = n4668 | n12903 ;
  assign n12932 = n12917 | n12931 ;
  assign n12933 = ~n12923 & n12932 ;
  assign n12934 = n12911 | n12914 ;
  assign n12935 = ( n4990 & ~n12908 ) | ( n4990 & n12934 ) | ( ~n12908 & n12934 ) ;
  assign n12936 = n4668 &  n12935 ;
  assign n12937 = n4353 | n12936 ;
  assign n12938 = n12933 | n12937 ;
  assign n12939 = n12930 &  n12938 ;
  assign n12918 = n12903 | n12917 ;
  assign n12924 = ( n4668 & ~n12923 ) | ( n4668 & n12918 ) | ( ~n12923 & n12918 ) ;
  assign n12925 = n4353 &  n12924 ;
  assign n12953 = n4053 | n12925 ;
  assign n12954 = n12939 | n12953 ;
  assign n12955 = ~n12945 & n12954 ;
  assign n12956 = n12933 | n12936 ;
  assign n12957 = ( n4353 & n12930 ) | ( n4353 & n12956 ) | ( n12930 & n12956 ) ;
  assign n12958 = n4053 &  n12957 ;
  assign n12959 = n3760 | n12958 ;
  assign n12960 = n12955 | n12959 ;
  assign n12961 = n12952 &  n12960 ;
  assign n12940 = n12925 | n12939 ;
  assign n12946 = ( n4053 & ~n12945 ) | ( n4053 & n12940 ) | ( ~n12945 & n12940 ) ;
  assign n12947 = n3760 &  n12946 ;
  assign n12975 = n3482 | n12947 ;
  assign n12976 = n12961 | n12975 ;
  assign n12977 = n12967 &  n12976 ;
  assign n12978 = n12955 | n12958 ;
  assign n12979 = ( n3760 & n12952 ) | ( n3760 & n12978 ) | ( n12952 & n12978 ) ;
  assign n12980 = n3482 &  n12979 ;
  assign n12981 = n3211 | n12980 ;
  assign n12982 = n12977 | n12981 ;
  assign n12983 = ~n12974 & n12982 ;
  assign n12962 = n12947 | n12961 ;
  assign n12968 = ( n3482 & n12962 ) | ( n3482 & n12967 ) | ( n12962 & n12967 ) ;
  assign n12969 = n3211 &  n12968 ;
  assign n12997 = n2955 | n12969 ;
  assign n12998 = n12983 | n12997 ;
  assign n12999 = ~n12989 & n12998 ;
  assign n13000 = n12977 | n12980 ;
  assign n13001 = ( n3211 & ~n12974 ) | ( n3211 & n13000 ) | ( ~n12974 & n13000 ) ;
  assign n13002 = n2955 &  n13001 ;
  assign n13003 = n2706 | n13002 ;
  assign n13004 = n12999 | n13003 ;
  assign n13005 = ~n12996 & n13004 ;
  assign n12984 = n12969 | n12983 ;
  assign n12990 = ( n2955 & ~n12989 ) | ( n2955 & n12984 ) | ( ~n12989 & n12984 ) ;
  assign n12991 = n2706 &  n12990 ;
  assign n13019 = n2472 | n12991 ;
  assign n13020 = n13005 | n13019 ;
  assign n13021 = ~n13011 & n13020 ;
  assign n13022 = n12999 | n13002 ;
  assign n13023 = ( n2706 & ~n12996 ) | ( n2706 & n13022 ) | ( ~n12996 & n13022 ) ;
  assign n13024 = n2472 &  n13023 ;
  assign n13025 = n2245 | n13024 ;
  assign n13026 = n13021 | n13025 ;
  assign n13027 = ~n13018 & n13026 ;
  assign n13006 = n12991 | n13005 ;
  assign n13012 = ( n2472 & ~n13011 ) | ( n2472 & n13006 ) | ( ~n13011 & n13006 ) ;
  assign n13013 = n2245 &  n13012 ;
  assign n13041 = ( n2033 & ~n13013 ) | ( n2033 & 1'b0 ) | ( ~n13013 & 1'b0 ) ;
  assign n13042 = ~n13027 & n13041 ;
  assign n13044 = n13021 | n13024 ;
  assign n13045 = ( n2245 & ~n13018 ) | ( n2245 & n13044 ) | ( ~n13018 & n13044 ) ;
  assign n13046 = ~n2033 & n13045 ;
  assign n13204 = n12653 | n12707 ;
  assign n13205 = ( n12653 & ~n12666 ) | ( n12653 & n12658 ) | ( ~n12666 & n12658 ) ;
  assign n13206 = ( n12666 & n13204 ) | ( n12666 & n13205 ) | ( n13204 & n13205 ) ;
  assign n13207 = ( n12653 & ~n13205 ) | ( n12653 & n13204 ) | ( ~n13205 & n13204 ) ;
  assign n13208 = ( n12658 & ~n13206 ) | ( n12658 & n13207 ) | ( ~n13206 & n13207 ) ;
  assign n13138 = ~n12600 & n12707 ;
  assign n13139 = ( n12587 & ~n13138 ) | ( n12587 & n12707 ) | ( ~n13138 & n12707 ) ;
  assign n13140 = ( n12592 & ~n12587 ) | ( n12592 & n13139 ) | ( ~n12587 & n13139 ) ;
  assign n13141 = ( n12587 & ~n13139 ) | ( n12587 & n12592 ) | ( ~n13139 & n12592 ) ;
  assign n13142 = ( n13140 & ~n12592 ) | ( n13140 & n13141 ) | ( ~n12592 & n13141 ) ;
  assign n13094 = n12556 &  n12707 ;
  assign n13095 = ( n12543 & n12548 ) | ( n12543 & n12707 ) | ( n12548 & n12707 ) ;
  assign n13097 = ( n13094 & ~n12543 ) | ( n13094 & n13095 ) | ( ~n12543 & n13095 ) ;
  assign n13096 = ( n12707 & ~n13095 ) | ( n12707 & n13094 ) | ( ~n13095 & n13094 ) ;
  assign n13098 = ( n12548 & ~n13097 ) | ( n12548 & n13096 ) | ( ~n13097 & n13096 ) ;
  assign n13028 = n13013 | n13027 ;
  assign n13034 = ( n13028 & ~n2033 ) | ( n13028 & n13033 ) | ( ~n2033 & n13033 ) ;
  assign n13035 = n1827 &  n13034 ;
  assign n13036 = n12506 | n12707 ;
  assign n13037 = ( n12498 & ~n12506 ) | ( n12498 & n12502 ) | ( ~n12506 & n12502 ) ;
  assign n13039 = ( n12506 & n13036 ) | ( n12506 & n13037 ) | ( n13036 & n13037 ) ;
  assign n13038 = ( n12502 & ~n13037 ) | ( n12502 & n13036 ) | ( ~n13037 & n13036 ) ;
  assign n13040 = ( n12498 & ~n13039 ) | ( n12498 & n13038 ) | ( ~n13039 & n13038 ) ;
  assign n13043 = ( n13033 & ~n13042 ) | ( n13033 & 1'b0 ) | ( ~n13042 & 1'b0 ) ;
  assign n13047 = n1827 | n13046 ;
  assign n13048 = n13043 | n13047 ;
  assign n13049 = ~n13040 & n13048 ;
  assign n13050 = n13035 | n13049 ;
  assign n13051 = ( n12500 & ~n12508 ) | ( n12500 & n12512 ) | ( ~n12508 & n12512 ) ;
  assign n13052 = ( n12508 & n12707 ) | ( n12508 & n13051 ) | ( n12707 & n13051 ) ;
  assign n13053 = ( n12500 & ~n13051 ) | ( n12500 & n12707 ) | ( ~n13051 & n12707 ) ;
  assign n13054 = ( n12512 & ~n13052 ) | ( n12512 & n13053 ) | ( ~n13052 & n13053 ) ;
  assign n13055 = ( n1636 & ~n13050 ) | ( n1636 & n13054 ) | ( ~n13050 & n13054 ) ;
  assign n13056 = n1452 | n13055 ;
  assign n13058 = ( n12528 & ~n12519 ) | ( n12528 & n12532 ) | ( ~n12519 & n12532 ) ;
  assign n13057 = ( n12532 & ~n12707 ) | ( n12532 & 1'b0 ) | ( ~n12707 & 1'b0 ) ;
  assign n13060 = ( n12532 & ~n13058 ) | ( n12532 & n13057 ) | ( ~n13058 & n13057 ) ;
  assign n13059 = ( n13057 & ~n12528 ) | ( n13057 & n13058 ) | ( ~n12528 & n13058 ) ;
  assign n13061 = ( n12519 & ~n13060 ) | ( n12519 & n13059 ) | ( ~n13060 & n13059 ) ;
  assign n13062 = ( n1636 & ~n13035 ) | ( n1636 & 1'b0 ) | ( ~n13035 & 1'b0 ) ;
  assign n13063 = ~n13049 & n13062 ;
  assign n13064 = n13054 | n13063 ;
  assign n13065 = n13043 | n13046 ;
  assign n13066 = ( n1827 & ~n13040 ) | ( n1827 & n13065 ) | ( ~n13040 & n13065 ) ;
  assign n13067 = ~n1636 & n13066 ;
  assign n13068 = ( n1452 & ~n13067 ) | ( n1452 & 1'b0 ) | ( ~n13067 & 1'b0 ) ;
  assign n13069 = n13064 &  n13068 ;
  assign n13070 = ( n13061 & ~n13069 ) | ( n13061 & 1'b0 ) | ( ~n13069 & 1'b0 ) ;
  assign n13071 = ( n13056 & ~n13070 ) | ( n13056 & 1'b0 ) | ( ~n13070 & 1'b0 ) ;
  assign n13072 = n12534 &  n12707 ;
  assign n13073 = ( n12526 & ~n12521 ) | ( n12526 & n12707 ) | ( ~n12521 & n12707 ) ;
  assign n13075 = ( n12521 & n13072 ) | ( n12521 & n13073 ) | ( n13072 & n13073 ) ;
  assign n13074 = ( n12707 & ~n13073 ) | ( n12707 & n13072 ) | ( ~n13073 & n13072 ) ;
  assign n13076 = ( n12526 & ~n13075 ) | ( n12526 & n13074 ) | ( ~n13075 & n13074 ) ;
  assign n13077 = ( n13071 & ~n1283 ) | ( n13071 & n13076 ) | ( ~n1283 & n13076 ) ;
  assign n13078 = n1122 | n13077 ;
  assign n13079 = n12554 | n12707 ;
  assign n13080 = ( n12541 & ~n12550 ) | ( n12541 & n12554 ) | ( ~n12550 & n12554 ) ;
  assign n13081 = ( n12550 & n13079 ) | ( n12550 & n13080 ) | ( n13079 & n13080 ) ;
  assign n13082 = ( n12554 & ~n13080 ) | ( n12554 & n13079 ) | ( ~n13080 & n13079 ) ;
  assign n13083 = ( n12541 & ~n13081 ) | ( n12541 & n13082 ) | ( ~n13081 & n13082 ) ;
  assign n13084 = ~n1283 & n13056 ;
  assign n13085 = ~n13070 & n13084 ;
  assign n13086 = n13076 | n13085 ;
  assign n13087 = ( n13064 & ~n13067 ) | ( n13064 & 1'b0 ) | ( ~n13067 & 1'b0 ) ;
  assign n13088 = ( n1452 & ~n13061 ) | ( n1452 & n13087 ) | ( ~n13061 & n13087 ) ;
  assign n13089 = ( n1283 & ~n13088 ) | ( n1283 & 1'b0 ) | ( ~n13088 & 1'b0 ) ;
  assign n13090 = ( n1122 & ~n13089 ) | ( n1122 & 1'b0 ) | ( ~n13089 & 1'b0 ) ;
  assign n13091 = n13086 &  n13090 ;
  assign n13092 = ( n13083 & ~n13091 ) | ( n13083 & 1'b0 ) | ( ~n13091 & 1'b0 ) ;
  assign n13093 = ( n13078 & ~n13092 ) | ( n13078 & 1'b0 ) | ( ~n13092 & 1'b0 ) ;
  assign n13099 = ( n976 & ~n13098 ) | ( n976 & n13093 ) | ( ~n13098 & n13093 ) ;
  assign n13100 = ( n837 & ~n13099 ) | ( n837 & 1'b0 ) | ( ~n13099 & 1'b0 ) ;
  assign n13101 = n12576 | n12707 ;
  assign n13102 = ( n12563 & ~n12576 ) | ( n12563 & n12572 ) | ( ~n12576 & n12572 ) ;
  assign n13104 = ( n12576 & n13101 ) | ( n12576 & n13102 ) | ( n13101 & n13102 ) ;
  assign n13103 = ( n12572 & ~n13102 ) | ( n12572 & n13101 ) | ( ~n13102 & n13101 ) ;
  assign n13105 = ( n12563 & ~n13104 ) | ( n12563 & n13103 ) | ( ~n13104 & n13103 ) ;
  assign n13106 = n976 &  n13078 ;
  assign n13107 = ~n13092 & n13106 ;
  assign n13108 = ( n13098 & ~n13107 ) | ( n13098 & 1'b0 ) | ( ~n13107 & 1'b0 ) ;
  assign n13109 = ( n13086 & ~n13089 ) | ( n13086 & 1'b0 ) | ( ~n13089 & 1'b0 ) ;
  assign n13110 = ( n1122 & ~n13083 ) | ( n1122 & n13109 ) | ( ~n13083 & n13109 ) ;
  assign n13111 = n976 | n13110 ;
  assign n13112 = ~n837 & n13111 ;
  assign n13113 = ~n13108 & n13112 ;
  assign n13114 = n13105 | n13113 ;
  assign n13115 = ~n13100 & n13114 ;
  assign n13116 = n12578 &  n12707 ;
  assign n13117 = ( n12565 & n12570 ) | ( n12565 & n12707 ) | ( n12570 & n12707 ) ;
  assign n13119 = ( n13116 & ~n12565 ) | ( n13116 & n13117 ) | ( ~n12565 & n13117 ) ;
  assign n13118 = ( n12707 & ~n13117 ) | ( n12707 & n13116 ) | ( ~n13117 & n13116 ) ;
  assign n13120 = ( n12570 & ~n13119 ) | ( n12570 & n13118 ) | ( ~n13119 & n13118 ) ;
  assign n13121 = ( n713 & ~n13115 ) | ( n713 & n13120 ) | ( ~n13115 & n13120 ) ;
  assign n13122 = n595 &  n13121 ;
  assign n13124 = ( n12594 & ~n12585 ) | ( n12594 & n12598 ) | ( ~n12585 & n12598 ) ;
  assign n13123 = n12598 | n12707 ;
  assign n13126 = ( n12598 & ~n13124 ) | ( n12598 & n13123 ) | ( ~n13124 & n13123 ) ;
  assign n13125 = ( n13123 & ~n12594 ) | ( n13123 & n13124 ) | ( ~n12594 & n13124 ) ;
  assign n13127 = ( n12585 & ~n13126 ) | ( n12585 & n13125 ) | ( ~n13126 & n13125 ) ;
  assign n13128 = n713 | n13100 ;
  assign n13129 = ( n13114 & ~n13128 ) | ( n13114 & 1'b0 ) | ( ~n13128 & 1'b0 ) ;
  assign n13130 = ( n13120 & ~n13129 ) | ( n13120 & 1'b0 ) | ( ~n13129 & 1'b0 ) ;
  assign n13131 = ~n13108 & n13111 ;
  assign n13132 = ( n13105 & ~n837 ) | ( n13105 & n13131 ) | ( ~n837 & n13131 ) ;
  assign n13133 = ( n713 & ~n13132 ) | ( n713 & 1'b0 ) | ( ~n13132 & 1'b0 ) ;
  assign n13134 = n595 | n13133 ;
  assign n13135 = n13130 | n13134 ;
  assign n13136 = ~n13127 & n13135 ;
  assign n13137 = n13122 | n13136 ;
  assign n13143 = ( n492 & ~n13142 ) | ( n492 & n13137 ) | ( ~n13142 & n13137 ) ;
  assign n13144 = n396 &  n13143 ;
  assign n13145 = n12620 | n12707 ;
  assign n13146 = ( n12607 & n12616 ) | ( n12607 & n12620 ) | ( n12616 & n12620 ) ;
  assign n13147 = ( n13145 & ~n12616 ) | ( n13145 & n13146 ) | ( ~n12616 & n13146 ) ;
  assign n13148 = ( n12620 & ~n13146 ) | ( n12620 & n13145 ) | ( ~n13146 & n13145 ) ;
  assign n13149 = ( n12607 & ~n13147 ) | ( n12607 & n13148 ) | ( ~n13147 & n13148 ) ;
  assign n13150 = n492 | n13122 ;
  assign n13151 = n13136 | n13150 ;
  assign n13152 = ~n13142 & n13151 ;
  assign n13153 = n13130 | n13133 ;
  assign n13154 = ( n595 & ~n13127 ) | ( n595 & n13153 ) | ( ~n13127 & n13153 ) ;
  assign n13155 = n492 &  n13154 ;
  assign n13156 = n396 | n13155 ;
  assign n13157 = n13152 | n13156 ;
  assign n13158 = n13149 &  n13157 ;
  assign n13159 = n13144 | n13158 ;
  assign n13160 = ~n12622 & n12707 ;
  assign n13161 = ( n12609 & n12614 ) | ( n12609 & n12707 ) | ( n12614 & n12707 ) ;
  assign n13163 = ( n13160 & ~n12609 ) | ( n13160 & n13161 ) | ( ~n12609 & n13161 ) ;
  assign n13162 = ( n12707 & ~n13161 ) | ( n12707 & n13160 ) | ( ~n13161 & n13160 ) ;
  assign n13164 = ( n12614 & ~n13163 ) | ( n12614 & n13162 ) | ( ~n13163 & n13162 ) ;
  assign n13165 = ( n315 & n13159 ) | ( n315 & n13164 ) | ( n13159 & n13164 ) ;
  assign n13166 = n240 &  n13165 ;
  assign n13168 = ( n12638 & ~n12629 ) | ( n12638 & n12642 ) | ( ~n12629 & n12642 ) ;
  assign n13167 = n12642 | n12707 ;
  assign n13170 = ( n12642 & ~n13168 ) | ( n12642 & n13167 ) | ( ~n13168 & n13167 ) ;
  assign n13169 = ( n13167 & ~n12638 ) | ( n13167 & n13168 ) | ( ~n12638 & n13168 ) ;
  assign n13171 = ( n12629 & ~n13170 ) | ( n12629 & n13169 ) | ( ~n13170 & n13169 ) ;
  assign n13172 = n315 | n13144 ;
  assign n13173 = n13158 | n13172 ;
  assign n13174 = n13164 &  n13173 ;
  assign n13175 = n13152 | n13155 ;
  assign n13176 = ( n396 & n13149 ) | ( n396 & n13175 ) | ( n13149 & n13175 ) ;
  assign n13177 = n315 &  n13176 ;
  assign n13178 = n240 | n13177 ;
  assign n13179 = n13174 | n13178 ;
  assign n13180 = ~n13171 & n13179 ;
  assign n13181 = n13166 | n13180 ;
  assign n13183 = ( n12631 & ~n12636 ) | ( n12631 & n12707 ) | ( ~n12636 & n12707 ) ;
  assign n13182 = ~n12644 & n12707 ;
  assign n13184 = ( n12707 & ~n13183 ) | ( n12707 & n13182 ) | ( ~n13183 & n13182 ) ;
  assign n13185 = ( n13182 & ~n12631 ) | ( n13182 & n13183 ) | ( ~n12631 & n13183 ) ;
  assign n13186 = ( n12636 & ~n13184 ) | ( n12636 & n13185 ) | ( ~n13184 & n13185 ) ;
  assign n13187 = ( n181 & n13181 ) | ( n181 & n13186 ) | ( n13181 & n13186 ) ;
  assign n13188 = ~n145 & n13187 ;
  assign n13190 = ( n12660 & ~n12651 ) | ( n12660 & n12664 ) | ( ~n12651 & n12664 ) ;
  assign n13189 = n12664 | n12707 ;
  assign n13192 = ( n12664 & ~n13190 ) | ( n12664 & n13189 ) | ( ~n13190 & n13189 ) ;
  assign n13191 = ( n13189 & ~n12660 ) | ( n13189 & n13190 ) | ( ~n12660 & n13190 ) ;
  assign n13193 = ( n12651 & ~n13192 ) | ( n12651 & n13191 ) | ( ~n13192 & n13191 ) ;
  assign n13194 = n181 | n13166 ;
  assign n13195 = n13180 | n13194 ;
  assign n13196 = n13186 &  n13195 ;
  assign n13197 = n13174 | n13177 ;
  assign n13198 = ( n240 & ~n13171 ) | ( n240 & n13197 ) | ( ~n13171 & n13197 ) ;
  assign n13199 = n181 &  n13198 ;
  assign n13200 = ( n145 & ~n13199 ) | ( n145 & 1'b0 ) | ( ~n13199 & 1'b0 ) ;
  assign n13201 = ~n13196 & n13200 ;
  assign n13202 = ( n13193 & ~n13201 ) | ( n13193 & 1'b0 ) | ( ~n13201 & 1'b0 ) ;
  assign n13203 = n13188 | n13202 ;
  assign n13209 = ( n150 & ~n13208 ) | ( n150 & n13203 ) | ( ~n13208 & n13203 ) ;
  assign n13210 = n12673 | n12689 ;
  assign n13211 = ( n12692 & ~n13210 ) | ( n12692 & n12707 ) | ( ~n13210 & n12707 ) ;
  assign n13212 = ~n12692 & n13211 ;
  assign n13213 = n12689 | n12692 ;
  assign n13214 = n12707 | n13213 ;
  assign n13215 = ( n12673 & ~n13214 ) | ( n12673 & n13213 ) | ( ~n13214 & n13213 ) ;
  assign n13216 = n13212 | n13215 ;
  assign n13217 = ( n12674 & ~n12681 ) | ( n12674 & 1'b0 ) | ( ~n12681 & 1'b0 ) ;
  assign n13218 = ~n12707 & n13217 ;
  assign n13219 = ( n12695 & ~n13218 ) | ( n12695 & n13217 ) | ( ~n13218 & n13217 ) ;
  assign n13220 = ( n13216 & ~n13219 ) | ( n13216 & 1'b0 ) | ( ~n13219 & 1'b0 ) ;
  assign n13221 = ~n13209 & n13220 ;
  assign n13222 = ( n133 & ~n13221 ) | ( n133 & n13220 ) | ( ~n13221 & n13220 ) ;
  assign n13223 = n150 | n13188 ;
  assign n13224 = n13202 | n13223 ;
  assign n13229 = n13224 | n13208 ;
  assign n13225 = n13196 | n13199 ;
  assign n13226 = ( n13193 & ~n145 ) | ( n13193 & n13225 ) | ( ~n145 & n13225 ) ;
  assign n13227 = n150 &  n13226 ;
  assign n13228 = n13216 | n13227 ;
  assign n13230 = ( n13229 & ~n13208 ) | ( n13229 & n13228 ) | ( ~n13208 & n13228 ) ;
  assign n13232 = ( n133 & ~n12681 ) | ( n133 & n12674 ) | ( ~n12681 & n12674 ) ;
  assign n13231 = ( n12681 & ~n12674 ) | ( n12681 & n12707 ) | ( ~n12674 & n12707 ) ;
  assign n13233 = ~n12681 & n13231 ;
  assign n13234 = ( n12681 & n13232 ) | ( n12681 & n13233 ) | ( n13232 & n13233 ) ;
  assign n13235 = n12677 | n12704 ;
  assign n13236 = ( n12680 & n12699 ) | ( n12680 & n13235 ) | ( n12699 & n13235 ) ;
  assign n13237 = ( n12680 & ~n13236 ) | ( n12680 & 1'b0 ) | ( ~n13236 & 1'b0 ) ;
  assign n13238 = ( n12687 & ~n13237 ) | ( n12687 & n12695 ) | ( ~n13237 & n12695 ) ;
  assign n13239 = ( n12687 & ~n13238 ) | ( n12687 & 1'b0 ) | ( ~n13238 & 1'b0 ) ;
  assign n13240 = n13234 | n13239 ;
  assign n13241 = ( n13230 & ~n13240 ) | ( n13230 & 1'b0 ) | ( ~n13240 & 1'b0 ) ;
  assign n13242 = ~n13222 | ~n13241 ;
  assign n13578 = n13046 | n13242 ;
  assign n13579 = ( n13033 & ~n13042 ) | ( n13033 & n13046 ) | ( ~n13042 & n13046 ) ;
  assign n13580 = ( n13042 & n13578 ) | ( n13042 & n13579 ) | ( n13578 & n13579 ) ;
  assign n13581 = ( n13046 & ~n13579 ) | ( n13046 & n13578 ) | ( ~n13579 & n13578 ) ;
  assign n13582 = ( n13033 & ~n13580 ) | ( n13033 & n13581 ) | ( ~n13580 & n13581 ) ;
  assign n13724 = ~n13179 & n13242 ;
  assign n13725 = ( n13166 & ~n13724 ) | ( n13166 & n13242 ) | ( ~n13724 & n13242 ) ;
  assign n13726 = ( n13171 & ~n13166 ) | ( n13171 & n13725 ) | ( ~n13166 & n13725 ) ;
  assign n13727 = ( n13166 & ~n13725 ) | ( n13166 & n13171 ) | ( ~n13725 & n13171 ) ;
  assign n13728 = ( n13726 & ~n13171 ) | ( n13726 & n13727 ) | ( ~n13171 & n13727 ) ;
  assign n13680 = ~n13135 & n13242 ;
  assign n13681 = ( n13122 & ~n13680 ) | ( n13122 & n13242 ) | ( ~n13680 & n13242 ) ;
  assign n13682 = ( n13127 & ~n13122 ) | ( n13127 & n13681 ) | ( ~n13122 & n13681 ) ;
  assign n13683 = ( n13122 & ~n13681 ) | ( n13122 & n13127 ) | ( ~n13681 & n13127 ) ;
  assign n13684 = ( n13682 & ~n13127 ) | ( n13682 & n13683 ) | ( ~n13127 & n13683 ) ;
  assign n13659 = ( n13100 & ~n13105 ) | ( n13100 & n13242 ) | ( ~n13105 & n13242 ) ;
  assign n13658 = n13113 &  n13242 ;
  assign n13660 = ( n13242 & ~n13659 ) | ( n13242 & n13658 ) | ( ~n13659 & n13658 ) ;
  assign n13661 = ( n13658 & ~n13100 ) | ( n13658 & n13659 ) | ( ~n13100 & n13659 ) ;
  assign n13662 = ( n13105 & ~n13660 ) | ( n13105 & n13661 ) | ( ~n13660 & n13661 ) ;
  assign n13636 = n13091 &  n13242 ;
  assign n13637 = ( n13078 & ~n13242 ) | ( n13078 & n13636 ) | ( ~n13242 & n13636 ) ;
  assign n13638 = ( n13083 & ~n13078 ) | ( n13083 & n13637 ) | ( ~n13078 & n13637 ) ;
  assign n13639 = ( n13078 & ~n13637 ) | ( n13078 & n13083 ) | ( ~n13637 & n13083 ) ;
  assign n13640 = ( n13638 & ~n13083 ) | ( n13638 & n13639 ) | ( ~n13083 & n13639 ) ;
  assign n13549 = ~n13004 & n13242 ;
  assign n13550 = ( n12991 & n12996 ) | ( n12991 & n13242 ) | ( n12996 & n13242 ) ;
  assign n13552 = ( n13549 & ~n12991 ) | ( n13549 & n13550 ) | ( ~n12991 & n13550 ) ;
  assign n13551 = ( n13242 & ~n13550 ) | ( n13242 & n13549 ) | ( ~n13550 & n13549 ) ;
  assign n13553 = ( n12996 & ~n13552 ) | ( n12996 & n13551 ) | ( ~n13552 & n13551 ) ;
  assign n13528 = ( n12969 & ~n12974 ) | ( n12969 & n12982 ) | ( ~n12974 & n12982 ) ;
  assign n13527 = n12969 | n13242 ;
  assign n13530 = ( n12969 & ~n13528 ) | ( n12969 & n13527 ) | ( ~n13528 & n13527 ) ;
  assign n13529 = ( n13527 & ~n12982 ) | ( n13527 & n13528 ) | ( ~n12982 & n13528 ) ;
  assign n13531 = ( n12974 & ~n13530 ) | ( n12974 & n13529 ) | ( ~n13530 & n13529 ) ;
  assign n13462 = ( n12903 & ~n12908 ) | ( n12903 & n12916 ) | ( ~n12908 & n12916 ) ;
  assign n13461 = n12903 | n13242 ;
  assign n13464 = ( n12903 & ~n13462 ) | ( n12903 & n13461 ) | ( ~n13462 & n13461 ) ;
  assign n13463 = ( n13461 & ~n12916 ) | ( n13461 & n13462 ) | ( ~n12916 & n13462 ) ;
  assign n13465 = ( n12908 & ~n13464 ) | ( n12908 & n13463 ) | ( ~n13464 & n13463 ) ;
  assign n12708 = x30 | x31 ;
  assign n12709 = x32 | n12708 ;
  assign n13243 = x32 &  n13242 ;
  assign n13244 = ( n12707 & ~n12709 ) | ( n12707 & n13243 ) | ( ~n12709 & n13243 ) ;
  assign n13245 = ( x32 & ~n13242 ) | ( x32 & x33 ) | ( ~n13242 & x33 ) ;
  assign n13251 = ( x32 & ~x33 ) | ( x32 & 1'b0 ) | ( ~x33 & 1'b0 ) ;
  assign n13246 = ~x32 & n12708 ;
  assign n13247 = ( x32 & ~n12705 ) | ( x32 & n13246 ) | ( ~n12705 & n13246 ) ;
  assign n13248 = ( n12687 & ~n13247 ) | ( n12687 & n12695 ) | ( ~n13247 & n12695 ) ;
  assign n13249 = ( n12687 & ~n13248 ) | ( n12687 & 1'b0 ) | ( ~n13248 & 1'b0 ) ;
  assign n13250 = ( n13242 & ~x33 ) | ( n13242 & n13249 ) | ( ~x33 & n13249 ) ;
  assign n13252 = ( n13245 & ~n13251 ) | ( n13245 & n13250 ) | ( ~n13251 & n13250 ) ;
  assign n13253 = ~n13244 & n13252 ;
  assign n13255 = ( n12707 & ~n13239 ) | ( n12707 & 1'b0 ) | ( ~n13239 & 1'b0 ) ;
  assign n13256 = ( n13230 & ~n13255 ) | ( n13230 & n13234 ) | ( ~n13255 & n13234 ) ;
  assign n13257 = ( n13230 & ~n13256 ) | ( n13230 & 1'b0 ) | ( ~n13256 & 1'b0 ) ;
  assign n13258 = n13222 &  n13257 ;
  assign n13254 = ~n12710 & n13242 ;
  assign n13259 = ( n13254 & ~n13258 ) | ( n13254 & 1'b0 ) | ( ~n13258 & 1'b0 ) ;
  assign n13260 = ( x34 & n13258 ) | ( x34 & n13259 ) | ( n13258 & n13259 ) ;
  assign n13261 = x34 | n13258 ;
  assign n13262 = n13254 | n13261 ;
  assign n13263 = ~n13260 & n13262 ;
  assign n13264 = ( n13253 & ~n12187 ) | ( n13253 & n13263 ) | ( ~n12187 & n13263 ) ;
  assign n13265 = ( n11674 & ~n13264 ) | ( n11674 & 1'b0 ) | ( ~n13264 & 1'b0 ) ;
  assign n13269 = ~x34 & n12707 ;
  assign n13270 = ( x35 & ~n13269 ) | ( x35 & 1'b0 ) | ( ~n13269 & 1'b0 ) ;
  assign n13271 = n12726 | n13270 ;
  assign n13266 = ( n12707 & ~x34 ) | ( n12707 & n12718 ) | ( ~x34 & n12718 ) ;
  assign n13267 = x34 &  n13266 ;
  assign n13268 = ( n12713 & ~n13267 ) | ( n12713 & n12718 ) | ( ~n13267 & n12718 ) ;
  assign n13272 = ( n13242 & ~n13271 ) | ( n13242 & n13268 ) | ( ~n13271 & n13268 ) ;
  assign n13274 = ( n13242 & ~n13272 ) | ( n13242 & 1'b0 ) | ( ~n13272 & 1'b0 ) ;
  assign n13273 = ~n13268 & n13272 ;
  assign n13275 = ( n13271 & ~n13274 ) | ( n13271 & n13273 ) | ( ~n13274 & n13273 ) ;
  assign n13276 = n12187 | n13244 ;
  assign n13277 = ( n13252 & ~n13276 ) | ( n13252 & 1'b0 ) | ( ~n13276 & 1'b0 ) ;
  assign n13278 = n13263 | n13277 ;
  assign n13279 = n13244 &  n13252 ;
  assign n13280 = ( n12187 & ~n13252 ) | ( n12187 & n13279 ) | ( ~n13252 & n13279 ) ;
  assign n13281 = n11674 | n13280 ;
  assign n13282 = ( n13278 & ~n13281 ) | ( n13278 & 1'b0 ) | ( ~n13281 & 1'b0 ) ;
  assign n13283 = n13275 | n13282 ;
  assign n13284 = ~n13265 & n13283 ;
  assign n13285 = ( n12723 & ~n12725 ) | ( n12723 & 1'b0 ) | ( ~n12725 & 1'b0 ) ;
  assign n13286 = ( n12725 & ~n13285 ) | ( n12725 & n12735 ) | ( ~n13285 & n12735 ) ;
  assign n13288 = ( n13242 & n13285 ) | ( n13242 & n13286 ) | ( n13285 & n13286 ) ;
  assign n13287 = ( n12725 & ~n13286 ) | ( n12725 & n13242 ) | ( ~n13286 & n13242 ) ;
  assign n13289 = ( n12735 & ~n13288 ) | ( n12735 & n13287 ) | ( ~n13288 & n13287 ) ;
  assign n13290 = ( n13284 & ~n11176 ) | ( n13284 & n13289 ) | ( ~n11176 & n13289 ) ;
  assign n13291 = ( n10685 & ~n13290 ) | ( n10685 & 1'b0 ) | ( ~n13290 & 1'b0 ) ;
  assign n13292 = n12760 | n13242 ;
  assign n13293 = ( n12747 & ~n12756 ) | ( n12747 & n12760 ) | ( ~n12756 & n12760 ) ;
  assign n13294 = ( n12756 & n13292 ) | ( n12756 & n13293 ) | ( n13292 & n13293 ) ;
  assign n13295 = ( n12760 & ~n13293 ) | ( n12760 & n13292 ) | ( ~n13293 & n13292 ) ;
  assign n13296 = ( n12747 & ~n13294 ) | ( n12747 & n13295 ) | ( ~n13294 & n13295 ) ;
  assign n13297 = n11176 | n13265 ;
  assign n13298 = ( n13283 & ~n13297 ) | ( n13283 & 1'b0 ) | ( ~n13297 & 1'b0 ) ;
  assign n13299 = n13289 | n13298 ;
  assign n13300 = ( n13278 & ~n13280 ) | ( n13278 & 1'b0 ) | ( ~n13280 & 1'b0 ) ;
  assign n13301 = ( n13275 & ~n11674 ) | ( n13275 & n13300 ) | ( ~n11674 & n13300 ) ;
  assign n13302 = ( n11176 & ~n13301 ) | ( n11176 & 1'b0 ) | ( ~n13301 & 1'b0 ) ;
  assign n13303 = n10685 | n13302 ;
  assign n13304 = ( n13299 & ~n13303 ) | ( n13299 & 1'b0 ) | ( ~n13303 & 1'b0 ) ;
  assign n13305 = n13296 | n13304 ;
  assign n13306 = ~n13291 & n13305 ;
  assign n13307 = n12749 | n13242 ;
  assign n13308 = ( n12754 & ~n12749 ) | ( n12754 & n12762 ) | ( ~n12749 & n12762 ) ;
  assign n13310 = ( n12749 & n13307 ) | ( n12749 & n13308 ) | ( n13307 & n13308 ) ;
  assign n13309 = ( n12762 & ~n13308 ) | ( n12762 & n13307 ) | ( ~n13308 & n13307 ) ;
  assign n13311 = ( n12754 & ~n13310 ) | ( n12754 & n13309 ) | ( ~n13310 & n13309 ) ;
  assign n13312 = ( n13306 & ~n10209 ) | ( n13306 & n13311 ) | ( ~n10209 & n13311 ) ;
  assign n13313 = n9740 | n13312 ;
  assign n13314 = n12782 | n13242 ;
  assign n13315 = ( n12769 & ~n12778 ) | ( n12769 & n12782 ) | ( ~n12778 & n12782 ) ;
  assign n13316 = ( n12778 & n13314 ) | ( n12778 & n13315 ) | ( n13314 & n13315 ) ;
  assign n13317 = ( n12782 & ~n13315 ) | ( n12782 & n13314 ) | ( ~n13315 & n13314 ) ;
  assign n13318 = ( n12769 & ~n13316 ) | ( n12769 & n13317 ) | ( ~n13316 & n13317 ) ;
  assign n13319 = n10209 | n13291 ;
  assign n13320 = ( n13305 & ~n13319 ) | ( n13305 & 1'b0 ) | ( ~n13319 & 1'b0 ) ;
  assign n13321 = n13311 | n13320 ;
  assign n13322 = ( n13299 & ~n13302 ) | ( n13299 & 1'b0 ) | ( ~n13302 & 1'b0 ) ;
  assign n13323 = ( n13296 & ~n10685 ) | ( n13296 & n13322 ) | ( ~n10685 & n13322 ) ;
  assign n13324 = ( n10209 & ~n13323 ) | ( n10209 & 1'b0 ) | ( ~n13323 & 1'b0 ) ;
  assign n13325 = ( n9740 & ~n13324 ) | ( n9740 & 1'b0 ) | ( ~n13324 & 1'b0 ) ;
  assign n13326 = n13321 &  n13325 ;
  assign n13327 = n13318 | n13326 ;
  assign n13328 = n13313 &  n13327 ;
  assign n13330 = ( n12771 & ~n12776 ) | ( n12771 & n12784 ) | ( ~n12776 & n12784 ) ;
  assign n13329 = ( n12771 & ~n13242 ) | ( n12771 & 1'b0 ) | ( ~n13242 & 1'b0 ) ;
  assign n13332 = ( n12771 & ~n13330 ) | ( n12771 & n13329 ) | ( ~n13330 & n13329 ) ;
  assign n13331 = ( n13329 & ~n12784 ) | ( n13329 & n13330 ) | ( ~n12784 & n13330 ) ;
  assign n13333 = ( n12776 & ~n13332 ) | ( n12776 & n13331 ) | ( ~n13332 & n13331 ) ;
  assign n13334 = ( n13328 & ~n9286 ) | ( n13328 & n13333 ) | ( ~n9286 & n13333 ) ;
  assign n13335 = ( n8839 & ~n13334 ) | ( n8839 & 1'b0 ) | ( ~n13334 & 1'b0 ) ;
  assign n13336 = n12804 | n13242 ;
  assign n13337 = ( n12791 & ~n12804 ) | ( n12791 & n12800 ) | ( ~n12804 & n12800 ) ;
  assign n13339 = ( n12804 & n13336 ) | ( n12804 & n13337 ) | ( n13336 & n13337 ) ;
  assign n13338 = ( n12800 & ~n13337 ) | ( n12800 & n13336 ) | ( ~n13337 & n13336 ) ;
  assign n13340 = ( n12791 & ~n13339 ) | ( n12791 & n13338 ) | ( ~n13339 & n13338 ) ;
  assign n13341 = ~n9286 & n13313 ;
  assign n13342 = n13327 &  n13341 ;
  assign n13343 = n13333 | n13342 ;
  assign n13344 = ( n13321 & ~n13324 ) | ( n13321 & 1'b0 ) | ( ~n13324 & 1'b0 ) ;
  assign n13345 = ( n9740 & n13318 ) | ( n9740 & n13344 ) | ( n13318 & n13344 ) ;
  assign n13346 = ( n9286 & ~n13345 ) | ( n9286 & 1'b0 ) | ( ~n13345 & 1'b0 ) ;
  assign n13347 = n8839 | n13346 ;
  assign n13348 = ( n13343 & ~n13347 ) | ( n13343 & 1'b0 ) | ( ~n13347 & 1'b0 ) ;
  assign n13349 = n13340 | n13348 ;
  assign n13350 = ~n13335 & n13349 ;
  assign n13351 = n12806 &  n13242 ;
  assign n13352 = ( n12793 & n12798 ) | ( n12793 & n13242 ) | ( n12798 & n13242 ) ;
  assign n13354 = ( n13351 & ~n12793 ) | ( n13351 & n13352 ) | ( ~n12793 & n13352 ) ;
  assign n13353 = ( n13242 & ~n13352 ) | ( n13242 & n13351 ) | ( ~n13352 & n13351 ) ;
  assign n13355 = ( n12798 & ~n13354 ) | ( n12798 & n13353 ) | ( ~n13354 & n13353 ) ;
  assign n13356 = ( n13350 & ~n8407 ) | ( n13350 & n13355 ) | ( ~n8407 & n13355 ) ;
  assign n13357 = ( n7982 & ~n13356 ) | ( n7982 & 1'b0 ) | ( ~n13356 & 1'b0 ) ;
  assign n13358 = n12826 | n13242 ;
  assign n13359 = ( n12813 & ~n12822 ) | ( n12813 & n12826 ) | ( ~n12822 & n12826 ) ;
  assign n13360 = ( n12822 & n13358 ) | ( n12822 & n13359 ) | ( n13358 & n13359 ) ;
  assign n13361 = ( n12826 & ~n13359 ) | ( n12826 & n13358 ) | ( ~n13359 & n13358 ) ;
  assign n13362 = ( n12813 & ~n13360 ) | ( n12813 & n13361 ) | ( ~n13360 & n13361 ) ;
  assign n13363 = n8407 | n13335 ;
  assign n13364 = ( n13349 & ~n13363 ) | ( n13349 & 1'b0 ) | ( ~n13363 & 1'b0 ) ;
  assign n13365 = n13355 | n13364 ;
  assign n13366 = ( n13343 & ~n13346 ) | ( n13343 & 1'b0 ) | ( ~n13346 & 1'b0 ) ;
  assign n13367 = ( n13340 & ~n8839 ) | ( n13340 & n13366 ) | ( ~n8839 & n13366 ) ;
  assign n13368 = ( n8407 & ~n13367 ) | ( n8407 & 1'b0 ) | ( ~n13367 & 1'b0 ) ;
  assign n13369 = n7982 | n13368 ;
  assign n13370 = ( n13365 & ~n13369 ) | ( n13365 & 1'b0 ) | ( ~n13369 & 1'b0 ) ;
  assign n13371 = n13362 | n13370 ;
  assign n13372 = ~n13357 & n13371 ;
  assign n13373 = n12815 | n13242 ;
  assign n13374 = ( n12820 & ~n12815 ) | ( n12820 & n12828 ) | ( ~n12815 & n12828 ) ;
  assign n13376 = ( n12815 & n13373 ) | ( n12815 & n13374 ) | ( n13373 & n13374 ) ;
  assign n13375 = ( n12828 & ~n13374 ) | ( n12828 & n13373 ) | ( ~n13374 & n13373 ) ;
  assign n13377 = ( n12820 & ~n13376 ) | ( n12820 & n13375 ) | ( ~n13376 & n13375 ) ;
  assign n13378 = ( n7572 & n13372 ) | ( n7572 & n13377 ) | ( n13372 & n13377 ) ;
  assign n13379 = n7169 | n13378 ;
  assign n13381 = ( n12844 & ~n12835 ) | ( n12844 & n12848 ) | ( ~n12835 & n12848 ) ;
  assign n13380 = ( n12848 & ~n13242 ) | ( n12848 & 1'b0 ) | ( ~n13242 & 1'b0 ) ;
  assign n13383 = ( n12848 & ~n13381 ) | ( n12848 & n13380 ) | ( ~n13381 & n13380 ) ;
  assign n13382 = ( n13380 & ~n12844 ) | ( n13380 & n13381 ) | ( ~n12844 & n13381 ) ;
  assign n13384 = ( n12835 & ~n13383 ) | ( n12835 & n13382 ) | ( ~n13383 & n13382 ) ;
  assign n13385 = ( n7572 & ~n13357 ) | ( n7572 & 1'b0 ) | ( ~n13357 & 1'b0 ) ;
  assign n13386 = n13371 &  n13385 ;
  assign n13387 = n13377 | n13386 ;
  assign n13388 = ( n13365 & ~n13368 ) | ( n13365 & 1'b0 ) | ( ~n13368 & 1'b0 ) ;
  assign n13389 = ( n13362 & ~n7982 ) | ( n13362 & n13388 ) | ( ~n7982 & n13388 ) ;
  assign n13390 = n7572 | n13389 ;
  assign n13391 = n7169 &  n13390 ;
  assign n13392 = n13387 &  n13391 ;
  assign n13393 = n13384 | n13392 ;
  assign n13394 = n13379 &  n13393 ;
  assign n13395 = ( n12837 & ~n13242 ) | ( n12837 & 1'b0 ) | ( ~n13242 & 1'b0 ) ;
  assign n13396 = ( n12837 & n12842 ) | ( n12837 & n12850 ) | ( n12842 & n12850 ) ;
  assign n13397 = ( n13395 & ~n12850 ) | ( n13395 & n13396 ) | ( ~n12850 & n13396 ) ;
  assign n13398 = ( n12837 & ~n13396 ) | ( n12837 & n13395 ) | ( ~n13396 & n13395 ) ;
  assign n13399 = ( n12842 & ~n13397 ) | ( n12842 & n13398 ) | ( ~n13397 & n13398 ) ;
  assign n13400 = ( n13394 & ~n6781 ) | ( n13394 & n13399 ) | ( ~n6781 & n13399 ) ;
  assign n13401 = n6399 | n13400 ;
  assign n13402 = n12870 | n13242 ;
  assign n13403 = ( n12857 & ~n12870 ) | ( n12857 & n12866 ) | ( ~n12870 & n12866 ) ;
  assign n13405 = ( n12870 & n13402 ) | ( n12870 & n13403 ) | ( n13402 & n13403 ) ;
  assign n13404 = ( n12866 & ~n13403 ) | ( n12866 & n13402 ) | ( ~n13403 & n13402 ) ;
  assign n13406 = ( n12857 & ~n13405 ) | ( n12857 & n13404 ) | ( ~n13405 & n13404 ) ;
  assign n13407 = ~n6781 & n13379 ;
  assign n13408 = n13393 &  n13407 ;
  assign n13409 = n13399 | n13408 ;
  assign n13410 = n13387 &  n13390 ;
  assign n13411 = ( n7169 & n13384 ) | ( n7169 & n13410 ) | ( n13384 & n13410 ) ;
  assign n13412 = ( n6781 & ~n13411 ) | ( n6781 & 1'b0 ) | ( ~n13411 & 1'b0 ) ;
  assign n13413 = ( n6399 & ~n13412 ) | ( n6399 & 1'b0 ) | ( ~n13412 & 1'b0 ) ;
  assign n13414 = n13409 &  n13413 ;
  assign n13415 = ( n13406 & ~n13414 ) | ( n13406 & 1'b0 ) | ( ~n13414 & 1'b0 ) ;
  assign n13416 = ( n13401 & ~n13415 ) | ( n13401 & 1'b0 ) | ( ~n13415 & 1'b0 ) ;
  assign n13417 = n12859 | n13242 ;
  assign n13418 = ( n12859 & ~n12872 ) | ( n12859 & n12864 ) | ( ~n12872 & n12864 ) ;
  assign n13419 = ( n12872 & n13417 ) | ( n12872 & n13418 ) | ( n13417 & n13418 ) ;
  assign n13420 = ( n12859 & ~n13418 ) | ( n12859 & n13417 ) | ( ~n13418 & n13417 ) ;
  assign n13421 = ( n12864 & ~n13419 ) | ( n12864 & n13420 ) | ( ~n13419 & n13420 ) ;
  assign n13422 = ( n6032 & ~n13416 ) | ( n6032 & n13421 ) | ( ~n13416 & n13421 ) ;
  assign n13423 = ~n5672 & n13422 ;
  assign n13425 = ( n12888 & ~n12879 ) | ( n12888 & n12892 ) | ( ~n12879 & n12892 ) ;
  assign n13424 = n12892 | n13242 ;
  assign n13427 = ( n12892 & ~n13425 ) | ( n12892 & n13424 ) | ( ~n13425 & n13424 ) ;
  assign n13426 = ( n13424 & ~n12888 ) | ( n13424 & n13425 ) | ( ~n12888 & n13425 ) ;
  assign n13428 = ( n12879 & ~n13427 ) | ( n12879 & n13426 ) | ( ~n13427 & n13426 ) ;
  assign n13429 = ~n6032 & n13401 ;
  assign n13430 = ~n13415 & n13429 ;
  assign n13431 = ( n13421 & ~n13430 ) | ( n13421 & 1'b0 ) | ( ~n13430 & 1'b0 ) ;
  assign n13432 = ( n13409 & ~n13412 ) | ( n13409 & 1'b0 ) | ( ~n13412 & 1'b0 ) ;
  assign n13433 = ( n6399 & ~n13406 ) | ( n6399 & n13432 ) | ( ~n13406 & n13432 ) ;
  assign n13434 = ( n6032 & ~n13433 ) | ( n6032 & 1'b0 ) | ( ~n13433 & 1'b0 ) ;
  assign n13435 = ( n5672 & ~n13434 ) | ( n5672 & 1'b0 ) | ( ~n13434 & 1'b0 ) ;
  assign n13436 = ~n13431 & n13435 ;
  assign n13437 = ( n13428 & ~n13436 ) | ( n13428 & 1'b0 ) | ( ~n13436 & 1'b0 ) ;
  assign n13438 = n13423 | n13437 ;
  assign n13439 = n12881 | n13242 ;
  assign n13440 = ( n12881 & ~n12894 ) | ( n12881 & n12886 ) | ( ~n12894 & n12886 ) ;
  assign n13441 = ( n12894 & n13439 ) | ( n12894 & n13440 ) | ( n13439 & n13440 ) ;
  assign n13442 = ( n12881 & ~n13440 ) | ( n12881 & n13439 ) | ( ~n13440 & n13439 ) ;
  assign n13443 = ( n12886 & ~n13441 ) | ( n12886 & n13442 ) | ( ~n13441 & n13442 ) ;
  assign n13444 = ( n5327 & n13438 ) | ( n5327 & n13443 ) | ( n13438 & n13443 ) ;
  assign n13445 = n4990 &  n13444 ;
  assign n13447 = ( n12910 & ~n12901 ) | ( n12910 & n12914 ) | ( ~n12901 & n12914 ) ;
  assign n13446 = n12914 | n13242 ;
  assign n13449 = ( n12914 & ~n13447 ) | ( n12914 & n13446 ) | ( ~n13447 & n13446 ) ;
  assign n13448 = ( n13446 & ~n12910 ) | ( n13446 & n13447 ) | ( ~n12910 & n13447 ) ;
  assign n13450 = ( n12901 & ~n13449 ) | ( n12901 & n13448 ) | ( ~n13449 & n13448 ) ;
  assign n13451 = n5327 | n13423 ;
  assign n13452 = n13437 | n13451 ;
  assign n13453 = n13443 &  n13452 ;
  assign n13454 = n13431 | n13434 ;
  assign n13455 = ( n13428 & ~n5672 ) | ( n13428 & n13454 ) | ( ~n5672 & n13454 ) ;
  assign n13456 = n5327 &  n13455 ;
  assign n13457 = n4990 | n13456 ;
  assign n13458 = n13453 | n13457 ;
  assign n13459 = n13450 &  n13458 ;
  assign n13460 = n13445 | n13459 ;
  assign n13466 = ( n4668 & ~n13465 ) | ( n4668 & n13460 ) | ( ~n13465 & n13460 ) ;
  assign n13467 = n4353 &  n13466 ;
  assign n13468 = n12936 | n13242 ;
  assign n13469 = ( n12923 & n12932 ) | ( n12923 & n12936 ) | ( n12932 & n12936 ) ;
  assign n13470 = ( n13468 & ~n12932 ) | ( n13468 & n13469 ) | ( ~n12932 & n13469 ) ;
  assign n13471 = ( n12936 & ~n13469 ) | ( n12936 & n13468 ) | ( ~n13469 & n13468 ) ;
  assign n13472 = ( n12923 & ~n13470 ) | ( n12923 & n13471 ) | ( ~n13470 & n13471 ) ;
  assign n13473 = n4668 | n13445 ;
  assign n13474 = n13459 | n13473 ;
  assign n13475 = ~n13465 & n13474 ;
  assign n13476 = n13453 | n13456 ;
  assign n13477 = ( n4990 & n13450 ) | ( n4990 & n13476 ) | ( n13450 & n13476 ) ;
  assign n13478 = n4668 &  n13477 ;
  assign n13479 = n4353 | n13478 ;
  assign n13480 = n13475 | n13479 ;
  assign n13481 = ~n13472 & n13480 ;
  assign n13482 = n13467 | n13481 ;
  assign n13483 = n12925 | n13242 ;
  assign n13484 = ( n12925 & n12930 ) | ( n12925 & n12938 ) | ( n12930 & n12938 ) ;
  assign n13485 = ( n13483 & ~n12938 ) | ( n13483 & n13484 ) | ( ~n12938 & n13484 ) ;
  assign n13486 = ( n12925 & ~n13484 ) | ( n12925 & n13483 ) | ( ~n13484 & n13483 ) ;
  assign n13487 = ( n12930 & ~n13485 ) | ( n12930 & n13486 ) | ( ~n13485 & n13486 ) ;
  assign n13488 = ( n4053 & n13482 ) | ( n4053 & n13487 ) | ( n13482 & n13487 ) ;
  assign n13489 = n3760 &  n13488 ;
  assign n13490 = n12958 | n13242 ;
  assign n13491 = ( n12945 & n12954 ) | ( n12945 & n12958 ) | ( n12954 & n12958 ) ;
  assign n13492 = ( n13490 & ~n12954 ) | ( n13490 & n13491 ) | ( ~n12954 & n13491 ) ;
  assign n13493 = ( n12958 & ~n13491 ) | ( n12958 & n13490 ) | ( ~n13491 & n13490 ) ;
  assign n13494 = ( n12945 & ~n13492 ) | ( n12945 & n13493 ) | ( ~n13492 & n13493 ) ;
  assign n13495 = n4053 | n13467 ;
  assign n13496 = n13481 | n13495 ;
  assign n13497 = n13487 &  n13496 ;
  assign n13498 = n13475 | n13478 ;
  assign n13499 = ( n4353 & ~n13472 ) | ( n4353 & n13498 ) | ( ~n13472 & n13498 ) ;
  assign n13500 = n4053 &  n13499 ;
  assign n13501 = n3760 | n13500 ;
  assign n13502 = n13497 | n13501 ;
  assign n13503 = ~n13494 & n13502 ;
  assign n13504 = n13489 | n13503 ;
  assign n13505 = n12947 | n13242 ;
  assign n13506 = ( n12947 & n12952 ) | ( n12947 & n12960 ) | ( n12952 & n12960 ) ;
  assign n13507 = ( n13505 & ~n12960 ) | ( n13505 & n13506 ) | ( ~n12960 & n13506 ) ;
  assign n13508 = ( n12947 & ~n13506 ) | ( n12947 & n13505 ) | ( ~n13506 & n13505 ) ;
  assign n13509 = ( n12952 & ~n13507 ) | ( n12952 & n13508 ) | ( ~n13507 & n13508 ) ;
  assign n13510 = ( n3482 & n13504 ) | ( n3482 & n13509 ) | ( n13504 & n13509 ) ;
  assign n13511 = n3211 &  n13510 ;
  assign n13513 = ( n12976 & ~n12967 ) | ( n12976 & n12980 ) | ( ~n12967 & n12980 ) ;
  assign n13512 = n12980 | n13242 ;
  assign n13515 = ( n12980 & ~n13513 ) | ( n12980 & n13512 ) | ( ~n13513 & n13512 ) ;
  assign n13514 = ( n13512 & ~n12976 ) | ( n13512 & n13513 ) | ( ~n12976 & n13513 ) ;
  assign n13516 = ( n12967 & ~n13515 ) | ( n12967 & n13514 ) | ( ~n13515 & n13514 ) ;
  assign n13517 = n3482 | n13489 ;
  assign n13518 = n13503 | n13517 ;
  assign n13519 = n13509 &  n13518 ;
  assign n13520 = n13497 | n13500 ;
  assign n13521 = ( n3760 & ~n13494 ) | ( n3760 & n13520 ) | ( ~n13494 & n13520 ) ;
  assign n13522 = n3482 &  n13521 ;
  assign n13523 = n3211 | n13522 ;
  assign n13524 = n13519 | n13523 ;
  assign n13525 = n13516 &  n13524 ;
  assign n13526 = n13511 | n13525 ;
  assign n13532 = ( n2955 & ~n13531 ) | ( n2955 & n13526 ) | ( ~n13531 & n13526 ) ;
  assign n13533 = n2706 &  n13532 ;
  assign n13535 = ( n12998 & ~n12989 ) | ( n12998 & n13002 ) | ( ~n12989 & n13002 ) ;
  assign n13534 = n13002 | n13242 ;
  assign n13537 = ( n13002 & ~n13535 ) | ( n13002 & n13534 ) | ( ~n13535 & n13534 ) ;
  assign n13536 = ( n13534 & ~n12998 ) | ( n13534 & n13535 ) | ( ~n12998 & n13535 ) ;
  assign n13538 = ( n12989 & ~n13537 ) | ( n12989 & n13536 ) | ( ~n13537 & n13536 ) ;
  assign n13539 = n2955 | n13511 ;
  assign n13540 = n13525 | n13539 ;
  assign n13541 = ~n13531 & n13540 ;
  assign n13542 = n13519 | n13522 ;
  assign n13543 = ( n3211 & n13516 ) | ( n3211 & n13542 ) | ( n13516 & n13542 ) ;
  assign n13544 = n2955 &  n13543 ;
  assign n13545 = n2706 | n13544 ;
  assign n13546 = n13541 | n13545 ;
  assign n13547 = ~n13538 & n13546 ;
  assign n13548 = n13533 | n13547 ;
  assign n13554 = ( n2472 & ~n13553 ) | ( n2472 & n13548 ) | ( ~n13553 & n13548 ) ;
  assign n13555 = n2245 &  n13554 ;
  assign n13557 = ( n13020 & ~n13011 ) | ( n13020 & n13024 ) | ( ~n13011 & n13024 ) ;
  assign n13556 = n13024 | n13242 ;
  assign n13559 = ( n13024 & ~n13557 ) | ( n13024 & n13556 ) | ( ~n13557 & n13556 ) ;
  assign n13558 = ( n13556 & ~n13020 ) | ( n13556 & n13557 ) | ( ~n13020 & n13557 ) ;
  assign n13560 = ( n13011 & ~n13559 ) | ( n13011 & n13558 ) | ( ~n13559 & n13558 ) ;
  assign n13561 = n2472 | n13533 ;
  assign n13562 = n13547 | n13561 ;
  assign n13563 = ~n13553 & n13562 ;
  assign n13564 = n13541 | n13544 ;
  assign n13565 = ( n2706 & ~n13538 ) | ( n2706 & n13564 ) | ( ~n13538 & n13564 ) ;
  assign n13566 = n2472 &  n13565 ;
  assign n13567 = n2245 | n13566 ;
  assign n13568 = n13563 | n13567 ;
  assign n13569 = ~n13560 & n13568 ;
  assign n13570 = n13555 | n13569 ;
  assign n13571 = ~n13026 & n13242 ;
  assign n13572 = ( n13013 & ~n13571 ) | ( n13013 & n13242 ) | ( ~n13571 & n13242 ) ;
  assign n13573 = ( n13018 & ~n13013 ) | ( n13018 & n13572 ) | ( ~n13013 & n13572 ) ;
  assign n13574 = ( n13013 & ~n13572 ) | ( n13013 & n13018 ) | ( ~n13572 & n13018 ) ;
  assign n13575 = ( n13573 & ~n13018 ) | ( n13573 & n13574 ) | ( ~n13018 & n13574 ) ;
  assign n13576 = ( n2033 & ~n13570 ) | ( n2033 & n13575 ) | ( ~n13570 & n13575 ) ;
  assign n13577 = ( n1827 & ~n13576 ) | ( n1827 & 1'b0 ) | ( ~n13576 & 1'b0 ) ;
  assign n13583 = ( n2033 & ~n13555 ) | ( n2033 & 1'b0 ) | ( ~n13555 & 1'b0 ) ;
  assign n13584 = ~n13569 & n13583 ;
  assign n13585 = n13575 | n13584 ;
  assign n13586 = n13563 | n13566 ;
  assign n13587 = ( n2245 & ~n13560 ) | ( n2245 & n13586 ) | ( ~n13560 & n13586 ) ;
  assign n13588 = ~n2033 & n13587 ;
  assign n13589 = n1827 | n13588 ;
  assign n13590 = ( n13585 & ~n13589 ) | ( n13585 & 1'b0 ) | ( ~n13589 & 1'b0 ) ;
  assign n13591 = ( n13582 & ~n13590 ) | ( n13582 & 1'b0 ) | ( ~n13590 & 1'b0 ) ;
  assign n13592 = n13577 | n13591 ;
  assign n13594 = ( n13035 & ~n13040 ) | ( n13035 & n13242 ) | ( ~n13040 & n13242 ) ;
  assign n13593 = ~n13048 & n13242 ;
  assign n13595 = ( n13242 & ~n13594 ) | ( n13242 & n13593 ) | ( ~n13594 & n13593 ) ;
  assign n13596 = ( n13593 & ~n13035 ) | ( n13593 & n13594 ) | ( ~n13035 & n13594 ) ;
  assign n13597 = ( n13040 & ~n13595 ) | ( n13040 & n13596 ) | ( ~n13595 & n13596 ) ;
  assign n13598 = ( n1636 & ~n13592 ) | ( n1636 & n13597 ) | ( ~n13592 & n13597 ) ;
  assign n13599 = n1452 | n13598 ;
  assign n13600 = ( n1636 & ~n13577 ) | ( n1636 & 1'b0 ) | ( ~n13577 & 1'b0 ) ;
  assign n13601 = ~n13591 & n13600 ;
  assign n13602 = n13597 | n13601 ;
  assign n13603 = ( n13585 & ~n13588 ) | ( n13585 & 1'b0 ) | ( ~n13588 & 1'b0 ) ;
  assign n13604 = ( n1827 & ~n13603 ) | ( n1827 & n13582 ) | ( ~n13603 & n13582 ) ;
  assign n13605 = ~n1636 & n13604 ;
  assign n13606 = ( n1452 & ~n13605 ) | ( n1452 & 1'b0 ) | ( ~n13605 & 1'b0 ) ;
  assign n13607 = n13602 &  n13606 ;
  assign n13608 = ( n13054 & ~n13063 ) | ( n13054 & n13067 ) | ( ~n13063 & n13067 ) ;
  assign n13609 = ( n13063 & n13242 ) | ( n13063 & n13608 ) | ( n13242 & n13608 ) ;
  assign n13610 = ( n13067 & ~n13608 ) | ( n13067 & n13242 ) | ( ~n13608 & n13242 ) ;
  assign n13611 = ( n13054 & ~n13609 ) | ( n13054 & n13610 ) | ( ~n13609 & n13610 ) ;
  assign n13612 = n13607 | n13611 ;
  assign n13613 = n13599 &  n13612 ;
  assign n13614 = n13069 &  n13242 ;
  assign n13615 = ( n13056 & ~n13242 ) | ( n13056 & n13614 ) | ( ~n13242 & n13614 ) ;
  assign n13616 = ( n13061 & ~n13056 ) | ( n13061 & n13615 ) | ( ~n13056 & n13615 ) ;
  assign n13617 = ( n13056 & ~n13615 ) | ( n13056 & n13061 ) | ( ~n13615 & n13061 ) ;
  assign n13618 = ( n13616 & ~n13061 ) | ( n13616 & n13617 ) | ( ~n13061 & n13617 ) ;
  assign n13619 = ( n1283 & ~n13613 ) | ( n1283 & n13618 ) | ( ~n13613 & n13618 ) ;
  assign n13620 = ~n1122 & n13619 ;
  assign n13621 = n13089 | n13242 ;
  assign n13622 = ( n13076 & ~n13089 ) | ( n13076 & n13085 ) | ( ~n13089 & n13085 ) ;
  assign n13624 = ( n13089 & n13621 ) | ( n13089 & n13622 ) | ( n13621 & n13622 ) ;
  assign n13623 = ( n13085 & ~n13622 ) | ( n13085 & n13621 ) | ( ~n13622 & n13621 ) ;
  assign n13625 = ( n13076 & ~n13624 ) | ( n13076 & n13623 ) | ( ~n13624 & n13623 ) ;
  assign n13626 = ~n1283 & n13599 ;
  assign n13627 = n13612 &  n13626 ;
  assign n13628 = ( n13618 & ~n13627 ) | ( n13618 & 1'b0 ) | ( ~n13627 & 1'b0 ) ;
  assign n13629 = ( n13602 & ~n13605 ) | ( n13602 & 1'b0 ) | ( ~n13605 & 1'b0 ) ;
  assign n13630 = ( n1452 & n13611 ) | ( n1452 & n13629 ) | ( n13611 & n13629 ) ;
  assign n13631 = ( n1283 & ~n13630 ) | ( n1283 & 1'b0 ) | ( ~n13630 & 1'b0 ) ;
  assign n13632 = ( n1122 & ~n13631 ) | ( n1122 & 1'b0 ) | ( ~n13631 & 1'b0 ) ;
  assign n13633 = ~n13628 & n13632 ;
  assign n13634 = n13625 | n13633 ;
  assign n13635 = ~n13620 & n13634 ;
  assign n13641 = ( n976 & ~n13640 ) | ( n976 & n13635 ) | ( ~n13640 & n13635 ) ;
  assign n13642 = ( n837 & ~n13641 ) | ( n837 & 1'b0 ) | ( ~n13641 & 1'b0 ) ;
  assign n13644 = ( n13107 & ~n13098 ) | ( n13107 & n13111 ) | ( ~n13098 & n13111 ) ;
  assign n13643 = ( n13111 & ~n13242 ) | ( n13111 & 1'b0 ) | ( ~n13242 & 1'b0 ) ;
  assign n13646 = ( n13111 & ~n13644 ) | ( n13111 & n13643 ) | ( ~n13644 & n13643 ) ;
  assign n13645 = ( n13643 & ~n13107 ) | ( n13643 & n13644 ) | ( ~n13107 & n13644 ) ;
  assign n13647 = ( n13098 & ~n13646 ) | ( n13098 & n13645 ) | ( ~n13646 & n13645 ) ;
  assign n13648 = ( n976 & ~n13620 ) | ( n976 & 1'b0 ) | ( ~n13620 & 1'b0 ) ;
  assign n13649 = n13634 &  n13648 ;
  assign n13650 = ( n13640 & ~n13649 ) | ( n13640 & 1'b0 ) | ( ~n13649 & 1'b0 ) ;
  assign n13651 = n13628 | n13631 ;
  assign n13652 = ( n1122 & ~n13651 ) | ( n1122 & n13625 ) | ( ~n13651 & n13625 ) ;
  assign n13653 = n976 | n13652 ;
  assign n13654 = ~n837 & n13653 ;
  assign n13655 = ~n13650 & n13654 ;
  assign n13656 = ( n13647 & ~n13655 ) | ( n13647 & 1'b0 ) | ( ~n13655 & 1'b0 ) ;
  assign n13657 = n13642 | n13656 ;
  assign n13663 = ( n713 & ~n13662 ) | ( n713 & n13657 ) | ( ~n13662 & n13657 ) ;
  assign n13664 = n595 &  n13663 ;
  assign n13665 = n13133 | n13242 ;
  assign n13666 = ( n13120 & ~n13129 ) | ( n13120 & n13133 ) | ( ~n13129 & n13133 ) ;
  assign n13667 = ( n13129 & n13665 ) | ( n13129 & n13666 ) | ( n13665 & n13666 ) ;
  assign n13668 = ( n13133 & ~n13666 ) | ( n13133 & n13665 ) | ( ~n13666 & n13665 ) ;
  assign n13669 = ( n13120 & ~n13667 ) | ( n13120 & n13668 ) | ( ~n13667 & n13668 ) ;
  assign n13670 = n713 | n13642 ;
  assign n13671 = n13656 | n13670 ;
  assign n13672 = ~n13662 & n13671 ;
  assign n13673 = ~n13650 & n13653 ;
  assign n13674 = ( n837 & ~n13673 ) | ( n837 & n13647 ) | ( ~n13673 & n13647 ) ;
  assign n13675 = n713 &  n13674 ;
  assign n13676 = n595 | n13675 ;
  assign n13677 = n13672 | n13676 ;
  assign n13678 = n13669 &  n13677 ;
  assign n13679 = n13664 | n13678 ;
  assign n13685 = ( n492 & ~n13684 ) | ( n492 & n13679 ) | ( ~n13684 & n13679 ) ;
  assign n13686 = n396 &  n13685 ;
  assign n13688 = ( n13151 & ~n13142 ) | ( n13151 & n13155 ) | ( ~n13142 & n13155 ) ;
  assign n13687 = n13155 | n13242 ;
  assign n13690 = ( n13155 & ~n13688 ) | ( n13155 & n13687 ) | ( ~n13688 & n13687 ) ;
  assign n13689 = ( n13687 & ~n13151 ) | ( n13687 & n13688 ) | ( ~n13151 & n13688 ) ;
  assign n13691 = ( n13142 & ~n13690 ) | ( n13142 & n13689 ) | ( ~n13690 & n13689 ) ;
  assign n13692 = n492 | n13664 ;
  assign n13693 = n13678 | n13692 ;
  assign n13694 = ~n13684 & n13693 ;
  assign n13695 = n13672 | n13675 ;
  assign n13696 = ( n595 & n13669 ) | ( n595 & n13695 ) | ( n13669 & n13695 ) ;
  assign n13697 = n492 &  n13696 ;
  assign n13698 = n396 | n13697 ;
  assign n13699 = n13694 | n13698 ;
  assign n13700 = ~n13691 & n13699 ;
  assign n13701 = n13686 | n13700 ;
  assign n13702 = ~n13157 & n13242 ;
  assign n13703 = ( n13144 & ~n13702 ) | ( n13144 & n13242 ) | ( ~n13702 & n13242 ) ;
  assign n13704 = ( n13144 & ~n13703 ) | ( n13144 & n13149 ) | ( ~n13703 & n13149 ) ;
  assign n13705 = ( n13149 & ~n13144 ) | ( n13149 & n13703 ) | ( ~n13144 & n13703 ) ;
  assign n13706 = ( n13704 & ~n13149 ) | ( n13704 & n13705 ) | ( ~n13149 & n13705 ) ;
  assign n13707 = ( n315 & n13701 ) | ( n315 & n13706 ) | ( n13701 & n13706 ) ;
  assign n13708 = n240 &  n13707 ;
  assign n13709 = n13177 | n13242 ;
  assign n13710 = ( n13164 & n13173 ) | ( n13164 & n13177 ) | ( n13173 & n13177 ) ;
  assign n13711 = ( n13709 & ~n13173 ) | ( n13709 & n13710 ) | ( ~n13173 & n13710 ) ;
  assign n13712 = ( n13177 & ~n13710 ) | ( n13177 & n13709 ) | ( ~n13710 & n13709 ) ;
  assign n13713 = ( n13164 & ~n13711 ) | ( n13164 & n13712 ) | ( ~n13711 & n13712 ) ;
  assign n13714 = n315 | n13686 ;
  assign n13715 = n13700 | n13714 ;
  assign n13716 = n13706 &  n13715 ;
  assign n13717 = n13694 | n13697 ;
  assign n13718 = ( n396 & ~n13691 ) | ( n396 & n13717 ) | ( ~n13691 & n13717 ) ;
  assign n13719 = n315 &  n13718 ;
  assign n13720 = n240 | n13719 ;
  assign n13721 = n13716 | n13720 ;
  assign n13722 = n13713 &  n13721 ;
  assign n13723 = n13708 | n13722 ;
  assign n13729 = ( n181 & ~n13728 ) | ( n181 & n13723 ) | ( ~n13728 & n13723 ) ;
  assign n13730 = ~n145 & n13729 ;
  assign n13732 = ( n13195 & ~n13186 ) | ( n13195 & n13199 ) | ( ~n13186 & n13199 ) ;
  assign n13731 = n13199 | n13242 ;
  assign n13734 = ( n13199 & ~n13732 ) | ( n13199 & n13731 ) | ( ~n13732 & n13731 ) ;
  assign n13733 = ( n13731 & ~n13195 ) | ( n13731 & n13732 ) | ( ~n13195 & n13732 ) ;
  assign n13735 = ( n13186 & ~n13734 ) | ( n13186 & n13733 ) | ( ~n13734 & n13733 ) ;
  assign n13736 = n181 | n13708 ;
  assign n13737 = n13722 | n13736 ;
  assign n13738 = ~n13728 & n13737 ;
  assign n13739 = n13716 | n13719 ;
  assign n13740 = ( n240 & n13713 ) | ( n240 & n13739 ) | ( n13713 & n13739 ) ;
  assign n13741 = n181 &  n13740 ;
  assign n13742 = ( n145 & ~n13741 ) | ( n145 & 1'b0 ) | ( ~n13741 & 1'b0 ) ;
  assign n13743 = ~n13738 & n13742 ;
  assign n13744 = ( n13735 & ~n13743 ) | ( n13735 & 1'b0 ) | ( ~n13743 & 1'b0 ) ;
  assign n13745 = n13730 | n13744 ;
  assign n13746 = n13188 | n13242 ;
  assign n13747 = ( n13193 & ~n13188 ) | ( n13193 & n13201 ) | ( ~n13188 & n13201 ) ;
  assign n13749 = ( n13188 & n13746 ) | ( n13188 & n13747 ) | ( n13746 & n13747 ) ;
  assign n13748 = ( n13201 & ~n13747 ) | ( n13201 & n13746 ) | ( ~n13747 & n13746 ) ;
  assign n13750 = ( n13193 & ~n13749 ) | ( n13193 & n13748 ) | ( ~n13749 & n13748 ) ;
  assign n13751 = ( n150 & n13745 ) | ( n150 & n13750 ) | ( n13745 & n13750 ) ;
  assign n13752 = ( n13208 & ~n13227 ) | ( n13208 & 1'b0 ) | ( ~n13227 & 1'b0 ) ;
  assign n13753 = ( n13242 & ~n13224 ) | ( n13242 & n13752 ) | ( ~n13224 & n13752 ) ;
  assign n13754 = n13224 &  n13753 ;
  assign n13755 = ( n13224 & ~n13227 ) | ( n13224 & 1'b0 ) | ( ~n13227 & 1'b0 ) ;
  assign n13756 = ~n13242 & n13755 ;
  assign n13757 = ( n13208 & ~n13756 ) | ( n13208 & n13755 ) | ( ~n13756 & n13755 ) ;
  assign n13758 = ~n13754 & n13757 ;
  assign n13759 = n13209 &  n13216 ;
  assign n13760 = ~n13242 & n13759 ;
  assign n13761 = ( n13230 & ~n13759 ) | ( n13230 & n13760 ) | ( ~n13759 & n13760 ) ;
  assign n13762 = ~n13758 & n13761 ;
  assign n13763 = ~n13751 & n13762 ;
  assign n13764 = ( n133 & ~n13763 ) | ( n133 & n13762 ) | ( ~n13763 & n13762 ) ;
  assign n13767 = n13738 | n13741 ;
  assign n13768 = ( n13735 & ~n145 ) | ( n13735 & n13767 ) | ( ~n145 & n13767 ) ;
  assign n13769 = n150 &  n13768 ;
  assign n13770 = ( n13758 & ~n13769 ) | ( n13758 & 1'b0 ) | ( ~n13769 & 1'b0 ) ;
  assign n13765 = n150 | n13730 ;
  assign n13766 = n13744 | n13765 ;
  assign n13771 = ( n13750 & ~n13766 ) | ( n13750 & 1'b0 ) | ( ~n13766 & 1'b0 ) ;
  assign n13772 = ( n13770 & ~n13750 ) | ( n13770 & n13771 ) | ( ~n13750 & n13771 ) ;
  assign n13774 = ( n133 & n13209 ) | ( n133 & n13216 ) | ( n13209 & n13216 ) ;
  assign n13773 = ( n13209 & ~n13242 ) | ( n13209 & n13216 ) | ( ~n13242 & n13216 ) ;
  assign n13775 = ( n13216 & ~n13773 ) | ( n13216 & 1'b0 ) | ( ~n13773 & 1'b0 ) ;
  assign n13776 = ( n13774 & ~n13216 ) | ( n13774 & n13775 ) | ( ~n13216 & n13775 ) ;
  assign n13777 = n13212 | n13239 ;
  assign n13778 = ( n13234 & ~n13215 ) | ( n13234 & n13777 ) | ( ~n13215 & n13777 ) ;
  assign n13779 = n13215 | n13778 ;
  assign n13780 = ( n13222 & ~n13230 ) | ( n13222 & n13779 ) | ( ~n13230 & n13779 ) ;
  assign n13781 = ( n13222 & ~n13780 ) | ( n13222 & 1'b0 ) | ( ~n13780 & 1'b0 ) ;
  assign n13782 = n13776 | n13781 ;
  assign n13783 = n13772 | n13782 ;
  assign n13784 = ~n13764 |  n13783 ;
  assign n14151 = ( n13577 & ~n13582 ) | ( n13577 & n13784 ) | ( ~n13582 & n13784 ) ;
  assign n14150 = n13590 &  n13784 ;
  assign n14152 = ( n13784 & ~n14151 ) | ( n13784 & n14150 ) | ( ~n14151 & n14150 ) ;
  assign n14153 = ( n14150 & ~n13577 ) | ( n14150 & n14151 ) | ( ~n13577 & n14151 ) ;
  assign n14154 = ( n13582 & ~n14152 ) | ( n13582 & n14153 ) | ( ~n14152 & n14153 ) ;
  assign n14107 = ( n13533 & ~n13538 ) | ( n13533 & n13546 ) | ( ~n13538 & n13546 ) ;
  assign n14106 = n13533 | n13784 ;
  assign n14109 = ( n13533 & ~n14107 ) | ( n13533 & n14106 ) | ( ~n14107 & n14106 ) ;
  assign n14108 = ( n14106 & ~n13546 ) | ( n14106 & n14107 ) | ( ~n13546 & n14107 ) ;
  assign n14110 = ( n13538 & ~n14109 ) | ( n13538 & n14108 ) | ( ~n14109 & n14108 ) ;
  assign n14063 = ( n13489 & ~n13494 ) | ( n13489 & n13502 ) | ( ~n13494 & n13502 ) ;
  assign n14062 = n13489 | n13784 ;
  assign n14065 = ( n13489 & ~n14063 ) | ( n13489 & n14062 ) | ( ~n14063 & n14062 ) ;
  assign n14064 = ( n14062 & ~n13502 ) | ( n14062 & n14063 ) | ( ~n13502 & n14063 ) ;
  assign n14066 = ( n13494 & ~n14065 ) | ( n13494 & n14064 ) | ( ~n14065 & n14064 ) ;
  assign n14041 = ( n13467 & ~n13472 ) | ( n13467 & n13480 ) | ( ~n13472 & n13480 ) ;
  assign n14040 = n13467 | n13784 ;
  assign n14043 = ( n13467 & ~n14041 ) | ( n13467 & n14040 ) | ( ~n14041 & n14040 ) ;
  assign n14042 = ( n14040 & ~n13480 ) | ( n14040 & n14041 ) | ( ~n13480 & n14041 ) ;
  assign n14044 = ( n13472 & ~n14043 ) | ( n13472 & n14042 ) | ( ~n14043 & n14042 ) ;
  assign n13791 = ( x30 & ~n13784 ) | ( x30 & x31 ) | ( ~n13784 & x31 ) ;
  assign n13797 = ( x30 & ~x31 ) | ( x30 & 1'b0 ) | ( ~x31 & 1'b0 ) ;
  assign n13787 = x28 | x29 ;
  assign n13792 = ~x30 & n13787 ;
  assign n13793 = ( x30 & ~n13240 ) | ( x30 & n13792 ) | ( ~n13240 & n13792 ) ;
  assign n13794 = ( n13230 & ~n13222 ) | ( n13230 & n13793 ) | ( ~n13222 & n13793 ) ;
  assign n13795 = n13222 &  n13794 ;
  assign n13796 = ( n13784 & ~x31 ) | ( n13784 & n13795 ) | ( ~x31 & n13795 ) ;
  assign n13798 = ( n13791 & ~n13797 ) | ( n13791 & n13796 ) | ( ~n13797 & n13796 ) ;
  assign n13788 = x30 | n13787 ;
  assign n13789 = x30 &  n13784 ;
  assign n13790 = ( n13242 & ~n13788 ) | ( n13242 & n13789 ) | ( ~n13788 & n13789 ) ;
  assign n13799 = n13790 &  n13798 ;
  assign n13800 = ( n12707 & ~n13798 ) | ( n12707 & n13799 ) | ( ~n13798 & n13799 ) ;
  assign n13801 = n12707 | n13790 ;
  assign n13802 = ( n13798 & ~n13801 ) | ( n13798 & 1'b0 ) | ( ~n13801 & 1'b0 ) ;
  assign n13804 = ( n13242 & ~n13781 ) | ( n13242 & 1'b0 ) | ( ~n13781 & 1'b0 ) ;
  assign n13805 = ( n13772 & ~n13776 ) | ( n13772 & n13804 ) | ( ~n13776 & n13804 ) ;
  assign n13806 = ~n13772 & n13805 ;
  assign n13807 = n13764 &  n13806 ;
  assign n13803 = ~n12708 & n13784 ;
  assign n13808 = ( n13803 & ~n13807 ) | ( n13803 & 1'b0 ) | ( ~n13807 & 1'b0 ) ;
  assign n13809 = ( x32 & n13807 ) | ( x32 & n13808 ) | ( n13807 & n13808 ) ;
  assign n13810 = x32 | n13807 ;
  assign n13811 = n13803 | n13810 ;
  assign n13812 = ~n13809 & n13811 ;
  assign n13813 = n13802 | n13812 ;
  assign n13814 = ~n13800 & n13813 ;
  assign n13818 = ~x32 & n13242 ;
  assign n13819 = ( x33 & ~n13818 ) | ( x33 & 1'b0 ) | ( ~n13818 & 1'b0 ) ;
  assign n13820 = n13254 | n13819 ;
  assign n13815 = ( n13242 & ~x32 ) | ( n13242 & n13249 ) | ( ~x32 & n13249 ) ;
  assign n13816 = x32 &  n13815 ;
  assign n13817 = ( n13244 & ~n13816 ) | ( n13244 & n13249 ) | ( ~n13816 & n13249 ) ;
  assign n13821 = ( n13784 & ~n13820 ) | ( n13784 & n13817 ) | ( ~n13820 & n13817 ) ;
  assign n13823 = ( n13784 & ~n13821 ) | ( n13784 & 1'b0 ) | ( ~n13821 & 1'b0 ) ;
  assign n13822 = ~n13817 & n13821 ;
  assign n13824 = ( n13820 & ~n13823 ) | ( n13820 & n13822 ) | ( ~n13823 & n13822 ) ;
  assign n13825 = ( n13814 & ~n12187 ) | ( n13814 & n13824 ) | ( ~n12187 & n13824 ) ;
  assign n13826 = ( n11674 & ~n13825 ) | ( n11674 & 1'b0 ) | ( ~n13825 & 1'b0 ) ;
  assign n13827 = ~n13277 & n13280 ;
  assign n13828 = ( n13263 & ~n13827 ) | ( n13263 & n13277 ) | ( ~n13827 & n13277 ) ;
  assign n13829 = ( n13784 & n13827 ) | ( n13784 & n13828 ) | ( n13827 & n13828 ) ;
  assign n13830 = ( n13277 & ~n13828 ) | ( n13277 & n13784 ) | ( ~n13828 & n13784 ) ;
  assign n13831 = ( n13263 & ~n13829 ) | ( n13263 & n13830 ) | ( ~n13829 & n13830 ) ;
  assign n13832 = n12187 | n13800 ;
  assign n13833 = ( n13813 & ~n13832 ) | ( n13813 & 1'b0 ) | ( ~n13832 & 1'b0 ) ;
  assign n13834 = n13824 | n13833 ;
  assign n13835 = ~n13790 & n13798 ;
  assign n13836 = ( n13812 & ~n12707 ) | ( n13812 & n13835 ) | ( ~n12707 & n13835 ) ;
  assign n13837 = ( n12187 & ~n13836 ) | ( n12187 & 1'b0 ) | ( ~n13836 & 1'b0 ) ;
  assign n13838 = n11674 | n13837 ;
  assign n13839 = ( n13834 & ~n13838 ) | ( n13834 & 1'b0 ) | ( ~n13838 & 1'b0 ) ;
  assign n13840 = n13831 | n13839 ;
  assign n13841 = ~n13826 & n13840 ;
  assign n13842 = n13265 | n13784 ;
  assign n13843 = ( n13265 & ~n13282 ) | ( n13265 & n13275 ) | ( ~n13282 & n13275 ) ;
  assign n13844 = ( n13282 & n13842 ) | ( n13282 & n13843 ) | ( n13842 & n13843 ) ;
  assign n13845 = ( n13265 & ~n13843 ) | ( n13265 & n13842 ) | ( ~n13843 & n13842 ) ;
  assign n13846 = ( n13275 & ~n13844 ) | ( n13275 & n13845 ) | ( ~n13844 & n13845 ) ;
  assign n13847 = ( n13841 & ~n11176 ) | ( n13841 & n13846 ) | ( ~n11176 & n13846 ) ;
  assign n13848 = ( n10685 & ~n13847 ) | ( n10685 & 1'b0 ) | ( ~n13847 & 1'b0 ) ;
  assign n13849 = n13302 | n13784 ;
  assign n13850 = ( n13289 & ~n13302 ) | ( n13289 & n13298 ) | ( ~n13302 & n13298 ) ;
  assign n13852 = ( n13302 & n13849 ) | ( n13302 & n13850 ) | ( n13849 & n13850 ) ;
  assign n13851 = ( n13298 & ~n13850 ) | ( n13298 & n13849 ) | ( ~n13850 & n13849 ) ;
  assign n13853 = ( n13289 & ~n13852 ) | ( n13289 & n13851 ) | ( ~n13852 & n13851 ) ;
  assign n13854 = n11176 | n13826 ;
  assign n13855 = ( n13840 & ~n13854 ) | ( n13840 & 1'b0 ) | ( ~n13854 & 1'b0 ) ;
  assign n13856 = n13846 | n13855 ;
  assign n13857 = ( n13834 & ~n13837 ) | ( n13834 & 1'b0 ) | ( ~n13837 & 1'b0 ) ;
  assign n13858 = ( n13831 & ~n11674 ) | ( n13831 & n13857 ) | ( ~n11674 & n13857 ) ;
  assign n13859 = ( n11176 & ~n13858 ) | ( n11176 & 1'b0 ) | ( ~n13858 & 1'b0 ) ;
  assign n13860 = n10685 | n13859 ;
  assign n13861 = ( n13856 & ~n13860 ) | ( n13856 & 1'b0 ) | ( ~n13860 & 1'b0 ) ;
  assign n13862 = n13853 | n13861 ;
  assign n13863 = ~n13848 & n13862 ;
  assign n13865 = ( n13291 & ~n13296 ) | ( n13291 & n13784 ) | ( ~n13296 & n13784 ) ;
  assign n13864 = n13304 &  n13784 ;
  assign n13866 = ( n13784 & ~n13865 ) | ( n13784 & n13864 ) | ( ~n13865 & n13864 ) ;
  assign n13867 = ( n13864 & ~n13291 ) | ( n13864 & n13865 ) | ( ~n13291 & n13865 ) ;
  assign n13868 = ( n13296 & ~n13866 ) | ( n13296 & n13867 ) | ( ~n13866 & n13867 ) ;
  assign n13869 = ( n13863 & ~n10209 ) | ( n13863 & n13868 ) | ( ~n10209 & n13868 ) ;
  assign n13870 = n9740 | n13869 ;
  assign n13871 = n13324 | n13784 ;
  assign n13872 = ( n13311 & ~n13320 ) | ( n13311 & n13324 ) | ( ~n13320 & n13324 ) ;
  assign n13873 = ( n13320 & n13871 ) | ( n13320 & n13872 ) | ( n13871 & n13872 ) ;
  assign n13874 = ( n13324 & ~n13872 ) | ( n13324 & n13871 ) | ( ~n13872 & n13871 ) ;
  assign n13875 = ( n13311 & ~n13873 ) | ( n13311 & n13874 ) | ( ~n13873 & n13874 ) ;
  assign n13876 = n10209 | n13848 ;
  assign n13877 = ( n13862 & ~n13876 ) | ( n13862 & 1'b0 ) | ( ~n13876 & 1'b0 ) ;
  assign n13878 = n13868 | n13877 ;
  assign n13879 = ( n13856 & ~n13859 ) | ( n13856 & 1'b0 ) | ( ~n13859 & 1'b0 ) ;
  assign n13880 = ( n13853 & ~n10685 ) | ( n13853 & n13879 ) | ( ~n10685 & n13879 ) ;
  assign n13881 = ( n10209 & ~n13880 ) | ( n10209 & 1'b0 ) | ( ~n13880 & 1'b0 ) ;
  assign n13882 = ( n9740 & ~n13881 ) | ( n9740 & 1'b0 ) | ( ~n13881 & 1'b0 ) ;
  assign n13883 = n13878 &  n13882 ;
  assign n13884 = n13875 | n13883 ;
  assign n13885 = n13870 &  n13884 ;
  assign n13886 = ( n13313 & ~n13784 ) | ( n13313 & 1'b0 ) | ( ~n13784 & 1'b0 ) ;
  assign n13887 = ( n13313 & n13318 ) | ( n13313 & n13326 ) | ( n13318 & n13326 ) ;
  assign n13888 = ( n13886 & ~n13326 ) | ( n13886 & n13887 ) | ( ~n13326 & n13887 ) ;
  assign n13889 = ( n13313 & ~n13887 ) | ( n13313 & n13886 ) | ( ~n13887 & n13886 ) ;
  assign n13890 = ( n13318 & ~n13888 ) | ( n13318 & n13889 ) | ( ~n13888 & n13889 ) ;
  assign n13891 = ( n13885 & ~n9286 ) | ( n13885 & n13890 ) | ( ~n9286 & n13890 ) ;
  assign n13892 = ( n8839 & ~n13891 ) | ( n8839 & 1'b0 ) | ( ~n13891 & 1'b0 ) ;
  assign n13893 = n13346 | n13784 ;
  assign n13894 = ( n13333 & ~n13342 ) | ( n13333 & n13346 ) | ( ~n13342 & n13346 ) ;
  assign n13895 = ( n13342 & n13893 ) | ( n13342 & n13894 ) | ( n13893 & n13894 ) ;
  assign n13896 = ( n13346 & ~n13894 ) | ( n13346 & n13893 ) | ( ~n13894 & n13893 ) ;
  assign n13897 = ( n13333 & ~n13895 ) | ( n13333 & n13896 ) | ( ~n13895 & n13896 ) ;
  assign n13898 = ~n9286 & n13870 ;
  assign n13899 = n13884 &  n13898 ;
  assign n13900 = n13890 | n13899 ;
  assign n13901 = ( n13878 & ~n13881 ) | ( n13878 & 1'b0 ) | ( ~n13881 & 1'b0 ) ;
  assign n13902 = ( n9740 & n13875 ) | ( n9740 & n13901 ) | ( n13875 & n13901 ) ;
  assign n13903 = ( n9286 & ~n13902 ) | ( n9286 & 1'b0 ) | ( ~n13902 & 1'b0 ) ;
  assign n13904 = n8839 | n13903 ;
  assign n13905 = ( n13900 & ~n13904 ) | ( n13900 & 1'b0 ) | ( ~n13904 & 1'b0 ) ;
  assign n13906 = n13897 | n13905 ;
  assign n13907 = ~n13892 & n13906 ;
  assign n13908 = n13335 | n13784 ;
  assign n13909 = ( n13335 & ~n13348 ) | ( n13335 & n13340 ) | ( ~n13348 & n13340 ) ;
  assign n13910 = ( n13348 & n13908 ) | ( n13348 & n13909 ) | ( n13908 & n13909 ) ;
  assign n13911 = ( n13335 & ~n13909 ) | ( n13335 & n13908 ) | ( ~n13909 & n13908 ) ;
  assign n13912 = ( n13340 & ~n13910 ) | ( n13340 & n13911 ) | ( ~n13910 & n13911 ) ;
  assign n13913 = ( n13907 & ~n8407 ) | ( n13907 & n13912 ) | ( ~n8407 & n13912 ) ;
  assign n13914 = ( n7982 & ~n13913 ) | ( n7982 & 1'b0 ) | ( ~n13913 & 1'b0 ) ;
  assign n13915 = n13368 | n13784 ;
  assign n13916 = ( n13355 & ~n13368 ) | ( n13355 & n13364 ) | ( ~n13368 & n13364 ) ;
  assign n13918 = ( n13368 & n13915 ) | ( n13368 & n13916 ) | ( n13915 & n13916 ) ;
  assign n13917 = ( n13364 & ~n13916 ) | ( n13364 & n13915 ) | ( ~n13916 & n13915 ) ;
  assign n13919 = ( n13355 & ~n13918 ) | ( n13355 & n13917 ) | ( ~n13918 & n13917 ) ;
  assign n13920 = n8407 | n13892 ;
  assign n13921 = ( n13906 & ~n13920 ) | ( n13906 & 1'b0 ) | ( ~n13920 & 1'b0 ) ;
  assign n13922 = n13912 | n13921 ;
  assign n13923 = ( n13900 & ~n13903 ) | ( n13900 & 1'b0 ) | ( ~n13903 & 1'b0 ) ;
  assign n13924 = ( n13897 & ~n8839 ) | ( n13897 & n13923 ) | ( ~n8839 & n13923 ) ;
  assign n13925 = ( n8407 & ~n13924 ) | ( n8407 & 1'b0 ) | ( ~n13924 & 1'b0 ) ;
  assign n13926 = n7982 | n13925 ;
  assign n13927 = ( n13922 & ~n13926 ) | ( n13922 & 1'b0 ) | ( ~n13926 & 1'b0 ) ;
  assign n13928 = n13919 | n13927 ;
  assign n13929 = ~n13914 & n13928 ;
  assign n13930 = n13357 | n13784 ;
  assign n13931 = ( n13362 & ~n13357 ) | ( n13362 & n13370 ) | ( ~n13357 & n13370 ) ;
  assign n13933 = ( n13357 & n13930 ) | ( n13357 & n13931 ) | ( n13930 & n13931 ) ;
  assign n13932 = ( n13370 & ~n13931 ) | ( n13370 & n13930 ) | ( ~n13931 & n13930 ) ;
  assign n13934 = ( n13362 & ~n13933 ) | ( n13362 & n13932 ) | ( ~n13933 & n13932 ) ;
  assign n13935 = ( n7572 & n13929 ) | ( n7572 & n13934 ) | ( n13929 & n13934 ) ;
  assign n13936 = n7169 | n13935 ;
  assign n13938 = ( n13386 & ~n13377 ) | ( n13386 & n13390 ) | ( ~n13377 & n13390 ) ;
  assign n13937 = ( n13390 & ~n13784 ) | ( n13390 & 1'b0 ) | ( ~n13784 & 1'b0 ) ;
  assign n13940 = ( n13390 & ~n13938 ) | ( n13390 & n13937 ) | ( ~n13938 & n13937 ) ;
  assign n13939 = ( n13937 & ~n13386 ) | ( n13937 & n13938 ) | ( ~n13386 & n13938 ) ;
  assign n13941 = ( n13377 & ~n13940 ) | ( n13377 & n13939 ) | ( ~n13940 & n13939 ) ;
  assign n13942 = ( n7572 & ~n13914 ) | ( n7572 & 1'b0 ) | ( ~n13914 & 1'b0 ) ;
  assign n13943 = n13928 &  n13942 ;
  assign n13944 = n13934 | n13943 ;
  assign n13945 = ( n13922 & ~n13925 ) | ( n13922 & 1'b0 ) | ( ~n13925 & 1'b0 ) ;
  assign n13946 = ( n13919 & ~n7982 ) | ( n13919 & n13945 ) | ( ~n7982 & n13945 ) ;
  assign n13947 = n7572 | n13946 ;
  assign n13948 = n7169 &  n13947 ;
  assign n13949 = n13944 &  n13948 ;
  assign n13950 = n13941 | n13949 ;
  assign n13951 = n13936 &  n13950 ;
  assign n13952 = ( n13379 & ~n13784 ) | ( n13379 & 1'b0 ) | ( ~n13784 & 1'b0 ) ;
  assign n13953 = ( n13379 & n13384 ) | ( n13379 & n13392 ) | ( n13384 & n13392 ) ;
  assign n13954 = ( n13952 & ~n13392 ) | ( n13952 & n13953 ) | ( ~n13392 & n13953 ) ;
  assign n13955 = ( n13379 & ~n13953 ) | ( n13379 & n13952 ) | ( ~n13953 & n13952 ) ;
  assign n13956 = ( n13384 & ~n13954 ) | ( n13384 & n13955 ) | ( ~n13954 & n13955 ) ;
  assign n13957 = ( n13951 & ~n6781 ) | ( n13951 & n13956 ) | ( ~n6781 & n13956 ) ;
  assign n13958 = n6399 | n13957 ;
  assign n13959 = n13412 | n13784 ;
  assign n13960 = ( n13399 & ~n13408 ) | ( n13399 & n13412 ) | ( ~n13408 & n13412 ) ;
  assign n13961 = ( n13408 & n13959 ) | ( n13408 & n13960 ) | ( n13959 & n13960 ) ;
  assign n13962 = ( n13412 & ~n13960 ) | ( n13412 & n13959 ) | ( ~n13960 & n13959 ) ;
  assign n13963 = ( n13399 & ~n13961 ) | ( n13399 & n13962 ) | ( ~n13961 & n13962 ) ;
  assign n13964 = ~n6781 & n13936 ;
  assign n13965 = n13950 &  n13964 ;
  assign n13966 = n13956 | n13965 ;
  assign n13967 = n13944 &  n13947 ;
  assign n13968 = ( n7169 & n13941 ) | ( n7169 & n13967 ) | ( n13941 & n13967 ) ;
  assign n13969 = ( n6781 & ~n13968 ) | ( n6781 & 1'b0 ) | ( ~n13968 & 1'b0 ) ;
  assign n13970 = ( n6399 & ~n13969 ) | ( n6399 & 1'b0 ) | ( ~n13969 & 1'b0 ) ;
  assign n13971 = n13966 &  n13970 ;
  assign n13972 = n13963 | n13971 ;
  assign n13973 = n13958 &  n13972 ;
  assign n13975 = ( n13401 & ~n13406 ) | ( n13401 & n13414 ) | ( ~n13406 & n13414 ) ;
  assign n13974 = ( n13401 & ~n13784 ) | ( n13401 & 1'b0 ) | ( ~n13784 & 1'b0 ) ;
  assign n13977 = ( n13401 & ~n13975 ) | ( n13401 & n13974 ) | ( ~n13975 & n13974 ) ;
  assign n13976 = ( n13974 & ~n13414 ) | ( n13974 & n13975 ) | ( ~n13414 & n13975 ) ;
  assign n13978 = ( n13406 & ~n13977 ) | ( n13406 & n13976 ) | ( ~n13977 & n13976 ) ;
  assign n13979 = ( n6032 & ~n13973 ) | ( n6032 & n13978 ) | ( ~n13973 & n13978 ) ;
  assign n13980 = ~n5672 & n13979 ;
  assign n13981 = n13434 | n13784 ;
  assign n13982 = ( n13421 & ~n13434 ) | ( n13421 & n13430 ) | ( ~n13434 & n13430 ) ;
  assign n13984 = ( n13434 & n13981 ) | ( n13434 & n13982 ) | ( n13981 & n13982 ) ;
  assign n13983 = ( n13430 & ~n13982 ) | ( n13430 & n13981 ) | ( ~n13982 & n13981 ) ;
  assign n13985 = ( n13421 & ~n13984 ) | ( n13421 & n13983 ) | ( ~n13984 & n13983 ) ;
  assign n13986 = ~n6032 & n13958 ;
  assign n13987 = n13972 &  n13986 ;
  assign n13988 = ( n13978 & ~n13987 ) | ( n13978 & 1'b0 ) | ( ~n13987 & 1'b0 ) ;
  assign n13989 = ( n13966 & ~n13969 ) | ( n13966 & 1'b0 ) | ( ~n13969 & 1'b0 ) ;
  assign n13990 = ( n6399 & n13963 ) | ( n6399 & n13989 ) | ( n13963 & n13989 ) ;
  assign n13991 = ( n6032 & ~n13990 ) | ( n6032 & 1'b0 ) | ( ~n13990 & 1'b0 ) ;
  assign n13992 = ( n5672 & ~n13991 ) | ( n5672 & 1'b0 ) | ( ~n13991 & 1'b0 ) ;
  assign n13993 = ~n13988 & n13992 ;
  assign n13994 = ( n13985 & ~n13993 ) | ( n13985 & 1'b0 ) | ( ~n13993 & 1'b0 ) ;
  assign n13995 = n13980 | n13994 ;
  assign n13996 = n13423 | n13784 ;
  assign n13997 = ( n13423 & ~n13436 ) | ( n13423 & n13428 ) | ( ~n13436 & n13428 ) ;
  assign n13998 = ( n13436 & n13996 ) | ( n13436 & n13997 ) | ( n13996 & n13997 ) ;
  assign n13999 = ( n13423 & ~n13997 ) | ( n13423 & n13996 ) | ( ~n13997 & n13996 ) ;
  assign n14000 = ( n13428 & ~n13998 ) | ( n13428 & n13999 ) | ( ~n13998 & n13999 ) ;
  assign n14001 = ( n5327 & n13995 ) | ( n5327 & n14000 ) | ( n13995 & n14000 ) ;
  assign n14002 = n4990 &  n14001 ;
  assign n14004 = ( n13452 & ~n13443 ) | ( n13452 & n13456 ) | ( ~n13443 & n13456 ) ;
  assign n14003 = n13456 | n13784 ;
  assign n14006 = ( n13456 & ~n14004 ) | ( n13456 & n14003 ) | ( ~n14004 & n14003 ) ;
  assign n14005 = ( n14003 & ~n13452 ) | ( n14003 & n14004 ) | ( ~n13452 & n14004 ) ;
  assign n14007 = ( n13443 & ~n14006 ) | ( n13443 & n14005 ) | ( ~n14006 & n14005 ) ;
  assign n14008 = n5327 | n13980 ;
  assign n14009 = n13994 | n14008 ;
  assign n14010 = n14000 &  n14009 ;
  assign n14011 = n13988 | n13991 ;
  assign n14012 = ( n13985 & ~n5672 ) | ( n13985 & n14011 ) | ( ~n5672 & n14011 ) ;
  assign n14013 = n5327 &  n14012 ;
  assign n14014 = n4990 | n14013 ;
  assign n14015 = n14010 | n14014 ;
  assign n14016 = n14007 &  n14015 ;
  assign n14017 = n14002 | n14016 ;
  assign n14018 = n13445 | n13784 ;
  assign n14019 = ( n13445 & n13450 ) | ( n13445 & n13458 ) | ( n13450 & n13458 ) ;
  assign n14020 = ( n14018 & ~n13458 ) | ( n14018 & n14019 ) | ( ~n13458 & n14019 ) ;
  assign n14021 = ( n13445 & ~n14019 ) | ( n13445 & n14018 ) | ( ~n14019 & n14018 ) ;
  assign n14022 = ( n13450 & ~n14020 ) | ( n13450 & n14021 ) | ( ~n14020 & n14021 ) ;
  assign n14023 = ( n4668 & n14017 ) | ( n4668 & n14022 ) | ( n14017 & n14022 ) ;
  assign n14024 = n4353 &  n14023 ;
  assign n14025 = n13478 | n13784 ;
  assign n14026 = ( n13465 & n13474 ) | ( n13465 & n13478 ) | ( n13474 & n13478 ) ;
  assign n14027 = ( n14025 & ~n13474 ) | ( n14025 & n14026 ) | ( ~n13474 & n14026 ) ;
  assign n14028 = ( n13478 & ~n14026 ) | ( n13478 & n14025 ) | ( ~n14026 & n14025 ) ;
  assign n14029 = ( n13465 & ~n14027 ) | ( n13465 & n14028 ) | ( ~n14027 & n14028 ) ;
  assign n14030 = n4668 | n14002 ;
  assign n14031 = n14016 | n14030 ;
  assign n14032 = n14022 &  n14031 ;
  assign n14033 = n14010 | n14013 ;
  assign n14034 = ( n4990 & n14007 ) | ( n4990 & n14033 ) | ( n14007 & n14033 ) ;
  assign n14035 = n4668 &  n14034 ;
  assign n14036 = n4353 | n14035 ;
  assign n14037 = n14032 | n14036 ;
  assign n14038 = ~n14029 & n14037 ;
  assign n14039 = n14024 | n14038 ;
  assign n14045 = ( n4053 & ~n14044 ) | ( n4053 & n14039 ) | ( ~n14044 & n14039 ) ;
  assign n14046 = n3760 &  n14045 ;
  assign n14048 = ( n13496 & ~n13487 ) | ( n13496 & n13500 ) | ( ~n13487 & n13500 ) ;
  assign n14047 = n13500 | n13784 ;
  assign n14050 = ( n13500 & ~n14048 ) | ( n13500 & n14047 ) | ( ~n14048 & n14047 ) ;
  assign n14049 = ( n14047 & ~n13496 ) | ( n14047 & n14048 ) | ( ~n13496 & n14048 ) ;
  assign n14051 = ( n13487 & ~n14050 ) | ( n13487 & n14049 ) | ( ~n14050 & n14049 ) ;
  assign n14052 = n4053 | n14024 ;
  assign n14053 = n14038 | n14052 ;
  assign n14054 = ~n14044 & n14053 ;
  assign n14055 = n14032 | n14035 ;
  assign n14056 = ( n4353 & ~n14029 ) | ( n4353 & n14055 ) | ( ~n14029 & n14055 ) ;
  assign n14057 = n4053 &  n14056 ;
  assign n14058 = n3760 | n14057 ;
  assign n14059 = n14054 | n14058 ;
  assign n14060 = n14051 &  n14059 ;
  assign n14061 = n14046 | n14060 ;
  assign n14067 = ( n3482 & ~n14066 ) | ( n3482 & n14061 ) | ( ~n14066 & n14061 ) ;
  assign n14068 = n3211 &  n14067 ;
  assign n14070 = ( n13518 & ~n13509 ) | ( n13518 & n13522 ) | ( ~n13509 & n13522 ) ;
  assign n14069 = n13522 | n13784 ;
  assign n14072 = ( n13522 & ~n14070 ) | ( n13522 & n14069 ) | ( ~n14070 & n14069 ) ;
  assign n14071 = ( n14069 & ~n13518 ) | ( n14069 & n14070 ) | ( ~n13518 & n14070 ) ;
  assign n14073 = ( n13509 & ~n14072 ) | ( n13509 & n14071 ) | ( ~n14072 & n14071 ) ;
  assign n14074 = n3482 | n14046 ;
  assign n14075 = n14060 | n14074 ;
  assign n14076 = ~n14066 & n14075 ;
  assign n14077 = n14054 | n14057 ;
  assign n14078 = ( n3760 & n14051 ) | ( n3760 & n14077 ) | ( n14051 & n14077 ) ;
  assign n14079 = n3482 &  n14078 ;
  assign n14080 = n3211 | n14079 ;
  assign n14081 = n14076 | n14080 ;
  assign n14082 = n14073 &  n14081 ;
  assign n14083 = n14068 | n14082 ;
  assign n14084 = n13511 | n13784 ;
  assign n14085 = ( n13511 & n13516 ) | ( n13511 & n13524 ) | ( n13516 & n13524 ) ;
  assign n14086 = ( n14084 & ~n13524 ) | ( n14084 & n14085 ) | ( ~n13524 & n14085 ) ;
  assign n14087 = ( n13511 & ~n14085 ) | ( n13511 & n14084 ) | ( ~n14085 & n14084 ) ;
  assign n14088 = ( n13516 & ~n14086 ) | ( n13516 & n14087 ) | ( ~n14086 & n14087 ) ;
  assign n14089 = ( n2955 & n14083 ) | ( n2955 & n14088 ) | ( n14083 & n14088 ) ;
  assign n14090 = n2706 &  n14089 ;
  assign n14091 = n13544 | n13784 ;
  assign n14092 = ( n13531 & n13540 ) | ( n13531 & n13544 ) | ( n13540 & n13544 ) ;
  assign n14093 = ( n14091 & ~n13540 ) | ( n14091 & n14092 ) | ( ~n13540 & n14092 ) ;
  assign n14094 = ( n13544 & ~n14092 ) | ( n13544 & n14091 ) | ( ~n14092 & n14091 ) ;
  assign n14095 = ( n13531 & ~n14093 ) | ( n13531 & n14094 ) | ( ~n14093 & n14094 ) ;
  assign n14096 = n2955 | n14068 ;
  assign n14097 = n14082 | n14096 ;
  assign n14098 = n14088 &  n14097 ;
  assign n14099 = n14076 | n14079 ;
  assign n14100 = ( n3211 & n14073 ) | ( n3211 & n14099 ) | ( n14073 & n14099 ) ;
  assign n14101 = n2955 &  n14100 ;
  assign n14102 = n2706 | n14101 ;
  assign n14103 = n14098 | n14102 ;
  assign n14104 = ~n14095 & n14103 ;
  assign n14105 = n14090 | n14104 ;
  assign n14111 = ( n2472 & ~n14110 ) | ( n2472 & n14105 ) | ( ~n14110 & n14105 ) ;
  assign n14112 = n2245 &  n14111 ;
  assign n14114 = ( n13562 & ~n13553 ) | ( n13562 & n13566 ) | ( ~n13553 & n13566 ) ;
  assign n14113 = n13566 | n13784 ;
  assign n14116 = ( n13566 & ~n14114 ) | ( n13566 & n14113 ) | ( ~n14114 & n14113 ) ;
  assign n14115 = ( n14113 & ~n13562 ) | ( n14113 & n14114 ) | ( ~n13562 & n14114 ) ;
  assign n14117 = ( n13553 & ~n14116 ) | ( n13553 & n14115 ) | ( ~n14116 & n14115 ) ;
  assign n14118 = n2472 | n14090 ;
  assign n14119 = n14104 | n14118 ;
  assign n14120 = ~n14110 & n14119 ;
  assign n14121 = n14098 | n14101 ;
  assign n14122 = ( n2706 & ~n14095 ) | ( n2706 & n14121 ) | ( ~n14095 & n14121 ) ;
  assign n14123 = n2472 &  n14122 ;
  assign n14124 = n2245 | n14123 ;
  assign n14125 = n14120 | n14124 ;
  assign n14126 = ~n14117 & n14125 ;
  assign n14127 = n14112 | n14126 ;
  assign n14128 = ~n13568 & n13784 ;
  assign n14129 = ( n13555 & ~n14128 ) | ( n13555 & n13784 ) | ( ~n14128 & n13784 ) ;
  assign n14130 = ( n13560 & ~n13555 ) | ( n13560 & n14129 ) | ( ~n13555 & n14129 ) ;
  assign n14131 = ( n13555 & ~n14129 ) | ( n13555 & n13560 ) | ( ~n14129 & n13560 ) ;
  assign n14132 = ( n14130 & ~n13560 ) | ( n14130 & n14131 ) | ( ~n13560 & n14131 ) ;
  assign n14133 = ( n2033 & ~n14127 ) | ( n2033 & n14132 ) | ( ~n14127 & n14132 ) ;
  assign n14134 = ( n1827 & ~n14133 ) | ( n1827 & 1'b0 ) | ( ~n14133 & 1'b0 ) ;
  assign n14135 = n13588 | n13784 ;
  assign n14136 = ( n13575 & ~n13588 ) | ( n13575 & n13584 ) | ( ~n13588 & n13584 ) ;
  assign n14138 = ( n13588 & n14135 ) | ( n13588 & n14136 ) | ( n14135 & n14136 ) ;
  assign n14137 = ( n13584 & ~n14136 ) | ( n13584 & n14135 ) | ( ~n14136 & n14135 ) ;
  assign n14139 = ( n13575 & ~n14138 ) | ( n13575 & n14137 ) | ( ~n14138 & n14137 ) ;
  assign n14140 = ( n2033 & ~n14112 ) | ( n2033 & 1'b0 ) | ( ~n14112 & 1'b0 ) ;
  assign n14141 = ~n14126 & n14140 ;
  assign n14142 = n14132 | n14141 ;
  assign n14143 = n14120 | n14123 ;
  assign n14144 = ( n2245 & ~n14117 ) | ( n2245 & n14143 ) | ( ~n14117 & n14143 ) ;
  assign n14145 = ~n2033 & n14144 ;
  assign n14146 = n1827 | n14145 ;
  assign n14147 = ( n14142 & ~n14146 ) | ( n14142 & 1'b0 ) | ( ~n14146 & 1'b0 ) ;
  assign n14148 = n14139 | n14147 ;
  assign n14149 = ~n14134 & n14148 ;
  assign n14155 = ( n1636 & ~n14154 ) | ( n1636 & n14149 ) | ( ~n14154 & n14149 ) ;
  assign n14156 = n1452 | n14155 ;
  assign n14259 = ~n13699 & n13784 ;
  assign n14260 = ( n13686 & n13691 ) | ( n13686 & n13784 ) | ( n13691 & n13784 ) ;
  assign n14262 = ( n14259 & ~n13686 ) | ( n14259 & n14260 ) | ( ~n13686 & n14260 ) ;
  assign n14261 = ( n13784 & ~n14260 ) | ( n13784 & n14259 ) | ( ~n14260 & n14259 ) ;
  assign n14263 = ( n13691 & ~n14262 ) | ( n13691 & n14261 ) | ( ~n14262 & n14261 ) ;
  assign n14157 = n13605 | n13784 ;
  assign n14158 = ( n13597 & ~n13605 ) | ( n13597 & n13601 ) | ( ~n13605 & n13601 ) ;
  assign n14160 = ( n13605 & n14157 ) | ( n13605 & n14158 ) | ( n14157 & n14158 ) ;
  assign n14159 = ( n13601 & ~n14158 ) | ( n13601 & n14157 ) | ( ~n14158 & n14157 ) ;
  assign n14161 = ( n13597 & ~n14160 ) | ( n13597 & n14159 ) | ( ~n14160 & n14159 ) ;
  assign n14162 = ( n1636 & ~n14134 ) | ( n1636 & 1'b0 ) | ( ~n14134 & 1'b0 ) ;
  assign n14163 = n14148 &  n14162 ;
  assign n14164 = ( n14154 & ~n14163 ) | ( n14154 & 1'b0 ) | ( ~n14163 & 1'b0 ) ;
  assign n14165 = ( n14142 & ~n14145 ) | ( n14142 & 1'b0 ) | ( ~n14145 & 1'b0 ) ;
  assign n14166 = ( n14139 & ~n1827 ) | ( n14139 & n14165 ) | ( ~n1827 & n14165 ) ;
  assign n14167 = n1636 | n14166 ;
  assign n14168 = n1452 &  n14167 ;
  assign n14169 = ~n14164 & n14168 ;
  assign n14170 = n14161 | n14169 ;
  assign n14171 = n14156 &  n14170 ;
  assign n14172 = ( n13599 & ~n13611 ) | ( n13599 & n13607 ) | ( ~n13611 & n13607 ) ;
  assign n14173 = ( n13607 & ~n14172 ) | ( n13607 & n13784 ) | ( ~n14172 & n13784 ) ;
  assign n14174 = ( n13784 & ~n13599 ) | ( n13784 & n14172 ) | ( ~n13599 & n14172 ) ;
  assign n14175 = ( n13611 & ~n14173 ) | ( n13611 & n14174 ) | ( ~n14173 & n14174 ) ;
  assign n14176 = ( n14171 & ~n1283 ) | ( n14171 & n14175 ) | ( ~n1283 & n14175 ) ;
  assign n14177 = n1122 | n14176 ;
  assign n14178 = n13631 | n13784 ;
  assign n14179 = ( n13618 & ~n13627 ) | ( n13618 & n13631 ) | ( ~n13627 & n13631 ) ;
  assign n14180 = ( n13627 & n14178 ) | ( n13627 & n14179 ) | ( n14178 & n14179 ) ;
  assign n14181 = ( n13631 & ~n14179 ) | ( n13631 & n14178 ) | ( ~n14179 & n14178 ) ;
  assign n14182 = ( n13618 & ~n14180 ) | ( n13618 & n14181 ) | ( ~n14180 & n14181 ) ;
  assign n14183 = ~n1283 & n14156 ;
  assign n14184 = n14170 &  n14183 ;
  assign n14185 = n14175 | n14184 ;
  assign n14186 = ~n14164 & n14167 ;
  assign n14187 = ( n1452 & n14161 ) | ( n1452 & n14186 ) | ( n14161 & n14186 ) ;
  assign n14188 = ( n1283 & ~n14187 ) | ( n1283 & 1'b0 ) | ( ~n14187 & 1'b0 ) ;
  assign n14189 = ( n1122 & ~n14188 ) | ( n1122 & 1'b0 ) | ( ~n14188 & 1'b0 ) ;
  assign n14190 = n14185 &  n14189 ;
  assign n14191 = ( n14182 & ~n14190 ) | ( n14182 & 1'b0 ) | ( ~n14190 & 1'b0 ) ;
  assign n14192 = ( n14177 & ~n14191 ) | ( n14177 & 1'b0 ) | ( ~n14191 & 1'b0 ) ;
  assign n14193 = n13633 &  n13784 ;
  assign n14194 = ( n13620 & ~n14193 ) | ( n13620 & n13784 ) | ( ~n14193 & n13784 ) ;
  assign n14195 = ( n13625 & ~n13620 ) | ( n13625 & n14194 ) | ( ~n13620 & n14194 ) ;
  assign n14196 = ( n13620 & ~n14194 ) | ( n13620 & n13625 ) | ( ~n14194 & n13625 ) ;
  assign n14197 = ( n14195 & ~n13625 ) | ( n14195 & n14196 ) | ( ~n13625 & n14196 ) ;
  assign n14198 = ( n976 & n14192 ) | ( n976 & n14197 ) | ( n14192 & n14197 ) ;
  assign n14199 = ( n837 & ~n14198 ) | ( n837 & 1'b0 ) | ( ~n14198 & 1'b0 ) ;
  assign n14201 = ( n13649 & ~n13640 ) | ( n13649 & n13653 ) | ( ~n13640 & n13653 ) ;
  assign n14200 = ( n13653 & ~n13784 ) | ( n13653 & 1'b0 ) | ( ~n13784 & 1'b0 ) ;
  assign n14203 = ( n13653 & ~n14201 ) | ( n13653 & n14200 ) | ( ~n14201 & n14200 ) ;
  assign n14202 = ( n14200 & ~n13649 ) | ( n14200 & n14201 ) | ( ~n13649 & n14201 ) ;
  assign n14204 = ( n13640 & ~n14203 ) | ( n13640 & n14202 ) | ( ~n14203 & n14202 ) ;
  assign n14205 = n976 &  n14177 ;
  assign n14206 = ~n14191 & n14205 ;
  assign n14207 = n14197 | n14206 ;
  assign n14208 = ( n14185 & ~n14188 ) | ( n14185 & 1'b0 ) | ( ~n14188 & 1'b0 ) ;
  assign n14209 = ( n1122 & ~n14182 ) | ( n1122 & n14208 ) | ( ~n14182 & n14208 ) ;
  assign n14210 = n976 | n14209 ;
  assign n14211 = ~n837 & n14210 ;
  assign n14212 = n14207 &  n14211 ;
  assign n14213 = ( n14204 & ~n14212 ) | ( n14204 & 1'b0 ) | ( ~n14212 & 1'b0 ) ;
  assign n14214 = n14199 | n14213 ;
  assign n14215 = n13655 &  n13784 ;
  assign n14216 = ( n13642 & n13647 ) | ( n13642 & n13784 ) | ( n13647 & n13784 ) ;
  assign n14218 = ( n14215 & ~n13642 ) | ( n14215 & n14216 ) | ( ~n13642 & n14216 ) ;
  assign n14217 = ( n13784 & ~n14216 ) | ( n13784 & n14215 ) | ( ~n14216 & n14215 ) ;
  assign n14219 = ( n13647 & ~n14218 ) | ( n13647 & n14217 ) | ( ~n14218 & n14217 ) ;
  assign n14220 = ( n713 & n14214 ) | ( n713 & n14219 ) | ( n14214 & n14219 ) ;
  assign n14221 = n595 &  n14220 ;
  assign n14223 = ( n13671 & ~n13662 ) | ( n13671 & n13675 ) | ( ~n13662 & n13675 ) ;
  assign n14222 = n13675 | n13784 ;
  assign n14225 = ( n13675 & ~n14223 ) | ( n13675 & n14222 ) | ( ~n14223 & n14222 ) ;
  assign n14224 = ( n14222 & ~n13671 ) | ( n14222 & n14223 ) | ( ~n13671 & n14223 ) ;
  assign n14226 = ( n13662 & ~n14225 ) | ( n13662 & n14224 ) | ( ~n14225 & n14224 ) ;
  assign n14227 = n713 | n14199 ;
  assign n14228 = n14213 | n14227 ;
  assign n14229 = n14219 &  n14228 ;
  assign n14230 = n14207 &  n14210 ;
  assign n14231 = ( n837 & ~n14230 ) | ( n837 & n14204 ) | ( ~n14230 & n14204 ) ;
  assign n14232 = n713 &  n14231 ;
  assign n14233 = n595 | n14232 ;
  assign n14234 = n14229 | n14233 ;
  assign n14235 = ~n14226 & n14234 ;
  assign n14236 = n14221 | n14235 ;
  assign n14237 = ~n13677 & n13784 ;
  assign n14238 = ( n13664 & ~n14237 ) | ( n13664 & n13784 ) | ( ~n14237 & n13784 ) ;
  assign n14239 = ( n13664 & ~n14238 ) | ( n13664 & n13669 ) | ( ~n14238 & n13669 ) ;
  assign n14240 = ( n13669 & ~n13664 ) | ( n13669 & n14238 ) | ( ~n13664 & n14238 ) ;
  assign n14241 = ( n14239 & ~n13669 ) | ( n14239 & n14240 ) | ( ~n13669 & n14240 ) ;
  assign n14242 = ( n492 & n14236 ) | ( n492 & n14241 ) | ( n14236 & n14241 ) ;
  assign n14243 = n396 &  n14242 ;
  assign n14245 = ( n13693 & ~n13684 ) | ( n13693 & n13697 ) | ( ~n13684 & n13697 ) ;
  assign n14244 = n13697 | n13784 ;
  assign n14247 = ( n13697 & ~n14245 ) | ( n13697 & n14244 ) | ( ~n14245 & n14244 ) ;
  assign n14246 = ( n14244 & ~n13693 ) | ( n14244 & n14245 ) | ( ~n13693 & n14245 ) ;
  assign n14248 = ( n13684 & ~n14247 ) | ( n13684 & n14246 ) | ( ~n14247 & n14246 ) ;
  assign n14249 = n492 | n14221 ;
  assign n14250 = n14235 | n14249 ;
  assign n14251 = n14241 &  n14250 ;
  assign n14252 = n14229 | n14232 ;
  assign n14253 = ( n595 & ~n14226 ) | ( n595 & n14252 ) | ( ~n14226 & n14252 ) ;
  assign n14254 = n492 &  n14253 ;
  assign n14255 = n396 | n14254 ;
  assign n14256 = n14251 | n14255 ;
  assign n14257 = ~n14248 & n14256 ;
  assign n14258 = n14243 | n14257 ;
  assign n14264 = ( n315 & ~n14263 ) | ( n315 & n14258 ) | ( ~n14263 & n14258 ) ;
  assign n14265 = n240 &  n14264 ;
  assign n14266 = n13719 | n13784 ;
  assign n14267 = ( n13706 & n13715 ) | ( n13706 & n13719 ) | ( n13715 & n13719 ) ;
  assign n14268 = ( n14266 & ~n13715 ) | ( n14266 & n14267 ) | ( ~n13715 & n14267 ) ;
  assign n14269 = ( n13719 & ~n14267 ) | ( n13719 & n14266 ) | ( ~n14267 & n14266 ) ;
  assign n14270 = ( n13706 & ~n14268 ) | ( n13706 & n14269 ) | ( ~n14268 & n14269 ) ;
  assign n14271 = n315 | n14243 ;
  assign n14272 = n14257 | n14271 ;
  assign n14273 = ~n14263 & n14272 ;
  assign n14274 = n14251 | n14254 ;
  assign n14275 = ( n396 & ~n14248 ) | ( n396 & n14274 ) | ( ~n14248 & n14274 ) ;
  assign n14276 = n315 &  n14275 ;
  assign n14277 = n240 | n14276 ;
  assign n14278 = n14273 | n14277 ;
  assign n14279 = n14270 &  n14278 ;
  assign n14280 = n14265 | n14279 ;
  assign n14281 = ~n13721 & n13784 ;
  assign n14282 = ( n13708 & ~n14281 ) | ( n13708 & n13784 ) | ( ~n14281 & n13784 ) ;
  assign n14283 = ( n13708 & ~n14282 ) | ( n13708 & n13713 ) | ( ~n14282 & n13713 ) ;
  assign n14284 = ( n13713 & ~n13708 ) | ( n13713 & n14282 ) | ( ~n13708 & n14282 ) ;
  assign n14285 = ( n14283 & ~n13713 ) | ( n14283 & n14284 ) | ( ~n13713 & n14284 ) ;
  assign n14286 = ( n181 & n14280 ) | ( n181 & n14285 ) | ( n14280 & n14285 ) ;
  assign n14287 = ~n145 & n14286 ;
  assign n14288 = n13741 | n13784 ;
  assign n14289 = ( n13728 & n13737 ) | ( n13728 & n13741 ) | ( n13737 & n13741 ) ;
  assign n14290 = ( n14288 & ~n13737 ) | ( n14288 & n14289 ) | ( ~n13737 & n14289 ) ;
  assign n14291 = ( n13741 & ~n14289 ) | ( n13741 & n14288 ) | ( ~n14289 & n14288 ) ;
  assign n14292 = ( n13728 & ~n14290 ) | ( n13728 & n14291 ) | ( ~n14290 & n14291 ) ;
  assign n14293 = n181 | n14265 ;
  assign n14294 = n14279 | n14293 ;
  assign n14295 = n14285 &  n14294 ;
  assign n14296 = n14273 | n14276 ;
  assign n14297 = ( n240 & n14270 ) | ( n240 & n14296 ) | ( n14270 & n14296 ) ;
  assign n14298 = n181 &  n14297 ;
  assign n14299 = ( n145 & ~n14298 ) | ( n145 & 1'b0 ) | ( ~n14298 & 1'b0 ) ;
  assign n14300 = ~n14295 & n14299 ;
  assign n14301 = n14292 | n14300 ;
  assign n14302 = ~n14287 & n14301 ;
  assign n14303 = n13730 | n13784 ;
  assign n14304 = ( n13735 & ~n13730 ) | ( n13735 & n13743 ) | ( ~n13730 & n13743 ) ;
  assign n14306 = ( n13730 & n14303 ) | ( n13730 & n14304 ) | ( n14303 & n14304 ) ;
  assign n14305 = ( n13743 & ~n14304 ) | ( n13743 & n14303 ) | ( ~n14304 & n14303 ) ;
  assign n14307 = ( n13735 & ~n14306 ) | ( n13735 & n14305 ) | ( ~n14306 & n14305 ) ;
  assign n14308 = ( n150 & ~n14302 ) | ( n150 & n14307 ) | ( ~n14302 & n14307 ) ;
  assign n14309 = ~n13750 & n13766 ;
  assign n14310 = ( n13769 & n13784 ) | ( n13769 & n14309 ) | ( n13784 & n14309 ) ;
  assign n14311 = ~n13769 & n14310 ;
  assign n14312 = ( n13766 & ~n13769 ) | ( n13766 & 1'b0 ) | ( ~n13769 & 1'b0 ) ;
  assign n14313 = ~n13784 & n14312 ;
  assign n14314 = ( n13750 & ~n14312 ) | ( n13750 & n14313 ) | ( ~n14312 & n14313 ) ;
  assign n14315 = n14311 | n14314 ;
  assign n14316 = ( n13751 & ~n13758 ) | ( n13751 & 1'b0 ) | ( ~n13758 & 1'b0 ) ;
  assign n14317 = ~n13784 & n14316 ;
  assign n14318 = ( n13772 & ~n14317 ) | ( n13772 & n14316 ) | ( ~n14317 & n14316 ) ;
  assign n14319 = ( n14315 & ~n14318 ) | ( n14315 & 1'b0 ) | ( ~n14318 & 1'b0 ) ;
  assign n14320 = ~n14308 & n14319 ;
  assign n14321 = ( n133 & ~n14320 ) | ( n133 & n14319 ) | ( ~n14320 & n14319 ) ;
  assign n14322 = n150 | n14287 ;
  assign n14323 = ( n14301 & ~n14322 ) | ( n14301 & 1'b0 ) | ( ~n14322 & 1'b0 ) ;
  assign n14328 = n14307 &  n14323 ;
  assign n14324 = n14295 | n14298 ;
  assign n14325 = ( n145 & ~n14324 ) | ( n145 & n14292 ) | ( ~n14324 & n14292 ) ;
  assign n14326 = ( n150 & ~n14325 ) | ( n150 & 1'b0 ) | ( ~n14325 & 1'b0 ) ;
  assign n14327 = n14315 | n14326 ;
  assign n14329 = ( n14307 & ~n14328 ) | ( n14307 & n14327 ) | ( ~n14328 & n14327 ) ;
  assign n14331 = ( n133 & ~n13758 ) | ( n133 & n13751 ) | ( ~n13758 & n13751 ) ;
  assign n14330 = ( n13758 & ~n13751 ) | ( n13758 & n13784 ) | ( ~n13751 & n13784 ) ;
  assign n14332 = ~n13758 & n14330 ;
  assign n14333 = ( n13758 & n14331 ) | ( n13758 & n14332 ) | ( n14331 & n14332 ) ;
  assign n14334 = n13754 | n13781 ;
  assign n14335 = ( n13757 & n13776 ) | ( n13757 & n14334 ) | ( n13776 & n14334 ) ;
  assign n14336 = ( n13757 & ~n14335 ) | ( n13757 & 1'b0 ) | ( ~n14335 & 1'b0 ) ;
  assign n14337 = ( n13764 & ~n14336 ) | ( n13764 & n13772 ) | ( ~n14336 & n13772 ) ;
  assign n14338 = ( n13764 & ~n14337 ) | ( n13764 & 1'b0 ) | ( ~n14337 & 1'b0 ) ;
  assign n14339 = n14333 | n14338 ;
  assign n14340 = ( n14329 & ~n14339 ) | ( n14329 & 1'b0 ) | ( ~n14339 & 1'b0 ) ;
  assign n14341 = ~n14321 | ~n14340 ;
  assign n14736 = n14169 &  n14341 ;
  assign n14737 = ( n14156 & ~n14341 ) | ( n14156 & n14736 ) | ( ~n14341 & n14736 ) ;
  assign n14738 = ( n14156 & ~n14737 ) | ( n14156 & n14161 ) | ( ~n14737 & n14161 ) ;
  assign n14739 = ( n14161 & ~n14156 ) | ( n14161 & n14737 ) | ( ~n14156 & n14737 ) ;
  assign n14740 = ( n14738 & ~n14161 ) | ( n14738 & n14739 ) | ( ~n14161 & n14739 ) ;
  assign n14722 = ( n14163 & ~n14154 ) | ( n14163 & n14167 ) | ( ~n14154 & n14167 ) ;
  assign n14721 = ( n14167 & ~n14341 ) | ( n14167 & 1'b0 ) | ( ~n14341 & 1'b0 ) ;
  assign n14724 = ( n14167 & ~n14722 ) | ( n14167 & n14721 ) | ( ~n14722 & n14721 ) ;
  assign n14723 = ( n14721 & ~n14163 ) | ( n14721 & n14722 ) | ( ~n14163 & n14722 ) ;
  assign n14725 = ( n14154 & ~n14724 ) | ( n14154 & n14723 ) | ( ~n14724 & n14723 ) ;
  assign n14714 = n14147 &  n14341 ;
  assign n14715 = ( n14134 & n14139 ) | ( n14134 & n14341 ) | ( n14139 & n14341 ) ;
  assign n14717 = ( n14714 & ~n14134 ) | ( n14714 & n14715 ) | ( ~n14134 & n14715 ) ;
  assign n14716 = ( n14341 & ~n14715 ) | ( n14341 & n14714 ) | ( ~n14715 & n14714 ) ;
  assign n14718 = ( n14139 & ~n14717 ) | ( n14139 & n14716 ) | ( ~n14717 & n14716 ) ;
  assign n14699 = n14145 | n14341 ;
  assign n14700 = ( n14132 & ~n14145 ) | ( n14132 & n14141 ) | ( ~n14145 & n14141 ) ;
  assign n14702 = ( n14145 & n14699 ) | ( n14145 & n14700 ) | ( n14699 & n14700 ) ;
  assign n14701 = ( n14141 & ~n14700 ) | ( n14141 & n14699 ) | ( ~n14700 & n14699 ) ;
  assign n14703 = ( n14132 & ~n14702 ) | ( n14132 & n14701 ) | ( ~n14702 & n14701 ) ;
  assign n14693 = ( n14112 & ~n14117 ) | ( n14112 & n14125 ) | ( ~n14117 & n14125 ) ;
  assign n14692 = n14112 | n14341 ;
  assign n14695 = ( n14112 & ~n14693 ) | ( n14112 & n14692 ) | ( ~n14693 & n14692 ) ;
  assign n14694 = ( n14692 & ~n14125 ) | ( n14692 & n14693 ) | ( ~n14125 & n14693 ) ;
  assign n14696 = ( n14117 & ~n14695 ) | ( n14117 & n14694 ) | ( ~n14695 & n14694 ) ;
  assign n14677 = n14123 | n14341 ;
  assign n14678 = ( n14110 & n14119 ) | ( n14110 & n14123 ) | ( n14119 & n14123 ) ;
  assign n14679 = ( n14677 & ~n14119 ) | ( n14677 & n14678 ) | ( ~n14119 & n14678 ) ;
  assign n14680 = ( n14123 & ~n14678 ) | ( n14123 & n14677 ) | ( ~n14678 & n14677 ) ;
  assign n14681 = ( n14110 & ~n14679 ) | ( n14110 & n14680 ) | ( ~n14679 & n14680 ) ;
  assign n14671 = ( n14090 & ~n14095 ) | ( n14090 & n14103 ) | ( ~n14095 & n14103 ) ;
  assign n14670 = n14090 | n14341 ;
  assign n14673 = ( n14090 & ~n14671 ) | ( n14090 & n14670 ) | ( ~n14671 & n14670 ) ;
  assign n14672 = ( n14670 & ~n14103 ) | ( n14670 & n14671 ) | ( ~n14103 & n14671 ) ;
  assign n14674 = ( n14095 & ~n14673 ) | ( n14095 & n14672 ) | ( ~n14673 & n14672 ) ;
  assign n14656 = ( n14097 & ~n14088 ) | ( n14097 & n14101 ) | ( ~n14088 & n14101 ) ;
  assign n14655 = n14101 | n14341 ;
  assign n14658 = ( n14101 & ~n14656 ) | ( n14101 & n14655 ) | ( ~n14656 & n14655 ) ;
  assign n14657 = ( n14655 & ~n14097 ) | ( n14655 & n14656 ) | ( ~n14097 & n14656 ) ;
  assign n14659 = ( n14088 & ~n14658 ) | ( n14088 & n14657 ) | ( ~n14658 & n14657 ) ;
  assign n14648 = n14068 | n14341 ;
  assign n14649 = ( n14068 & n14073 ) | ( n14068 & n14081 ) | ( n14073 & n14081 ) ;
  assign n14650 = ( n14648 & ~n14081 ) | ( n14648 & n14649 ) | ( ~n14081 & n14649 ) ;
  assign n14651 = ( n14068 & ~n14649 ) | ( n14068 & n14648 ) | ( ~n14649 & n14648 ) ;
  assign n14652 = ( n14073 & ~n14650 ) | ( n14073 & n14651 ) | ( ~n14650 & n14651 ) ;
  assign n14633 = n14079 | n14341 ;
  assign n14634 = ( n14066 & n14075 ) | ( n14066 & n14079 ) | ( n14075 & n14079 ) ;
  assign n14635 = ( n14633 & ~n14075 ) | ( n14633 & n14634 ) | ( ~n14075 & n14634 ) ;
  assign n14636 = ( n14079 & ~n14634 ) | ( n14079 & n14633 ) | ( ~n14634 & n14633 ) ;
  assign n14637 = ( n14066 & ~n14635 ) | ( n14066 & n14636 ) | ( ~n14635 & n14636 ) ;
  assign n14626 = n14046 | n14341 ;
  assign n14627 = ( n14046 & n14051 ) | ( n14046 & n14059 ) | ( n14051 & n14059 ) ;
  assign n14628 = ( n14626 & ~n14059 ) | ( n14626 & n14627 ) | ( ~n14059 & n14627 ) ;
  assign n14629 = ( n14046 & ~n14627 ) | ( n14046 & n14626 ) | ( ~n14627 & n14626 ) ;
  assign n14630 = ( n14051 & ~n14628 ) | ( n14051 & n14629 ) | ( ~n14628 & n14629 ) ;
  assign n14611 = n14057 | n14341 ;
  assign n14612 = ( n14044 & n14053 ) | ( n14044 & n14057 ) | ( n14053 & n14057 ) ;
  assign n14613 = ( n14611 & ~n14053 ) | ( n14611 & n14612 ) | ( ~n14053 & n14612 ) ;
  assign n14614 = ( n14057 & ~n14612 ) | ( n14057 & n14611 ) | ( ~n14612 & n14611 ) ;
  assign n14615 = ( n14044 & ~n14613 ) | ( n14044 & n14614 ) | ( ~n14613 & n14614 ) ;
  assign n14605 = ( n14024 & ~n14029 ) | ( n14024 & n14037 ) | ( ~n14029 & n14037 ) ;
  assign n14604 = n14024 | n14341 ;
  assign n14607 = ( n14024 & ~n14605 ) | ( n14024 & n14604 ) | ( ~n14605 & n14604 ) ;
  assign n14606 = ( n14604 & ~n14037 ) | ( n14604 & n14605 ) | ( ~n14037 & n14605 ) ;
  assign n14608 = ( n14029 & ~n14607 ) | ( n14029 & n14606 ) | ( ~n14607 & n14606 ) ;
  assign n14590 = ( n14031 & ~n14022 ) | ( n14031 & n14035 ) | ( ~n14022 & n14035 ) ;
  assign n14589 = n14035 | n14341 ;
  assign n14592 = ( n14035 & ~n14590 ) | ( n14035 & n14589 ) | ( ~n14590 & n14589 ) ;
  assign n14591 = ( n14589 & ~n14031 ) | ( n14589 & n14590 ) | ( ~n14031 & n14590 ) ;
  assign n14593 = ( n14022 & ~n14592 ) | ( n14022 & n14591 ) | ( ~n14592 & n14591 ) ;
  assign n14582 = n14002 | n14341 ;
  assign n14583 = ( n14002 & n14007 ) | ( n14002 & n14015 ) | ( n14007 & n14015 ) ;
  assign n14584 = ( n14582 & ~n14015 ) | ( n14582 & n14583 ) | ( ~n14015 & n14583 ) ;
  assign n14585 = ( n14002 & ~n14583 ) | ( n14002 & n14582 ) | ( ~n14583 & n14582 ) ;
  assign n14586 = ( n14007 & ~n14584 ) | ( n14007 & n14585 ) | ( ~n14584 & n14585 ) ;
  assign n14568 = ( n14009 & ~n14000 ) | ( n14009 & n14013 ) | ( ~n14000 & n14013 ) ;
  assign n14567 = n14013 | n14341 ;
  assign n14570 = ( n14013 & ~n14568 ) | ( n14013 & n14567 ) | ( ~n14568 & n14567 ) ;
  assign n14569 = ( n14567 & ~n14009 ) | ( n14567 & n14568 ) | ( ~n14009 & n14568 ) ;
  assign n14571 = ( n14000 & ~n14570 ) | ( n14000 & n14569 ) | ( ~n14570 & n14569 ) ;
  assign n14560 = n13980 | n14341 ;
  assign n14561 = ( n13980 & ~n13993 ) | ( n13980 & n13985 ) | ( ~n13993 & n13985 ) ;
  assign n14562 = ( n13993 & n14560 ) | ( n13993 & n14561 ) | ( n14560 & n14561 ) ;
  assign n14563 = ( n13980 & ~n14561 ) | ( n13980 & n14560 ) | ( ~n14561 & n14560 ) ;
  assign n14564 = ( n13985 & ~n14562 ) | ( n13985 & n14563 ) | ( ~n14562 & n14563 ) ;
  assign n14545 = n13991 | n14341 ;
  assign n14546 = ( n13978 & ~n13991 ) | ( n13978 & n13987 ) | ( ~n13991 & n13987 ) ;
  assign n14548 = ( n13991 & n14545 ) | ( n13991 & n14546 ) | ( n14545 & n14546 ) ;
  assign n14547 = ( n13987 & ~n14546 ) | ( n13987 & n14545 ) | ( ~n14546 & n14545 ) ;
  assign n14549 = ( n13978 & ~n14548 ) | ( n13978 & n14547 ) | ( ~n14548 & n14547 ) ;
  assign n14538 = ( n13958 & ~n14341 ) | ( n13958 & 1'b0 ) | ( ~n14341 & 1'b0 ) ;
  assign n14539 = ( n13958 & n13963 ) | ( n13958 & n13971 ) | ( n13963 & n13971 ) ;
  assign n14540 = ( n14538 & ~n13971 ) | ( n14538 & n14539 ) | ( ~n13971 & n14539 ) ;
  assign n14541 = ( n13958 & ~n14539 ) | ( n13958 & n14538 ) | ( ~n14539 & n14538 ) ;
  assign n14542 = ( n13963 & ~n14540 ) | ( n13963 & n14541 ) | ( ~n14540 & n14541 ) ;
  assign n14523 = n13969 | n14341 ;
  assign n14524 = ( n13956 & ~n13965 ) | ( n13956 & n13969 ) | ( ~n13965 & n13969 ) ;
  assign n14525 = ( n13965 & n14523 ) | ( n13965 & n14524 ) | ( n14523 & n14524 ) ;
  assign n14526 = ( n13969 & ~n14524 ) | ( n13969 & n14523 ) | ( ~n14524 & n14523 ) ;
  assign n14527 = ( n13956 & ~n14525 ) | ( n13956 & n14526 ) | ( ~n14525 & n14526 ) ;
  assign n14516 = ( n13936 & ~n14341 ) | ( n13936 & 1'b0 ) | ( ~n14341 & 1'b0 ) ;
  assign n14517 = ( n13936 & n13941 ) | ( n13936 & n13949 ) | ( n13941 & n13949 ) ;
  assign n14518 = ( n14516 & ~n13949 ) | ( n14516 & n14517 ) | ( ~n13949 & n14517 ) ;
  assign n14519 = ( n13936 & ~n14517 ) | ( n13936 & n14516 ) | ( ~n14517 & n14516 ) ;
  assign n14520 = ( n13941 & ~n14518 ) | ( n13941 & n14519 ) | ( ~n14518 & n14519 ) ;
  assign n14502 = ( n13943 & ~n13934 ) | ( n13943 & n13947 ) | ( ~n13934 & n13947 ) ;
  assign n14501 = ( n13947 & ~n14341 ) | ( n13947 & 1'b0 ) | ( ~n14341 & 1'b0 ) ;
  assign n14504 = ( n13947 & ~n14502 ) | ( n13947 & n14501 ) | ( ~n14502 & n14501 ) ;
  assign n14503 = ( n14501 & ~n13943 ) | ( n14501 & n14502 ) | ( ~n13943 & n14502 ) ;
  assign n14505 = ( n13934 & ~n14504 ) | ( n13934 & n14503 ) | ( ~n14504 & n14503 ) ;
  assign n14494 = n13914 | n14341 ;
  assign n14495 = ( n13919 & ~n13914 ) | ( n13919 & n13927 ) | ( ~n13914 & n13927 ) ;
  assign n14497 = ( n13914 & n14494 ) | ( n13914 & n14495 ) | ( n14494 & n14495 ) ;
  assign n14496 = ( n13927 & ~n14495 ) | ( n13927 & n14494 ) | ( ~n14495 & n14494 ) ;
  assign n14498 = ( n13919 & ~n14497 ) | ( n13919 & n14496 ) | ( ~n14497 & n14496 ) ;
  assign n14479 = n13925 | n14341 ;
  assign n14480 = ( n13912 & ~n13921 ) | ( n13912 & n13925 ) | ( ~n13921 & n13925 ) ;
  assign n14481 = ( n13921 & n14479 ) | ( n13921 & n14480 ) | ( n14479 & n14480 ) ;
  assign n14482 = ( n13925 & ~n14480 ) | ( n13925 & n14479 ) | ( ~n14480 & n14479 ) ;
  assign n14483 = ( n13912 & ~n14481 ) | ( n13912 & n14482 ) | ( ~n14481 & n14482 ) ;
  assign n14472 = n13892 | n14341 ;
  assign n14473 = ( n13897 & ~n13892 ) | ( n13897 & n13905 ) | ( ~n13892 & n13905 ) ;
  assign n14475 = ( n13892 & n14472 ) | ( n13892 & n14473 ) | ( n14472 & n14473 ) ;
  assign n14474 = ( n13905 & ~n14473 ) | ( n13905 & n14472 ) | ( ~n14473 & n14472 ) ;
  assign n14476 = ( n13897 & ~n14475 ) | ( n13897 & n14474 ) | ( ~n14475 & n14474 ) ;
  assign n14457 = n13903 | n14341 ;
  assign n14458 = ( n13890 & ~n13899 ) | ( n13890 & n13903 ) | ( ~n13899 & n13903 ) ;
  assign n14459 = ( n13899 & n14457 ) | ( n13899 & n14458 ) | ( n14457 & n14458 ) ;
  assign n14460 = ( n13903 & ~n14458 ) | ( n13903 & n14457 ) | ( ~n14458 & n14457 ) ;
  assign n14461 = ( n13890 & ~n14459 ) | ( n13890 & n14460 ) | ( ~n14459 & n14460 ) ;
  assign n14450 = n13883 &  n14341 ;
  assign n14451 = ( n13875 & ~n13870 ) | ( n13875 & n14341 ) | ( ~n13870 & n14341 ) ;
  assign n14453 = ( n14450 & n13870 ) | ( n14450 & n14451 ) | ( n13870 & n14451 ) ;
  assign n14452 = ( n14341 & ~n14451 ) | ( n14341 & n14450 ) | ( ~n14451 & n14450 ) ;
  assign n14454 = ( n13875 & ~n14453 ) | ( n13875 & n14452 ) | ( ~n14453 & n14452 ) ;
  assign n14435 = n13881 | n14341 ;
  assign n14436 = ( n13868 & ~n13881 ) | ( n13868 & n13877 ) | ( ~n13881 & n13877 ) ;
  assign n14438 = ( n13881 & n14435 ) | ( n13881 & n14436 ) | ( n14435 & n14436 ) ;
  assign n14437 = ( n13877 & ~n14436 ) | ( n13877 & n14435 ) | ( ~n14436 & n14435 ) ;
  assign n14439 = ( n13868 & ~n14438 ) | ( n13868 & n14437 ) | ( ~n14438 & n14437 ) ;
  assign n14428 = n13848 | n14341 ;
  assign n14429 = ( n13848 & ~n13861 ) | ( n13848 & n13853 ) | ( ~n13861 & n13853 ) ;
  assign n14430 = ( n13861 & n14428 ) | ( n13861 & n14429 ) | ( n14428 & n14429 ) ;
  assign n14431 = ( n13848 & ~n14429 ) | ( n13848 & n14428 ) | ( ~n14429 & n14428 ) ;
  assign n14432 = ( n13853 & ~n14430 ) | ( n13853 & n14431 ) | ( ~n14430 & n14431 ) ;
  assign n14413 = n13859 | n14341 ;
  assign n14414 = ( n13846 & ~n13855 ) | ( n13846 & n13859 ) | ( ~n13855 & n13859 ) ;
  assign n14415 = ( n13855 & n14413 ) | ( n13855 & n14414 ) | ( n14413 & n14414 ) ;
  assign n14416 = ( n13859 & ~n14414 ) | ( n13859 & n14413 ) | ( ~n14414 & n14413 ) ;
  assign n14417 = ( n13846 & ~n14415 ) | ( n13846 & n14416 ) | ( ~n14415 & n14416 ) ;
  assign n14406 = n13826 | n14341 ;
  assign n14407 = ( n13831 & ~n13826 ) | ( n13831 & n13839 ) | ( ~n13826 & n13839 ) ;
  assign n14409 = ( n13826 & n14406 ) | ( n13826 & n14407 ) | ( n14406 & n14407 ) ;
  assign n14408 = ( n13839 & ~n14407 ) | ( n13839 & n14406 ) | ( ~n14407 & n14406 ) ;
  assign n14410 = ( n13831 & ~n14409 ) | ( n13831 & n14408 ) | ( ~n14409 & n14408 ) ;
  assign n14391 = n13837 | n14341 ;
  assign n14392 = ( n13824 & ~n13833 ) | ( n13824 & n13837 ) | ( ~n13833 & n13837 ) ;
  assign n14393 = ( n13833 & n14391 ) | ( n13833 & n14392 ) | ( n14391 & n14392 ) ;
  assign n14394 = ( n13837 & ~n14392 ) | ( n13837 & n14391 ) | ( ~n14392 & n14391 ) ;
  assign n14395 = ( n13824 & ~n14393 ) | ( n13824 & n14394 ) | ( ~n14393 & n14394 ) ;
  assign n14384 = ( n13800 & ~n13802 ) | ( n13800 & 1'b0 ) | ( ~n13802 & 1'b0 ) ;
  assign n14385 = ( n13802 & ~n14384 ) | ( n13802 & n13812 ) | ( ~n14384 & n13812 ) ;
  assign n14387 = ( n14341 & n14384 ) | ( n14341 & n14385 ) | ( n14384 & n14385 ) ;
  assign n14386 = ( n13802 & ~n14385 ) | ( n13802 & n14341 ) | ( ~n14385 & n14341 ) ;
  assign n14388 = ( n13812 & ~n14387 ) | ( n13812 & n14386 ) | ( ~n14387 & n14386 ) ;
  assign n14368 = ~x30 & n13784 ;
  assign n14369 = ( x31 & ~n14368 ) | ( x31 & 1'b0 ) | ( ~n14368 & 1'b0 ) ;
  assign n14370 = n13803 | n14369 ;
  assign n14365 = ( n13784 & ~x30 ) | ( n13784 & n13795 ) | ( ~x30 & n13795 ) ;
  assign n14366 = x30 &  n14365 ;
  assign n14367 = ( n13790 & ~n14366 ) | ( n13790 & n13795 ) | ( ~n14366 & n13795 ) ;
  assign n14371 = ( n14341 & ~n14370 ) | ( n14341 & n14367 ) | ( ~n14370 & n14367 ) ;
  assign n14373 = ( n14341 & ~n14371 ) | ( n14341 & 1'b0 ) | ( ~n14371 & 1'b0 ) ;
  assign n14372 = ~n14367 & n14371 ;
  assign n14374 = ( n14370 & ~n14373 ) | ( n14370 & n14372 ) | ( ~n14373 & n14372 ) ;
  assign n14354 = ( n13784 & ~n14338 ) | ( n13784 & 1'b0 ) | ( ~n14338 & 1'b0 ) ;
  assign n14355 = ( n14329 & ~n14354 ) | ( n14329 & n14333 ) | ( ~n14354 & n14333 ) ;
  assign n14356 = ( n14329 & ~n14355 ) | ( n14329 & 1'b0 ) | ( ~n14355 & 1'b0 ) ;
  assign n14357 = n14321 &  n14356 ;
  assign n14353 = ~n13787 & n14341 ;
  assign n14358 = ( n14353 & ~n14357 ) | ( n14353 & 1'b0 ) | ( ~n14357 & 1'b0 ) ;
  assign n14359 = ( x30 & n14357 ) | ( x30 & n14358 ) | ( n14357 & n14358 ) ;
  assign n14360 = x30 | n14357 ;
  assign n14361 = n14353 | n14360 ;
  assign n14362 = ~n14359 & n14361 ;
  assign n14344 = ( x28 & ~n14341 ) | ( x28 & x29 ) | ( ~n14341 & x29 ) ;
  assign n14350 = ( x28 & ~x29 ) | ( x28 & 1'b0 ) | ( ~x29 & 1'b0 ) ;
  assign n13785 = x26 | x27 ;
  assign n14345 = ~x28 & n13785 ;
  assign n14346 = ( x28 & ~n13782 ) | ( x28 & n14345 ) | ( ~n13782 & n14345 ) ;
  assign n14347 = ( n13764 & ~n14346 ) | ( n13764 & n13772 ) | ( ~n14346 & n13772 ) ;
  assign n14348 = ( n13764 & ~n14347 ) | ( n13764 & 1'b0 ) | ( ~n14347 & 1'b0 ) ;
  assign n14349 = ( n14341 & ~x29 ) | ( n14341 & n14348 ) | ( ~x29 & n14348 ) ;
  assign n14351 = ( n14344 & ~n14350 ) | ( n14344 & n14349 ) | ( ~n14350 & n14349 ) ;
  assign n13786 = x28 | n13785 ;
  assign n14342 = x28 &  n14341 ;
  assign n14343 = ( n13784 & ~n13786 ) | ( n13784 & n14342 ) | ( ~n13786 & n14342 ) ;
  assign n14375 = n13242 | n14343 ;
  assign n14376 = ( n14351 & ~n14375 ) | ( n14351 & 1'b0 ) | ( ~n14375 & 1'b0 ) ;
  assign n14377 = n14362 | n14376 ;
  assign n14378 = n14343 &  n14351 ;
  assign n14379 = ( n13242 & ~n14351 ) | ( n13242 & n14378 ) | ( ~n14351 & n14378 ) ;
  assign n14380 = n12707 | n14379 ;
  assign n14381 = ( n14377 & ~n14380 ) | ( n14377 & 1'b0 ) | ( ~n14380 & 1'b0 ) ;
  assign n14382 = n14374 | n14381 ;
  assign n14352 = ~n14343 & n14351 ;
  assign n14363 = ( n14352 & ~n13242 ) | ( n14352 & n14362 ) | ( ~n13242 & n14362 ) ;
  assign n14364 = ( n12707 & ~n14363 ) | ( n12707 & 1'b0 ) | ( ~n14363 & 1'b0 ) ;
  assign n14396 = n12187 | n14364 ;
  assign n14397 = ( n14382 & ~n14396 ) | ( n14382 & 1'b0 ) | ( ~n14396 & 1'b0 ) ;
  assign n14398 = n14388 | n14397 ;
  assign n14399 = ( n14377 & ~n14379 ) | ( n14377 & 1'b0 ) | ( ~n14379 & 1'b0 ) ;
  assign n14400 = ( n14374 & ~n12707 ) | ( n14374 & n14399 ) | ( ~n12707 & n14399 ) ;
  assign n14401 = ( n12187 & ~n14400 ) | ( n12187 & 1'b0 ) | ( ~n14400 & 1'b0 ) ;
  assign n14402 = n11674 | n14401 ;
  assign n14403 = ( n14398 & ~n14402 ) | ( n14398 & 1'b0 ) | ( ~n14402 & 1'b0 ) ;
  assign n14404 = n14395 | n14403 ;
  assign n14383 = ~n14364 & n14382 ;
  assign n14389 = ( n14383 & ~n12187 ) | ( n14383 & n14388 ) | ( ~n12187 & n14388 ) ;
  assign n14390 = ( n11674 & ~n14389 ) | ( n11674 & 1'b0 ) | ( ~n14389 & 1'b0 ) ;
  assign n14418 = n11176 | n14390 ;
  assign n14419 = ( n14404 & ~n14418 ) | ( n14404 & 1'b0 ) | ( ~n14418 & 1'b0 ) ;
  assign n14420 = n14410 | n14419 ;
  assign n14421 = ( n14398 & ~n14401 ) | ( n14398 & 1'b0 ) | ( ~n14401 & 1'b0 ) ;
  assign n14422 = ( n14395 & ~n11674 ) | ( n14395 & n14421 ) | ( ~n11674 & n14421 ) ;
  assign n14423 = ( n11176 & ~n14422 ) | ( n11176 & 1'b0 ) | ( ~n14422 & 1'b0 ) ;
  assign n14424 = n10685 | n14423 ;
  assign n14425 = ( n14420 & ~n14424 ) | ( n14420 & 1'b0 ) | ( ~n14424 & 1'b0 ) ;
  assign n14426 = n14417 | n14425 ;
  assign n14405 = ~n14390 & n14404 ;
  assign n14411 = ( n14405 & ~n11176 ) | ( n14405 & n14410 ) | ( ~n11176 & n14410 ) ;
  assign n14412 = ( n10685 & ~n14411 ) | ( n10685 & 1'b0 ) | ( ~n14411 & 1'b0 ) ;
  assign n14440 = n10209 | n14412 ;
  assign n14441 = ( n14426 & ~n14440 ) | ( n14426 & 1'b0 ) | ( ~n14440 & 1'b0 ) ;
  assign n14442 = n14432 | n14441 ;
  assign n14443 = ( n14420 & ~n14423 ) | ( n14420 & 1'b0 ) | ( ~n14423 & 1'b0 ) ;
  assign n14444 = ( n14417 & ~n10685 ) | ( n14417 & n14443 ) | ( ~n10685 & n14443 ) ;
  assign n14445 = ( n10209 & ~n14444 ) | ( n10209 & 1'b0 ) | ( ~n14444 & 1'b0 ) ;
  assign n14446 = ( n9740 & ~n14445 ) | ( n9740 & 1'b0 ) | ( ~n14445 & 1'b0 ) ;
  assign n14447 = n14442 &  n14446 ;
  assign n14448 = n14439 | n14447 ;
  assign n14427 = ~n14412 & n14426 ;
  assign n14433 = ( n14427 & ~n10209 ) | ( n14427 & n14432 ) | ( ~n10209 & n14432 ) ;
  assign n14434 = n9740 | n14433 ;
  assign n14462 = ~n9286 & n14434 ;
  assign n14463 = n14448 &  n14462 ;
  assign n14464 = n14454 | n14463 ;
  assign n14465 = ( n14442 & ~n14445 ) | ( n14442 & 1'b0 ) | ( ~n14445 & 1'b0 ) ;
  assign n14466 = ( n9740 & n14439 ) | ( n9740 & n14465 ) | ( n14439 & n14465 ) ;
  assign n14467 = ( n9286 & ~n14466 ) | ( n9286 & 1'b0 ) | ( ~n14466 & 1'b0 ) ;
  assign n14468 = n8839 | n14467 ;
  assign n14469 = ( n14464 & ~n14468 ) | ( n14464 & 1'b0 ) | ( ~n14468 & 1'b0 ) ;
  assign n14470 = n14461 | n14469 ;
  assign n14449 = n14434 &  n14448 ;
  assign n14455 = ( n14449 & ~n9286 ) | ( n14449 & n14454 ) | ( ~n9286 & n14454 ) ;
  assign n14456 = ( n8839 & ~n14455 ) | ( n8839 & 1'b0 ) | ( ~n14455 & 1'b0 ) ;
  assign n14484 = n8407 | n14456 ;
  assign n14485 = ( n14470 & ~n14484 ) | ( n14470 & 1'b0 ) | ( ~n14484 & 1'b0 ) ;
  assign n14486 = n14476 | n14485 ;
  assign n14487 = ( n14464 & ~n14467 ) | ( n14464 & 1'b0 ) | ( ~n14467 & 1'b0 ) ;
  assign n14488 = ( n14461 & ~n8839 ) | ( n14461 & n14487 ) | ( ~n8839 & n14487 ) ;
  assign n14489 = ( n8407 & ~n14488 ) | ( n8407 & 1'b0 ) | ( ~n14488 & 1'b0 ) ;
  assign n14490 = n7982 | n14489 ;
  assign n14491 = ( n14486 & ~n14490 ) | ( n14486 & 1'b0 ) | ( ~n14490 & 1'b0 ) ;
  assign n14492 = n14483 | n14491 ;
  assign n14471 = ~n14456 & n14470 ;
  assign n14477 = ( n14471 & ~n8407 ) | ( n14471 & n14476 ) | ( ~n8407 & n14476 ) ;
  assign n14478 = ( n7982 & ~n14477 ) | ( n7982 & 1'b0 ) | ( ~n14477 & 1'b0 ) ;
  assign n14506 = ( n7572 & ~n14478 ) | ( n7572 & 1'b0 ) | ( ~n14478 & 1'b0 ) ;
  assign n14507 = n14492 &  n14506 ;
  assign n14508 = n14498 | n14507 ;
  assign n14509 = ( n14486 & ~n14489 ) | ( n14486 & 1'b0 ) | ( ~n14489 & 1'b0 ) ;
  assign n14510 = ( n14483 & ~n7982 ) | ( n14483 & n14509 ) | ( ~n7982 & n14509 ) ;
  assign n14511 = n7572 | n14510 ;
  assign n14512 = n7169 &  n14511 ;
  assign n14513 = n14508 &  n14512 ;
  assign n14514 = n14505 | n14513 ;
  assign n14493 = ~n14478 & n14492 ;
  assign n14499 = ( n7572 & n14493 ) | ( n7572 & n14498 ) | ( n14493 & n14498 ) ;
  assign n14500 = n7169 | n14499 ;
  assign n14528 = ~n6781 & n14500 ;
  assign n14529 = n14514 &  n14528 ;
  assign n14530 = n14520 | n14529 ;
  assign n14531 = n14508 &  n14511 ;
  assign n14532 = ( n7169 & n14505 ) | ( n7169 & n14531 ) | ( n14505 & n14531 ) ;
  assign n14533 = ( n6781 & ~n14532 ) | ( n6781 & 1'b0 ) | ( ~n14532 & 1'b0 ) ;
  assign n14534 = ( n6399 & ~n14533 ) | ( n6399 & 1'b0 ) | ( ~n14533 & 1'b0 ) ;
  assign n14535 = n14530 &  n14534 ;
  assign n14536 = n14527 | n14535 ;
  assign n14515 = n14500 &  n14514 ;
  assign n14521 = ( n14515 & ~n6781 ) | ( n14515 & n14520 ) | ( ~n6781 & n14520 ) ;
  assign n14522 = n6399 | n14521 ;
  assign n14550 = ~n6032 & n14522 ;
  assign n14551 = n14536 &  n14550 ;
  assign n14552 = n14542 | n14551 ;
  assign n14553 = ( n14530 & ~n14533 ) | ( n14530 & 1'b0 ) | ( ~n14533 & 1'b0 ) ;
  assign n14554 = ( n6399 & n14527 ) | ( n6399 & n14553 ) | ( n14527 & n14553 ) ;
  assign n14555 = ( n6032 & ~n14554 ) | ( n6032 & 1'b0 ) | ( ~n14554 & 1'b0 ) ;
  assign n14556 = ( n5672 & ~n14555 ) | ( n5672 & 1'b0 ) | ( ~n14555 & 1'b0 ) ;
  assign n14557 = n14552 &  n14556 ;
  assign n14558 = ( n14549 & ~n14557 ) | ( n14549 & 1'b0 ) | ( ~n14557 & 1'b0 ) ;
  assign n14537 = n14522 &  n14536 ;
  assign n14543 = ( n14537 & ~n6032 ) | ( n14537 & n14542 ) | ( ~n6032 & n14542 ) ;
  assign n14544 = n5672 | n14543 ;
  assign n14572 = ~n5327 & n14544 ;
  assign n14573 = ~n14558 & n14572 ;
  assign n14574 = ( n14564 & ~n14573 ) | ( n14564 & 1'b0 ) | ( ~n14573 & 1'b0 ) ;
  assign n14575 = ( n14552 & ~n14555 ) | ( n14552 & 1'b0 ) | ( ~n14555 & 1'b0 ) ;
  assign n14576 = ( n5672 & ~n14549 ) | ( n5672 & n14575 ) | ( ~n14549 & n14575 ) ;
  assign n14577 = ( n5327 & ~n14576 ) | ( n5327 & 1'b0 ) | ( ~n14576 & 1'b0 ) ;
  assign n14578 = n4990 | n14577 ;
  assign n14579 = n14574 | n14578 ;
  assign n14580 = n14571 &  n14579 ;
  assign n14559 = ( n14544 & ~n14558 ) | ( n14544 & 1'b0 ) | ( ~n14558 & 1'b0 ) ;
  assign n14565 = ( n5327 & ~n14559 ) | ( n5327 & n14564 ) | ( ~n14559 & n14564 ) ;
  assign n14566 = n4990 &  n14565 ;
  assign n14594 = n4668 | n14566 ;
  assign n14595 = n14580 | n14594 ;
  assign n14596 = n14586 &  n14595 ;
  assign n14597 = n14574 | n14577 ;
  assign n14598 = ( n4990 & n14571 ) | ( n4990 & n14597 ) | ( n14571 & n14597 ) ;
  assign n14599 = n4668 &  n14598 ;
  assign n14600 = n4353 | n14599 ;
  assign n14601 = n14596 | n14600 ;
  assign n14602 = n14593 &  n14601 ;
  assign n14581 = n14566 | n14580 ;
  assign n14587 = ( n4668 & n14581 ) | ( n4668 & n14586 ) | ( n14581 & n14586 ) ;
  assign n14588 = n4353 &  n14587 ;
  assign n14616 = n4053 | n14588 ;
  assign n14617 = n14602 | n14616 ;
  assign n14618 = ~n14608 & n14617 ;
  assign n14619 = n14596 | n14599 ;
  assign n14620 = ( n4353 & n14593 ) | ( n4353 & n14619 ) | ( n14593 & n14619 ) ;
  assign n14621 = n4053 &  n14620 ;
  assign n14622 = n3760 | n14621 ;
  assign n14623 = n14618 | n14622 ;
  assign n14624 = ~n14615 & n14623 ;
  assign n14603 = n14588 | n14602 ;
  assign n14609 = ( n4053 & ~n14608 ) | ( n4053 & n14603 ) | ( ~n14608 & n14603 ) ;
  assign n14610 = n3760 &  n14609 ;
  assign n14638 = n3482 | n14610 ;
  assign n14639 = n14624 | n14638 ;
  assign n14640 = n14630 &  n14639 ;
  assign n14641 = n14618 | n14621 ;
  assign n14642 = ( n3760 & ~n14615 ) | ( n3760 & n14641 ) | ( ~n14615 & n14641 ) ;
  assign n14643 = n3482 &  n14642 ;
  assign n14644 = n3211 | n14643 ;
  assign n14645 = n14640 | n14644 ;
  assign n14646 = ~n14637 & n14645 ;
  assign n14625 = n14610 | n14624 ;
  assign n14631 = ( n3482 & n14625 ) | ( n3482 & n14630 ) | ( n14625 & n14630 ) ;
  assign n14632 = n3211 &  n14631 ;
  assign n14660 = n2955 | n14632 ;
  assign n14661 = n14646 | n14660 ;
  assign n14662 = n14652 &  n14661 ;
  assign n14663 = n14640 | n14643 ;
  assign n14664 = ( n3211 & ~n14637 ) | ( n3211 & n14663 ) | ( ~n14637 & n14663 ) ;
  assign n14665 = n2955 &  n14664 ;
  assign n14666 = n2706 | n14665 ;
  assign n14667 = n14662 | n14666 ;
  assign n14668 = n14659 &  n14667 ;
  assign n14647 = n14632 | n14646 ;
  assign n14653 = ( n2955 & n14647 ) | ( n2955 & n14652 ) | ( n14647 & n14652 ) ;
  assign n14654 = n2706 &  n14653 ;
  assign n14682 = n2472 | n14654 ;
  assign n14683 = n14668 | n14682 ;
  assign n14684 = ~n14674 & n14683 ;
  assign n14685 = n14662 | n14665 ;
  assign n14686 = ( n2706 & n14659 ) | ( n2706 & n14685 ) | ( n14659 & n14685 ) ;
  assign n14687 = n2472 &  n14686 ;
  assign n14688 = n2245 | n14687 ;
  assign n14689 = n14684 | n14688 ;
  assign n14690 = ~n14681 & n14689 ;
  assign n14669 = n14654 | n14668 ;
  assign n14675 = ( n2472 & ~n14674 ) | ( n2472 & n14669 ) | ( ~n14674 & n14669 ) ;
  assign n14676 = n2245 &  n14675 ;
  assign n14704 = ( n2033 & ~n14676 ) | ( n2033 & 1'b0 ) | ( ~n14676 & 1'b0 ) ;
  assign n14705 = ~n14690 & n14704 ;
  assign n14706 = n14696 | n14705 ;
  assign n14707 = n14684 | n14687 ;
  assign n14708 = ( n2245 & ~n14681 ) | ( n2245 & n14707 ) | ( ~n14681 & n14707 ) ;
  assign n14709 = ~n2033 & n14708 ;
  assign n14710 = n1827 | n14709 ;
  assign n14711 = ( n14706 & ~n14710 ) | ( n14706 & 1'b0 ) | ( ~n14710 & 1'b0 ) ;
  assign n14712 = n14703 | n14711 ;
  assign n14691 = n14676 | n14690 ;
  assign n14697 = ( n2033 & ~n14691 ) | ( n2033 & n14696 ) | ( ~n14691 & n14696 ) ;
  assign n14698 = ( n1827 & ~n14697 ) | ( n1827 & 1'b0 ) | ( ~n14697 & 1'b0 ) ;
  assign n14726 = ( n1636 & ~n14698 ) | ( n1636 & 1'b0 ) | ( ~n14698 & 1'b0 ) ;
  assign n14727 = n14712 &  n14726 ;
  assign n14728 = n14718 | n14727 ;
  assign n14729 = ( n14706 & ~n14709 ) | ( n14706 & 1'b0 ) | ( ~n14709 & 1'b0 ) ;
  assign n14730 = ( n14703 & ~n1827 ) | ( n14703 & n14729 ) | ( ~n1827 & n14729 ) ;
  assign n14731 = n1636 | n14730 ;
  assign n14746 = n14728 &  n14731 ;
  assign n14747 = ( n1452 & ~n14725 ) | ( n1452 & n14746 ) | ( ~n14725 & n14746 ) ;
  assign n14748 = ( n1283 & ~n14747 ) | ( n1283 & 1'b0 ) | ( ~n14747 & 1'b0 ) ;
  assign n14867 = n14287 | n14341 ;
  assign n14868 = ( n14287 & ~n14300 ) | ( n14287 & n14292 ) | ( ~n14300 & n14292 ) ;
  assign n14869 = ( n14300 & n14867 ) | ( n14300 & n14868 ) | ( n14867 & n14868 ) ;
  assign n14870 = ( n14287 & ~n14868 ) | ( n14287 & n14867 ) | ( ~n14868 & n14867 ) ;
  assign n14871 = ( n14292 & ~n14869 ) | ( n14292 & n14870 ) | ( ~n14869 & n14870 ) ;
  assign n14823 = ~n14256 & n14341 ;
  assign n14824 = ( n14243 & ~n14823 ) | ( n14243 & n14341 ) | ( ~n14823 & n14341 ) ;
  assign n14825 = ( n14248 & ~n14243 ) | ( n14248 & n14824 ) | ( ~n14243 & n14824 ) ;
  assign n14826 = ( n14243 & ~n14824 ) | ( n14243 & n14248 ) | ( ~n14824 & n14248 ) ;
  assign n14827 = ( n14825 & ~n14248 ) | ( n14825 & n14826 ) | ( ~n14248 & n14826 ) ;
  assign n14802 = ( n14221 & ~n14226 ) | ( n14221 & n14341 ) | ( ~n14226 & n14341 ) ;
  assign n14801 = ~n14234 & n14341 ;
  assign n14803 = ( n14341 & ~n14802 ) | ( n14341 & n14801 ) | ( ~n14802 & n14801 ) ;
  assign n14804 = ( n14801 & ~n14221 ) | ( n14801 & n14802 ) | ( ~n14221 & n14802 ) ;
  assign n14805 = ( n14226 & ~n14803 ) | ( n14226 & n14804 ) | ( ~n14803 & n14804 ) ;
  assign n14757 = n14190 &  n14341 ;
  assign n14758 = ( n14182 & ~n14177 ) | ( n14182 & n14341 ) | ( ~n14177 & n14341 ) ;
  assign n14760 = ( n14177 & n14757 ) | ( n14177 & n14758 ) | ( n14757 & n14758 ) ;
  assign n14759 = ( n14341 & ~n14758 ) | ( n14341 & n14757 ) | ( ~n14758 & n14757 ) ;
  assign n14761 = ( n14182 & ~n14760 ) | ( n14182 & n14759 ) | ( ~n14760 & n14759 ) ;
  assign n14713 = ~n14698 & n14712 ;
  assign n14719 = ( n1636 & n14713 ) | ( n1636 & n14718 ) | ( n14713 & n14718 ) ;
  assign n14720 = n1452 | n14719 ;
  assign n14732 = n1452 &  n14731 ;
  assign n14733 = n14728 &  n14732 ;
  assign n14734 = ( n14725 & ~n14733 ) | ( n14725 & 1'b0 ) | ( ~n14733 & 1'b0 ) ;
  assign n14735 = ( n14720 & ~n14734 ) | ( n14720 & 1'b0 ) | ( ~n14734 & 1'b0 ) ;
  assign n14741 = ( n14735 & ~n1283 ) | ( n14735 & n14740 ) | ( ~n1283 & n14740 ) ;
  assign n14742 = n1122 | n14741 ;
  assign n14743 = ~n1283 & n14720 ;
  assign n14744 = ~n14734 & n14743 ;
  assign n14745 = n14740 | n14744 ;
  assign n14749 = ( n1122 & ~n14748 ) | ( n1122 & 1'b0 ) | ( ~n14748 & 1'b0 ) ;
  assign n14750 = n14745 &  n14749 ;
  assign n14751 = ( n14175 & ~n14188 ) | ( n14175 & n14184 ) | ( ~n14188 & n14184 ) ;
  assign n14753 = ( n14188 & n14341 ) | ( n14188 & n14751 ) | ( n14341 & n14751 ) ;
  assign n14752 = ( n14184 & ~n14751 ) | ( n14184 & n14341 ) | ( ~n14751 & n14341 ) ;
  assign n14754 = ( n14175 & ~n14753 ) | ( n14175 & n14752 ) | ( ~n14753 & n14752 ) ;
  assign n14755 = n14750 | n14754 ;
  assign n14756 = n14742 &  n14755 ;
  assign n14762 = ( n976 & ~n14761 ) | ( n976 & n14756 ) | ( ~n14761 & n14756 ) ;
  assign n14763 = ( n837 & ~n14762 ) | ( n837 & 1'b0 ) | ( ~n14762 & 1'b0 ) ;
  assign n14764 = ( n14210 & ~n14341 ) | ( n14210 & 1'b0 ) | ( ~n14341 & 1'b0 ) ;
  assign n14765 = ( n14197 & n14206 ) | ( n14197 & n14210 ) | ( n14206 & n14210 ) ;
  assign n14766 = ( n14764 & ~n14206 ) | ( n14764 & n14765 ) | ( ~n14206 & n14765 ) ;
  assign n14767 = ( n14210 & ~n14765 ) | ( n14210 & n14764 ) | ( ~n14765 & n14764 ) ;
  assign n14768 = ( n14197 & ~n14766 ) | ( n14197 & n14767 ) | ( ~n14766 & n14767 ) ;
  assign n14769 = n976 &  n14742 ;
  assign n14770 = n14755 &  n14769 ;
  assign n14771 = ( n14761 & ~n14770 ) | ( n14761 & 1'b0 ) | ( ~n14770 & 1'b0 ) ;
  assign n14772 = ( n14745 & ~n14748 ) | ( n14745 & 1'b0 ) | ( ~n14748 & 1'b0 ) ;
  assign n14773 = ( n1122 & n14754 ) | ( n1122 & n14772 ) | ( n14754 & n14772 ) ;
  assign n14774 = n976 | n14773 ;
  assign n14775 = ~n837 & n14774 ;
  assign n14776 = ~n14771 & n14775 ;
  assign n14777 = n14768 | n14776 ;
  assign n14778 = ~n14763 & n14777 ;
  assign n14779 = n14212 &  n14341 ;
  assign n14780 = ( n14199 & n14204 ) | ( n14199 & n14341 ) | ( n14204 & n14341 ) ;
  assign n14782 = ( n14779 & ~n14199 ) | ( n14779 & n14780 ) | ( ~n14199 & n14780 ) ;
  assign n14781 = ( n14341 & ~n14780 ) | ( n14341 & n14779 ) | ( ~n14780 & n14779 ) ;
  assign n14783 = ( n14204 & ~n14782 ) | ( n14204 & n14781 ) | ( ~n14782 & n14781 ) ;
  assign n14784 = ( n713 & ~n14778 ) | ( n713 & n14783 ) | ( ~n14778 & n14783 ) ;
  assign n14785 = n595 &  n14784 ;
  assign n14786 = n14232 | n14341 ;
  assign n14787 = ( n14219 & n14228 ) | ( n14219 & n14232 ) | ( n14228 & n14232 ) ;
  assign n14788 = ( n14786 & ~n14228 ) | ( n14786 & n14787 ) | ( ~n14228 & n14787 ) ;
  assign n14789 = ( n14232 & ~n14787 ) | ( n14232 & n14786 ) | ( ~n14787 & n14786 ) ;
  assign n14790 = ( n14219 & ~n14788 ) | ( n14219 & n14789 ) | ( ~n14788 & n14789 ) ;
  assign n14791 = n713 | n14763 ;
  assign n14792 = ( n14777 & ~n14791 ) | ( n14777 & 1'b0 ) | ( ~n14791 & 1'b0 ) ;
  assign n14793 = ( n14783 & ~n14792 ) | ( n14783 & 1'b0 ) | ( ~n14792 & 1'b0 ) ;
  assign n14794 = ~n14771 & n14774 ;
  assign n14795 = ( n14768 & ~n837 ) | ( n14768 & n14794 ) | ( ~n837 & n14794 ) ;
  assign n14796 = ( n713 & ~n14795 ) | ( n713 & 1'b0 ) | ( ~n14795 & 1'b0 ) ;
  assign n14797 = n595 | n14796 ;
  assign n14798 = n14793 | n14797 ;
  assign n14799 = n14790 &  n14798 ;
  assign n14800 = n14785 | n14799 ;
  assign n14806 = ( n492 & ~n14805 ) | ( n492 & n14800 ) | ( ~n14805 & n14800 ) ;
  assign n14807 = n396 &  n14806 ;
  assign n14808 = n14254 | n14341 ;
  assign n14809 = ( n14241 & n14250 ) | ( n14241 & n14254 ) | ( n14250 & n14254 ) ;
  assign n14810 = ( n14808 & ~n14250 ) | ( n14808 & n14809 ) | ( ~n14250 & n14809 ) ;
  assign n14811 = ( n14254 & ~n14809 ) | ( n14254 & n14808 ) | ( ~n14809 & n14808 ) ;
  assign n14812 = ( n14241 & ~n14810 ) | ( n14241 & n14811 ) | ( ~n14810 & n14811 ) ;
  assign n14813 = n492 | n14785 ;
  assign n14814 = n14799 | n14813 ;
  assign n14815 = ~n14805 & n14814 ;
  assign n14816 = n14793 | n14796 ;
  assign n14817 = ( n595 & n14790 ) | ( n595 & n14816 ) | ( n14790 & n14816 ) ;
  assign n14818 = n492 &  n14817 ;
  assign n14819 = n396 | n14818 ;
  assign n14820 = n14815 | n14819 ;
  assign n14821 = n14812 &  n14820 ;
  assign n14822 = n14807 | n14821 ;
  assign n14828 = ( n315 & ~n14827 ) | ( n315 & n14822 ) | ( ~n14827 & n14822 ) ;
  assign n14829 = n240 &  n14828 ;
  assign n14831 = ( n14272 & ~n14263 ) | ( n14272 & n14276 ) | ( ~n14263 & n14276 ) ;
  assign n14830 = n14276 | n14341 ;
  assign n14833 = ( n14276 & ~n14831 ) | ( n14276 & n14830 ) | ( ~n14831 & n14830 ) ;
  assign n14832 = ( n14830 & ~n14272 ) | ( n14830 & n14831 ) | ( ~n14272 & n14831 ) ;
  assign n14834 = ( n14263 & ~n14833 ) | ( n14263 & n14832 ) | ( ~n14833 & n14832 ) ;
  assign n14835 = n315 | n14807 ;
  assign n14836 = n14821 | n14835 ;
  assign n14837 = ~n14827 & n14836 ;
  assign n14838 = n14815 | n14818 ;
  assign n14839 = ( n396 & n14812 ) | ( n396 & n14838 ) | ( n14812 & n14838 ) ;
  assign n14840 = n315 &  n14839 ;
  assign n14841 = n240 | n14840 ;
  assign n14842 = n14837 | n14841 ;
  assign n14843 = ~n14834 & n14842 ;
  assign n14844 = n14829 | n14843 ;
  assign n14845 = ~n14278 & n14341 ;
  assign n14846 = ( n14265 & n14270 ) | ( n14265 & n14341 ) | ( n14270 & n14341 ) ;
  assign n14848 = ( n14845 & ~n14265 ) | ( n14845 & n14846 ) | ( ~n14265 & n14846 ) ;
  assign n14847 = ( n14341 & ~n14846 ) | ( n14341 & n14845 ) | ( ~n14846 & n14845 ) ;
  assign n14849 = ( n14270 & ~n14848 ) | ( n14270 & n14847 ) | ( ~n14848 & n14847 ) ;
  assign n14850 = ( n181 & n14844 ) | ( n181 & n14849 ) | ( n14844 & n14849 ) ;
  assign n14851 = ~n145 & n14850 ;
  assign n14853 = ( n14294 & ~n14285 ) | ( n14294 & n14298 ) | ( ~n14285 & n14298 ) ;
  assign n14852 = n14298 | n14341 ;
  assign n14855 = ( n14298 & ~n14853 ) | ( n14298 & n14852 ) | ( ~n14853 & n14852 ) ;
  assign n14854 = ( n14852 & ~n14294 ) | ( n14852 & n14853 ) | ( ~n14294 & n14853 ) ;
  assign n14856 = ( n14285 & ~n14855 ) | ( n14285 & n14854 ) | ( ~n14855 & n14854 ) ;
  assign n14857 = n181 | n14829 ;
  assign n14858 = n14843 | n14857 ;
  assign n14859 = n14849 &  n14858 ;
  assign n14860 = n14837 | n14840 ;
  assign n14861 = ( n240 & ~n14834 ) | ( n240 & n14860 ) | ( ~n14834 & n14860 ) ;
  assign n14862 = n181 &  n14861 ;
  assign n14863 = ( n145 & ~n14862 ) | ( n145 & 1'b0 ) | ( ~n14862 & 1'b0 ) ;
  assign n14864 = ~n14859 & n14863 ;
  assign n14865 = ( n14856 & ~n14864 ) | ( n14856 & 1'b0 ) | ( ~n14864 & 1'b0 ) ;
  assign n14866 = n14851 | n14865 ;
  assign n14872 = ( n150 & ~n14871 ) | ( n150 & n14866 ) | ( ~n14871 & n14866 ) ;
  assign n14873 = n14307 | n14326 ;
  assign n14874 = ( n14323 & ~n14873 ) | ( n14323 & n14341 ) | ( ~n14873 & n14341 ) ;
  assign n14875 = ~n14323 & n14874 ;
  assign n14876 = n14323 | n14326 ;
  assign n14877 = n14341 | n14876 ;
  assign n14878 = ( n14307 & ~n14877 ) | ( n14307 & n14876 ) | ( ~n14877 & n14876 ) ;
  assign n14879 = n14875 | n14878 ;
  assign n14880 = n14308 &  n14315 ;
  assign n14881 = ~n14341 & n14880 ;
  assign n14882 = ( n14329 & ~n14880 ) | ( n14329 & n14881 ) | ( ~n14880 & n14881 ) ;
  assign n14883 = n14879 &  n14882 ;
  assign n14884 = ~n14872 & n14883 ;
  assign n14885 = ( n133 & ~n14884 ) | ( n133 & n14883 ) | ( ~n14884 & n14883 ) ;
  assign n14888 = n14859 | n14862 ;
  assign n14889 = ( n14856 & ~n145 ) | ( n14856 & n14888 ) | ( ~n145 & n14888 ) ;
  assign n14890 = n150 &  n14889 ;
  assign n14891 = n14879 | n14890 ;
  assign n14886 = n150 | n14851 ;
  assign n14887 = n14865 | n14886 ;
  assign n14892 = n14871 | n14887 ;
  assign n14893 = ( n14891 & ~n14871 ) | ( n14891 & n14892 ) | ( ~n14871 & n14892 ) ;
  assign n14895 = ( n133 & n14308 ) | ( n133 & n14315 ) | ( n14308 & n14315 ) ;
  assign n14894 = ( n14308 & ~n14341 ) | ( n14308 & n14315 ) | ( ~n14341 & n14315 ) ;
  assign n14896 = ( n14315 & ~n14894 ) | ( n14315 & 1'b0 ) | ( ~n14894 & 1'b0 ) ;
  assign n14897 = ( n14895 & ~n14315 ) | ( n14895 & n14896 ) | ( ~n14315 & n14896 ) ;
  assign n14898 = n14311 | n14338 ;
  assign n14899 = ( n14333 & ~n14314 ) | ( n14333 & n14898 ) | ( ~n14314 & n14898 ) ;
  assign n14900 = n14314 | n14899 ;
  assign n14901 = ( n14321 & ~n14329 ) | ( n14321 & n14900 ) | ( ~n14329 & n14900 ) ;
  assign n14902 = ( n14321 & ~n14901 ) | ( n14321 & 1'b0 ) | ( ~n14901 & 1'b0 ) ;
  assign n14903 = n14897 | n14902 ;
  assign n14904 = ( n14893 & ~n14903 ) | ( n14893 & 1'b0 ) | ( ~n14903 & 1'b0 ) ;
  assign n14905 = ~n14885 | ~n14904 ;
  assign n15322 = n14748 | n14905 ;
  assign n15323 = ( n14740 & ~n14748 ) | ( n14740 & n14744 ) | ( ~n14748 & n14744 ) ;
  assign n15325 = ( n14748 & n15322 ) | ( n14748 & n15323 ) | ( n15322 & n15323 ) ;
  assign n15324 = ( n14744 & ~n15323 ) | ( n14744 & n15322 ) | ( ~n15323 & n15322 ) ;
  assign n15326 = ( n14740 & ~n15325 ) | ( n14740 & n15324 ) | ( ~n15325 & n15324 ) ;
  assign n15425 = ( n14829 & ~n14834 ) | ( n14829 & n14905 ) | ( ~n14834 & n14905 ) ;
  assign n15424 = ~n14842 & n14905 ;
  assign n15426 = ( n14905 & ~n15425 ) | ( n14905 & n15424 ) | ( ~n15425 & n15424 ) ;
  assign n15427 = ( n15424 & ~n14829 ) | ( n15424 & n15425 ) | ( ~n14829 & n15425 ) ;
  assign n15428 = ( n14834 & ~n15426 ) | ( n14834 & n15427 ) | ( ~n15426 & n15427 ) ;
  assign n15359 = ( n14763 & ~n14768 ) | ( n14763 & n14905 ) | ( ~n14768 & n14905 ) ;
  assign n15358 = n14776 &  n14905 ;
  assign n15360 = ( n14905 & ~n15359 ) | ( n14905 & n15358 ) | ( ~n15359 & n15358 ) ;
  assign n15361 = ( n15358 & ~n14763 ) | ( n15358 & n15359 ) | ( ~n14763 & n15359 ) ;
  assign n15362 = ( n14768 & ~n15360 ) | ( n14768 & n15361 ) | ( ~n15360 & n15361 ) ;
  assign n15228 = ( n14632 & ~n14637 ) | ( n14632 & n14645 ) | ( ~n14637 & n14645 ) ;
  assign n15227 = n14632 | n14905 ;
  assign n15230 = ( n14632 & ~n15228 ) | ( n14632 & n15227 ) | ( ~n15228 & n15227 ) ;
  assign n15229 = ( n15227 & ~n14645 ) | ( n15227 & n15228 ) | ( ~n14645 & n15228 ) ;
  assign n15231 = ( n14637 & ~n15230 ) | ( n14637 & n15229 ) | ( ~n15230 & n15229 ) ;
  assign n15206 = ( n14610 & ~n14615 ) | ( n14610 & n14623 ) | ( ~n14615 & n14623 ) ;
  assign n15205 = n14610 | n14905 ;
  assign n15208 = ( n14610 & ~n15206 ) | ( n14610 & n15205 ) | ( ~n15206 & n15205 ) ;
  assign n15207 = ( n15205 & ~n14623 ) | ( n15205 & n15206 ) | ( ~n14623 & n15206 ) ;
  assign n15209 = ( n14615 & ~n15208 ) | ( n14615 & n15207 ) | ( ~n15208 & n15207 ) ;
  assign n14912 = ( x26 & ~n14905 ) | ( x26 & x27 ) | ( ~n14905 & x27 ) ;
  assign n14918 = ( x26 & ~x27 ) | ( x26 & 1'b0 ) | ( ~x27 & 1'b0 ) ;
  assign n14908 = x24 | x25 ;
  assign n14913 = ~x26 & n14908 ;
  assign n14914 = ( x26 & ~n14339 ) | ( x26 & n14913 ) | ( ~n14339 & n14913 ) ;
  assign n14915 = ( n14329 & ~n14321 ) | ( n14329 & n14914 ) | ( ~n14321 & n14914 ) ;
  assign n14916 = n14321 &  n14915 ;
  assign n14917 = ( n14905 & ~x27 ) | ( n14905 & n14916 ) | ( ~x27 & n14916 ) ;
  assign n14919 = ( n14912 & ~n14918 ) | ( n14912 & n14917 ) | ( ~n14918 & n14917 ) ;
  assign n14909 = x26 | n14908 ;
  assign n14910 = x26 &  n14905 ;
  assign n14911 = ( n14341 & ~n14909 ) | ( n14341 & n14910 ) | ( ~n14909 & n14910 ) ;
  assign n14920 = n14911 &  n14919 ;
  assign n14921 = ( n13784 & ~n14919 ) | ( n13784 & n14920 ) | ( ~n14919 & n14920 ) ;
  assign n14922 = n13784 | n14911 ;
  assign n14923 = ( n14919 & ~n14922 ) | ( n14919 & 1'b0 ) | ( ~n14922 & 1'b0 ) ;
  assign n14925 = ( n14341 & ~n14902 ) | ( n14341 & 1'b0 ) | ( ~n14902 & 1'b0 ) ;
  assign n14926 = ( n14893 & ~n14925 ) | ( n14893 & n14897 ) | ( ~n14925 & n14897 ) ;
  assign n14927 = ( n14893 & ~n14926 ) | ( n14893 & 1'b0 ) | ( ~n14926 & 1'b0 ) ;
  assign n14928 = n14885 &  n14927 ;
  assign n14924 = ~n13785 & n14905 ;
  assign n14929 = ( n14924 & ~n14928 ) | ( n14924 & 1'b0 ) | ( ~n14928 & 1'b0 ) ;
  assign n14930 = ( x28 & n14928 ) | ( x28 & n14929 ) | ( n14928 & n14929 ) ;
  assign n14931 = x28 | n14928 ;
  assign n14932 = n14924 | n14931 ;
  assign n14933 = ~n14930 & n14932 ;
  assign n14934 = n14923 | n14933 ;
  assign n14935 = ~n14921 & n14934 ;
  assign n14939 = ~x28 & n14341 ;
  assign n14940 = ( x29 & ~n14939 ) | ( x29 & 1'b0 ) | ( ~n14939 & 1'b0 ) ;
  assign n14941 = n14353 | n14940 ;
  assign n14936 = ( n14341 & ~x28 ) | ( n14341 & n14348 ) | ( ~x28 & n14348 ) ;
  assign n14937 = x28 &  n14936 ;
  assign n14938 = ( n14343 & ~n14937 ) | ( n14343 & n14348 ) | ( ~n14937 & n14348 ) ;
  assign n14942 = ( n14905 & ~n14941 ) | ( n14905 & n14938 ) | ( ~n14941 & n14938 ) ;
  assign n14944 = ( n14905 & ~n14942 ) | ( n14905 & 1'b0 ) | ( ~n14942 & 1'b0 ) ;
  assign n14943 = ~n14938 & n14942 ;
  assign n14945 = ( n14941 & ~n14944 ) | ( n14941 & n14943 ) | ( ~n14944 & n14943 ) ;
  assign n14946 = ( n14935 & ~n13242 ) | ( n14935 & n14945 ) | ( ~n13242 & n14945 ) ;
  assign n14947 = ( n12707 & ~n14946 ) | ( n12707 & 1'b0 ) | ( ~n14946 & 1'b0 ) ;
  assign n14948 = ~n14376 & n14379 ;
  assign n14949 = ( n14362 & ~n14376 ) | ( n14362 & n14948 ) | ( ~n14376 & n14948 ) ;
  assign n14951 = ( n14905 & n14376 ) | ( n14905 & n14949 ) | ( n14376 & n14949 ) ;
  assign n14950 = ( n14905 & ~n14949 ) | ( n14905 & n14948 ) | ( ~n14949 & n14948 ) ;
  assign n14952 = ( n14362 & ~n14951 ) | ( n14362 & n14950 ) | ( ~n14951 & n14950 ) ;
  assign n14953 = n13242 | n14921 ;
  assign n14954 = ( n14934 & ~n14953 ) | ( n14934 & 1'b0 ) | ( ~n14953 & 1'b0 ) ;
  assign n14955 = n14945 | n14954 ;
  assign n14956 = ~n14911 & n14919 ;
  assign n14957 = ( n14933 & ~n13784 ) | ( n14933 & n14956 ) | ( ~n13784 & n14956 ) ;
  assign n14958 = ( n13242 & ~n14957 ) | ( n13242 & 1'b0 ) | ( ~n14957 & 1'b0 ) ;
  assign n14959 = n12707 | n14958 ;
  assign n14960 = ( n14955 & ~n14959 ) | ( n14955 & 1'b0 ) | ( ~n14959 & 1'b0 ) ;
  assign n14961 = n14952 | n14960 ;
  assign n14962 = ~n14947 & n14961 ;
  assign n14963 = n14364 | n14905 ;
  assign n14964 = ( n14364 & ~n14381 ) | ( n14364 & n14374 ) | ( ~n14381 & n14374 ) ;
  assign n14965 = ( n14381 & n14963 ) | ( n14381 & n14964 ) | ( n14963 & n14964 ) ;
  assign n14966 = ( n14364 & ~n14964 ) | ( n14364 & n14963 ) | ( ~n14964 & n14963 ) ;
  assign n14967 = ( n14374 & ~n14965 ) | ( n14374 & n14966 ) | ( ~n14965 & n14966 ) ;
  assign n14968 = ( n14962 & ~n12187 ) | ( n14962 & n14967 ) | ( ~n12187 & n14967 ) ;
  assign n14969 = ( n11674 & ~n14968 ) | ( n11674 & 1'b0 ) | ( ~n14968 & 1'b0 ) ;
  assign n14970 = n14401 | n14905 ;
  assign n14971 = ( n14388 & ~n14401 ) | ( n14388 & n14397 ) | ( ~n14401 & n14397 ) ;
  assign n14973 = ( n14401 & n14970 ) | ( n14401 & n14971 ) | ( n14970 & n14971 ) ;
  assign n14972 = ( n14397 & ~n14971 ) | ( n14397 & n14970 ) | ( ~n14971 & n14970 ) ;
  assign n14974 = ( n14388 & ~n14973 ) | ( n14388 & n14972 ) | ( ~n14973 & n14972 ) ;
  assign n14975 = n12187 | n14947 ;
  assign n14976 = ( n14961 & ~n14975 ) | ( n14961 & 1'b0 ) | ( ~n14975 & 1'b0 ) ;
  assign n14977 = n14967 | n14976 ;
  assign n14978 = ( n14955 & ~n14958 ) | ( n14955 & 1'b0 ) | ( ~n14958 & 1'b0 ) ;
  assign n14979 = ( n14952 & ~n12707 ) | ( n14952 & n14978 ) | ( ~n12707 & n14978 ) ;
  assign n14980 = ( n12187 & ~n14979 ) | ( n12187 & 1'b0 ) | ( ~n14979 & 1'b0 ) ;
  assign n14981 = n11674 | n14980 ;
  assign n14982 = ( n14977 & ~n14981 ) | ( n14977 & 1'b0 ) | ( ~n14981 & 1'b0 ) ;
  assign n14983 = n14974 | n14982 ;
  assign n14984 = ~n14969 & n14983 ;
  assign n14985 = n14403 &  n14905 ;
  assign n14986 = ( n14390 & n14395 ) | ( n14390 & n14905 ) | ( n14395 & n14905 ) ;
  assign n14988 = ( n14985 & ~n14390 ) | ( n14985 & n14986 ) | ( ~n14390 & n14986 ) ;
  assign n14987 = ( n14905 & ~n14986 ) | ( n14905 & n14985 ) | ( ~n14986 & n14985 ) ;
  assign n14989 = ( n14395 & ~n14988 ) | ( n14395 & n14987 ) | ( ~n14988 & n14987 ) ;
  assign n14990 = ( n14984 & ~n11176 ) | ( n14984 & n14989 ) | ( ~n11176 & n14989 ) ;
  assign n14991 = ( n10685 & ~n14990 ) | ( n10685 & 1'b0 ) | ( ~n14990 & 1'b0 ) ;
  assign n14992 = n14423 | n14905 ;
  assign n14993 = ( n14410 & ~n14419 ) | ( n14410 & n14423 ) | ( ~n14419 & n14423 ) ;
  assign n14994 = ( n14419 & n14992 ) | ( n14419 & n14993 ) | ( n14992 & n14993 ) ;
  assign n14995 = ( n14423 & ~n14993 ) | ( n14423 & n14992 ) | ( ~n14993 & n14992 ) ;
  assign n14996 = ( n14410 & ~n14994 ) | ( n14410 & n14995 ) | ( ~n14994 & n14995 ) ;
  assign n14997 = n11176 | n14969 ;
  assign n14998 = ( n14983 & ~n14997 ) | ( n14983 & 1'b0 ) | ( ~n14997 & 1'b0 ) ;
  assign n14999 = n14989 | n14998 ;
  assign n15000 = ( n14977 & ~n14980 ) | ( n14977 & 1'b0 ) | ( ~n14980 & 1'b0 ) ;
  assign n15001 = ( n14974 & ~n11674 ) | ( n14974 & n15000 ) | ( ~n11674 & n15000 ) ;
  assign n15002 = ( n11176 & ~n15001 ) | ( n11176 & 1'b0 ) | ( ~n15001 & 1'b0 ) ;
  assign n15003 = n10685 | n15002 ;
  assign n15004 = ( n14999 & ~n15003 ) | ( n14999 & 1'b0 ) | ( ~n15003 & 1'b0 ) ;
  assign n15005 = n14996 | n15004 ;
  assign n15006 = ~n14991 & n15005 ;
  assign n15007 = n14412 | n14905 ;
  assign n15008 = ( n14417 & ~n14412 ) | ( n14417 & n14425 ) | ( ~n14412 & n14425 ) ;
  assign n15010 = ( n14412 & n15007 ) | ( n14412 & n15008 ) | ( n15007 & n15008 ) ;
  assign n15009 = ( n14425 & ~n15008 ) | ( n14425 & n15007 ) | ( ~n15008 & n15007 ) ;
  assign n15011 = ( n14417 & ~n15010 ) | ( n14417 & n15009 ) | ( ~n15010 & n15009 ) ;
  assign n15012 = ( n15006 & ~n10209 ) | ( n15006 & n15011 ) | ( ~n10209 & n15011 ) ;
  assign n15013 = n9740 | n15012 ;
  assign n15014 = n14445 | n14905 ;
  assign n15015 = ( n14432 & ~n14441 ) | ( n14432 & n14445 ) | ( ~n14441 & n14445 ) ;
  assign n15016 = ( n14441 & n15014 ) | ( n14441 & n15015 ) | ( n15014 & n15015 ) ;
  assign n15017 = ( n14445 & ~n15015 ) | ( n14445 & n15014 ) | ( ~n15015 & n15014 ) ;
  assign n15018 = ( n14432 & ~n15016 ) | ( n14432 & n15017 ) | ( ~n15016 & n15017 ) ;
  assign n15019 = n10209 | n14991 ;
  assign n15020 = ( n15005 & ~n15019 ) | ( n15005 & 1'b0 ) | ( ~n15019 & 1'b0 ) ;
  assign n15021 = n15011 | n15020 ;
  assign n15022 = ( n14999 & ~n15002 ) | ( n14999 & 1'b0 ) | ( ~n15002 & 1'b0 ) ;
  assign n15023 = ( n14996 & ~n10685 ) | ( n14996 & n15022 ) | ( ~n10685 & n15022 ) ;
  assign n15024 = ( n10209 & ~n15023 ) | ( n10209 & 1'b0 ) | ( ~n15023 & 1'b0 ) ;
  assign n15025 = ( n9740 & ~n15024 ) | ( n9740 & 1'b0 ) | ( ~n15024 & 1'b0 ) ;
  assign n15026 = n15021 &  n15025 ;
  assign n15027 = n15018 | n15026 ;
  assign n15028 = n15013 &  n15027 ;
  assign n15030 = ( n14434 & ~n14439 ) | ( n14434 & n14447 ) | ( ~n14439 & n14447 ) ;
  assign n15029 = ( n14434 & ~n14905 ) | ( n14434 & 1'b0 ) | ( ~n14905 & 1'b0 ) ;
  assign n15032 = ( n14434 & ~n15030 ) | ( n14434 & n15029 ) | ( ~n15030 & n15029 ) ;
  assign n15031 = ( n15029 & ~n14447 ) | ( n15029 & n15030 ) | ( ~n14447 & n15030 ) ;
  assign n15033 = ( n14439 & ~n15032 ) | ( n14439 & n15031 ) | ( ~n15032 & n15031 ) ;
  assign n15034 = ( n15028 & ~n9286 ) | ( n15028 & n15033 ) | ( ~n9286 & n15033 ) ;
  assign n15035 = ( n8839 & ~n15034 ) | ( n8839 & 1'b0 ) | ( ~n15034 & 1'b0 ) ;
  assign n15036 = n14467 | n14905 ;
  assign n15037 = ( n14454 & ~n14467 ) | ( n14454 & n14463 ) | ( ~n14467 & n14463 ) ;
  assign n15039 = ( n14467 & n15036 ) | ( n14467 & n15037 ) | ( n15036 & n15037 ) ;
  assign n15038 = ( n14463 & ~n15037 ) | ( n14463 & n15036 ) | ( ~n15037 & n15036 ) ;
  assign n15040 = ( n14454 & ~n15039 ) | ( n14454 & n15038 ) | ( ~n15039 & n15038 ) ;
  assign n15041 = ~n9286 & n15013 ;
  assign n15042 = n15027 &  n15041 ;
  assign n15043 = n15033 | n15042 ;
  assign n15044 = ( n15021 & ~n15024 ) | ( n15021 & 1'b0 ) | ( ~n15024 & 1'b0 ) ;
  assign n15045 = ( n9740 & n15018 ) | ( n9740 & n15044 ) | ( n15018 & n15044 ) ;
  assign n15046 = ( n9286 & ~n15045 ) | ( n9286 & 1'b0 ) | ( ~n15045 & 1'b0 ) ;
  assign n15047 = n8839 | n15046 ;
  assign n15048 = ( n15043 & ~n15047 ) | ( n15043 & 1'b0 ) | ( ~n15047 & 1'b0 ) ;
  assign n15049 = n15040 | n15048 ;
  assign n15050 = ~n15035 & n15049 ;
  assign n15051 = n14469 &  n14905 ;
  assign n15052 = ( n14456 & n14461 ) | ( n14456 & n14905 ) | ( n14461 & n14905 ) ;
  assign n15054 = ( n15051 & ~n14456 ) | ( n15051 & n15052 ) | ( ~n14456 & n15052 ) ;
  assign n15053 = ( n14905 & ~n15052 ) | ( n14905 & n15051 ) | ( ~n15052 & n15051 ) ;
  assign n15055 = ( n14461 & ~n15054 ) | ( n14461 & n15053 ) | ( ~n15054 & n15053 ) ;
  assign n15056 = ( n15050 & ~n8407 ) | ( n15050 & n15055 ) | ( ~n8407 & n15055 ) ;
  assign n15057 = ( n7982 & ~n15056 ) | ( n7982 & 1'b0 ) | ( ~n15056 & 1'b0 ) ;
  assign n15058 = n14489 | n14905 ;
  assign n15059 = ( n14476 & ~n14485 ) | ( n14476 & n14489 ) | ( ~n14485 & n14489 ) ;
  assign n15060 = ( n14485 & n15058 ) | ( n14485 & n15059 ) | ( n15058 & n15059 ) ;
  assign n15061 = ( n14489 & ~n15059 ) | ( n14489 & n15058 ) | ( ~n15059 & n15058 ) ;
  assign n15062 = ( n14476 & ~n15060 ) | ( n14476 & n15061 ) | ( ~n15060 & n15061 ) ;
  assign n15063 = n8407 | n15035 ;
  assign n15064 = ( n15049 & ~n15063 ) | ( n15049 & 1'b0 ) | ( ~n15063 & 1'b0 ) ;
  assign n15065 = n15055 | n15064 ;
  assign n15066 = ( n15043 & ~n15046 ) | ( n15043 & 1'b0 ) | ( ~n15046 & 1'b0 ) ;
  assign n15067 = ( n15040 & ~n8839 ) | ( n15040 & n15066 ) | ( ~n8839 & n15066 ) ;
  assign n15068 = ( n8407 & ~n15067 ) | ( n8407 & 1'b0 ) | ( ~n15067 & 1'b0 ) ;
  assign n15069 = n7982 | n15068 ;
  assign n15070 = ( n15065 & ~n15069 ) | ( n15065 & 1'b0 ) | ( ~n15069 & 1'b0 ) ;
  assign n15071 = n15062 | n15070 ;
  assign n15072 = ~n15057 & n15071 ;
  assign n15073 = n14478 | n14905 ;
  assign n15074 = ( n14483 & ~n14478 ) | ( n14483 & n14491 ) | ( ~n14478 & n14491 ) ;
  assign n15076 = ( n14478 & n15073 ) | ( n14478 & n15074 ) | ( n15073 & n15074 ) ;
  assign n15075 = ( n14491 & ~n15074 ) | ( n14491 & n15073 ) | ( ~n15074 & n15073 ) ;
  assign n15077 = ( n14483 & ~n15076 ) | ( n14483 & n15075 ) | ( ~n15076 & n15075 ) ;
  assign n15078 = ( n7572 & n15072 ) | ( n7572 & n15077 ) | ( n15072 & n15077 ) ;
  assign n15079 = n7169 | n15078 ;
  assign n15081 = ( n14507 & ~n14498 ) | ( n14507 & n14511 ) | ( ~n14498 & n14511 ) ;
  assign n15080 = ( n14511 & ~n14905 ) | ( n14511 & 1'b0 ) | ( ~n14905 & 1'b0 ) ;
  assign n15083 = ( n14511 & ~n15081 ) | ( n14511 & n15080 ) | ( ~n15081 & n15080 ) ;
  assign n15082 = ( n15080 & ~n14507 ) | ( n15080 & n15081 ) | ( ~n14507 & n15081 ) ;
  assign n15084 = ( n14498 & ~n15083 ) | ( n14498 & n15082 ) | ( ~n15083 & n15082 ) ;
  assign n15085 = ( n7572 & ~n15057 ) | ( n7572 & 1'b0 ) | ( ~n15057 & 1'b0 ) ;
  assign n15086 = n15071 &  n15085 ;
  assign n15087 = n15077 | n15086 ;
  assign n15088 = ( n15065 & ~n15068 ) | ( n15065 & 1'b0 ) | ( ~n15068 & 1'b0 ) ;
  assign n15089 = ( n15062 & ~n7982 ) | ( n15062 & n15088 ) | ( ~n7982 & n15088 ) ;
  assign n15090 = n7572 | n15089 ;
  assign n15091 = n7169 &  n15090 ;
  assign n15092 = n15087 &  n15091 ;
  assign n15093 = n15084 | n15092 ;
  assign n15094 = n15079 &  n15093 ;
  assign n15095 = ( n14500 & ~n14905 ) | ( n14500 & 1'b0 ) | ( ~n14905 & 1'b0 ) ;
  assign n15096 = ( n14500 & n14505 ) | ( n14500 & n14513 ) | ( n14505 & n14513 ) ;
  assign n15097 = ( n15095 & ~n14513 ) | ( n15095 & n15096 ) | ( ~n14513 & n15096 ) ;
  assign n15098 = ( n14500 & ~n15096 ) | ( n14500 & n15095 ) | ( ~n15096 & n15095 ) ;
  assign n15099 = ( n14505 & ~n15097 ) | ( n14505 & n15098 ) | ( ~n15097 & n15098 ) ;
  assign n15100 = ( n15094 & ~n6781 ) | ( n15094 & n15099 ) | ( ~n6781 & n15099 ) ;
  assign n15101 = n6399 | n15100 ;
  assign n15102 = n14533 | n14905 ;
  assign n15103 = ( n14520 & ~n14529 ) | ( n14520 & n14533 ) | ( ~n14529 & n14533 ) ;
  assign n15104 = ( n14529 & n15102 ) | ( n14529 & n15103 ) | ( n15102 & n15103 ) ;
  assign n15105 = ( n14533 & ~n15103 ) | ( n14533 & n15102 ) | ( ~n15103 & n15102 ) ;
  assign n15106 = ( n14520 & ~n15104 ) | ( n14520 & n15105 ) | ( ~n15104 & n15105 ) ;
  assign n15107 = ~n6781 & n15079 ;
  assign n15108 = n15093 &  n15107 ;
  assign n15109 = n15099 | n15108 ;
  assign n15110 = n15087 &  n15090 ;
  assign n15111 = ( n7169 & n15084 ) | ( n7169 & n15110 ) | ( n15084 & n15110 ) ;
  assign n15112 = ( n6781 & ~n15111 ) | ( n6781 & 1'b0 ) | ( ~n15111 & 1'b0 ) ;
  assign n15113 = ( n6399 & ~n15112 ) | ( n6399 & 1'b0 ) | ( ~n15112 & 1'b0 ) ;
  assign n15114 = n15109 &  n15113 ;
  assign n15115 = n15106 | n15114 ;
  assign n15116 = n15101 &  n15115 ;
  assign n15117 = ( n14522 & ~n14905 ) | ( n14522 & 1'b0 ) | ( ~n14905 & 1'b0 ) ;
  assign n15118 = ( n14522 & n14527 ) | ( n14522 & n14535 ) | ( n14527 & n14535 ) ;
  assign n15119 = ( n15117 & ~n14535 ) | ( n15117 & n15118 ) | ( ~n14535 & n15118 ) ;
  assign n15120 = ( n14522 & ~n15118 ) | ( n14522 & n15117 ) | ( ~n15118 & n15117 ) ;
  assign n15121 = ( n14527 & ~n15119 ) | ( n14527 & n15120 ) | ( ~n15119 & n15120 ) ;
  assign n15122 = ( n15116 & ~n6032 ) | ( n15116 & n15121 ) | ( ~n6032 & n15121 ) ;
  assign n15123 = n5672 | n15122 ;
  assign n15124 = n14555 | n14905 ;
  assign n15125 = ( n14542 & ~n14551 ) | ( n14542 & n14555 ) | ( ~n14551 & n14555 ) ;
  assign n15126 = ( n14551 & n15124 ) | ( n14551 & n15125 ) | ( n15124 & n15125 ) ;
  assign n15127 = ( n14555 & ~n15125 ) | ( n14555 & n15124 ) | ( ~n15125 & n15124 ) ;
  assign n15128 = ( n14542 & ~n15126 ) | ( n14542 & n15127 ) | ( ~n15126 & n15127 ) ;
  assign n15129 = ~n6032 & n15101 ;
  assign n15130 = n15115 &  n15129 ;
  assign n15131 = n15121 | n15130 ;
  assign n15132 = ( n15109 & ~n15112 ) | ( n15109 & 1'b0 ) | ( ~n15112 & 1'b0 ) ;
  assign n15133 = ( n6399 & n15106 ) | ( n6399 & n15132 ) | ( n15106 & n15132 ) ;
  assign n15134 = ( n6032 & ~n15133 ) | ( n6032 & 1'b0 ) | ( ~n15133 & 1'b0 ) ;
  assign n15135 = ( n5672 & ~n15134 ) | ( n5672 & 1'b0 ) | ( ~n15134 & 1'b0 ) ;
  assign n15136 = n15131 &  n15135 ;
  assign n15137 = n15128 | n15136 ;
  assign n15138 = n15123 &  n15137 ;
  assign n15140 = ( n14544 & ~n14549 ) | ( n14544 & n14557 ) | ( ~n14549 & n14557 ) ;
  assign n15139 = ( n14544 & ~n14905 ) | ( n14544 & 1'b0 ) | ( ~n14905 & 1'b0 ) ;
  assign n15142 = ( n14544 & ~n15140 ) | ( n14544 & n15139 ) | ( ~n15140 & n15139 ) ;
  assign n15141 = ( n15139 & ~n14557 ) | ( n15139 & n15140 ) | ( ~n14557 & n15140 ) ;
  assign n15143 = ( n14549 & ~n15142 ) | ( n14549 & n15141 ) | ( ~n15142 & n15141 ) ;
  assign n15144 = ( n5327 & ~n15138 ) | ( n5327 & n15143 ) | ( ~n15138 & n15143 ) ;
  assign n15145 = n4990 &  n15144 ;
  assign n15146 = n14577 | n14905 ;
  assign n15147 = ( n14564 & ~n14577 ) | ( n14564 & n14573 ) | ( ~n14577 & n14573 ) ;
  assign n15149 = ( n14577 & n15146 ) | ( n14577 & n15147 ) | ( n15146 & n15147 ) ;
  assign n15148 = ( n14573 & ~n15147 ) | ( n14573 & n15146 ) | ( ~n15147 & n15146 ) ;
  assign n15150 = ( n14564 & ~n15149 ) | ( n14564 & n15148 ) | ( ~n15149 & n15148 ) ;
  assign n15151 = ~n5327 & n15123 ;
  assign n15152 = n15137 &  n15151 ;
  assign n15153 = ( n15143 & ~n15152 ) | ( n15143 & 1'b0 ) | ( ~n15152 & 1'b0 ) ;
  assign n15154 = ( n15131 & ~n15134 ) | ( n15131 & 1'b0 ) | ( ~n15134 & 1'b0 ) ;
  assign n15155 = ( n5672 & n15128 ) | ( n5672 & n15154 ) | ( n15128 & n15154 ) ;
  assign n15156 = ( n5327 & ~n15155 ) | ( n5327 & 1'b0 ) | ( ~n15155 & 1'b0 ) ;
  assign n15157 = n4990 | n15156 ;
  assign n15158 = n15153 | n15157 ;
  assign n15159 = n15150 &  n15158 ;
  assign n15160 = n15145 | n15159 ;
  assign n15161 = n14566 | n14905 ;
  assign n15162 = ( n14566 & n14571 ) | ( n14566 & n14579 ) | ( n14571 & n14579 ) ;
  assign n15163 = ( n15161 & ~n14579 ) | ( n15161 & n15162 ) | ( ~n14579 & n15162 ) ;
  assign n15164 = ( n14566 & ~n15162 ) | ( n14566 & n15161 ) | ( ~n15162 & n15161 ) ;
  assign n15165 = ( n14571 & ~n15163 ) | ( n14571 & n15164 ) | ( ~n15163 & n15164 ) ;
  assign n15166 = ( n4668 & n15160 ) | ( n4668 & n15165 ) | ( n15160 & n15165 ) ;
  assign n15167 = n4353 &  n15166 ;
  assign n15169 = ( n14595 & ~n14586 ) | ( n14595 & n14599 ) | ( ~n14586 & n14599 ) ;
  assign n15168 = n14599 | n14905 ;
  assign n15171 = ( n14599 & ~n15169 ) | ( n14599 & n15168 ) | ( ~n15169 & n15168 ) ;
  assign n15170 = ( n15168 & ~n14595 ) | ( n15168 & n15169 ) | ( ~n14595 & n15169 ) ;
  assign n15172 = ( n14586 & ~n15171 ) | ( n14586 & n15170 ) | ( ~n15171 & n15170 ) ;
  assign n15173 = n4668 | n15145 ;
  assign n15174 = n15159 | n15173 ;
  assign n15175 = n15165 &  n15174 ;
  assign n15176 = n15153 | n15156 ;
  assign n15177 = ( n4990 & n15150 ) | ( n4990 & n15176 ) | ( n15150 & n15176 ) ;
  assign n15178 = n4668 &  n15177 ;
  assign n15179 = n4353 | n15178 ;
  assign n15180 = n15175 | n15179 ;
  assign n15181 = n15172 &  n15180 ;
  assign n15182 = n15167 | n15181 ;
  assign n15183 = n14588 | n14905 ;
  assign n15184 = ( n14588 & n14593 ) | ( n14588 & n14601 ) | ( n14593 & n14601 ) ;
  assign n15185 = ( n15183 & ~n14601 ) | ( n15183 & n15184 ) | ( ~n14601 & n15184 ) ;
  assign n15186 = ( n14588 & ~n15184 ) | ( n14588 & n15183 ) | ( ~n15184 & n15183 ) ;
  assign n15187 = ( n14593 & ~n15185 ) | ( n14593 & n15186 ) | ( ~n15185 & n15186 ) ;
  assign n15188 = ( n4053 & n15182 ) | ( n4053 & n15187 ) | ( n15182 & n15187 ) ;
  assign n15189 = n3760 &  n15188 ;
  assign n15190 = n14621 | n14905 ;
  assign n15191 = ( n14608 & n14617 ) | ( n14608 & n14621 ) | ( n14617 & n14621 ) ;
  assign n15192 = ( n15190 & ~n14617 ) | ( n15190 & n15191 ) | ( ~n14617 & n15191 ) ;
  assign n15193 = ( n14621 & ~n15191 ) | ( n14621 & n15190 ) | ( ~n15191 & n15190 ) ;
  assign n15194 = ( n14608 & ~n15192 ) | ( n14608 & n15193 ) | ( ~n15192 & n15193 ) ;
  assign n15195 = n4053 | n15167 ;
  assign n15196 = n15181 | n15195 ;
  assign n15197 = n15187 &  n15196 ;
  assign n15198 = n15175 | n15178 ;
  assign n15199 = ( n4353 & n15172 ) | ( n4353 & n15198 ) | ( n15172 & n15198 ) ;
  assign n15200 = n4053 &  n15199 ;
  assign n15201 = n3760 | n15200 ;
  assign n15202 = n15197 | n15201 ;
  assign n15203 = ~n15194 & n15202 ;
  assign n15204 = n15189 | n15203 ;
  assign n15210 = ( n3482 & ~n15209 ) | ( n3482 & n15204 ) | ( ~n15209 & n15204 ) ;
  assign n15211 = n3211 &  n15210 ;
  assign n15213 = ( n14639 & ~n14630 ) | ( n14639 & n14643 ) | ( ~n14630 & n14643 ) ;
  assign n15212 = n14643 | n14905 ;
  assign n15215 = ( n14643 & ~n15213 ) | ( n14643 & n15212 ) | ( ~n15213 & n15212 ) ;
  assign n15214 = ( n15212 & ~n14639 ) | ( n15212 & n15213 ) | ( ~n14639 & n15213 ) ;
  assign n15216 = ( n14630 & ~n15215 ) | ( n14630 & n15214 ) | ( ~n15215 & n15214 ) ;
  assign n15217 = n3482 | n15189 ;
  assign n15218 = n15203 | n15217 ;
  assign n15219 = ~n15209 & n15218 ;
  assign n15220 = n15197 | n15200 ;
  assign n15221 = ( n3760 & ~n15194 ) | ( n3760 & n15220 ) | ( ~n15194 & n15220 ) ;
  assign n15222 = n3482 &  n15221 ;
  assign n15223 = n3211 | n15222 ;
  assign n15224 = n15219 | n15223 ;
  assign n15225 = n15216 &  n15224 ;
  assign n15226 = n15211 | n15225 ;
  assign n15232 = ( n2955 & ~n15231 ) | ( n2955 & n15226 ) | ( ~n15231 & n15226 ) ;
  assign n15233 = n2706 &  n15232 ;
  assign n15235 = ( n14661 & ~n14652 ) | ( n14661 & n14665 ) | ( ~n14652 & n14665 ) ;
  assign n15234 = n14665 | n14905 ;
  assign n15237 = ( n14665 & ~n15235 ) | ( n14665 & n15234 ) | ( ~n15235 & n15234 ) ;
  assign n15236 = ( n15234 & ~n14661 ) | ( n15234 & n15235 ) | ( ~n14661 & n15235 ) ;
  assign n15238 = ( n14652 & ~n15237 ) | ( n14652 & n15236 ) | ( ~n15237 & n15236 ) ;
  assign n15239 = n2955 | n15211 ;
  assign n15240 = n15225 | n15239 ;
  assign n15241 = ~n15231 & n15240 ;
  assign n15242 = n15219 | n15222 ;
  assign n15243 = ( n3211 & n15216 ) | ( n3211 & n15242 ) | ( n15216 & n15242 ) ;
  assign n15244 = n2955 &  n15243 ;
  assign n15245 = n2706 | n15244 ;
  assign n15246 = n15241 | n15245 ;
  assign n15247 = n15238 &  n15246 ;
  assign n15248 = n15233 | n15247 ;
  assign n15249 = n14654 | n14905 ;
  assign n15250 = ( n14654 & n14659 ) | ( n14654 & n14667 ) | ( n14659 & n14667 ) ;
  assign n15251 = ( n15249 & ~n14667 ) | ( n15249 & n15250 ) | ( ~n14667 & n15250 ) ;
  assign n15252 = ( n14654 & ~n15250 ) | ( n14654 & n15249 ) | ( ~n15250 & n15249 ) ;
  assign n15253 = ( n14659 & ~n15251 ) | ( n14659 & n15252 ) | ( ~n15251 & n15252 ) ;
  assign n15254 = ( n2472 & n15248 ) | ( n2472 & n15253 ) | ( n15248 & n15253 ) ;
  assign n15255 = n2245 &  n15254 ;
  assign n15256 = n14687 | n14905 ;
  assign n15257 = ( n14674 & n14683 ) | ( n14674 & n14687 ) | ( n14683 & n14687 ) ;
  assign n15258 = ( n15256 & ~n14683 ) | ( n15256 & n15257 ) | ( ~n14683 & n15257 ) ;
  assign n15259 = ( n14687 & ~n15257 ) | ( n14687 & n15256 ) | ( ~n15257 & n15256 ) ;
  assign n15260 = ( n14674 & ~n15258 ) | ( n14674 & n15259 ) | ( ~n15258 & n15259 ) ;
  assign n15261 = n2472 | n15233 ;
  assign n15262 = n15247 | n15261 ;
  assign n15263 = n15253 &  n15262 ;
  assign n15264 = n15241 | n15244 ;
  assign n15265 = ( n2706 & n15238 ) | ( n2706 & n15264 ) | ( n15238 & n15264 ) ;
  assign n15266 = n2472 &  n15265 ;
  assign n15267 = n2245 | n15266 ;
  assign n15268 = n15263 | n15267 ;
  assign n15269 = ~n15260 & n15268 ;
  assign n15270 = n15255 | n15269 ;
  assign n15272 = ( n14676 & ~n14681 ) | ( n14676 & n14689 ) | ( ~n14681 & n14689 ) ;
  assign n15271 = n14676 | n14905 ;
  assign n15274 = ( n14676 & ~n15272 ) | ( n14676 & n15271 ) | ( ~n15272 & n15271 ) ;
  assign n15273 = ( n15271 & ~n14689 ) | ( n15271 & n15272 ) | ( ~n14689 & n15272 ) ;
  assign n15275 = ( n14681 & ~n15274 ) | ( n14681 & n15273 ) | ( ~n15274 & n15273 ) ;
  assign n15276 = ( n2033 & ~n15270 ) | ( n2033 & n15275 ) | ( ~n15270 & n15275 ) ;
  assign n15277 = ( n1827 & ~n15276 ) | ( n1827 & 1'b0 ) | ( ~n15276 & 1'b0 ) ;
  assign n15278 = n14709 | n14905 ;
  assign n15279 = ( n14696 & ~n14705 ) | ( n14696 & n14709 ) | ( ~n14705 & n14709 ) ;
  assign n15280 = ( n14705 & n15278 ) | ( n14705 & n15279 ) | ( n15278 & n15279 ) ;
  assign n15281 = ( n14709 & ~n15279 ) | ( n14709 & n15278 ) | ( ~n15279 & n15278 ) ;
  assign n15282 = ( n14696 & ~n15280 ) | ( n14696 & n15281 ) | ( ~n15280 & n15281 ) ;
  assign n15283 = ( n2033 & ~n15255 ) | ( n2033 & 1'b0 ) | ( ~n15255 & 1'b0 ) ;
  assign n15284 = ~n15269 & n15283 ;
  assign n15285 = n15275 | n15284 ;
  assign n15286 = n15263 | n15266 ;
  assign n15287 = ( n2245 & ~n15260 ) | ( n2245 & n15286 ) | ( ~n15260 & n15286 ) ;
  assign n15288 = ~n2033 & n15287 ;
  assign n15289 = n1827 | n15288 ;
  assign n15290 = ( n15285 & ~n15289 ) | ( n15285 & 1'b0 ) | ( ~n15289 & 1'b0 ) ;
  assign n15291 = n15282 | n15290 ;
  assign n15292 = ~n15277 & n15291 ;
  assign n15293 = n14698 | n14905 ;
  assign n15294 = ( n14703 & ~n14698 ) | ( n14703 & n14711 ) | ( ~n14698 & n14711 ) ;
  assign n15296 = ( n14698 & n15293 ) | ( n14698 & n15294 ) | ( n15293 & n15294 ) ;
  assign n15295 = ( n14711 & ~n15294 ) | ( n14711 & n15293 ) | ( ~n15294 & n15293 ) ;
  assign n15297 = ( n14703 & ~n15296 ) | ( n14703 & n15295 ) | ( ~n15296 & n15295 ) ;
  assign n15298 = ( n1636 & n15292 ) | ( n1636 & n15297 ) | ( n15292 & n15297 ) ;
  assign n15299 = n1452 | n15298 ;
  assign n15300 = ( n14731 & ~n14905 ) | ( n14731 & 1'b0 ) | ( ~n14905 & 1'b0 ) ;
  assign n15301 = ( n14718 & n14727 ) | ( n14718 & n14731 ) | ( n14727 & n14731 ) ;
  assign n15302 = ( n15300 & ~n14727 ) | ( n15300 & n15301 ) | ( ~n14727 & n15301 ) ;
  assign n15303 = ( n14731 & ~n15301 ) | ( n14731 & n15300 ) | ( ~n15301 & n15300 ) ;
  assign n15304 = ( n14718 & ~n15302 ) | ( n14718 & n15303 ) | ( ~n15302 & n15303 ) ;
  assign n15305 = ( n1636 & ~n15277 ) | ( n1636 & 1'b0 ) | ( ~n15277 & 1'b0 ) ;
  assign n15306 = n15291 &  n15305 ;
  assign n15307 = n15297 | n15306 ;
  assign n15308 = ( n15285 & ~n15288 ) | ( n15285 & 1'b0 ) | ( ~n15288 & 1'b0 ) ;
  assign n15309 = ( n15282 & ~n1827 ) | ( n15282 & n15308 ) | ( ~n1827 & n15308 ) ;
  assign n15310 = n1636 | n15309 ;
  assign n15311 = n1452 &  n15310 ;
  assign n15312 = n15307 &  n15311 ;
  assign n15313 = n15304 | n15312 ;
  assign n15314 = n15299 &  n15313 ;
  assign n15315 = n14733 &  n14905 ;
  assign n15316 = ( n14725 & ~n14720 ) | ( n14725 & n14905 ) | ( ~n14720 & n14905 ) ;
  assign n15318 = ( n14720 & n15315 ) | ( n14720 & n15316 ) | ( n15315 & n15316 ) ;
  assign n15317 = ( n14905 & ~n15316 ) | ( n14905 & n15315 ) | ( ~n15316 & n15315 ) ;
  assign n15319 = ( n14725 & ~n15318 ) | ( n14725 & n15317 ) | ( ~n15318 & n15317 ) ;
  assign n15320 = ( n1283 & ~n15314 ) | ( n1283 & n15319 ) | ( ~n15314 & n15319 ) ;
  assign n15321 = ~n1122 & n15320 ;
  assign n15327 = ~n1283 & n15299 ;
  assign n15328 = n15313 &  n15327 ;
  assign n15329 = ( n15319 & ~n15328 ) | ( n15319 & 1'b0 ) | ( ~n15328 & 1'b0 ) ;
  assign n15330 = n15307 &  n15310 ;
  assign n15331 = ( n1452 & n15304 ) | ( n1452 & n15330 ) | ( n15304 & n15330 ) ;
  assign n15332 = ( n1283 & ~n15331 ) | ( n1283 & 1'b0 ) | ( ~n15331 & 1'b0 ) ;
  assign n15333 = ( n1122 & ~n15332 ) | ( n1122 & 1'b0 ) | ( ~n15332 & 1'b0 ) ;
  assign n15334 = ~n15329 & n15333 ;
  assign n15335 = n15326 | n15334 ;
  assign n15336 = ~n15321 & n15335 ;
  assign n15337 = ( n14742 & ~n14754 ) | ( n14742 & n14750 ) | ( ~n14754 & n14750 ) ;
  assign n15338 = ( n14750 & ~n15337 ) | ( n14750 & n14905 ) | ( ~n15337 & n14905 ) ;
  assign n15339 = ( n14905 & ~n14742 ) | ( n14905 & n15337 ) | ( ~n14742 & n15337 ) ;
  assign n15340 = ( n14754 & ~n15338 ) | ( n14754 & n15339 ) | ( ~n15338 & n15339 ) ;
  assign n15341 = ( n976 & n15336 ) | ( n976 & n15340 ) | ( n15336 & n15340 ) ;
  assign n15342 = ( n837 & ~n15341 ) | ( n837 & 1'b0 ) | ( ~n15341 & 1'b0 ) ;
  assign n15344 = ( n14770 & ~n14761 ) | ( n14770 & n14774 ) | ( ~n14761 & n14774 ) ;
  assign n15343 = ( n14774 & ~n14905 ) | ( n14774 & 1'b0 ) | ( ~n14905 & 1'b0 ) ;
  assign n15346 = ( n14774 & ~n15344 ) | ( n14774 & n15343 ) | ( ~n15344 & n15343 ) ;
  assign n15345 = ( n15343 & ~n14770 ) | ( n15343 & n15344 ) | ( ~n14770 & n15344 ) ;
  assign n15347 = ( n14761 & ~n15346 ) | ( n14761 & n15345 ) | ( ~n15346 & n15345 ) ;
  assign n15348 = ( n976 & ~n15321 ) | ( n976 & 1'b0 ) | ( ~n15321 & 1'b0 ) ;
  assign n15349 = n15335 &  n15348 ;
  assign n15350 = n15340 | n15349 ;
  assign n15351 = n15329 | n15332 ;
  assign n15352 = ( n1122 & ~n15351 ) | ( n1122 & n15326 ) | ( ~n15351 & n15326 ) ;
  assign n15353 = n976 | n15352 ;
  assign n15354 = ~n837 & n15353 ;
  assign n15355 = n15350 &  n15354 ;
  assign n15356 = ( n15347 & ~n15355 ) | ( n15347 & 1'b0 ) | ( ~n15355 & 1'b0 ) ;
  assign n15357 = n15342 | n15356 ;
  assign n15363 = ( n713 & ~n15362 ) | ( n713 & n15357 ) | ( ~n15362 & n15357 ) ;
  assign n15364 = n595 &  n15363 ;
  assign n15365 = n14796 | n14905 ;
  assign n15366 = ( n14783 & ~n14792 ) | ( n14783 & n14796 ) | ( ~n14792 & n14796 ) ;
  assign n15367 = ( n14792 & n15365 ) | ( n14792 & n15366 ) | ( n15365 & n15366 ) ;
  assign n15368 = ( n14796 & ~n15366 ) | ( n14796 & n15365 ) | ( ~n15366 & n15365 ) ;
  assign n15369 = ( n14783 & ~n15367 ) | ( n14783 & n15368 ) | ( ~n15367 & n15368 ) ;
  assign n15370 = n713 | n15342 ;
  assign n15371 = n15356 | n15370 ;
  assign n15372 = ~n15362 & n15371 ;
  assign n15373 = n15350 &  n15353 ;
  assign n15374 = ( n837 & ~n15373 ) | ( n837 & n15347 ) | ( ~n15373 & n15347 ) ;
  assign n15375 = n713 &  n15374 ;
  assign n15376 = n595 | n15375 ;
  assign n15377 = n15372 | n15376 ;
  assign n15378 = n15369 &  n15377 ;
  assign n15379 = n15364 | n15378 ;
  assign n15380 = ~n14798 & n14905 ;
  assign n15381 = ( n14785 & n14790 ) | ( n14785 & n14905 ) | ( n14790 & n14905 ) ;
  assign n15383 = ( n15380 & ~n14785 ) | ( n15380 & n15381 ) | ( ~n14785 & n15381 ) ;
  assign n15382 = ( n14905 & ~n15381 ) | ( n14905 & n15380 ) | ( ~n15381 & n15380 ) ;
  assign n15384 = ( n14790 & ~n15383 ) | ( n14790 & n15382 ) | ( ~n15383 & n15382 ) ;
  assign n15385 = ( n492 & n15379 ) | ( n492 & n15384 ) | ( n15379 & n15384 ) ;
  assign n15386 = n396 &  n15385 ;
  assign n15388 = ( n14814 & ~n14805 ) | ( n14814 & n14818 ) | ( ~n14805 & n14818 ) ;
  assign n15387 = n14818 | n14905 ;
  assign n15390 = ( n14818 & ~n15388 ) | ( n14818 & n15387 ) | ( ~n15388 & n15387 ) ;
  assign n15389 = ( n15387 & ~n14814 ) | ( n15387 & n15388 ) | ( ~n14814 & n15388 ) ;
  assign n15391 = ( n14805 & ~n15390 ) | ( n14805 & n15389 ) | ( ~n15390 & n15389 ) ;
  assign n15392 = n492 | n15364 ;
  assign n15393 = n15378 | n15392 ;
  assign n15394 = n15384 &  n15393 ;
  assign n15395 = n15372 | n15375 ;
  assign n15396 = ( n595 & n15369 ) | ( n595 & n15395 ) | ( n15369 & n15395 ) ;
  assign n15397 = n492 &  n15396 ;
  assign n15398 = n396 | n15397 ;
  assign n15399 = n15394 | n15398 ;
  assign n15400 = ~n15391 & n15399 ;
  assign n15401 = n15386 | n15400 ;
  assign n15403 = ( n14807 & ~n14812 ) | ( n14807 & n14905 ) | ( ~n14812 & n14905 ) ;
  assign n15402 = ~n14820 & n14905 ;
  assign n15404 = ( n14905 & ~n15403 ) | ( n14905 & n15402 ) | ( ~n15403 & n15402 ) ;
  assign n15405 = ( n15402 & ~n14807 ) | ( n15402 & n15403 ) | ( ~n14807 & n15403 ) ;
  assign n15406 = ( n14812 & ~n15404 ) | ( n14812 & n15405 ) | ( ~n15404 & n15405 ) ;
  assign n15407 = ( n315 & n15401 ) | ( n315 & n15406 ) | ( n15401 & n15406 ) ;
  assign n15408 = n240 &  n15407 ;
  assign n15410 = ( n14836 & ~n14827 ) | ( n14836 & n14840 ) | ( ~n14827 & n14840 ) ;
  assign n15409 = n14840 | n14905 ;
  assign n15412 = ( n14840 & ~n15410 ) | ( n14840 & n15409 ) | ( ~n15410 & n15409 ) ;
  assign n15411 = ( n15409 & ~n14836 ) | ( n15409 & n15410 ) | ( ~n14836 & n15410 ) ;
  assign n15413 = ( n14827 & ~n15412 ) | ( n14827 & n15411 ) | ( ~n15412 & n15411 ) ;
  assign n15414 = n315 | n15386 ;
  assign n15415 = n15400 | n15414 ;
  assign n15416 = n15406 &  n15415 ;
  assign n15417 = n15394 | n15397 ;
  assign n15418 = ( n396 & ~n15391 ) | ( n396 & n15417 ) | ( ~n15391 & n15417 ) ;
  assign n15419 = n315 &  n15418 ;
  assign n15420 = n240 | n15419 ;
  assign n15421 = n15416 | n15420 ;
  assign n15422 = ~n15413 & n15421 ;
  assign n15423 = n15408 | n15422 ;
  assign n15429 = ( n181 & ~n15428 ) | ( n181 & n15423 ) | ( ~n15428 & n15423 ) ;
  assign n15430 = ~n145 & n15429 ;
  assign n15432 = ( n14858 & ~n14849 ) | ( n14858 & n14862 ) | ( ~n14849 & n14862 ) ;
  assign n15431 = n14862 | n14905 ;
  assign n15434 = ( n14862 & ~n15432 ) | ( n14862 & n15431 ) | ( ~n15432 & n15431 ) ;
  assign n15433 = ( n15431 & ~n14858 ) | ( n15431 & n15432 ) | ( ~n14858 & n15432 ) ;
  assign n15435 = ( n14849 & ~n15434 ) | ( n14849 & n15433 ) | ( ~n15434 & n15433 ) ;
  assign n15436 = n181 | n15408 ;
  assign n15437 = n15422 | n15436 ;
  assign n15438 = ~n15428 & n15437 ;
  assign n15439 = n15416 | n15419 ;
  assign n15440 = ( n240 & ~n15413 ) | ( n240 & n15439 ) | ( ~n15413 & n15439 ) ;
  assign n15441 = n181 &  n15440 ;
  assign n15442 = ( n145 & ~n15441 ) | ( n145 & 1'b0 ) | ( ~n15441 & 1'b0 ) ;
  assign n15443 = ~n15438 & n15442 ;
  assign n15444 = ( n15435 & ~n15443 ) | ( n15435 & 1'b0 ) | ( ~n15443 & 1'b0 ) ;
  assign n15445 = n15430 | n15444 ;
  assign n15446 = n14851 | n14905 ;
  assign n15447 = ( n14856 & ~n14851 ) | ( n14856 & n14864 ) | ( ~n14851 & n14864 ) ;
  assign n15449 = ( n14851 & n15446 ) | ( n14851 & n15447 ) | ( n15446 & n15447 ) ;
  assign n15448 = ( n14864 & ~n15447 ) | ( n14864 & n15446 ) | ( ~n15447 & n15446 ) ;
  assign n15450 = ( n14856 & ~n15449 ) | ( n14856 & n15448 ) | ( ~n15449 & n15448 ) ;
  assign n15451 = ( n150 & n15445 ) | ( n150 & n15450 ) | ( n15445 & n15450 ) ;
  assign n15452 = n14871 &  n14887 ;
  assign n15453 = ( n14890 & n14905 ) | ( n14890 & n15452 ) | ( n14905 & n15452 ) ;
  assign n15454 = ~n14890 & n15453 ;
  assign n15455 = ( n14887 & ~n14890 ) | ( n14887 & 1'b0 ) | ( ~n14890 & 1'b0 ) ;
  assign n15456 = ~n14905 & n15455 ;
  assign n15457 = ( n14871 & ~n15456 ) | ( n14871 & n15455 ) | ( ~n15456 & n15455 ) ;
  assign n15458 = ~n15454 & n15457 ;
  assign n15459 = n14872 &  n14879 ;
  assign n15460 = ~n14905 & n15459 ;
  assign n15461 = ( n14893 & ~n15459 ) | ( n14893 & n15460 ) | ( ~n15459 & n15460 ) ;
  assign n15462 = ~n15458 & n15461 ;
  assign n15463 = ~n15451 & n15462 ;
  assign n15464 = ( n133 & ~n15463 ) | ( n133 & n15462 ) | ( ~n15463 & n15462 ) ;
  assign n15467 = n15438 | n15441 ;
  assign n15468 = ( n15435 & ~n145 ) | ( n15435 & n15467 ) | ( ~n145 & n15467 ) ;
  assign n15469 = n150 &  n15468 ;
  assign n15470 = ( n15458 & ~n15469 ) | ( n15458 & 1'b0 ) | ( ~n15469 & 1'b0 ) ;
  assign n15465 = n150 | n15430 ;
  assign n15466 = n15444 | n15465 ;
  assign n15471 = ( n15450 & ~n15466 ) | ( n15450 & 1'b0 ) | ( ~n15466 & 1'b0 ) ;
  assign n15472 = ( n15470 & ~n15450 ) | ( n15470 & n15471 ) | ( ~n15450 & n15471 ) ;
  assign n15474 = ( n133 & n14872 ) | ( n133 & n14879 ) | ( n14872 & n14879 ) ;
  assign n15473 = ( n14872 & ~n14905 ) | ( n14872 & n14879 ) | ( ~n14905 & n14879 ) ;
  assign n15475 = ( n14879 & ~n15473 ) | ( n14879 & 1'b0 ) | ( ~n15473 & 1'b0 ) ;
  assign n15476 = ( n15474 & ~n14879 ) | ( n15474 & n15475 ) | ( ~n14879 & n15475 ) ;
  assign n15477 = n14875 | n14902 ;
  assign n15478 = ( n14897 & ~n14878 ) | ( n14897 & n15477 ) | ( ~n14878 & n15477 ) ;
  assign n15479 = n14878 | n15478 ;
  assign n15480 = ( n14885 & ~n14893 ) | ( n14885 & n15479 ) | ( ~n14893 & n15479 ) ;
  assign n15481 = ( n14885 & ~n15480 ) | ( n14885 & 1'b0 ) | ( ~n15480 & 1'b0 ) ;
  assign n15482 = n15476 | n15481 ;
  assign n15483 = n15472 | n15482 ;
  assign n15484 = ~n15464 |  n15483 ;
  assign n15924 = ( n15321 & ~n15326 ) | ( n15321 & n15484 ) | ( ~n15326 & n15484 ) ;
  assign n15923 = n15334 &  n15484 ;
  assign n15925 = ( n15484 & ~n15924 ) | ( n15484 & n15923 ) | ( ~n15924 & n15923 ) ;
  assign n15926 = ( n15923 & ~n15321 ) | ( n15923 & n15924 ) | ( ~n15321 & n15924 ) ;
  assign n15927 = ( n15326 & ~n15925 ) | ( n15326 & n15926 ) | ( ~n15925 & n15926 ) ;
  assign n15908 = n15332 | n15484 ;
  assign n15909 = ( n15319 & ~n15328 ) | ( n15319 & n15332 ) | ( ~n15328 & n15332 ) ;
  assign n15910 = ( n15328 & n15908 ) | ( n15328 & n15909 ) | ( n15908 & n15909 ) ;
  assign n15911 = ( n15332 & ~n15909 ) | ( n15332 & n15908 ) | ( ~n15909 & n15908 ) ;
  assign n15912 = ( n15319 & ~n15910 ) | ( n15319 & n15911 ) | ( ~n15910 & n15911 ) ;
  assign n15901 = ( n15299 & ~n15484 ) | ( n15299 & 1'b0 ) | ( ~n15484 & 1'b0 ) ;
  assign n15902 = ( n15299 & n15304 ) | ( n15299 & n15312 ) | ( n15304 & n15312 ) ;
  assign n15903 = ( n15901 & ~n15312 ) | ( n15901 & n15902 ) | ( ~n15312 & n15902 ) ;
  assign n15904 = ( n15299 & ~n15902 ) | ( n15299 & n15901 ) | ( ~n15902 & n15901 ) ;
  assign n15905 = ( n15304 & ~n15903 ) | ( n15304 & n15904 ) | ( ~n15903 & n15904 ) ;
  assign n15887 = ( n15306 & ~n15297 ) | ( n15306 & n15310 ) | ( ~n15297 & n15310 ) ;
  assign n15886 = ( n15310 & ~n15484 ) | ( n15310 & 1'b0 ) | ( ~n15484 & 1'b0 ) ;
  assign n15889 = ( n15310 & ~n15887 ) | ( n15310 & n15886 ) | ( ~n15887 & n15886 ) ;
  assign n15888 = ( n15886 & ~n15306 ) | ( n15886 & n15887 ) | ( ~n15306 & n15887 ) ;
  assign n15890 = ( n15297 & ~n15889 ) | ( n15297 & n15888 ) | ( ~n15889 & n15888 ) ;
  assign n15879 = n15277 | n15484 ;
  assign n15880 = ( n15282 & ~n15277 ) | ( n15282 & n15290 ) | ( ~n15277 & n15290 ) ;
  assign n15882 = ( n15277 & n15879 ) | ( n15277 & n15880 ) | ( n15879 & n15880 ) ;
  assign n15881 = ( n15290 & ~n15880 ) | ( n15290 & n15879 ) | ( ~n15880 & n15879 ) ;
  assign n15883 = ( n15282 & ~n15882 ) | ( n15282 & n15881 ) | ( ~n15882 & n15881 ) ;
  assign n15864 = n15288 | n15484 ;
  assign n15865 = ( n15275 & ~n15284 ) | ( n15275 & n15288 ) | ( ~n15284 & n15288 ) ;
  assign n15866 = ( n15284 & n15864 ) | ( n15284 & n15865 ) | ( n15864 & n15865 ) ;
  assign n15867 = ( n15288 & ~n15865 ) | ( n15288 & n15864 ) | ( ~n15865 & n15864 ) ;
  assign n15868 = ( n15275 & ~n15866 ) | ( n15275 & n15867 ) | ( ~n15866 & n15867 ) ;
  assign n15858 = ( n15255 & ~n15260 ) | ( n15255 & n15268 ) | ( ~n15260 & n15268 ) ;
  assign n15857 = n15255 | n15484 ;
  assign n15860 = ( n15255 & ~n15858 ) | ( n15255 & n15857 ) | ( ~n15858 & n15857 ) ;
  assign n15859 = ( n15857 & ~n15268 ) | ( n15857 & n15858 ) | ( ~n15268 & n15858 ) ;
  assign n15861 = ( n15260 & ~n15860 ) | ( n15260 & n15859 ) | ( ~n15860 & n15859 ) ;
  assign n15843 = ( n15262 & ~n15253 ) | ( n15262 & n15266 ) | ( ~n15253 & n15266 ) ;
  assign n15842 = n15266 | n15484 ;
  assign n15845 = ( n15266 & ~n15843 ) | ( n15266 & n15842 ) | ( ~n15843 & n15842 ) ;
  assign n15844 = ( n15842 & ~n15262 ) | ( n15842 & n15843 ) | ( ~n15262 & n15843 ) ;
  assign n15846 = ( n15253 & ~n15845 ) | ( n15253 & n15844 ) | ( ~n15845 & n15844 ) ;
  assign n15835 = n15233 | n15484 ;
  assign n15836 = ( n15233 & n15238 ) | ( n15233 & n15246 ) | ( n15238 & n15246 ) ;
  assign n15837 = ( n15835 & ~n15246 ) | ( n15835 & n15836 ) | ( ~n15246 & n15836 ) ;
  assign n15838 = ( n15233 & ~n15836 ) | ( n15233 & n15835 ) | ( ~n15836 & n15835 ) ;
  assign n15839 = ( n15238 & ~n15837 ) | ( n15238 & n15838 ) | ( ~n15837 & n15838 ) ;
  assign n15820 = n15244 | n15484 ;
  assign n15821 = ( n15231 & n15240 ) | ( n15231 & n15244 ) | ( n15240 & n15244 ) ;
  assign n15822 = ( n15820 & ~n15240 ) | ( n15820 & n15821 ) | ( ~n15240 & n15821 ) ;
  assign n15823 = ( n15244 & ~n15821 ) | ( n15244 & n15820 ) | ( ~n15821 & n15820 ) ;
  assign n15824 = ( n15231 & ~n15822 ) | ( n15231 & n15823 ) | ( ~n15822 & n15823 ) ;
  assign n15813 = n15211 | n15484 ;
  assign n15814 = ( n15211 & n15216 ) | ( n15211 & n15224 ) | ( n15216 & n15224 ) ;
  assign n15815 = ( n15813 & ~n15224 ) | ( n15813 & n15814 ) | ( ~n15224 & n15814 ) ;
  assign n15816 = ( n15211 & ~n15814 ) | ( n15211 & n15813 ) | ( ~n15814 & n15813 ) ;
  assign n15817 = ( n15216 & ~n15815 ) | ( n15216 & n15816 ) | ( ~n15815 & n15816 ) ;
  assign n15798 = n15222 | n15484 ;
  assign n15799 = ( n15209 & n15218 ) | ( n15209 & n15222 ) | ( n15218 & n15222 ) ;
  assign n15800 = ( n15798 & ~n15218 ) | ( n15798 & n15799 ) | ( ~n15218 & n15799 ) ;
  assign n15801 = ( n15222 & ~n15799 ) | ( n15222 & n15798 ) | ( ~n15799 & n15798 ) ;
  assign n15802 = ( n15209 & ~n15800 ) | ( n15209 & n15801 ) | ( ~n15800 & n15801 ) ;
  assign n15792 = ( n15189 & ~n15194 ) | ( n15189 & n15202 ) | ( ~n15194 & n15202 ) ;
  assign n15791 = n15189 | n15484 ;
  assign n15794 = ( n15189 & ~n15792 ) | ( n15189 & n15791 ) | ( ~n15792 & n15791 ) ;
  assign n15793 = ( n15791 & ~n15202 ) | ( n15791 & n15792 ) | ( ~n15202 & n15792 ) ;
  assign n15795 = ( n15194 & ~n15794 ) | ( n15194 & n15793 ) | ( ~n15794 & n15793 ) ;
  assign n15777 = ( n15196 & ~n15187 ) | ( n15196 & n15200 ) | ( ~n15187 & n15200 ) ;
  assign n15776 = n15200 | n15484 ;
  assign n15779 = ( n15200 & ~n15777 ) | ( n15200 & n15776 ) | ( ~n15777 & n15776 ) ;
  assign n15778 = ( n15776 & ~n15196 ) | ( n15776 & n15777 ) | ( ~n15196 & n15777 ) ;
  assign n15780 = ( n15187 & ~n15779 ) | ( n15187 & n15778 ) | ( ~n15779 & n15778 ) ;
  assign n15769 = n15167 | n15484 ;
  assign n15770 = ( n15167 & n15172 ) | ( n15167 & n15180 ) | ( n15172 & n15180 ) ;
  assign n15771 = ( n15769 & ~n15180 ) | ( n15769 & n15770 ) | ( ~n15180 & n15770 ) ;
  assign n15772 = ( n15167 & ~n15770 ) | ( n15167 & n15769 ) | ( ~n15770 & n15769 ) ;
  assign n15773 = ( n15172 & ~n15771 ) | ( n15172 & n15772 ) | ( ~n15771 & n15772 ) ;
  assign n15755 = ( n15174 & ~n15165 ) | ( n15174 & n15178 ) | ( ~n15165 & n15178 ) ;
  assign n15754 = n15178 | n15484 ;
  assign n15757 = ( n15178 & ~n15755 ) | ( n15178 & n15754 ) | ( ~n15755 & n15754 ) ;
  assign n15756 = ( n15754 & ~n15174 ) | ( n15754 & n15755 ) | ( ~n15174 & n15755 ) ;
  assign n15758 = ( n15165 & ~n15757 ) | ( n15165 & n15756 ) | ( ~n15757 & n15756 ) ;
  assign n15747 = n15145 | n15484 ;
  assign n15748 = ( n15145 & n15150 ) | ( n15145 & n15158 ) | ( n15150 & n15158 ) ;
  assign n15749 = ( n15747 & ~n15158 ) | ( n15747 & n15748 ) | ( ~n15158 & n15748 ) ;
  assign n15750 = ( n15145 & ~n15748 ) | ( n15145 & n15747 ) | ( ~n15748 & n15747 ) ;
  assign n15751 = ( n15150 & ~n15749 ) | ( n15150 & n15750 ) | ( ~n15749 & n15750 ) ;
  assign n15732 = n15156 | n15484 ;
  assign n15733 = ( n15143 & ~n15156 ) | ( n15143 & n15152 ) | ( ~n15156 & n15152 ) ;
  assign n15735 = ( n15156 & n15732 ) | ( n15156 & n15733 ) | ( n15732 & n15733 ) ;
  assign n15734 = ( n15152 & ~n15733 ) | ( n15152 & n15732 ) | ( ~n15733 & n15732 ) ;
  assign n15736 = ( n15143 & ~n15735 ) | ( n15143 & n15734 ) | ( ~n15735 & n15734 ) ;
  assign n15725 = ( n15123 & ~n15484 ) | ( n15123 & 1'b0 ) | ( ~n15484 & 1'b0 ) ;
  assign n15726 = ( n15123 & n15128 ) | ( n15123 & n15136 ) | ( n15128 & n15136 ) ;
  assign n15727 = ( n15725 & ~n15136 ) | ( n15725 & n15726 ) | ( ~n15136 & n15726 ) ;
  assign n15728 = ( n15123 & ~n15726 ) | ( n15123 & n15725 ) | ( ~n15726 & n15725 ) ;
  assign n15729 = ( n15128 & ~n15727 ) | ( n15128 & n15728 ) | ( ~n15727 & n15728 ) ;
  assign n15710 = n15134 | n15484 ;
  assign n15711 = ( n15121 & ~n15130 ) | ( n15121 & n15134 ) | ( ~n15130 & n15134 ) ;
  assign n15712 = ( n15130 & n15710 ) | ( n15130 & n15711 ) | ( n15710 & n15711 ) ;
  assign n15713 = ( n15134 & ~n15711 ) | ( n15134 & n15710 ) | ( ~n15711 & n15710 ) ;
  assign n15714 = ( n15121 & ~n15712 ) | ( n15121 & n15713 ) | ( ~n15712 & n15713 ) ;
  assign n15703 = ( n15101 & ~n15484 ) | ( n15101 & 1'b0 ) | ( ~n15484 & 1'b0 ) ;
  assign n15704 = ( n15101 & n15106 ) | ( n15101 & n15114 ) | ( n15106 & n15114 ) ;
  assign n15705 = ( n15703 & ~n15114 ) | ( n15703 & n15704 ) | ( ~n15114 & n15704 ) ;
  assign n15706 = ( n15101 & ~n15704 ) | ( n15101 & n15703 ) | ( ~n15704 & n15703 ) ;
  assign n15707 = ( n15106 & ~n15705 ) | ( n15106 & n15706 ) | ( ~n15705 & n15706 ) ;
  assign n15688 = n15112 | n15484 ;
  assign n15689 = ( n15099 & ~n15108 ) | ( n15099 & n15112 ) | ( ~n15108 & n15112 ) ;
  assign n15690 = ( n15108 & n15688 ) | ( n15108 & n15689 ) | ( n15688 & n15689 ) ;
  assign n15691 = ( n15112 & ~n15689 ) | ( n15112 & n15688 ) | ( ~n15689 & n15688 ) ;
  assign n15692 = ( n15099 & ~n15690 ) | ( n15099 & n15691 ) | ( ~n15690 & n15691 ) ;
  assign n15681 = ( n15079 & ~n15484 ) | ( n15079 & 1'b0 ) | ( ~n15484 & 1'b0 ) ;
  assign n15682 = ( n15079 & n15084 ) | ( n15079 & n15092 ) | ( n15084 & n15092 ) ;
  assign n15683 = ( n15681 & ~n15092 ) | ( n15681 & n15682 ) | ( ~n15092 & n15682 ) ;
  assign n15684 = ( n15079 & ~n15682 ) | ( n15079 & n15681 ) | ( ~n15682 & n15681 ) ;
  assign n15685 = ( n15084 & ~n15683 ) | ( n15084 & n15684 ) | ( ~n15683 & n15684 ) ;
  assign n15667 = ( n15086 & ~n15077 ) | ( n15086 & n15090 ) | ( ~n15077 & n15090 ) ;
  assign n15666 = ( n15090 & ~n15484 ) | ( n15090 & 1'b0 ) | ( ~n15484 & 1'b0 ) ;
  assign n15669 = ( n15090 & ~n15667 ) | ( n15090 & n15666 ) | ( ~n15667 & n15666 ) ;
  assign n15668 = ( n15666 & ~n15086 ) | ( n15666 & n15667 ) | ( ~n15086 & n15667 ) ;
  assign n15670 = ( n15077 & ~n15669 ) | ( n15077 & n15668 ) | ( ~n15669 & n15668 ) ;
  assign n15659 = n15057 | n15484 ;
  assign n15660 = ( n15062 & ~n15057 ) | ( n15062 & n15070 ) | ( ~n15057 & n15070 ) ;
  assign n15662 = ( n15057 & n15659 ) | ( n15057 & n15660 ) | ( n15659 & n15660 ) ;
  assign n15661 = ( n15070 & ~n15660 ) | ( n15070 & n15659 ) | ( ~n15660 & n15659 ) ;
  assign n15663 = ( n15062 & ~n15662 ) | ( n15062 & n15661 ) | ( ~n15662 & n15661 ) ;
  assign n15644 = n15068 | n15484 ;
  assign n15645 = ( n15055 & ~n15068 ) | ( n15055 & n15064 ) | ( ~n15068 & n15064 ) ;
  assign n15647 = ( n15068 & n15644 ) | ( n15068 & n15645 ) | ( n15644 & n15645 ) ;
  assign n15646 = ( n15064 & ~n15645 ) | ( n15064 & n15644 ) | ( ~n15645 & n15644 ) ;
  assign n15648 = ( n15055 & ~n15647 ) | ( n15055 & n15646 ) | ( ~n15647 & n15646 ) ;
  assign n15637 = n15035 | n15484 ;
  assign n15638 = ( n15035 & ~n15048 ) | ( n15035 & n15040 ) | ( ~n15048 & n15040 ) ;
  assign n15639 = ( n15048 & n15637 ) | ( n15048 & n15638 ) | ( n15637 & n15638 ) ;
  assign n15640 = ( n15035 & ~n15638 ) | ( n15035 & n15637 ) | ( ~n15638 & n15637 ) ;
  assign n15641 = ( n15040 & ~n15639 ) | ( n15040 & n15640 ) | ( ~n15639 & n15640 ) ;
  assign n15622 = n15046 | n15484 ;
  assign n15623 = ( n15033 & ~n15042 ) | ( n15033 & n15046 ) | ( ~n15042 & n15046 ) ;
  assign n15624 = ( n15042 & n15622 ) | ( n15042 & n15623 ) | ( n15622 & n15623 ) ;
  assign n15625 = ( n15046 & ~n15623 ) | ( n15046 & n15622 ) | ( ~n15623 & n15622 ) ;
  assign n15626 = ( n15033 & ~n15624 ) | ( n15033 & n15625 ) | ( ~n15624 & n15625 ) ;
  assign n15615 = ( n15013 & ~n15484 ) | ( n15013 & 1'b0 ) | ( ~n15484 & 1'b0 ) ;
  assign n15616 = ( n15013 & n15018 ) | ( n15013 & n15026 ) | ( n15018 & n15026 ) ;
  assign n15617 = ( n15615 & ~n15026 ) | ( n15615 & n15616 ) | ( ~n15026 & n15616 ) ;
  assign n15618 = ( n15013 & ~n15616 ) | ( n15013 & n15615 ) | ( ~n15616 & n15615 ) ;
  assign n15619 = ( n15018 & ~n15617 ) | ( n15018 & n15618 ) | ( ~n15617 & n15618 ) ;
  assign n15600 = n15024 | n15484 ;
  assign n15601 = ( n15011 & ~n15020 ) | ( n15011 & n15024 ) | ( ~n15020 & n15024 ) ;
  assign n15602 = ( n15020 & n15600 ) | ( n15020 & n15601 ) | ( n15600 & n15601 ) ;
  assign n15603 = ( n15024 & ~n15601 ) | ( n15024 & n15600 ) | ( ~n15601 & n15600 ) ;
  assign n15604 = ( n15011 & ~n15602 ) | ( n15011 & n15603 ) | ( ~n15602 & n15603 ) ;
  assign n15593 = n15004 &  n15484 ;
  assign n15594 = ( n14991 & n14996 ) | ( n14991 & n15484 ) | ( n14996 & n15484 ) ;
  assign n15596 = ( n15593 & ~n14991 ) | ( n15593 & n15594 ) | ( ~n14991 & n15594 ) ;
  assign n15595 = ( n15484 & ~n15594 ) | ( n15484 & n15593 ) | ( ~n15594 & n15593 ) ;
  assign n15597 = ( n14996 & ~n15596 ) | ( n14996 & n15595 ) | ( ~n15596 & n15595 ) ;
  assign n15578 = n15002 | n15484 ;
  assign n15579 = ( n14989 & ~n15002 ) | ( n14989 & n14998 ) | ( ~n15002 & n14998 ) ;
  assign n15581 = ( n15002 & n15578 ) | ( n15002 & n15579 ) | ( n15578 & n15579 ) ;
  assign n15580 = ( n14998 & ~n15579 ) | ( n14998 & n15578 ) | ( ~n15579 & n15578 ) ;
  assign n15582 = ( n14989 & ~n15581 ) | ( n14989 & n15580 ) | ( ~n15581 & n15580 ) ;
  assign n15571 = n14969 | n15484 ;
  assign n15572 = ( n14969 & ~n14982 ) | ( n14969 & n14974 ) | ( ~n14982 & n14974 ) ;
  assign n15573 = ( n14982 & n15571 ) | ( n14982 & n15572 ) | ( n15571 & n15572 ) ;
  assign n15574 = ( n14969 & ~n15572 ) | ( n14969 & n15571 ) | ( ~n15572 & n15571 ) ;
  assign n15575 = ( n14974 & ~n15573 ) | ( n14974 & n15574 ) | ( ~n15573 & n15574 ) ;
  assign n15556 = n14980 | n15484 ;
  assign n15557 = ( n14967 & ~n14976 ) | ( n14967 & n14980 ) | ( ~n14976 & n14980 ) ;
  assign n15558 = ( n14976 & n15556 ) | ( n14976 & n15557 ) | ( n15556 & n15557 ) ;
  assign n15559 = ( n14980 & ~n15557 ) | ( n14980 & n15556 ) | ( ~n15557 & n15556 ) ;
  assign n15560 = ( n14967 & ~n15558 ) | ( n14967 & n15559 ) | ( ~n15558 & n15559 ) ;
  assign n15549 = n14947 | n15484 ;
  assign n15550 = ( n14952 & ~n14947 ) | ( n14952 & n14960 ) | ( ~n14947 & n14960 ) ;
  assign n15552 = ( n14947 & n15549 ) | ( n14947 & n15550 ) | ( n15549 & n15550 ) ;
  assign n15551 = ( n14960 & ~n15550 ) | ( n14960 & n15549 ) | ( ~n15550 & n15549 ) ;
  assign n15553 = ( n14952 & ~n15552 ) | ( n14952 & n15551 ) | ( ~n15552 & n15551 ) ;
  assign n15534 = n14958 | n15484 ;
  assign n15535 = ( n14945 & ~n14954 ) | ( n14945 & n14958 ) | ( ~n14954 & n14958 ) ;
  assign n15536 = ( n14954 & n15534 ) | ( n14954 & n15535 ) | ( n15534 & n15535 ) ;
  assign n15537 = ( n14958 & ~n15535 ) | ( n14958 & n15534 ) | ( ~n15535 & n15534 ) ;
  assign n15538 = ( n14945 & ~n15536 ) | ( n14945 & n15537 ) | ( ~n15536 & n15537 ) ;
  assign n15527 = ( n14921 & ~n14923 ) | ( n14921 & 1'b0 ) | ( ~n14923 & 1'b0 ) ;
  assign n15528 = ( n14923 & ~n15527 ) | ( n14923 & n14933 ) | ( ~n15527 & n14933 ) ;
  assign n15530 = ( n15484 & n15527 ) | ( n15484 & n15528 ) | ( n15527 & n15528 ) ;
  assign n15529 = ( n14923 & ~n15528 ) | ( n14923 & n15484 ) | ( ~n15528 & n15484 ) ;
  assign n15531 = ( n14933 & ~n15530 ) | ( n14933 & n15529 ) | ( ~n15530 & n15529 ) ;
  assign n15511 = ~x26 & n14905 ;
  assign n15512 = ( x27 & ~n15511 ) | ( x27 & 1'b0 ) | ( ~n15511 & 1'b0 ) ;
  assign n15513 = n14924 | n15512 ;
  assign n15508 = ( n14905 & ~x26 ) | ( n14905 & n14916 ) | ( ~x26 & n14916 ) ;
  assign n15509 = x26 &  n15508 ;
  assign n15510 = ( n14911 & ~n15509 ) | ( n14911 & n14916 ) | ( ~n15509 & n14916 ) ;
  assign n15514 = ( n15484 & ~n15513 ) | ( n15484 & n15510 ) | ( ~n15513 & n15510 ) ;
  assign n15516 = ( n15484 & ~n15514 ) | ( n15484 & 1'b0 ) | ( ~n15514 & 1'b0 ) ;
  assign n15515 = ~n15510 & n15514 ;
  assign n15517 = ( n15513 & ~n15516 ) | ( n15513 & n15515 ) | ( ~n15516 & n15515 ) ;
  assign n15497 = ( n14905 & ~n15481 ) | ( n14905 & 1'b0 ) | ( ~n15481 & 1'b0 ) ;
  assign n15498 = ( n15472 & ~n15476 ) | ( n15472 & n15497 ) | ( ~n15476 & n15497 ) ;
  assign n15499 = ~n15472 & n15498 ;
  assign n15500 = n15464 &  n15499 ;
  assign n15496 = ~n14908 & n15484 ;
  assign n15501 = ( n15496 & ~n15500 ) | ( n15496 & 1'b0 ) | ( ~n15500 & 1'b0 ) ;
  assign n15502 = ( x26 & n15500 ) | ( x26 & n15501 ) | ( n15500 & n15501 ) ;
  assign n15503 = x26 | n15500 ;
  assign n15504 = n15496 | n15503 ;
  assign n15505 = ~n15502 & n15504 ;
  assign n15487 = ( x24 & ~n15484 ) | ( x24 & x25 ) | ( ~n15484 & x25 ) ;
  assign n15493 = ( x24 & ~x25 ) | ( x24 & 1'b0 ) | ( ~x25 & 1'b0 ) ;
  assign n14906 = x22 | x23 ;
  assign n15488 = ~x24 & n14906 ;
  assign n15489 = ( x24 & ~n14903 ) | ( x24 & n15488 ) | ( ~n14903 & n15488 ) ;
  assign n15490 = ( n14893 & ~n14885 ) | ( n14893 & n15489 ) | ( ~n14885 & n15489 ) ;
  assign n15491 = n14885 &  n15490 ;
  assign n15492 = ( n15484 & ~x25 ) | ( n15484 & n15491 ) | ( ~x25 & n15491 ) ;
  assign n15494 = ( n15487 & ~n15493 ) | ( n15487 & n15492 ) | ( ~n15493 & n15492 ) ;
  assign n14907 = x24 | n14906 ;
  assign n15485 = x24 &  n15484 ;
  assign n15486 = ( n14905 & ~n14907 ) | ( n14905 & n15485 ) | ( ~n14907 & n15485 ) ;
  assign n15518 = n14341 | n15486 ;
  assign n15519 = ( n15494 & ~n15518 ) | ( n15494 & 1'b0 ) | ( ~n15518 & 1'b0 ) ;
  assign n15520 = n15505 | n15519 ;
  assign n15521 = n15486 &  n15494 ;
  assign n15522 = ( n14341 & ~n15494 ) | ( n14341 & n15521 ) | ( ~n15494 & n15521 ) ;
  assign n15523 = n13784 | n15522 ;
  assign n15524 = ( n15520 & ~n15523 ) | ( n15520 & 1'b0 ) | ( ~n15523 & 1'b0 ) ;
  assign n15525 = n15517 | n15524 ;
  assign n15495 = ~n15486 & n15494 ;
  assign n15506 = ( n15495 & ~n14341 ) | ( n15495 & n15505 ) | ( ~n14341 & n15505 ) ;
  assign n15507 = ( n13784 & ~n15506 ) | ( n13784 & 1'b0 ) | ( ~n15506 & 1'b0 ) ;
  assign n15539 = n13242 | n15507 ;
  assign n15540 = ( n15525 & ~n15539 ) | ( n15525 & 1'b0 ) | ( ~n15539 & 1'b0 ) ;
  assign n15541 = n15531 | n15540 ;
  assign n15542 = ( n15520 & ~n15522 ) | ( n15520 & 1'b0 ) | ( ~n15522 & 1'b0 ) ;
  assign n15543 = ( n15517 & ~n13784 ) | ( n15517 & n15542 ) | ( ~n13784 & n15542 ) ;
  assign n15544 = ( n13242 & ~n15543 ) | ( n13242 & 1'b0 ) | ( ~n15543 & 1'b0 ) ;
  assign n15545 = n12707 | n15544 ;
  assign n15546 = ( n15541 & ~n15545 ) | ( n15541 & 1'b0 ) | ( ~n15545 & 1'b0 ) ;
  assign n15547 = n15538 | n15546 ;
  assign n15526 = ~n15507 & n15525 ;
  assign n15532 = ( n15526 & ~n13242 ) | ( n15526 & n15531 ) | ( ~n13242 & n15531 ) ;
  assign n15533 = ( n12707 & ~n15532 ) | ( n12707 & 1'b0 ) | ( ~n15532 & 1'b0 ) ;
  assign n15561 = n12187 | n15533 ;
  assign n15562 = ( n15547 & ~n15561 ) | ( n15547 & 1'b0 ) | ( ~n15561 & 1'b0 ) ;
  assign n15563 = n15553 | n15562 ;
  assign n15564 = ( n15541 & ~n15544 ) | ( n15541 & 1'b0 ) | ( ~n15544 & 1'b0 ) ;
  assign n15565 = ( n15538 & ~n12707 ) | ( n15538 & n15564 ) | ( ~n12707 & n15564 ) ;
  assign n15566 = ( n12187 & ~n15565 ) | ( n12187 & 1'b0 ) | ( ~n15565 & 1'b0 ) ;
  assign n15567 = n11674 | n15566 ;
  assign n15568 = ( n15563 & ~n15567 ) | ( n15563 & 1'b0 ) | ( ~n15567 & 1'b0 ) ;
  assign n15569 = n15560 | n15568 ;
  assign n15548 = ~n15533 & n15547 ;
  assign n15554 = ( n15548 & ~n12187 ) | ( n15548 & n15553 ) | ( ~n12187 & n15553 ) ;
  assign n15555 = ( n11674 & ~n15554 ) | ( n11674 & 1'b0 ) | ( ~n15554 & 1'b0 ) ;
  assign n15583 = n11176 | n15555 ;
  assign n15584 = ( n15569 & ~n15583 ) | ( n15569 & 1'b0 ) | ( ~n15583 & 1'b0 ) ;
  assign n15585 = n15575 | n15584 ;
  assign n15586 = ( n15563 & ~n15566 ) | ( n15563 & 1'b0 ) | ( ~n15566 & 1'b0 ) ;
  assign n15587 = ( n15560 & ~n11674 ) | ( n15560 & n15586 ) | ( ~n11674 & n15586 ) ;
  assign n15588 = ( n11176 & ~n15587 ) | ( n11176 & 1'b0 ) | ( ~n15587 & 1'b0 ) ;
  assign n15589 = n10685 | n15588 ;
  assign n15590 = ( n15585 & ~n15589 ) | ( n15585 & 1'b0 ) | ( ~n15589 & 1'b0 ) ;
  assign n15591 = n15582 | n15590 ;
  assign n15570 = ~n15555 & n15569 ;
  assign n15576 = ( n15570 & ~n11176 ) | ( n15570 & n15575 ) | ( ~n11176 & n15575 ) ;
  assign n15577 = ( n10685 & ~n15576 ) | ( n10685 & 1'b0 ) | ( ~n15576 & 1'b0 ) ;
  assign n15605 = n10209 | n15577 ;
  assign n15606 = ( n15591 & ~n15605 ) | ( n15591 & 1'b0 ) | ( ~n15605 & 1'b0 ) ;
  assign n15607 = n15597 | n15606 ;
  assign n15608 = ( n15585 & ~n15588 ) | ( n15585 & 1'b0 ) | ( ~n15588 & 1'b0 ) ;
  assign n15609 = ( n15582 & ~n10685 ) | ( n15582 & n15608 ) | ( ~n10685 & n15608 ) ;
  assign n15610 = ( n10209 & ~n15609 ) | ( n10209 & 1'b0 ) | ( ~n15609 & 1'b0 ) ;
  assign n15611 = ( n9740 & ~n15610 ) | ( n9740 & 1'b0 ) | ( ~n15610 & 1'b0 ) ;
  assign n15612 = n15607 &  n15611 ;
  assign n15613 = n15604 | n15612 ;
  assign n15592 = ~n15577 & n15591 ;
  assign n15598 = ( n15592 & ~n10209 ) | ( n15592 & n15597 ) | ( ~n10209 & n15597 ) ;
  assign n15599 = n9740 | n15598 ;
  assign n15627 = ~n9286 & n15599 ;
  assign n15628 = n15613 &  n15627 ;
  assign n15629 = n15619 | n15628 ;
  assign n15630 = ( n15607 & ~n15610 ) | ( n15607 & 1'b0 ) | ( ~n15610 & 1'b0 ) ;
  assign n15631 = ( n9740 & n15604 ) | ( n9740 & n15630 ) | ( n15604 & n15630 ) ;
  assign n15632 = ( n9286 & ~n15631 ) | ( n9286 & 1'b0 ) | ( ~n15631 & 1'b0 ) ;
  assign n15633 = n8839 | n15632 ;
  assign n15634 = ( n15629 & ~n15633 ) | ( n15629 & 1'b0 ) | ( ~n15633 & 1'b0 ) ;
  assign n15635 = n15626 | n15634 ;
  assign n15614 = n15599 &  n15613 ;
  assign n15620 = ( n15614 & ~n9286 ) | ( n15614 & n15619 ) | ( ~n9286 & n15619 ) ;
  assign n15621 = ( n8839 & ~n15620 ) | ( n8839 & 1'b0 ) | ( ~n15620 & 1'b0 ) ;
  assign n15649 = n8407 | n15621 ;
  assign n15650 = ( n15635 & ~n15649 ) | ( n15635 & 1'b0 ) | ( ~n15649 & 1'b0 ) ;
  assign n15651 = n15641 | n15650 ;
  assign n15652 = ( n15629 & ~n15632 ) | ( n15629 & 1'b0 ) | ( ~n15632 & 1'b0 ) ;
  assign n15653 = ( n15626 & ~n8839 ) | ( n15626 & n15652 ) | ( ~n8839 & n15652 ) ;
  assign n15654 = ( n8407 & ~n15653 ) | ( n8407 & 1'b0 ) | ( ~n15653 & 1'b0 ) ;
  assign n15655 = n7982 | n15654 ;
  assign n15656 = ( n15651 & ~n15655 ) | ( n15651 & 1'b0 ) | ( ~n15655 & 1'b0 ) ;
  assign n15657 = n15648 | n15656 ;
  assign n15636 = ~n15621 & n15635 ;
  assign n15642 = ( n15636 & ~n8407 ) | ( n15636 & n15641 ) | ( ~n8407 & n15641 ) ;
  assign n15643 = ( n7982 & ~n15642 ) | ( n7982 & 1'b0 ) | ( ~n15642 & 1'b0 ) ;
  assign n15671 = ( n7572 & ~n15643 ) | ( n7572 & 1'b0 ) | ( ~n15643 & 1'b0 ) ;
  assign n15672 = n15657 &  n15671 ;
  assign n15673 = n15663 | n15672 ;
  assign n15674 = ( n15651 & ~n15654 ) | ( n15651 & 1'b0 ) | ( ~n15654 & 1'b0 ) ;
  assign n15675 = ( n15648 & ~n7982 ) | ( n15648 & n15674 ) | ( ~n7982 & n15674 ) ;
  assign n15676 = n7572 | n15675 ;
  assign n15677 = n7169 &  n15676 ;
  assign n15678 = n15673 &  n15677 ;
  assign n15679 = n15670 | n15678 ;
  assign n15658 = ~n15643 & n15657 ;
  assign n15664 = ( n7572 & n15658 ) | ( n7572 & n15663 ) | ( n15658 & n15663 ) ;
  assign n15665 = n7169 | n15664 ;
  assign n15693 = ~n6781 & n15665 ;
  assign n15694 = n15679 &  n15693 ;
  assign n15695 = n15685 | n15694 ;
  assign n15696 = n15673 &  n15676 ;
  assign n15697 = ( n7169 & n15670 ) | ( n7169 & n15696 ) | ( n15670 & n15696 ) ;
  assign n15698 = ( n6781 & ~n15697 ) | ( n6781 & 1'b0 ) | ( ~n15697 & 1'b0 ) ;
  assign n15699 = ( n6399 & ~n15698 ) | ( n6399 & 1'b0 ) | ( ~n15698 & 1'b0 ) ;
  assign n15700 = n15695 &  n15699 ;
  assign n15701 = n15692 | n15700 ;
  assign n15680 = n15665 &  n15679 ;
  assign n15686 = ( n15680 & ~n6781 ) | ( n15680 & n15685 ) | ( ~n6781 & n15685 ) ;
  assign n15687 = n6399 | n15686 ;
  assign n15715 = ~n6032 & n15687 ;
  assign n15716 = n15701 &  n15715 ;
  assign n15717 = n15707 | n15716 ;
  assign n15718 = ( n15695 & ~n15698 ) | ( n15695 & 1'b0 ) | ( ~n15698 & 1'b0 ) ;
  assign n15719 = ( n6399 & n15692 ) | ( n6399 & n15718 ) | ( n15692 & n15718 ) ;
  assign n15720 = ( n6032 & ~n15719 ) | ( n6032 & 1'b0 ) | ( ~n15719 & 1'b0 ) ;
  assign n15721 = ( n5672 & ~n15720 ) | ( n5672 & 1'b0 ) | ( ~n15720 & 1'b0 ) ;
  assign n15722 = n15717 &  n15721 ;
  assign n15723 = n15714 | n15722 ;
  assign n15702 = n15687 &  n15701 ;
  assign n15708 = ( n15702 & ~n6032 ) | ( n15702 & n15707 ) | ( ~n6032 & n15707 ) ;
  assign n15709 = n5672 | n15708 ;
  assign n15737 = ~n5327 & n15709 ;
  assign n15738 = n15723 &  n15737 ;
  assign n15739 = n15729 | n15738 ;
  assign n15740 = ( n15717 & ~n15720 ) | ( n15717 & 1'b0 ) | ( ~n15720 & 1'b0 ) ;
  assign n15741 = ( n5672 & n15714 ) | ( n5672 & n15740 ) | ( n15714 & n15740 ) ;
  assign n15742 = ( n5327 & ~n15741 ) | ( n5327 & 1'b0 ) | ( ~n15741 & 1'b0 ) ;
  assign n15743 = n4990 | n15742 ;
  assign n15744 = ( n15739 & ~n15743 ) | ( n15739 & 1'b0 ) | ( ~n15743 & 1'b0 ) ;
  assign n15745 = ( n15736 & ~n15744 ) | ( n15736 & 1'b0 ) | ( ~n15744 & 1'b0 ) ;
  assign n15724 = n15709 &  n15723 ;
  assign n15730 = ( n15724 & ~n5327 ) | ( n15724 & n15729 ) | ( ~n5327 & n15729 ) ;
  assign n15731 = ( n4990 & ~n15730 ) | ( n4990 & 1'b0 ) | ( ~n15730 & 1'b0 ) ;
  assign n15759 = n4668 | n15731 ;
  assign n15760 = n15745 | n15759 ;
  assign n15761 = n15751 &  n15760 ;
  assign n15762 = ( n15739 & ~n15742 ) | ( n15739 & 1'b0 ) | ( ~n15742 & 1'b0 ) ;
  assign n15763 = ( n4990 & ~n15762 ) | ( n4990 & n15736 ) | ( ~n15762 & n15736 ) ;
  assign n15764 = n4668 &  n15763 ;
  assign n15765 = n4353 | n15764 ;
  assign n15766 = n15761 | n15765 ;
  assign n15767 = n15758 &  n15766 ;
  assign n15746 = n15731 | n15745 ;
  assign n15752 = ( n4668 & n15746 ) | ( n4668 & n15751 ) | ( n15746 & n15751 ) ;
  assign n15753 = n4353 &  n15752 ;
  assign n15781 = n4053 | n15753 ;
  assign n15782 = n15767 | n15781 ;
  assign n15783 = n15773 &  n15782 ;
  assign n15784 = n15761 | n15764 ;
  assign n15785 = ( n4353 & n15758 ) | ( n4353 & n15784 ) | ( n15758 & n15784 ) ;
  assign n15786 = n4053 &  n15785 ;
  assign n15787 = n3760 | n15786 ;
  assign n15788 = n15783 | n15787 ;
  assign n15789 = n15780 &  n15788 ;
  assign n15768 = n15753 | n15767 ;
  assign n15774 = ( n4053 & n15768 ) | ( n4053 & n15773 ) | ( n15768 & n15773 ) ;
  assign n15775 = n3760 &  n15774 ;
  assign n15803 = n3482 | n15775 ;
  assign n15804 = n15789 | n15803 ;
  assign n15805 = ~n15795 & n15804 ;
  assign n15806 = n15783 | n15786 ;
  assign n15807 = ( n3760 & n15780 ) | ( n3760 & n15806 ) | ( n15780 & n15806 ) ;
  assign n15808 = n3482 &  n15807 ;
  assign n15809 = n3211 | n15808 ;
  assign n15810 = n15805 | n15809 ;
  assign n15811 = ~n15802 & n15810 ;
  assign n15790 = n15775 | n15789 ;
  assign n15796 = ( n3482 & ~n15795 ) | ( n3482 & n15790 ) | ( ~n15795 & n15790 ) ;
  assign n15797 = n3211 &  n15796 ;
  assign n15825 = n2955 | n15797 ;
  assign n15826 = n15811 | n15825 ;
  assign n15827 = n15817 &  n15826 ;
  assign n15828 = n15805 | n15808 ;
  assign n15829 = ( n3211 & ~n15802 ) | ( n3211 & n15828 ) | ( ~n15802 & n15828 ) ;
  assign n15830 = n2955 &  n15829 ;
  assign n15831 = n2706 | n15830 ;
  assign n15832 = n15827 | n15831 ;
  assign n15833 = ~n15824 & n15832 ;
  assign n15812 = n15797 | n15811 ;
  assign n15818 = ( n2955 & n15812 ) | ( n2955 & n15817 ) | ( n15812 & n15817 ) ;
  assign n15819 = n2706 &  n15818 ;
  assign n15847 = n2472 | n15819 ;
  assign n15848 = n15833 | n15847 ;
  assign n15849 = n15839 &  n15848 ;
  assign n15850 = n15827 | n15830 ;
  assign n15851 = ( n2706 & ~n15824 ) | ( n2706 & n15850 ) | ( ~n15824 & n15850 ) ;
  assign n15852 = n2472 &  n15851 ;
  assign n15853 = n2245 | n15852 ;
  assign n15854 = n15849 | n15853 ;
  assign n15855 = n15846 &  n15854 ;
  assign n15834 = n15819 | n15833 ;
  assign n15840 = ( n2472 & n15834 ) | ( n2472 & n15839 ) | ( n15834 & n15839 ) ;
  assign n15841 = n2245 &  n15840 ;
  assign n15869 = ( n2033 & ~n15841 ) | ( n2033 & 1'b0 ) | ( ~n15841 & 1'b0 ) ;
  assign n15870 = ~n15855 & n15869 ;
  assign n15871 = n15861 | n15870 ;
  assign n15872 = n15849 | n15852 ;
  assign n15873 = ( n2245 & n15846 ) | ( n2245 & n15872 ) | ( n15846 & n15872 ) ;
  assign n15874 = ~n2033 & n15873 ;
  assign n15875 = n1827 | n15874 ;
  assign n15876 = ( n15871 & ~n15875 ) | ( n15871 & 1'b0 ) | ( ~n15875 & 1'b0 ) ;
  assign n15877 = n15868 | n15876 ;
  assign n15856 = n15841 | n15855 ;
  assign n15862 = ( n2033 & ~n15856 ) | ( n2033 & n15861 ) | ( ~n15856 & n15861 ) ;
  assign n15863 = ( n1827 & ~n15862 ) | ( n1827 & 1'b0 ) | ( ~n15862 & 1'b0 ) ;
  assign n15891 = ( n1636 & ~n15863 ) | ( n1636 & 1'b0 ) | ( ~n15863 & 1'b0 ) ;
  assign n15892 = n15877 &  n15891 ;
  assign n15893 = n15883 | n15892 ;
  assign n15894 = ( n15871 & ~n15874 ) | ( n15871 & 1'b0 ) | ( ~n15874 & 1'b0 ) ;
  assign n15895 = ( n15868 & ~n1827 ) | ( n15868 & n15894 ) | ( ~n1827 & n15894 ) ;
  assign n15896 = n1636 | n15895 ;
  assign n15897 = n1452 &  n15896 ;
  assign n15898 = n15893 &  n15897 ;
  assign n15899 = n15890 | n15898 ;
  assign n15878 = ~n15863 & n15877 ;
  assign n15884 = ( n1636 & n15878 ) | ( n1636 & n15883 ) | ( n15878 & n15883 ) ;
  assign n15885 = n1452 | n15884 ;
  assign n15913 = ~n1283 & n15885 ;
  assign n15914 = n15899 &  n15913 ;
  assign n15915 = n15905 | n15914 ;
  assign n15916 = n15893 &  n15896 ;
  assign n15917 = ( n1452 & n15890 ) | ( n1452 & n15916 ) | ( n15890 & n15916 ) ;
  assign n15918 = ( n1283 & ~n15917 ) | ( n1283 & 1'b0 ) | ( ~n15917 & 1'b0 ) ;
  assign n15933 = ( n15915 & ~n15918 ) | ( n15915 & 1'b0 ) | ( ~n15918 & 1'b0 ) ;
  assign n15934 = ( n1122 & ~n15912 ) | ( n1122 & n15933 ) | ( ~n15912 & n15933 ) ;
  assign n15935 = n976 | n15934 ;
  assign n16010 = ~n15421 & n15484 ;
  assign n16011 = ( n15408 & n15413 ) | ( n15408 & n15484 ) | ( n15413 & n15484 ) ;
  assign n16013 = ( n16010 & ~n15408 ) | ( n16010 & n16011 ) | ( ~n15408 & n16011 ) ;
  assign n16012 = ( n15484 & ~n16011 ) | ( n15484 & n16010 ) | ( ~n16011 & n16010 ) ;
  assign n16014 = ( n15413 & ~n16013 ) | ( n15413 & n16012 ) | ( ~n16013 & n16012 ) ;
  assign n15988 = ~n15399 & n15484 ;
  assign n15989 = ( n15386 & n15391 ) | ( n15386 & n15484 ) | ( n15391 & n15484 ) ;
  assign n15991 = ( n15988 & ~n15386 ) | ( n15988 & n15989 ) | ( ~n15386 & n15989 ) ;
  assign n15990 = ( n15484 & ~n15989 ) | ( n15484 & n15988 ) | ( ~n15989 & n15988 ) ;
  assign n15992 = ( n15391 & ~n15991 ) | ( n15391 & n15990 ) | ( ~n15991 & n15990 ) ;
  assign n15900 = n15885 &  n15899 ;
  assign n15906 = ( n15900 & ~n1283 ) | ( n15900 & n15905 ) | ( ~n1283 & n15905 ) ;
  assign n15907 = n1122 | n15906 ;
  assign n15919 = ( n1122 & ~n15918 ) | ( n1122 & 1'b0 ) | ( ~n15918 & 1'b0 ) ;
  assign n15920 = n15915 &  n15919 ;
  assign n15921 = ( n15912 & ~n15920 ) | ( n15912 & 1'b0 ) | ( ~n15920 & 1'b0 ) ;
  assign n15922 = ( n15907 & ~n15921 ) | ( n15907 & 1'b0 ) | ( ~n15921 & 1'b0 ) ;
  assign n15928 = ( n976 & n15922 ) | ( n976 & n15927 ) | ( n15922 & n15927 ) ;
  assign n15929 = ( n837 & ~n15928 ) | ( n837 & 1'b0 ) | ( ~n15928 & 1'b0 ) ;
  assign n15930 = n976 &  n15907 ;
  assign n15931 = ~n15921 & n15930 ;
  assign n15932 = n15927 | n15931 ;
  assign n15936 = ~n837 & n15935 ;
  assign n15937 = n15932 &  n15936 ;
  assign n15938 = ( n15349 & ~n15340 ) | ( n15349 & n15353 ) | ( ~n15340 & n15353 ) ;
  assign n15939 = ( n15349 & ~n15938 ) | ( n15349 & n15484 ) | ( ~n15938 & n15484 ) ;
  assign n15940 = ( n15484 & ~n15353 ) | ( n15484 & n15938 ) | ( ~n15353 & n15938 ) ;
  assign n15941 = ( n15340 & ~n15939 ) | ( n15340 & n15940 ) | ( ~n15939 & n15940 ) ;
  assign n15942 = n15937 | n15941 ;
  assign n15943 = ~n15929 & n15942 ;
  assign n15945 = ( n15342 & ~n15347 ) | ( n15342 & n15484 ) | ( ~n15347 & n15484 ) ;
  assign n15944 = n15355 &  n15484 ;
  assign n15946 = ( n15484 & ~n15945 ) | ( n15484 & n15944 ) | ( ~n15945 & n15944 ) ;
  assign n15947 = ( n15944 & ~n15342 ) | ( n15944 & n15945 ) | ( ~n15342 & n15945 ) ;
  assign n15948 = ( n15347 & ~n15946 ) | ( n15347 & n15947 ) | ( ~n15946 & n15947 ) ;
  assign n15949 = ( n713 & ~n15943 ) | ( n713 & n15948 ) | ( ~n15943 & n15948 ) ;
  assign n15950 = n595 &  n15949 ;
  assign n15952 = ( n15371 & ~n15362 ) | ( n15371 & n15375 ) | ( ~n15362 & n15375 ) ;
  assign n15951 = n15375 | n15484 ;
  assign n15954 = ( n15375 & ~n15952 ) | ( n15375 & n15951 ) | ( ~n15952 & n15951 ) ;
  assign n15953 = ( n15951 & ~n15371 ) | ( n15951 & n15952 ) | ( ~n15371 & n15952 ) ;
  assign n15955 = ( n15362 & ~n15954 ) | ( n15362 & n15953 ) | ( ~n15954 & n15953 ) ;
  assign n15956 = n713 | n15929 ;
  assign n15957 = ( n15942 & ~n15956 ) | ( n15942 & 1'b0 ) | ( ~n15956 & 1'b0 ) ;
  assign n15958 = ( n15948 & ~n15957 ) | ( n15948 & 1'b0 ) | ( ~n15957 & 1'b0 ) ;
  assign n15959 = n15932 &  n15935 ;
  assign n15960 = ( n15941 & ~n837 ) | ( n15941 & n15959 ) | ( ~n837 & n15959 ) ;
  assign n15961 = ( n713 & ~n15960 ) | ( n713 & 1'b0 ) | ( ~n15960 & 1'b0 ) ;
  assign n15962 = n595 | n15961 ;
  assign n15963 = n15958 | n15962 ;
  assign n15964 = ~n15955 & n15963 ;
  assign n15965 = n15950 | n15964 ;
  assign n15966 = ~n15377 & n15484 ;
  assign n15967 = ( n15364 & n15369 ) | ( n15364 & n15484 ) | ( n15369 & n15484 ) ;
  assign n15969 = ( n15966 & ~n15364 ) | ( n15966 & n15967 ) | ( ~n15364 & n15967 ) ;
  assign n15968 = ( n15484 & ~n15967 ) | ( n15484 & n15966 ) | ( ~n15967 & n15966 ) ;
  assign n15970 = ( n15369 & ~n15969 ) | ( n15369 & n15968 ) | ( ~n15969 & n15968 ) ;
  assign n15971 = ( n492 & n15965 ) | ( n492 & n15970 ) | ( n15965 & n15970 ) ;
  assign n15972 = n396 &  n15971 ;
  assign n15973 = n15397 | n15484 ;
  assign n15974 = ( n15384 & n15393 ) | ( n15384 & n15397 ) | ( n15393 & n15397 ) ;
  assign n15975 = ( n15973 & ~n15393 ) | ( n15973 & n15974 ) | ( ~n15393 & n15974 ) ;
  assign n15976 = ( n15397 & ~n15974 ) | ( n15397 & n15973 ) | ( ~n15974 & n15973 ) ;
  assign n15977 = ( n15384 & ~n15975 ) | ( n15384 & n15976 ) | ( ~n15975 & n15976 ) ;
  assign n15978 = n492 | n15950 ;
  assign n15979 = n15964 | n15978 ;
  assign n15980 = n15970 &  n15979 ;
  assign n15981 = n15958 | n15961 ;
  assign n15982 = ( n595 & ~n15955 ) | ( n595 & n15981 ) | ( ~n15955 & n15981 ) ;
  assign n15983 = n492 &  n15982 ;
  assign n15984 = n396 | n15983 ;
  assign n15985 = n15980 | n15984 ;
  assign n15986 = n15977 &  n15985 ;
  assign n15987 = n15972 | n15986 ;
  assign n15993 = ( n315 & ~n15992 ) | ( n315 & n15987 ) | ( ~n15992 & n15987 ) ;
  assign n15994 = n240 &  n15993 ;
  assign n15995 = n15419 | n15484 ;
  assign n15996 = ( n15406 & n15415 ) | ( n15406 & n15419 ) | ( n15415 & n15419 ) ;
  assign n15997 = ( n15995 & ~n15415 ) | ( n15995 & n15996 ) | ( ~n15415 & n15996 ) ;
  assign n15998 = ( n15419 & ~n15996 ) | ( n15419 & n15995 ) | ( ~n15996 & n15995 ) ;
  assign n15999 = ( n15406 & ~n15997 ) | ( n15406 & n15998 ) | ( ~n15997 & n15998 ) ;
  assign n16000 = n315 | n15972 ;
  assign n16001 = n15986 | n16000 ;
  assign n16002 = ~n15992 & n16001 ;
  assign n16003 = n15980 | n15983 ;
  assign n16004 = ( n396 & n15977 ) | ( n396 & n16003 ) | ( n15977 & n16003 ) ;
  assign n16005 = n315 &  n16004 ;
  assign n16006 = n240 | n16005 ;
  assign n16007 = n16002 | n16006 ;
  assign n16008 = n15999 &  n16007 ;
  assign n16009 = n15994 | n16008 ;
  assign n16015 = ( n181 & ~n16014 ) | ( n181 & n16009 ) | ( ~n16014 & n16009 ) ;
  assign n16016 = ~n145 & n16015 ;
  assign n16017 = n15441 | n15484 ;
  assign n16018 = ( n15428 & n15437 ) | ( n15428 & n15441 ) | ( n15437 & n15441 ) ;
  assign n16019 = ( n16017 & ~n15437 ) | ( n16017 & n16018 ) | ( ~n15437 & n16018 ) ;
  assign n16020 = ( n15441 & ~n16018 ) | ( n15441 & n16017 ) | ( ~n16018 & n16017 ) ;
  assign n16021 = ( n15428 & ~n16019 ) | ( n15428 & n16020 ) | ( ~n16019 & n16020 ) ;
  assign n16022 = n181 | n15994 ;
  assign n16023 = n16008 | n16022 ;
  assign n16024 = ~n16014 & n16023 ;
  assign n16025 = n16002 | n16005 ;
  assign n16026 = ( n240 & n15999 ) | ( n240 & n16025 ) | ( n15999 & n16025 ) ;
  assign n16027 = n181 &  n16026 ;
  assign n16028 = ( n145 & ~n16027 ) | ( n145 & 1'b0 ) | ( ~n16027 & 1'b0 ) ;
  assign n16029 = ~n16024 & n16028 ;
  assign n16030 = n16021 | n16029 ;
  assign n16031 = ~n16016 & n16030 ;
  assign n16032 = n15430 | n15484 ;
  assign n16033 = ( n15435 & ~n15430 ) | ( n15435 & n15443 ) | ( ~n15430 & n15443 ) ;
  assign n16035 = ( n15430 & n16032 ) | ( n15430 & n16033 ) | ( n16032 & n16033 ) ;
  assign n16034 = ( n15443 & ~n16033 ) | ( n15443 & n16032 ) | ( ~n16033 & n16032 ) ;
  assign n16036 = ( n15435 & ~n16035 ) | ( n15435 & n16034 ) | ( ~n16035 & n16034 ) ;
  assign n16037 = ( n150 & ~n16031 ) | ( n150 & n16036 ) | ( ~n16031 & n16036 ) ;
  assign n16038 = n15450 | n15469 ;
  assign n16039 = ( n15466 & ~n15484 ) | ( n15466 & n16038 ) | ( ~n15484 & n16038 ) ;
  assign n16040 = ( n15466 & ~n16039 ) | ( n15466 & 1'b0 ) | ( ~n16039 & 1'b0 ) ;
  assign n16041 = ( n15466 & ~n15469 ) | ( n15466 & 1'b0 ) | ( ~n15469 & 1'b0 ) ;
  assign n16042 = ~n15484 & n16041 ;
  assign n16043 = ( n15450 & ~n16041 ) | ( n15450 & n16042 ) | ( ~n16041 & n16042 ) ;
  assign n16044 = n16040 | n16043 ;
  assign n16045 = ( n15451 & ~n15458 ) | ( n15451 & 1'b0 ) | ( ~n15458 & 1'b0 ) ;
  assign n16046 = ~n15484 & n16045 ;
  assign n16047 = ( n15472 & ~n16046 ) | ( n15472 & n16045 ) | ( ~n16046 & n16045 ) ;
  assign n16048 = ( n16044 & ~n16047 ) | ( n16044 & 1'b0 ) | ( ~n16047 & 1'b0 ) ;
  assign n16049 = ~n16037 & n16048 ;
  assign n16050 = ( n133 & ~n16049 ) | ( n133 & n16048 ) | ( ~n16049 & n16048 ) ;
  assign n16051 = n150 | n16016 ;
  assign n16052 = ( n16030 & ~n16051 ) | ( n16030 & 1'b0 ) | ( ~n16051 & 1'b0 ) ;
  assign n16057 = n16036 &  n16052 ;
  assign n16053 = n16024 | n16027 ;
  assign n16054 = ( n145 & ~n16053 ) | ( n145 & n16021 ) | ( ~n16053 & n16021 ) ;
  assign n16055 = ( n150 & ~n16054 ) | ( n150 & 1'b0 ) | ( ~n16054 & 1'b0 ) ;
  assign n16056 = n16044 | n16055 ;
  assign n16058 = ( n16036 & ~n16057 ) | ( n16036 & n16056 ) | ( ~n16057 & n16056 ) ;
  assign n16060 = ( n133 & ~n15458 ) | ( n133 & n15451 ) | ( ~n15458 & n15451 ) ;
  assign n16059 = ( n15458 & ~n15451 ) | ( n15458 & n15484 ) | ( ~n15451 & n15484 ) ;
  assign n16061 = ~n15458 & n16059 ;
  assign n16062 = ( n15458 & n16060 ) | ( n15458 & n16061 ) | ( n16060 & n16061 ) ;
  assign n16063 = n15454 | n15481 ;
  assign n16064 = ( n15457 & n15476 ) | ( n15457 & n16063 ) | ( n15476 & n16063 ) ;
  assign n16065 = ( n15457 & ~n16064 ) | ( n15457 & 1'b0 ) | ( ~n16064 & 1'b0 ) ;
  assign n16066 = ( n15464 & ~n16065 ) | ( n15464 & n15472 ) | ( ~n16065 & n15472 ) ;
  assign n16067 = ( n15464 & ~n16066 ) | ( n15464 & 1'b0 ) | ( ~n16066 & 1'b0 ) ;
  assign n16068 = n16062 | n16067 ;
  assign n16069 = ( n16058 & ~n16068 ) | ( n16058 & 1'b0 ) | ( ~n16068 & 1'b0 ) ;
  assign n16070 = ~n16050 | ~n16069 ;
  assign n16531 = ( n15935 & ~n16070 ) | ( n15935 & 1'b0 ) | ( ~n16070 & 1'b0 ) ;
  assign n16532 = ( n15927 & n15931 ) | ( n15927 & n15935 ) | ( n15931 & n15935 ) ;
  assign n16533 = ( n16531 & ~n15931 ) | ( n16531 & n16532 ) | ( ~n15931 & n16532 ) ;
  assign n16534 = ( n15935 & ~n16532 ) | ( n15935 & n16531 ) | ( ~n16532 & n16531 ) ;
  assign n16535 = ( n15927 & ~n16533 ) | ( n15927 & n16534 ) | ( ~n16533 & n16534 ) ;
  assign n16525 = ( n15907 & ~n15912 ) | ( n15907 & n15920 ) | ( ~n15912 & n15920 ) ;
  assign n16524 = ( n15907 & ~n16070 ) | ( n15907 & 1'b0 ) | ( ~n16070 & 1'b0 ) ;
  assign n16527 = ( n15907 & ~n16525 ) | ( n15907 & n16524 ) | ( ~n16525 & n16524 ) ;
  assign n16526 = ( n16524 & ~n15920 ) | ( n16524 & n16525 ) | ( ~n15920 & n16525 ) ;
  assign n16528 = ( n15912 & ~n16527 ) | ( n15912 & n16526 ) | ( ~n16527 & n16526 ) ;
  assign n16437 = ( n15819 & ~n15824 ) | ( n15819 & n15832 ) | ( ~n15824 & n15832 ) ;
  assign n16436 = n15819 | n16070 ;
  assign n16439 = ( n15819 & ~n16437 ) | ( n15819 & n16436 ) | ( ~n16437 & n16436 ) ;
  assign n16438 = ( n16436 & ~n15832 ) | ( n16436 & n16437 ) | ( ~n15832 & n16437 ) ;
  assign n16440 = ( n15824 & ~n16439 ) | ( n15824 & n16438 ) | ( ~n16439 & n16438 ) ;
  assign n16415 = ( n15797 & ~n15802 ) | ( n15797 & n15810 ) | ( ~n15802 & n15810 ) ;
  assign n16414 = n15797 | n16070 ;
  assign n16417 = ( n15797 & ~n16415 ) | ( n15797 & n16414 ) | ( ~n16415 & n16414 ) ;
  assign n16416 = ( n16414 & ~n15810 ) | ( n16414 & n16415 ) | ( ~n15810 & n16415 ) ;
  assign n16418 = ( n15802 & ~n16417 ) | ( n15802 & n16416 ) | ( ~n16417 & n16416 ) ;
  assign n16077 = ( x22 & ~n16070 ) | ( x22 & x23 ) | ( ~n16070 & x23 ) ;
  assign n16083 = ( x22 & ~x23 ) | ( x22 & 1'b0 ) | ( ~x23 & 1'b0 ) ;
  assign n16073 = x20 | x21 ;
  assign n16078 = ~x22 & n16073 ;
  assign n16079 = ( x22 & ~n15482 ) | ( x22 & n16078 ) | ( ~n15482 & n16078 ) ;
  assign n16080 = ( n15464 & ~n16079 ) | ( n15464 & n15472 ) | ( ~n16079 & n15472 ) ;
  assign n16081 = ( n15464 & ~n16080 ) | ( n15464 & 1'b0 ) | ( ~n16080 & 1'b0 ) ;
  assign n16082 = ( n16070 & ~x23 ) | ( n16070 & n16081 ) | ( ~x23 & n16081 ) ;
  assign n16084 = ( n16077 & ~n16083 ) | ( n16077 & n16082 ) | ( ~n16083 & n16082 ) ;
  assign n16074 = x22 | n16073 ;
  assign n16075 = x22 &  n16070 ;
  assign n16076 = ( n15484 & ~n16074 ) | ( n15484 & n16075 ) | ( ~n16074 & n16075 ) ;
  assign n16085 = n16076 &  n16084 ;
  assign n16086 = ( n14905 & ~n16084 ) | ( n14905 & n16085 ) | ( ~n16084 & n16085 ) ;
  assign n16087 = n14905 | n16076 ;
  assign n16088 = ( n16084 & ~n16087 ) | ( n16084 & 1'b0 ) | ( ~n16087 & 1'b0 ) ;
  assign n16090 = ( n15484 & ~n16067 ) | ( n15484 & 1'b0 ) | ( ~n16067 & 1'b0 ) ;
  assign n16091 = ( n16058 & ~n16090 ) | ( n16058 & n16062 ) | ( ~n16090 & n16062 ) ;
  assign n16092 = ( n16058 & ~n16091 ) | ( n16058 & 1'b0 ) | ( ~n16091 & 1'b0 ) ;
  assign n16093 = n16050 &  n16092 ;
  assign n16089 = ~n14906 & n16070 ;
  assign n16094 = ( n16089 & ~n16093 ) | ( n16089 & 1'b0 ) | ( ~n16093 & 1'b0 ) ;
  assign n16095 = ( x24 & n16093 ) | ( x24 & n16094 ) | ( n16093 & n16094 ) ;
  assign n16096 = x24 | n16093 ;
  assign n16097 = n16089 | n16096 ;
  assign n16098 = ~n16095 & n16097 ;
  assign n16099 = n16088 | n16098 ;
  assign n16100 = ~n16086 & n16099 ;
  assign n16104 = ~x24 & n15484 ;
  assign n16105 = ( x25 & ~n16104 ) | ( x25 & 1'b0 ) | ( ~n16104 & 1'b0 ) ;
  assign n16106 = n15496 | n16105 ;
  assign n16101 = ( n15484 & ~x24 ) | ( n15484 & n15491 ) | ( ~x24 & n15491 ) ;
  assign n16102 = x24 &  n16101 ;
  assign n16103 = ( n15486 & ~n16102 ) | ( n15486 & n15491 ) | ( ~n16102 & n15491 ) ;
  assign n16107 = ( n16070 & ~n16106 ) | ( n16070 & n16103 ) | ( ~n16106 & n16103 ) ;
  assign n16109 = ( n16070 & ~n16107 ) | ( n16070 & 1'b0 ) | ( ~n16107 & 1'b0 ) ;
  assign n16108 = ~n16103 & n16107 ;
  assign n16110 = ( n16106 & ~n16109 ) | ( n16106 & n16108 ) | ( ~n16109 & n16108 ) ;
  assign n16111 = ( n16100 & ~n14341 ) | ( n16100 & n16110 ) | ( ~n14341 & n16110 ) ;
  assign n16112 = ( n13784 & ~n16111 ) | ( n13784 & 1'b0 ) | ( ~n16111 & 1'b0 ) ;
  assign n16113 = ~n15519 & n15522 ;
  assign n16114 = ( n15505 & ~n15519 ) | ( n15505 & n16113 ) | ( ~n15519 & n16113 ) ;
  assign n16116 = ( n15519 & n16070 ) | ( n15519 & n16114 ) | ( n16070 & n16114 ) ;
  assign n16115 = ( n16070 & ~n16114 ) | ( n16070 & n16113 ) | ( ~n16114 & n16113 ) ;
  assign n16117 = ( n15505 & ~n16116 ) | ( n15505 & n16115 ) | ( ~n16116 & n16115 ) ;
  assign n16118 = n14341 | n16086 ;
  assign n16119 = ( n16099 & ~n16118 ) | ( n16099 & 1'b0 ) | ( ~n16118 & 1'b0 ) ;
  assign n16120 = n16110 | n16119 ;
  assign n16121 = ~n16076 & n16084 ;
  assign n16122 = ( n16098 & ~n14905 ) | ( n16098 & n16121 ) | ( ~n14905 & n16121 ) ;
  assign n16123 = ( n14341 & ~n16122 ) | ( n14341 & 1'b0 ) | ( ~n16122 & 1'b0 ) ;
  assign n16124 = n13784 | n16123 ;
  assign n16125 = ( n16120 & ~n16124 ) | ( n16120 & 1'b0 ) | ( ~n16124 & 1'b0 ) ;
  assign n16126 = n16117 | n16125 ;
  assign n16127 = ~n16112 & n16126 ;
  assign n16128 = n15507 | n16070 ;
  assign n16129 = ( n15507 & ~n15524 ) | ( n15507 & n15517 ) | ( ~n15524 & n15517 ) ;
  assign n16130 = ( n15524 & n16128 ) | ( n15524 & n16129 ) | ( n16128 & n16129 ) ;
  assign n16131 = ( n15507 & ~n16129 ) | ( n15507 & n16128 ) | ( ~n16129 & n16128 ) ;
  assign n16132 = ( n15517 & ~n16130 ) | ( n15517 & n16131 ) | ( ~n16130 & n16131 ) ;
  assign n16133 = ( n16127 & ~n13242 ) | ( n16127 & n16132 ) | ( ~n13242 & n16132 ) ;
  assign n16134 = ( n12707 & ~n16133 ) | ( n12707 & 1'b0 ) | ( ~n16133 & 1'b0 ) ;
  assign n16135 = n15544 | n16070 ;
  assign n16136 = ( n15531 & ~n15544 ) | ( n15531 & n15540 ) | ( ~n15544 & n15540 ) ;
  assign n16138 = ( n15544 & n16135 ) | ( n15544 & n16136 ) | ( n16135 & n16136 ) ;
  assign n16137 = ( n15540 & ~n16136 ) | ( n15540 & n16135 ) | ( ~n16136 & n16135 ) ;
  assign n16139 = ( n15531 & ~n16138 ) | ( n15531 & n16137 ) | ( ~n16138 & n16137 ) ;
  assign n16140 = n13242 | n16112 ;
  assign n16141 = ( n16126 & ~n16140 ) | ( n16126 & 1'b0 ) | ( ~n16140 & 1'b0 ) ;
  assign n16142 = n16132 | n16141 ;
  assign n16143 = ( n16120 & ~n16123 ) | ( n16120 & 1'b0 ) | ( ~n16123 & 1'b0 ) ;
  assign n16144 = ( n16117 & ~n13784 ) | ( n16117 & n16143 ) | ( ~n13784 & n16143 ) ;
  assign n16145 = ( n13242 & ~n16144 ) | ( n13242 & 1'b0 ) | ( ~n16144 & 1'b0 ) ;
  assign n16146 = n12707 | n16145 ;
  assign n16147 = ( n16142 & ~n16146 ) | ( n16142 & 1'b0 ) | ( ~n16146 & 1'b0 ) ;
  assign n16148 = n16139 | n16147 ;
  assign n16149 = ~n16134 & n16148 ;
  assign n16150 = n15546 &  n16070 ;
  assign n16151 = ( n15533 & n15538 ) | ( n15533 & n16070 ) | ( n15538 & n16070 ) ;
  assign n16153 = ( n16150 & ~n15533 ) | ( n16150 & n16151 ) | ( ~n15533 & n16151 ) ;
  assign n16152 = ( n16070 & ~n16151 ) | ( n16070 & n16150 ) | ( ~n16151 & n16150 ) ;
  assign n16154 = ( n15538 & ~n16153 ) | ( n15538 & n16152 ) | ( ~n16153 & n16152 ) ;
  assign n16155 = ( n16149 & ~n12187 ) | ( n16149 & n16154 ) | ( ~n12187 & n16154 ) ;
  assign n16156 = ( n11674 & ~n16155 ) | ( n11674 & 1'b0 ) | ( ~n16155 & 1'b0 ) ;
  assign n16157 = n15566 | n16070 ;
  assign n16158 = ( n15553 & ~n15562 ) | ( n15553 & n15566 ) | ( ~n15562 & n15566 ) ;
  assign n16159 = ( n15562 & n16157 ) | ( n15562 & n16158 ) | ( n16157 & n16158 ) ;
  assign n16160 = ( n15566 & ~n16158 ) | ( n15566 & n16157 ) | ( ~n16158 & n16157 ) ;
  assign n16161 = ( n15553 & ~n16159 ) | ( n15553 & n16160 ) | ( ~n16159 & n16160 ) ;
  assign n16162 = n12187 | n16134 ;
  assign n16163 = ( n16148 & ~n16162 ) | ( n16148 & 1'b0 ) | ( ~n16162 & 1'b0 ) ;
  assign n16164 = n16154 | n16163 ;
  assign n16165 = ( n16142 & ~n16145 ) | ( n16142 & 1'b0 ) | ( ~n16145 & 1'b0 ) ;
  assign n16166 = ( n16139 & ~n12707 ) | ( n16139 & n16165 ) | ( ~n12707 & n16165 ) ;
  assign n16167 = ( n12187 & ~n16166 ) | ( n12187 & 1'b0 ) | ( ~n16166 & 1'b0 ) ;
  assign n16168 = n11674 | n16167 ;
  assign n16169 = ( n16164 & ~n16168 ) | ( n16164 & 1'b0 ) | ( ~n16168 & 1'b0 ) ;
  assign n16170 = n16161 | n16169 ;
  assign n16171 = ~n16156 & n16170 ;
  assign n16172 = n15555 | n16070 ;
  assign n16173 = ( n15560 & ~n15555 ) | ( n15560 & n15568 ) | ( ~n15555 & n15568 ) ;
  assign n16175 = ( n15555 & n16172 ) | ( n15555 & n16173 ) | ( n16172 & n16173 ) ;
  assign n16174 = ( n15568 & ~n16173 ) | ( n15568 & n16172 ) | ( ~n16173 & n16172 ) ;
  assign n16176 = ( n15560 & ~n16175 ) | ( n15560 & n16174 ) | ( ~n16175 & n16174 ) ;
  assign n16177 = ( n16171 & ~n11176 ) | ( n16171 & n16176 ) | ( ~n11176 & n16176 ) ;
  assign n16178 = ( n10685 & ~n16177 ) | ( n10685 & 1'b0 ) | ( ~n16177 & 1'b0 ) ;
  assign n16179 = n15588 | n16070 ;
  assign n16180 = ( n15575 & ~n15584 ) | ( n15575 & n15588 ) | ( ~n15584 & n15588 ) ;
  assign n16181 = ( n15584 & n16179 ) | ( n15584 & n16180 ) | ( n16179 & n16180 ) ;
  assign n16182 = ( n15588 & ~n16180 ) | ( n15588 & n16179 ) | ( ~n16180 & n16179 ) ;
  assign n16183 = ( n15575 & ~n16181 ) | ( n15575 & n16182 ) | ( ~n16181 & n16182 ) ;
  assign n16184 = n11176 | n16156 ;
  assign n16185 = ( n16170 & ~n16184 ) | ( n16170 & 1'b0 ) | ( ~n16184 & 1'b0 ) ;
  assign n16186 = n16176 | n16185 ;
  assign n16187 = ( n16164 & ~n16167 ) | ( n16164 & 1'b0 ) | ( ~n16167 & 1'b0 ) ;
  assign n16188 = ( n16161 & ~n11674 ) | ( n16161 & n16187 ) | ( ~n11674 & n16187 ) ;
  assign n16189 = ( n11176 & ~n16188 ) | ( n11176 & 1'b0 ) | ( ~n16188 & 1'b0 ) ;
  assign n16190 = n10685 | n16189 ;
  assign n16191 = ( n16186 & ~n16190 ) | ( n16186 & 1'b0 ) | ( ~n16190 & 1'b0 ) ;
  assign n16192 = n16183 | n16191 ;
  assign n16193 = ~n16178 & n16192 ;
  assign n16194 = n15577 | n16070 ;
  assign n16195 = ( n15577 & ~n15590 ) | ( n15577 & n15582 ) | ( ~n15590 & n15582 ) ;
  assign n16196 = ( n15590 & n16194 ) | ( n15590 & n16195 ) | ( n16194 & n16195 ) ;
  assign n16197 = ( n15577 & ~n16195 ) | ( n15577 & n16194 ) | ( ~n16195 & n16194 ) ;
  assign n16198 = ( n15582 & ~n16196 ) | ( n15582 & n16197 ) | ( ~n16196 & n16197 ) ;
  assign n16199 = ( n16193 & ~n10209 ) | ( n16193 & n16198 ) | ( ~n10209 & n16198 ) ;
  assign n16200 = n9740 | n16199 ;
  assign n16201 = n15610 | n16070 ;
  assign n16202 = ( n15597 & ~n15610 ) | ( n15597 & n15606 ) | ( ~n15610 & n15606 ) ;
  assign n16204 = ( n15610 & n16201 ) | ( n15610 & n16202 ) | ( n16201 & n16202 ) ;
  assign n16203 = ( n15606 & ~n16202 ) | ( n15606 & n16201 ) | ( ~n16202 & n16201 ) ;
  assign n16205 = ( n15597 & ~n16204 ) | ( n15597 & n16203 ) | ( ~n16204 & n16203 ) ;
  assign n16206 = n10209 | n16178 ;
  assign n16207 = ( n16192 & ~n16206 ) | ( n16192 & 1'b0 ) | ( ~n16206 & 1'b0 ) ;
  assign n16208 = n16198 | n16207 ;
  assign n16209 = ( n16186 & ~n16189 ) | ( n16186 & 1'b0 ) | ( ~n16189 & 1'b0 ) ;
  assign n16210 = ( n16183 & ~n10685 ) | ( n16183 & n16209 ) | ( ~n10685 & n16209 ) ;
  assign n16211 = ( n10209 & ~n16210 ) | ( n10209 & 1'b0 ) | ( ~n16210 & 1'b0 ) ;
  assign n16212 = ( n9740 & ~n16211 ) | ( n9740 & 1'b0 ) | ( ~n16211 & 1'b0 ) ;
  assign n16213 = n16208 &  n16212 ;
  assign n16214 = n16205 | n16213 ;
  assign n16215 = n16200 &  n16214 ;
  assign n16216 = n15612 &  n16070 ;
  assign n16217 = ( n15604 & ~n15599 ) | ( n15604 & n16070 ) | ( ~n15599 & n16070 ) ;
  assign n16219 = ( n16216 & n15599 ) | ( n16216 & n16217 ) | ( n15599 & n16217 ) ;
  assign n16218 = ( n16070 & ~n16217 ) | ( n16070 & n16216 ) | ( ~n16217 & n16216 ) ;
  assign n16220 = ( n15604 & ~n16219 ) | ( n15604 & n16218 ) | ( ~n16219 & n16218 ) ;
  assign n16221 = ( n16215 & ~n9286 ) | ( n16215 & n16220 ) | ( ~n9286 & n16220 ) ;
  assign n16222 = ( n8839 & ~n16221 ) | ( n8839 & 1'b0 ) | ( ~n16221 & 1'b0 ) ;
  assign n16223 = n15632 | n16070 ;
  assign n16224 = ( n15619 & ~n15628 ) | ( n15619 & n15632 ) | ( ~n15628 & n15632 ) ;
  assign n16225 = ( n15628 & n16223 ) | ( n15628 & n16224 ) | ( n16223 & n16224 ) ;
  assign n16226 = ( n15632 & ~n16224 ) | ( n15632 & n16223 ) | ( ~n16224 & n16223 ) ;
  assign n16227 = ( n15619 & ~n16225 ) | ( n15619 & n16226 ) | ( ~n16225 & n16226 ) ;
  assign n16228 = ~n9286 & n16200 ;
  assign n16229 = n16214 &  n16228 ;
  assign n16230 = n16220 | n16229 ;
  assign n16231 = ( n16208 & ~n16211 ) | ( n16208 & 1'b0 ) | ( ~n16211 & 1'b0 ) ;
  assign n16232 = ( n9740 & n16205 ) | ( n9740 & n16231 ) | ( n16205 & n16231 ) ;
  assign n16233 = ( n9286 & ~n16232 ) | ( n9286 & 1'b0 ) | ( ~n16232 & 1'b0 ) ;
  assign n16234 = n8839 | n16233 ;
  assign n16235 = ( n16230 & ~n16234 ) | ( n16230 & 1'b0 ) | ( ~n16234 & 1'b0 ) ;
  assign n16236 = n16227 | n16235 ;
  assign n16237 = ~n16222 & n16236 ;
  assign n16238 = n15621 | n16070 ;
  assign n16239 = ( n15626 & ~n15621 ) | ( n15626 & n15634 ) | ( ~n15621 & n15634 ) ;
  assign n16241 = ( n15621 & n16238 ) | ( n15621 & n16239 ) | ( n16238 & n16239 ) ;
  assign n16240 = ( n15634 & ~n16239 ) | ( n15634 & n16238 ) | ( ~n16239 & n16238 ) ;
  assign n16242 = ( n15626 & ~n16241 ) | ( n15626 & n16240 ) | ( ~n16241 & n16240 ) ;
  assign n16243 = ( n16237 & ~n8407 ) | ( n16237 & n16242 ) | ( ~n8407 & n16242 ) ;
  assign n16244 = ( n7982 & ~n16243 ) | ( n7982 & 1'b0 ) | ( ~n16243 & 1'b0 ) ;
  assign n16245 = n15654 | n16070 ;
  assign n16246 = ( n15641 & ~n15650 ) | ( n15641 & n15654 ) | ( ~n15650 & n15654 ) ;
  assign n16247 = ( n15650 & n16245 ) | ( n15650 & n16246 ) | ( n16245 & n16246 ) ;
  assign n16248 = ( n15654 & ~n16246 ) | ( n15654 & n16245 ) | ( ~n16246 & n16245 ) ;
  assign n16249 = ( n15641 & ~n16247 ) | ( n15641 & n16248 ) | ( ~n16247 & n16248 ) ;
  assign n16250 = n8407 | n16222 ;
  assign n16251 = ( n16236 & ~n16250 ) | ( n16236 & 1'b0 ) | ( ~n16250 & 1'b0 ) ;
  assign n16252 = n16242 | n16251 ;
  assign n16253 = ( n16230 & ~n16233 ) | ( n16230 & 1'b0 ) | ( ~n16233 & 1'b0 ) ;
  assign n16254 = ( n16227 & ~n8839 ) | ( n16227 & n16253 ) | ( ~n8839 & n16253 ) ;
  assign n16255 = ( n8407 & ~n16254 ) | ( n8407 & 1'b0 ) | ( ~n16254 & 1'b0 ) ;
  assign n16256 = n7982 | n16255 ;
  assign n16257 = ( n16252 & ~n16256 ) | ( n16252 & 1'b0 ) | ( ~n16256 & 1'b0 ) ;
  assign n16258 = n16249 | n16257 ;
  assign n16259 = ~n16244 & n16258 ;
  assign n16260 = n15643 | n16070 ;
  assign n16261 = ( n15648 & ~n15643 ) | ( n15648 & n15656 ) | ( ~n15643 & n15656 ) ;
  assign n16263 = ( n15643 & n16260 ) | ( n15643 & n16261 ) | ( n16260 & n16261 ) ;
  assign n16262 = ( n15656 & ~n16261 ) | ( n15656 & n16260 ) | ( ~n16261 & n16260 ) ;
  assign n16264 = ( n15648 & ~n16263 ) | ( n15648 & n16262 ) | ( ~n16263 & n16262 ) ;
  assign n16265 = ( n7572 & n16259 ) | ( n7572 & n16264 ) | ( n16259 & n16264 ) ;
  assign n16266 = n7169 | n16265 ;
  assign n16268 = ( n15672 & ~n15663 ) | ( n15672 & n15676 ) | ( ~n15663 & n15676 ) ;
  assign n16267 = ( n15676 & ~n16070 ) | ( n15676 & 1'b0 ) | ( ~n16070 & 1'b0 ) ;
  assign n16270 = ( n15676 & ~n16268 ) | ( n15676 & n16267 ) | ( ~n16268 & n16267 ) ;
  assign n16269 = ( n16267 & ~n15672 ) | ( n16267 & n16268 ) | ( ~n15672 & n16268 ) ;
  assign n16271 = ( n15663 & ~n16270 ) | ( n15663 & n16269 ) | ( ~n16270 & n16269 ) ;
  assign n16272 = ( n7572 & ~n16244 ) | ( n7572 & 1'b0 ) | ( ~n16244 & 1'b0 ) ;
  assign n16273 = n16258 &  n16272 ;
  assign n16274 = n16264 | n16273 ;
  assign n16275 = ( n16252 & ~n16255 ) | ( n16252 & 1'b0 ) | ( ~n16255 & 1'b0 ) ;
  assign n16276 = ( n16249 & ~n7982 ) | ( n16249 & n16275 ) | ( ~n7982 & n16275 ) ;
  assign n16277 = n7572 | n16276 ;
  assign n16278 = n7169 &  n16277 ;
  assign n16279 = n16274 &  n16278 ;
  assign n16280 = n16271 | n16279 ;
  assign n16281 = n16266 &  n16280 ;
  assign n16282 = ( n15665 & ~n16070 ) | ( n15665 & 1'b0 ) | ( ~n16070 & 1'b0 ) ;
  assign n16283 = ( n15665 & n15670 ) | ( n15665 & n15678 ) | ( n15670 & n15678 ) ;
  assign n16284 = ( n16282 & ~n15678 ) | ( n16282 & n16283 ) | ( ~n15678 & n16283 ) ;
  assign n16285 = ( n15665 & ~n16283 ) | ( n15665 & n16282 ) | ( ~n16283 & n16282 ) ;
  assign n16286 = ( n15670 & ~n16284 ) | ( n15670 & n16285 ) | ( ~n16284 & n16285 ) ;
  assign n16287 = ( n16281 & ~n6781 ) | ( n16281 & n16286 ) | ( ~n6781 & n16286 ) ;
  assign n16288 = n6399 | n16287 ;
  assign n16289 = n15698 | n16070 ;
  assign n16290 = ( n15685 & ~n15694 ) | ( n15685 & n15698 ) | ( ~n15694 & n15698 ) ;
  assign n16291 = ( n15694 & n16289 ) | ( n15694 & n16290 ) | ( n16289 & n16290 ) ;
  assign n16292 = ( n15698 & ~n16290 ) | ( n15698 & n16289 ) | ( ~n16290 & n16289 ) ;
  assign n16293 = ( n15685 & ~n16291 ) | ( n15685 & n16292 ) | ( ~n16291 & n16292 ) ;
  assign n16294 = ~n6781 & n16266 ;
  assign n16295 = n16280 &  n16294 ;
  assign n16296 = n16286 | n16295 ;
  assign n16297 = n16274 &  n16277 ;
  assign n16298 = ( n7169 & n16271 ) | ( n7169 & n16297 ) | ( n16271 & n16297 ) ;
  assign n16299 = ( n6781 & ~n16298 ) | ( n6781 & 1'b0 ) | ( ~n16298 & 1'b0 ) ;
  assign n16300 = ( n6399 & ~n16299 ) | ( n6399 & 1'b0 ) | ( ~n16299 & 1'b0 ) ;
  assign n16301 = n16296 &  n16300 ;
  assign n16302 = n16293 | n16301 ;
  assign n16303 = n16288 &  n16302 ;
  assign n16304 = ( n15687 & ~n16070 ) | ( n15687 & 1'b0 ) | ( ~n16070 & 1'b0 ) ;
  assign n16305 = ( n15687 & n15692 ) | ( n15687 & n15700 ) | ( n15692 & n15700 ) ;
  assign n16306 = ( n16304 & ~n15700 ) | ( n16304 & n16305 ) | ( ~n15700 & n16305 ) ;
  assign n16307 = ( n15687 & ~n16305 ) | ( n15687 & n16304 ) | ( ~n16305 & n16304 ) ;
  assign n16308 = ( n15692 & ~n16306 ) | ( n15692 & n16307 ) | ( ~n16306 & n16307 ) ;
  assign n16309 = ( n16303 & ~n6032 ) | ( n16303 & n16308 ) | ( ~n6032 & n16308 ) ;
  assign n16310 = n5672 | n16309 ;
  assign n16311 = n15720 | n16070 ;
  assign n16312 = ( n15707 & ~n15716 ) | ( n15707 & n15720 ) | ( ~n15716 & n15720 ) ;
  assign n16313 = ( n15716 & n16311 ) | ( n15716 & n16312 ) | ( n16311 & n16312 ) ;
  assign n16314 = ( n15720 & ~n16312 ) | ( n15720 & n16311 ) | ( ~n16312 & n16311 ) ;
  assign n16315 = ( n15707 & ~n16313 ) | ( n15707 & n16314 ) | ( ~n16313 & n16314 ) ;
  assign n16316 = ~n6032 & n16288 ;
  assign n16317 = n16302 &  n16316 ;
  assign n16318 = n16308 | n16317 ;
  assign n16319 = ( n16296 & ~n16299 ) | ( n16296 & 1'b0 ) | ( ~n16299 & 1'b0 ) ;
  assign n16320 = ( n6399 & n16293 ) | ( n6399 & n16319 ) | ( n16293 & n16319 ) ;
  assign n16321 = ( n6032 & ~n16320 ) | ( n6032 & 1'b0 ) | ( ~n16320 & 1'b0 ) ;
  assign n16322 = ( n5672 & ~n16321 ) | ( n5672 & 1'b0 ) | ( ~n16321 & 1'b0 ) ;
  assign n16323 = n16318 &  n16322 ;
  assign n16324 = n16315 | n16323 ;
  assign n16325 = n16310 &  n16324 ;
  assign n16326 = ( n15709 & ~n16070 ) | ( n15709 & 1'b0 ) | ( ~n16070 & 1'b0 ) ;
  assign n16327 = ( n15709 & n15714 ) | ( n15709 & n15722 ) | ( n15714 & n15722 ) ;
  assign n16328 = ( n16326 & ~n15722 ) | ( n16326 & n16327 ) | ( ~n15722 & n16327 ) ;
  assign n16329 = ( n15709 & ~n16327 ) | ( n15709 & n16326 ) | ( ~n16327 & n16326 ) ;
  assign n16330 = ( n15714 & ~n16328 ) | ( n15714 & n16329 ) | ( ~n16328 & n16329 ) ;
  assign n16331 = ( n16325 & ~n5327 ) | ( n16325 & n16330 ) | ( ~n5327 & n16330 ) ;
  assign n16332 = ( n4990 & ~n16331 ) | ( n4990 & 1'b0 ) | ( ~n16331 & 1'b0 ) ;
  assign n16333 = n15742 | n16070 ;
  assign n16334 = ( n15729 & ~n15738 ) | ( n15729 & n15742 ) | ( ~n15738 & n15742 ) ;
  assign n16335 = ( n15738 & n16333 ) | ( n15738 & n16334 ) | ( n16333 & n16334 ) ;
  assign n16336 = ( n15742 & ~n16334 ) | ( n15742 & n16333 ) | ( ~n16334 & n16333 ) ;
  assign n16337 = ( n15729 & ~n16335 ) | ( n15729 & n16336 ) | ( ~n16335 & n16336 ) ;
  assign n16338 = ~n5327 & n16310 ;
  assign n16339 = n16324 &  n16338 ;
  assign n16340 = n16330 | n16339 ;
  assign n16341 = ( n16318 & ~n16321 ) | ( n16318 & 1'b0 ) | ( ~n16321 & 1'b0 ) ;
  assign n16342 = ( n5672 & n16315 ) | ( n5672 & n16341 ) | ( n16315 & n16341 ) ;
  assign n16343 = ( n5327 & ~n16342 ) | ( n5327 & 1'b0 ) | ( ~n16342 & 1'b0 ) ;
  assign n16344 = n4990 | n16343 ;
  assign n16345 = ( n16340 & ~n16344 ) | ( n16340 & 1'b0 ) | ( ~n16344 & 1'b0 ) ;
  assign n16346 = n16337 | n16345 ;
  assign n16347 = ~n16332 & n16346 ;
  assign n16348 = n15731 | n16070 ;
  assign n16349 = ( n15731 & ~n15744 ) | ( n15731 & n15736 ) | ( ~n15744 & n15736 ) ;
  assign n16350 = ( n15744 & n16348 ) | ( n15744 & n16349 ) | ( n16348 & n16349 ) ;
  assign n16351 = ( n15731 & ~n16349 ) | ( n15731 & n16348 ) | ( ~n16349 & n16348 ) ;
  assign n16352 = ( n15736 & ~n16350 ) | ( n15736 & n16351 ) | ( ~n16350 & n16351 ) ;
  assign n16353 = ( n4668 & ~n16347 ) | ( n4668 & n16352 ) | ( ~n16347 & n16352 ) ;
  assign n16354 = n4353 &  n16353 ;
  assign n16356 = ( n15760 & ~n15751 ) | ( n15760 & n15764 ) | ( ~n15751 & n15764 ) ;
  assign n16355 = n15764 | n16070 ;
  assign n16358 = ( n15764 & ~n16356 ) | ( n15764 & n16355 ) | ( ~n16356 & n16355 ) ;
  assign n16357 = ( n16355 & ~n15760 ) | ( n16355 & n16356 ) | ( ~n15760 & n16356 ) ;
  assign n16359 = ( n15751 & ~n16358 ) | ( n15751 & n16357 ) | ( ~n16358 & n16357 ) ;
  assign n16360 = n4668 | n16332 ;
  assign n16361 = ( n16346 & ~n16360 ) | ( n16346 & 1'b0 ) | ( ~n16360 & 1'b0 ) ;
  assign n16362 = ( n16352 & ~n16361 ) | ( n16352 & 1'b0 ) | ( ~n16361 & 1'b0 ) ;
  assign n16363 = ( n16340 & ~n16343 ) | ( n16340 & 1'b0 ) | ( ~n16343 & 1'b0 ) ;
  assign n16364 = ( n16337 & ~n4990 ) | ( n16337 & n16363 ) | ( ~n4990 & n16363 ) ;
  assign n16365 = ( n4668 & ~n16364 ) | ( n4668 & 1'b0 ) | ( ~n16364 & 1'b0 ) ;
  assign n16366 = n4353 | n16365 ;
  assign n16367 = n16362 | n16366 ;
  assign n16368 = n16359 &  n16367 ;
  assign n16369 = n16354 | n16368 ;
  assign n16370 = n15753 | n16070 ;
  assign n16371 = ( n15753 & n15758 ) | ( n15753 & n15766 ) | ( n15758 & n15766 ) ;
  assign n16372 = ( n16370 & ~n15766 ) | ( n16370 & n16371 ) | ( ~n15766 & n16371 ) ;
  assign n16373 = ( n15753 & ~n16371 ) | ( n15753 & n16370 ) | ( ~n16371 & n16370 ) ;
  assign n16374 = ( n15758 & ~n16372 ) | ( n15758 & n16373 ) | ( ~n16372 & n16373 ) ;
  assign n16375 = ( n4053 & n16369 ) | ( n4053 & n16374 ) | ( n16369 & n16374 ) ;
  assign n16376 = n3760 &  n16375 ;
  assign n16378 = ( n15782 & ~n15773 ) | ( n15782 & n15786 ) | ( ~n15773 & n15786 ) ;
  assign n16377 = n15786 | n16070 ;
  assign n16380 = ( n15786 & ~n16378 ) | ( n15786 & n16377 ) | ( ~n16378 & n16377 ) ;
  assign n16379 = ( n16377 & ~n15782 ) | ( n16377 & n16378 ) | ( ~n15782 & n16378 ) ;
  assign n16381 = ( n15773 & ~n16380 ) | ( n15773 & n16379 ) | ( ~n16380 & n16379 ) ;
  assign n16382 = n4053 | n16354 ;
  assign n16383 = n16368 | n16382 ;
  assign n16384 = n16374 &  n16383 ;
  assign n16385 = n16362 | n16365 ;
  assign n16386 = ( n4353 & n16359 ) | ( n4353 & n16385 ) | ( n16359 & n16385 ) ;
  assign n16387 = n4053 &  n16386 ;
  assign n16388 = n3760 | n16387 ;
  assign n16389 = n16384 | n16388 ;
  assign n16390 = n16381 &  n16389 ;
  assign n16391 = n16376 | n16390 ;
  assign n16392 = n15775 | n16070 ;
  assign n16393 = ( n15775 & n15780 ) | ( n15775 & n15788 ) | ( n15780 & n15788 ) ;
  assign n16394 = ( n16392 & ~n15788 ) | ( n16392 & n16393 ) | ( ~n15788 & n16393 ) ;
  assign n16395 = ( n15775 & ~n16393 ) | ( n15775 & n16392 ) | ( ~n16393 & n16392 ) ;
  assign n16396 = ( n15780 & ~n16394 ) | ( n15780 & n16395 ) | ( ~n16394 & n16395 ) ;
  assign n16397 = ( n3482 & n16391 ) | ( n3482 & n16396 ) | ( n16391 & n16396 ) ;
  assign n16398 = n3211 &  n16397 ;
  assign n16399 = n15808 | n16070 ;
  assign n16400 = ( n15795 & n15804 ) | ( n15795 & n15808 ) | ( n15804 & n15808 ) ;
  assign n16401 = ( n16399 & ~n15804 ) | ( n16399 & n16400 ) | ( ~n15804 & n16400 ) ;
  assign n16402 = ( n15808 & ~n16400 ) | ( n15808 & n16399 ) | ( ~n16400 & n16399 ) ;
  assign n16403 = ( n15795 & ~n16401 ) | ( n15795 & n16402 ) | ( ~n16401 & n16402 ) ;
  assign n16404 = n3482 | n16376 ;
  assign n16405 = n16390 | n16404 ;
  assign n16406 = n16396 &  n16405 ;
  assign n16407 = n16384 | n16387 ;
  assign n16408 = ( n3760 & n16381 ) | ( n3760 & n16407 ) | ( n16381 & n16407 ) ;
  assign n16409 = n3482 &  n16408 ;
  assign n16410 = n3211 | n16409 ;
  assign n16411 = n16406 | n16410 ;
  assign n16412 = ~n16403 & n16411 ;
  assign n16413 = n16398 | n16412 ;
  assign n16419 = ( n2955 & ~n16418 ) | ( n2955 & n16413 ) | ( ~n16418 & n16413 ) ;
  assign n16420 = n2706 &  n16419 ;
  assign n16422 = ( n15826 & ~n15817 ) | ( n15826 & n15830 ) | ( ~n15817 & n15830 ) ;
  assign n16421 = n15830 | n16070 ;
  assign n16424 = ( n15830 & ~n16422 ) | ( n15830 & n16421 ) | ( ~n16422 & n16421 ) ;
  assign n16423 = ( n16421 & ~n15826 ) | ( n16421 & n16422 ) | ( ~n15826 & n16422 ) ;
  assign n16425 = ( n15817 & ~n16424 ) | ( n15817 & n16423 ) | ( ~n16424 & n16423 ) ;
  assign n16426 = n2955 | n16398 ;
  assign n16427 = n16412 | n16426 ;
  assign n16428 = ~n16418 & n16427 ;
  assign n16429 = n16406 | n16409 ;
  assign n16430 = ( n3211 & ~n16403 ) | ( n3211 & n16429 ) | ( ~n16403 & n16429 ) ;
  assign n16431 = n2955 &  n16430 ;
  assign n16432 = n2706 | n16431 ;
  assign n16433 = n16428 | n16432 ;
  assign n16434 = n16425 &  n16433 ;
  assign n16435 = n16420 | n16434 ;
  assign n16441 = ( n2472 & ~n16440 ) | ( n2472 & n16435 ) | ( ~n16440 & n16435 ) ;
  assign n16442 = n2245 &  n16441 ;
  assign n16444 = ( n15848 & ~n15839 ) | ( n15848 & n15852 ) | ( ~n15839 & n15852 ) ;
  assign n16443 = n15852 | n16070 ;
  assign n16446 = ( n15852 & ~n16444 ) | ( n15852 & n16443 ) | ( ~n16444 & n16443 ) ;
  assign n16445 = ( n16443 & ~n15848 ) | ( n16443 & n16444 ) | ( ~n15848 & n16444 ) ;
  assign n16447 = ( n15839 & ~n16446 ) | ( n15839 & n16445 ) | ( ~n16446 & n16445 ) ;
  assign n16448 = n2472 | n16420 ;
  assign n16449 = n16434 | n16448 ;
  assign n16450 = ~n16440 & n16449 ;
  assign n16451 = n16428 | n16431 ;
  assign n16452 = ( n2706 & n16425 ) | ( n2706 & n16451 ) | ( n16425 & n16451 ) ;
  assign n16453 = n2472 &  n16452 ;
  assign n16454 = n2245 | n16453 ;
  assign n16455 = n16450 | n16454 ;
  assign n16456 = n16447 &  n16455 ;
  assign n16457 = n16442 | n16456 ;
  assign n16458 = n15841 | n16070 ;
  assign n16459 = ( n15841 & n15846 ) | ( n15841 & n15854 ) | ( n15846 & n15854 ) ;
  assign n16460 = ( n16458 & ~n15854 ) | ( n16458 & n16459 ) | ( ~n15854 & n16459 ) ;
  assign n16461 = ( n15841 & ~n16459 ) | ( n15841 & n16458 ) | ( ~n16459 & n16458 ) ;
  assign n16462 = ( n15846 & ~n16460 ) | ( n15846 & n16461 ) | ( ~n16460 & n16461 ) ;
  assign n16463 = ( n16457 & ~n2033 ) | ( n16457 & n16462 ) | ( ~n2033 & n16462 ) ;
  assign n16464 = n1827 &  n16463 ;
  assign n16465 = n15874 | n16070 ;
  assign n16466 = ( n15861 & ~n15870 ) | ( n15861 & n15874 ) | ( ~n15870 & n15874 ) ;
  assign n16467 = ( n15870 & n16465 ) | ( n15870 & n16466 ) | ( n16465 & n16466 ) ;
  assign n16468 = ( n15874 & ~n16466 ) | ( n15874 & n16465 ) | ( ~n16466 & n16465 ) ;
  assign n16469 = ( n15861 & ~n16467 ) | ( n15861 & n16468 ) | ( ~n16467 & n16468 ) ;
  assign n16470 = ( n2033 & ~n16442 ) | ( n2033 & 1'b0 ) | ( ~n16442 & 1'b0 ) ;
  assign n16471 = ~n16456 & n16470 ;
  assign n16472 = ( n16462 & ~n16471 ) | ( n16462 & 1'b0 ) | ( ~n16471 & 1'b0 ) ;
  assign n16473 = n16450 | n16453 ;
  assign n16474 = ( n2245 & n16447 ) | ( n2245 & n16473 ) | ( n16447 & n16473 ) ;
  assign n16475 = ~n2033 & n16474 ;
  assign n16476 = n1827 | n16475 ;
  assign n16477 = n16472 | n16476 ;
  assign n16478 = ~n16469 & n16477 ;
  assign n16479 = n16464 | n16478 ;
  assign n16480 = n15863 | n16070 ;
  assign n16481 = ( n15868 & ~n15863 ) | ( n15868 & n15876 ) | ( ~n15863 & n15876 ) ;
  assign n16483 = ( n15863 & n16480 ) | ( n15863 & n16481 ) | ( n16480 & n16481 ) ;
  assign n16482 = ( n15876 & ~n16481 ) | ( n15876 & n16480 ) | ( ~n16481 & n16480 ) ;
  assign n16484 = ( n15868 & ~n16483 ) | ( n15868 & n16482 ) | ( ~n16483 & n16482 ) ;
  assign n16485 = ( n1636 & ~n16479 ) | ( n1636 & n16484 ) | ( ~n16479 & n16484 ) ;
  assign n16486 = n1452 | n16485 ;
  assign n16488 = ( n15892 & ~n15883 ) | ( n15892 & n15896 ) | ( ~n15883 & n15896 ) ;
  assign n16487 = ( n15896 & ~n16070 ) | ( n15896 & 1'b0 ) | ( ~n16070 & 1'b0 ) ;
  assign n16490 = ( n15896 & ~n16488 ) | ( n15896 & n16487 ) | ( ~n16488 & n16487 ) ;
  assign n16489 = ( n16487 & ~n15892 ) | ( n16487 & n16488 ) | ( ~n15892 & n16488 ) ;
  assign n16491 = ( n15883 & ~n16490 ) | ( n15883 & n16489 ) | ( ~n16490 & n16489 ) ;
  assign n16492 = ( n1636 & ~n16464 ) | ( n1636 & 1'b0 ) | ( ~n16464 & 1'b0 ) ;
  assign n16493 = ~n16478 & n16492 ;
  assign n16494 = n16484 | n16493 ;
  assign n16495 = n16472 | n16475 ;
  assign n16496 = ( n1827 & ~n16469 ) | ( n1827 & n16495 ) | ( ~n16469 & n16495 ) ;
  assign n16497 = ~n1636 & n16496 ;
  assign n16498 = ( n1452 & ~n16497 ) | ( n1452 & 1'b0 ) | ( ~n16497 & 1'b0 ) ;
  assign n16499 = n16494 &  n16498 ;
  assign n16500 = n16491 | n16499 ;
  assign n16501 = n16486 &  n16500 ;
  assign n16502 = ( n15885 & ~n16070 ) | ( n15885 & 1'b0 ) | ( ~n16070 & 1'b0 ) ;
  assign n16503 = ( n15885 & n15890 ) | ( n15885 & n15898 ) | ( n15890 & n15898 ) ;
  assign n16504 = ( n16502 & ~n15898 ) | ( n16502 & n16503 ) | ( ~n15898 & n16503 ) ;
  assign n16505 = ( n15885 & ~n16503 ) | ( n15885 & n16502 ) | ( ~n16503 & n16502 ) ;
  assign n16506 = ( n15890 & ~n16504 ) | ( n15890 & n16505 ) | ( ~n16504 & n16505 ) ;
  assign n16507 = ( n16501 & ~n1283 ) | ( n16501 & n16506 ) | ( ~n1283 & n16506 ) ;
  assign n16508 = n1122 | n16507 ;
  assign n16509 = n15918 | n16070 ;
  assign n16510 = ( n15905 & ~n15914 ) | ( n15905 & n15918 ) | ( ~n15914 & n15918 ) ;
  assign n16511 = ( n15914 & n16509 ) | ( n15914 & n16510 ) | ( n16509 & n16510 ) ;
  assign n16512 = ( n15918 & ~n16510 ) | ( n15918 & n16509 ) | ( ~n16510 & n16509 ) ;
  assign n16513 = ( n15905 & ~n16511 ) | ( n15905 & n16512 ) | ( ~n16511 & n16512 ) ;
  assign n16514 = ~n1283 & n16486 ;
  assign n16515 = n16500 &  n16514 ;
  assign n16516 = n16506 | n16515 ;
  assign n16517 = ( n16494 & ~n16497 ) | ( n16494 & 1'b0 ) | ( ~n16497 & 1'b0 ) ;
  assign n16518 = ( n1452 & n16491 ) | ( n1452 & n16517 ) | ( n16491 & n16517 ) ;
  assign n16519 = ( n1283 & ~n16518 ) | ( n1283 & 1'b0 ) | ( ~n16518 & 1'b0 ) ;
  assign n16520 = ( n1122 & ~n16519 ) | ( n1122 & 1'b0 ) | ( ~n16519 & 1'b0 ) ;
  assign n16521 = n16516 &  n16520 ;
  assign n16522 = n16513 | n16521 ;
  assign n16523 = n16508 &  n16522 ;
  assign n16529 = ( n976 & ~n16528 ) | ( n976 & n16523 ) | ( ~n16528 & n16523 ) ;
  assign n16530 = ( n837 & ~n16529 ) | ( n837 & 1'b0 ) | ( ~n16529 & 1'b0 ) ;
  assign n16568 = ( n15950 & ~n15955 ) | ( n15950 & n16070 ) | ( ~n15955 & n16070 ) ;
  assign n16567 = ~n15963 & n16070 ;
  assign n16569 = ( n16070 & ~n16568 ) | ( n16070 & n16567 ) | ( ~n16568 & n16567 ) ;
  assign n16570 = ( n16567 & ~n15950 ) | ( n16567 & n16568 ) | ( ~n15950 & n16568 ) ;
  assign n16571 = ( n15955 & ~n16569 ) | ( n15955 & n16570 ) | ( ~n16569 & n16570 ) ;
  assign n16536 = n976 &  n16508 ;
  assign n16537 = n16522 &  n16536 ;
  assign n16538 = ( n16528 & ~n16537 ) | ( n16528 & 1'b0 ) | ( ~n16537 & 1'b0 ) ;
  assign n16539 = ( n16516 & ~n16519 ) | ( n16516 & 1'b0 ) | ( ~n16519 & 1'b0 ) ;
  assign n16540 = ( n1122 & n16513 ) | ( n1122 & n16539 ) | ( n16513 & n16539 ) ;
  assign n16541 = n976 | n16540 ;
  assign n16542 = ~n837 & n16541 ;
  assign n16543 = ~n16538 & n16542 ;
  assign n16544 = n16535 | n16543 ;
  assign n16545 = ~n16530 & n16544 ;
  assign n16546 = ( n15929 & ~n15937 ) | ( n15929 & n15941 ) | ( ~n15937 & n15941 ) ;
  assign n16547 = ( n15937 & n16070 ) | ( n15937 & n16546 ) | ( n16070 & n16546 ) ;
  assign n16548 = ( n15929 & ~n16546 ) | ( n15929 & n16070 ) | ( ~n16546 & n16070 ) ;
  assign n16549 = ( n15941 & ~n16547 ) | ( n15941 & n16548 ) | ( ~n16547 & n16548 ) ;
  assign n16550 = ( n16545 & ~n713 ) | ( n16545 & n16549 ) | ( ~n713 & n16549 ) ;
  assign n16551 = ( n595 & ~n16550 ) | ( n595 & 1'b0 ) | ( ~n16550 & 1'b0 ) ;
  assign n16552 = n15961 | n16070 ;
  assign n16553 = ( n15948 & ~n15957 ) | ( n15948 & n15961 ) | ( ~n15957 & n15961 ) ;
  assign n16554 = ( n15957 & n16552 ) | ( n15957 & n16553 ) | ( n16552 & n16553 ) ;
  assign n16555 = ( n15961 & ~n16553 ) | ( n15961 & n16552 ) | ( ~n16553 & n16552 ) ;
  assign n16556 = ( n15948 & ~n16554 ) | ( n15948 & n16555 ) | ( ~n16554 & n16555 ) ;
  assign n16557 = n713 | n16530 ;
  assign n16558 = ( n16544 & ~n16557 ) | ( n16544 & 1'b0 ) | ( ~n16557 & 1'b0 ) ;
  assign n16559 = n16549 | n16558 ;
  assign n16560 = ~n16538 & n16541 ;
  assign n16561 = ( n16535 & ~n837 ) | ( n16535 & n16560 ) | ( ~n837 & n16560 ) ;
  assign n16562 = ( n713 & ~n16561 ) | ( n713 & 1'b0 ) | ( ~n16561 & 1'b0 ) ;
  assign n16563 = n595 | n16562 ;
  assign n16564 = ( n16559 & ~n16563 ) | ( n16559 & 1'b0 ) | ( ~n16563 & 1'b0 ) ;
  assign n16565 = ( n16556 & ~n16564 ) | ( n16556 & 1'b0 ) | ( ~n16564 & 1'b0 ) ;
  assign n16566 = n16551 | n16565 ;
  assign n16572 = ( n492 & ~n16571 ) | ( n492 & n16566 ) | ( ~n16571 & n16566 ) ;
  assign n16573 = n396 &  n16572 ;
  assign n16574 = n15983 | n16070 ;
  assign n16575 = ( n15970 & n15979 ) | ( n15970 & n15983 ) | ( n15979 & n15983 ) ;
  assign n16576 = ( n16574 & ~n15979 ) | ( n16574 & n16575 ) | ( ~n15979 & n16575 ) ;
  assign n16577 = ( n15983 & ~n16575 ) | ( n15983 & n16574 ) | ( ~n16575 & n16574 ) ;
  assign n16578 = ( n15970 & ~n16576 ) | ( n15970 & n16577 ) | ( ~n16576 & n16577 ) ;
  assign n16579 = n492 | n16551 ;
  assign n16580 = n16565 | n16579 ;
  assign n16581 = ~n16571 & n16580 ;
  assign n16582 = ( n16559 & ~n16562 ) | ( n16559 & 1'b0 ) | ( ~n16562 & 1'b0 ) ;
  assign n16583 = ( n595 & ~n16582 ) | ( n595 & n16556 ) | ( ~n16582 & n16556 ) ;
  assign n16584 = n492 &  n16583 ;
  assign n16585 = n396 | n16584 ;
  assign n16586 = n16581 | n16585 ;
  assign n16587 = n16578 &  n16586 ;
  assign n16588 = n16573 | n16587 ;
  assign n16590 = ( n15972 & ~n15977 ) | ( n15972 & n16070 ) | ( ~n15977 & n16070 ) ;
  assign n16589 = ~n15985 & n16070 ;
  assign n16591 = ( n16070 & ~n16590 ) | ( n16070 & n16589 ) | ( ~n16590 & n16589 ) ;
  assign n16592 = ( n16589 & ~n15972 ) | ( n16589 & n16590 ) | ( ~n15972 & n16590 ) ;
  assign n16593 = ( n15977 & ~n16591 ) | ( n15977 & n16592 ) | ( ~n16591 & n16592 ) ;
  assign n16594 = ( n315 & n16588 ) | ( n315 & n16593 ) | ( n16588 & n16593 ) ;
  assign n16595 = n240 &  n16594 ;
  assign n16597 = ( n16001 & ~n15992 ) | ( n16001 & n16005 ) | ( ~n15992 & n16005 ) ;
  assign n16596 = n16005 | n16070 ;
  assign n16599 = ( n16005 & ~n16597 ) | ( n16005 & n16596 ) | ( ~n16597 & n16596 ) ;
  assign n16598 = ( n16596 & ~n16001 ) | ( n16596 & n16597 ) | ( ~n16001 & n16597 ) ;
  assign n16600 = ( n15992 & ~n16599 ) | ( n15992 & n16598 ) | ( ~n16599 & n16598 ) ;
  assign n16601 = n315 | n16573 ;
  assign n16602 = n16587 | n16601 ;
  assign n16603 = n16593 &  n16602 ;
  assign n16604 = n16581 | n16584 ;
  assign n16605 = ( n396 & n16578 ) | ( n396 & n16604 ) | ( n16578 & n16604 ) ;
  assign n16606 = n315 &  n16605 ;
  assign n16607 = n240 | n16606 ;
  assign n16608 = n16603 | n16607 ;
  assign n16609 = ~n16600 & n16608 ;
  assign n16610 = n16595 | n16609 ;
  assign n16612 = ( n15994 & ~n15999 ) | ( n15994 & n16070 ) | ( ~n15999 & n16070 ) ;
  assign n16611 = ~n16007 & n16070 ;
  assign n16613 = ( n16070 & ~n16612 ) | ( n16070 & n16611 ) | ( ~n16612 & n16611 ) ;
  assign n16614 = ( n16611 & ~n15994 ) | ( n16611 & n16612 ) | ( ~n15994 & n16612 ) ;
  assign n16615 = ( n15999 & ~n16613 ) | ( n15999 & n16614 ) | ( ~n16613 & n16614 ) ;
  assign n16616 = ( n181 & n16610 ) | ( n181 & n16615 ) | ( n16610 & n16615 ) ;
  assign n16617 = ~n145 & n16616 ;
  assign n16618 = n16027 | n16070 ;
  assign n16619 = ( n16014 & n16023 ) | ( n16014 & n16027 ) | ( n16023 & n16027 ) ;
  assign n16620 = ( n16618 & ~n16023 ) | ( n16618 & n16619 ) | ( ~n16023 & n16619 ) ;
  assign n16621 = ( n16027 & ~n16619 ) | ( n16027 & n16618 ) | ( ~n16619 & n16618 ) ;
  assign n16622 = ( n16014 & ~n16620 ) | ( n16014 & n16621 ) | ( ~n16620 & n16621 ) ;
  assign n16623 = n181 | n16595 ;
  assign n16624 = n16609 | n16623 ;
  assign n16625 = n16615 &  n16624 ;
  assign n16626 = n16603 | n16606 ;
  assign n16627 = ( n240 & ~n16600 ) | ( n240 & n16626 ) | ( ~n16600 & n16626 ) ;
  assign n16628 = n181 &  n16627 ;
  assign n16629 = ( n145 & ~n16628 ) | ( n145 & 1'b0 ) | ( ~n16628 & 1'b0 ) ;
  assign n16630 = ~n16625 & n16629 ;
  assign n16631 = n16622 | n16630 ;
  assign n16632 = ~n16617 & n16631 ;
  assign n16633 = n16016 | n16070 ;
  assign n16634 = ( n16016 & ~n16029 ) | ( n16016 & n16021 ) | ( ~n16029 & n16021 ) ;
  assign n16635 = ( n16029 & n16633 ) | ( n16029 & n16634 ) | ( n16633 & n16634 ) ;
  assign n16636 = ( n16016 & ~n16634 ) | ( n16016 & n16633 ) | ( ~n16634 & n16633 ) ;
  assign n16637 = ( n16021 & ~n16635 ) | ( n16021 & n16636 ) | ( ~n16635 & n16636 ) ;
  assign n16638 = ( n16632 & ~n150 ) | ( n16632 & n16637 ) | ( ~n150 & n16637 ) ;
  assign n16639 = n16036 | n16052 ;
  assign n16640 = ( n16055 & ~n16639 ) | ( n16055 & n16070 ) | ( ~n16639 & n16070 ) ;
  assign n16641 = ~n16055 & n16640 ;
  assign n16642 = n16052 | n16055 ;
  assign n16643 = n16070 | n16642 ;
  assign n16644 = ( n16036 & ~n16643 ) | ( n16036 & n16642 ) | ( ~n16643 & n16642 ) ;
  assign n16645 = n16641 | n16644 ;
  assign n16646 = n16037 &  n16044 ;
  assign n16647 = ~n16070 & n16646 ;
  assign n16648 = ( n16058 & ~n16646 ) | ( n16058 & n16647 ) | ( ~n16646 & n16647 ) ;
  assign n16649 = n16645 &  n16648 ;
  assign n16650 = n16638 &  n16649 ;
  assign n16651 = ( n133 & ~n16650 ) | ( n133 & n16649 ) | ( ~n16650 & n16649 ) ;
  assign n16654 = n16625 | n16628 ;
  assign n16655 = ( n145 & ~n16654 ) | ( n145 & n16622 ) | ( ~n16654 & n16622 ) ;
  assign n16656 = ( n150 & ~n16655 ) | ( n150 & 1'b0 ) | ( ~n16655 & 1'b0 ) ;
  assign n16657 = n16645 | n16656 ;
  assign n16652 = n150 | n16617 ;
  assign n16653 = ( n16631 & ~n16652 ) | ( n16631 & 1'b0 ) | ( ~n16652 & 1'b0 ) ;
  assign n16658 = ~n16637 & n16653 ;
  assign n16659 = ( n16637 & ~n16657 ) | ( n16637 & n16658 ) | ( ~n16657 & n16658 ) ;
  assign n16661 = ( n133 & n16037 ) | ( n133 & n16044 ) | ( n16037 & n16044 ) ;
  assign n16660 = ( n16037 & ~n16070 ) | ( n16037 & n16044 ) | ( ~n16070 & n16044 ) ;
  assign n16662 = ( n16044 & ~n16660 ) | ( n16044 & 1'b0 ) | ( ~n16660 & 1'b0 ) ;
  assign n16663 = ( n16661 & ~n16044 ) | ( n16661 & n16662 ) | ( ~n16044 & n16662 ) ;
  assign n16664 = n16040 | n16067 ;
  assign n16665 = ( n16062 & ~n16043 ) | ( n16062 & n16664 ) | ( ~n16043 & n16664 ) ;
  assign n16666 = n16043 | n16665 ;
  assign n16667 = ( n16050 & ~n16058 ) | ( n16050 & n16666 ) | ( ~n16058 & n16666 ) ;
  assign n16668 = ( n16050 & ~n16667 ) | ( n16050 & 1'b0 ) | ( ~n16667 & 1'b0 ) ;
  assign n16669 = n16663 | n16668 ;
  assign n16670 = n16659 | n16669 ;
  assign n16671 = ~n16651 |  n16670 ;
  assign n17154 = n16530 | n16671 ;
  assign n17155 = ( n16535 & ~n16530 ) | ( n16535 & n16543 ) | ( ~n16530 & n16543 ) ;
  assign n17157 = ( n16530 & n17154 ) | ( n16530 & n17155 ) | ( n17154 & n17155 ) ;
  assign n17156 = ( n16543 & ~n17155 ) | ( n16543 & n17154 ) | ( ~n17155 & n17154 ) ;
  assign n17158 = ( n16535 & ~n17157 ) | ( n16535 & n17156 ) | ( ~n17157 & n17156 ) ;
  assign n17132 = ( n16508 & ~n16671 ) | ( n16508 & 1'b0 ) | ( ~n16671 & 1'b0 ) ;
  assign n17133 = ( n16508 & n16513 ) | ( n16508 & n16521 ) | ( n16513 & n16521 ) ;
  assign n17134 = ( n17132 & ~n16521 ) | ( n17132 & n17133 ) | ( ~n16521 & n17133 ) ;
  assign n17135 = ( n16508 & ~n17133 ) | ( n16508 & n17132 ) | ( ~n17133 & n17132 ) ;
  assign n17136 = ( n16513 & ~n17134 ) | ( n16513 & n17135 ) | ( ~n17134 & n17135 ) ;
  assign n17117 = n16519 | n16671 ;
  assign n17118 = ( n16506 & ~n16515 ) | ( n16506 & n16519 ) | ( ~n16515 & n16519 ) ;
  assign n17119 = ( n16515 & n17117 ) | ( n16515 & n17118 ) | ( n17117 & n17118 ) ;
  assign n17120 = ( n16519 & ~n17118 ) | ( n16519 & n17117 ) | ( ~n17118 & n17117 ) ;
  assign n17121 = ( n16506 & ~n17119 ) | ( n16506 & n17120 ) | ( ~n17119 & n17120 ) ;
  assign n17110 = ( n16486 & ~n16671 ) | ( n16486 & 1'b0 ) | ( ~n16671 & 1'b0 ) ;
  assign n17111 = ( n16486 & n16491 ) | ( n16486 & n16499 ) | ( n16491 & n16499 ) ;
  assign n17112 = ( n17110 & ~n16499 ) | ( n17110 & n17111 ) | ( ~n16499 & n17111 ) ;
  assign n17113 = ( n16486 & ~n17111 ) | ( n16486 & n17110 ) | ( ~n17111 & n17110 ) ;
  assign n17114 = ( n16491 & ~n17112 ) | ( n16491 & n17113 ) | ( ~n17112 & n17113 ) ;
  assign n17095 = n16497 | n16671 ;
  assign n17096 = ( n16484 & ~n16493 ) | ( n16484 & n16497 ) | ( ~n16493 & n16497 ) ;
  assign n17097 = ( n16493 & n17095 ) | ( n16493 & n17096 ) | ( n17095 & n17096 ) ;
  assign n17098 = ( n16497 & ~n17096 ) | ( n16497 & n17095 ) | ( ~n17096 & n17095 ) ;
  assign n17099 = ( n16484 & ~n17097 ) | ( n16484 & n17098 ) | ( ~n17097 & n17098 ) ;
  assign n17089 = ( n16464 & ~n16469 ) | ( n16464 & n16477 ) | ( ~n16469 & n16477 ) ;
  assign n17088 = n16464 | n16671 ;
  assign n17091 = ( n16464 & ~n17089 ) | ( n16464 & n17088 ) | ( ~n17089 & n17088 ) ;
  assign n17090 = ( n17088 & ~n16477 ) | ( n17088 & n17089 ) | ( ~n16477 & n17089 ) ;
  assign n17092 = ( n16469 & ~n17091 ) | ( n16469 & n17090 ) | ( ~n17091 & n17090 ) ;
  assign n17073 = n16475 | n16671 ;
  assign n17074 = ( n16462 & ~n16475 ) | ( n16462 & n16471 ) | ( ~n16475 & n16471 ) ;
  assign n17076 = ( n16475 & n17073 ) | ( n16475 & n17074 ) | ( n17073 & n17074 ) ;
  assign n17075 = ( n16471 & ~n17074 ) | ( n16471 & n17073 ) | ( ~n17074 & n17073 ) ;
  assign n17077 = ( n16462 & ~n17076 ) | ( n16462 & n17075 ) | ( ~n17076 & n17075 ) ;
  assign n17066 = n16442 | n16671 ;
  assign n17067 = ( n16442 & n16447 ) | ( n16442 & n16455 ) | ( n16447 & n16455 ) ;
  assign n17068 = ( n17066 & ~n16455 ) | ( n17066 & n17067 ) | ( ~n16455 & n17067 ) ;
  assign n17069 = ( n16442 & ~n17067 ) | ( n16442 & n17066 ) | ( ~n17067 & n17066 ) ;
  assign n17070 = ( n16447 & ~n17068 ) | ( n16447 & n17069 ) | ( ~n17068 & n17069 ) ;
  assign n17051 = n16453 | n16671 ;
  assign n17052 = ( n16440 & n16449 ) | ( n16440 & n16453 ) | ( n16449 & n16453 ) ;
  assign n17053 = ( n17051 & ~n16449 ) | ( n17051 & n17052 ) | ( ~n16449 & n17052 ) ;
  assign n17054 = ( n16453 & ~n17052 ) | ( n16453 & n17051 ) | ( ~n17052 & n17051 ) ;
  assign n17055 = ( n16440 & ~n17053 ) | ( n16440 & n17054 ) | ( ~n17053 & n17054 ) ;
  assign n17044 = n16420 | n16671 ;
  assign n17045 = ( n16420 & n16425 ) | ( n16420 & n16433 ) | ( n16425 & n16433 ) ;
  assign n17046 = ( n17044 & ~n16433 ) | ( n17044 & n17045 ) | ( ~n16433 & n17045 ) ;
  assign n17047 = ( n16420 & ~n17045 ) | ( n16420 & n17044 ) | ( ~n17045 & n17044 ) ;
  assign n17048 = ( n16425 & ~n17046 ) | ( n16425 & n17047 ) | ( ~n17046 & n17047 ) ;
  assign n17029 = n16431 | n16671 ;
  assign n17030 = ( n16418 & n16427 ) | ( n16418 & n16431 ) | ( n16427 & n16431 ) ;
  assign n17031 = ( n17029 & ~n16427 ) | ( n17029 & n17030 ) | ( ~n16427 & n17030 ) ;
  assign n17032 = ( n16431 & ~n17030 ) | ( n16431 & n17029 ) | ( ~n17030 & n17029 ) ;
  assign n17033 = ( n16418 & ~n17031 ) | ( n16418 & n17032 ) | ( ~n17031 & n17032 ) ;
  assign n17023 = ( n16398 & ~n16403 ) | ( n16398 & n16411 ) | ( ~n16403 & n16411 ) ;
  assign n17022 = n16398 | n16671 ;
  assign n17025 = ( n16398 & ~n17023 ) | ( n16398 & n17022 ) | ( ~n17023 & n17022 ) ;
  assign n17024 = ( n17022 & ~n16411 ) | ( n17022 & n17023 ) | ( ~n16411 & n17023 ) ;
  assign n17026 = ( n16403 & ~n17025 ) | ( n16403 & n17024 ) | ( ~n17025 & n17024 ) ;
  assign n17008 = ( n16405 & ~n16396 ) | ( n16405 & n16409 ) | ( ~n16396 & n16409 ) ;
  assign n17007 = n16409 | n16671 ;
  assign n17010 = ( n16409 & ~n17008 ) | ( n16409 & n17007 ) | ( ~n17008 & n17007 ) ;
  assign n17009 = ( n17007 & ~n16405 ) | ( n17007 & n17008 ) | ( ~n16405 & n17008 ) ;
  assign n17011 = ( n16396 & ~n17010 ) | ( n16396 & n17009 ) | ( ~n17010 & n17009 ) ;
  assign n17000 = n16376 | n16671 ;
  assign n17001 = ( n16376 & n16381 ) | ( n16376 & n16389 ) | ( n16381 & n16389 ) ;
  assign n17002 = ( n17000 & ~n16389 ) | ( n17000 & n17001 ) | ( ~n16389 & n17001 ) ;
  assign n17003 = ( n16376 & ~n17001 ) | ( n16376 & n17000 ) | ( ~n17001 & n17000 ) ;
  assign n17004 = ( n16381 & ~n17002 ) | ( n16381 & n17003 ) | ( ~n17002 & n17003 ) ;
  assign n16986 = ( n16383 & ~n16374 ) | ( n16383 & n16387 ) | ( ~n16374 & n16387 ) ;
  assign n16985 = n16387 | n16671 ;
  assign n16988 = ( n16387 & ~n16986 ) | ( n16387 & n16985 ) | ( ~n16986 & n16985 ) ;
  assign n16987 = ( n16985 & ~n16383 ) | ( n16985 & n16986 ) | ( ~n16383 & n16986 ) ;
  assign n16989 = ( n16374 & ~n16988 ) | ( n16374 & n16987 ) | ( ~n16988 & n16987 ) ;
  assign n16978 = n16354 | n16671 ;
  assign n16979 = ( n16354 & n16359 ) | ( n16354 & n16367 ) | ( n16359 & n16367 ) ;
  assign n16980 = ( n16978 & ~n16367 ) | ( n16978 & n16979 ) | ( ~n16367 & n16979 ) ;
  assign n16981 = ( n16354 & ~n16979 ) | ( n16354 & n16978 ) | ( ~n16979 & n16978 ) ;
  assign n16982 = ( n16359 & ~n16980 ) | ( n16359 & n16981 ) | ( ~n16980 & n16981 ) ;
  assign n16963 = n16365 | n16671 ;
  assign n16964 = ( n16352 & ~n16365 ) | ( n16352 & n16361 ) | ( ~n16365 & n16361 ) ;
  assign n16966 = ( n16365 & n16963 ) | ( n16365 & n16964 ) | ( n16963 & n16964 ) ;
  assign n16965 = ( n16361 & ~n16964 ) | ( n16361 & n16963 ) | ( ~n16964 & n16963 ) ;
  assign n16967 = ( n16352 & ~n16966 ) | ( n16352 & n16965 ) | ( ~n16966 & n16965 ) ;
  assign n16956 = n16332 | n16671 ;
  assign n16957 = ( n16337 & ~n16332 ) | ( n16337 & n16345 ) | ( ~n16332 & n16345 ) ;
  assign n16959 = ( n16332 & n16956 ) | ( n16332 & n16957 ) | ( n16956 & n16957 ) ;
  assign n16958 = ( n16345 & ~n16957 ) | ( n16345 & n16956 ) | ( ~n16957 & n16956 ) ;
  assign n16960 = ( n16337 & ~n16959 ) | ( n16337 & n16958 ) | ( ~n16959 & n16958 ) ;
  assign n16941 = n16343 | n16671 ;
  assign n16942 = ( n16330 & ~n16339 ) | ( n16330 & n16343 ) | ( ~n16339 & n16343 ) ;
  assign n16943 = ( n16339 & n16941 ) | ( n16339 & n16942 ) | ( n16941 & n16942 ) ;
  assign n16944 = ( n16343 & ~n16942 ) | ( n16343 & n16941 ) | ( ~n16942 & n16941 ) ;
  assign n16945 = ( n16330 & ~n16943 ) | ( n16330 & n16944 ) | ( ~n16943 & n16944 ) ;
  assign n16934 = ( n16310 & ~n16671 ) | ( n16310 & 1'b0 ) | ( ~n16671 & 1'b0 ) ;
  assign n16935 = ( n16310 & n16315 ) | ( n16310 & n16323 ) | ( n16315 & n16323 ) ;
  assign n16936 = ( n16934 & ~n16323 ) | ( n16934 & n16935 ) | ( ~n16323 & n16935 ) ;
  assign n16937 = ( n16310 & ~n16935 ) | ( n16310 & n16934 ) | ( ~n16935 & n16934 ) ;
  assign n16938 = ( n16315 & ~n16936 ) | ( n16315 & n16937 ) | ( ~n16936 & n16937 ) ;
  assign n16919 = n16321 | n16671 ;
  assign n16920 = ( n16308 & ~n16317 ) | ( n16308 & n16321 ) | ( ~n16317 & n16321 ) ;
  assign n16921 = ( n16317 & n16919 ) | ( n16317 & n16920 ) | ( n16919 & n16920 ) ;
  assign n16922 = ( n16321 & ~n16920 ) | ( n16321 & n16919 ) | ( ~n16920 & n16919 ) ;
  assign n16923 = ( n16308 & ~n16921 ) | ( n16308 & n16922 ) | ( ~n16921 & n16922 ) ;
  assign n16912 = ( n16288 & ~n16671 ) | ( n16288 & 1'b0 ) | ( ~n16671 & 1'b0 ) ;
  assign n16913 = ( n16288 & n16293 ) | ( n16288 & n16301 ) | ( n16293 & n16301 ) ;
  assign n16914 = ( n16912 & ~n16301 ) | ( n16912 & n16913 ) | ( ~n16301 & n16913 ) ;
  assign n16915 = ( n16288 & ~n16913 ) | ( n16288 & n16912 ) | ( ~n16913 & n16912 ) ;
  assign n16916 = ( n16293 & ~n16914 ) | ( n16293 & n16915 ) | ( ~n16914 & n16915 ) ;
  assign n16897 = n16299 | n16671 ;
  assign n16898 = ( n16286 & ~n16295 ) | ( n16286 & n16299 ) | ( ~n16295 & n16299 ) ;
  assign n16899 = ( n16295 & n16897 ) | ( n16295 & n16898 ) | ( n16897 & n16898 ) ;
  assign n16900 = ( n16299 & ~n16898 ) | ( n16299 & n16897 ) | ( ~n16898 & n16897 ) ;
  assign n16901 = ( n16286 & ~n16899 ) | ( n16286 & n16900 ) | ( ~n16899 & n16900 ) ;
  assign n16890 = ( n16266 & ~n16671 ) | ( n16266 & 1'b0 ) | ( ~n16671 & 1'b0 ) ;
  assign n16891 = ( n16266 & n16271 ) | ( n16266 & n16279 ) | ( n16271 & n16279 ) ;
  assign n16892 = ( n16890 & ~n16279 ) | ( n16890 & n16891 ) | ( ~n16279 & n16891 ) ;
  assign n16893 = ( n16266 & ~n16891 ) | ( n16266 & n16890 ) | ( ~n16891 & n16890 ) ;
  assign n16894 = ( n16271 & ~n16892 ) | ( n16271 & n16893 ) | ( ~n16892 & n16893 ) ;
  assign n16876 = ( n16273 & ~n16264 ) | ( n16273 & n16277 ) | ( ~n16264 & n16277 ) ;
  assign n16875 = ( n16277 & ~n16671 ) | ( n16277 & 1'b0 ) | ( ~n16671 & 1'b0 ) ;
  assign n16878 = ( n16277 & ~n16876 ) | ( n16277 & n16875 ) | ( ~n16876 & n16875 ) ;
  assign n16877 = ( n16875 & ~n16273 ) | ( n16875 & n16876 ) | ( ~n16273 & n16876 ) ;
  assign n16879 = ( n16264 & ~n16878 ) | ( n16264 & n16877 ) | ( ~n16878 & n16877 ) ;
  assign n16868 = n16244 | n16671 ;
  assign n16869 = ( n16249 & ~n16244 ) | ( n16249 & n16257 ) | ( ~n16244 & n16257 ) ;
  assign n16871 = ( n16244 & n16868 ) | ( n16244 & n16869 ) | ( n16868 & n16869 ) ;
  assign n16870 = ( n16257 & ~n16869 ) | ( n16257 & n16868 ) | ( ~n16869 & n16868 ) ;
  assign n16872 = ( n16249 & ~n16871 ) | ( n16249 & n16870 ) | ( ~n16871 & n16870 ) ;
  assign n16853 = n16255 | n16671 ;
  assign n16854 = ( n16242 & ~n16251 ) | ( n16242 & n16255 ) | ( ~n16251 & n16255 ) ;
  assign n16855 = ( n16251 & n16853 ) | ( n16251 & n16854 ) | ( n16853 & n16854 ) ;
  assign n16856 = ( n16255 & ~n16854 ) | ( n16255 & n16853 ) | ( ~n16854 & n16853 ) ;
  assign n16857 = ( n16242 & ~n16855 ) | ( n16242 & n16856 ) | ( ~n16855 & n16856 ) ;
  assign n16846 = n16235 &  n16671 ;
  assign n16847 = ( n16222 & n16227 ) | ( n16222 & n16671 ) | ( n16227 & n16671 ) ;
  assign n16849 = ( n16846 & ~n16222 ) | ( n16846 & n16847 ) | ( ~n16222 & n16847 ) ;
  assign n16848 = ( n16671 & ~n16847 ) | ( n16671 & n16846 ) | ( ~n16847 & n16846 ) ;
  assign n16850 = ( n16227 & ~n16849 ) | ( n16227 & n16848 ) | ( ~n16849 & n16848 ) ;
  assign n16831 = n16233 | n16671 ;
  assign n16832 = ( n16220 & ~n16233 ) | ( n16220 & n16229 ) | ( ~n16233 & n16229 ) ;
  assign n16834 = ( n16233 & n16831 ) | ( n16233 & n16832 ) | ( n16831 & n16832 ) ;
  assign n16833 = ( n16229 & ~n16832 ) | ( n16229 & n16831 ) | ( ~n16832 & n16831 ) ;
  assign n16835 = ( n16220 & ~n16834 ) | ( n16220 & n16833 ) | ( ~n16834 & n16833 ) ;
  assign n16825 = ( n16200 & ~n16205 ) | ( n16200 & n16213 ) | ( ~n16205 & n16213 ) ;
  assign n16824 = ( n16200 & ~n16671 ) | ( n16200 & 1'b0 ) | ( ~n16671 & 1'b0 ) ;
  assign n16827 = ( n16200 & ~n16825 ) | ( n16200 & n16824 ) | ( ~n16825 & n16824 ) ;
  assign n16826 = ( n16824 & ~n16213 ) | ( n16824 & n16825 ) | ( ~n16213 & n16825 ) ;
  assign n16828 = ( n16205 & ~n16827 ) | ( n16205 & n16826 ) | ( ~n16827 & n16826 ) ;
  assign n16809 = n16211 | n16671 ;
  assign n16810 = ( n16198 & ~n16207 ) | ( n16198 & n16211 ) | ( ~n16207 & n16211 ) ;
  assign n16811 = ( n16207 & n16809 ) | ( n16207 & n16810 ) | ( n16809 & n16810 ) ;
  assign n16812 = ( n16211 & ~n16810 ) | ( n16211 & n16809 ) | ( ~n16810 & n16809 ) ;
  assign n16813 = ( n16198 & ~n16811 ) | ( n16198 & n16812 ) | ( ~n16811 & n16812 ) ;
  assign n16802 = n16178 | n16671 ;
  assign n16803 = ( n16183 & ~n16178 ) | ( n16183 & n16191 ) | ( ~n16178 & n16191 ) ;
  assign n16805 = ( n16178 & n16802 ) | ( n16178 & n16803 ) | ( n16802 & n16803 ) ;
  assign n16804 = ( n16191 & ~n16803 ) | ( n16191 & n16802 ) | ( ~n16803 & n16802 ) ;
  assign n16806 = ( n16183 & ~n16805 ) | ( n16183 & n16804 ) | ( ~n16805 & n16804 ) ;
  assign n16787 = n16189 | n16671 ;
  assign n16788 = ( n16176 & ~n16185 ) | ( n16176 & n16189 ) | ( ~n16185 & n16189 ) ;
  assign n16789 = ( n16185 & n16787 ) | ( n16185 & n16788 ) | ( n16787 & n16788 ) ;
  assign n16790 = ( n16189 & ~n16788 ) | ( n16189 & n16787 ) | ( ~n16788 & n16787 ) ;
  assign n16791 = ( n16176 & ~n16789 ) | ( n16176 & n16790 ) | ( ~n16789 & n16790 ) ;
  assign n16780 = n16169 &  n16671 ;
  assign n16781 = ( n16156 & n16161 ) | ( n16156 & n16671 ) | ( n16161 & n16671 ) ;
  assign n16783 = ( n16780 & ~n16156 ) | ( n16780 & n16781 ) | ( ~n16156 & n16781 ) ;
  assign n16782 = ( n16671 & ~n16781 ) | ( n16671 & n16780 ) | ( ~n16781 & n16780 ) ;
  assign n16784 = ( n16161 & ~n16783 ) | ( n16161 & n16782 ) | ( ~n16783 & n16782 ) ;
  assign n16765 = n16167 | n16671 ;
  assign n16766 = ( n16154 & ~n16167 ) | ( n16154 & n16163 ) | ( ~n16167 & n16163 ) ;
  assign n16768 = ( n16167 & n16765 ) | ( n16167 & n16766 ) | ( n16765 & n16766 ) ;
  assign n16767 = ( n16163 & ~n16766 ) | ( n16163 & n16765 ) | ( ~n16766 & n16765 ) ;
  assign n16769 = ( n16154 & ~n16768 ) | ( n16154 & n16767 ) | ( ~n16768 & n16767 ) ;
  assign n16758 = n16134 | n16671 ;
  assign n16759 = ( n16134 & ~n16147 ) | ( n16134 & n16139 ) | ( ~n16147 & n16139 ) ;
  assign n16760 = ( n16147 & n16758 ) | ( n16147 & n16759 ) | ( n16758 & n16759 ) ;
  assign n16761 = ( n16134 & ~n16759 ) | ( n16134 & n16758 ) | ( ~n16759 & n16758 ) ;
  assign n16762 = ( n16139 & ~n16760 ) | ( n16139 & n16761 ) | ( ~n16760 & n16761 ) ;
  assign n16743 = n16145 | n16671 ;
  assign n16744 = ( n16132 & ~n16141 ) | ( n16132 & n16145 ) | ( ~n16141 & n16145 ) ;
  assign n16745 = ( n16141 & n16743 ) | ( n16141 & n16744 ) | ( n16743 & n16744 ) ;
  assign n16746 = ( n16145 & ~n16744 ) | ( n16145 & n16743 ) | ( ~n16744 & n16743 ) ;
  assign n16747 = ( n16132 & ~n16745 ) | ( n16132 & n16746 ) | ( ~n16745 & n16746 ) ;
  assign n16736 = n16112 | n16671 ;
  assign n16737 = ( n16117 & ~n16112 ) | ( n16117 & n16125 ) | ( ~n16112 & n16125 ) ;
  assign n16739 = ( n16112 & n16736 ) | ( n16112 & n16737 ) | ( n16736 & n16737 ) ;
  assign n16738 = ( n16125 & ~n16737 ) | ( n16125 & n16736 ) | ( ~n16737 & n16736 ) ;
  assign n16740 = ( n16117 & ~n16739 ) | ( n16117 & n16738 ) | ( ~n16739 & n16738 ) ;
  assign n16721 = n16123 | n16671 ;
  assign n16722 = ( n16110 & ~n16119 ) | ( n16110 & n16123 ) | ( ~n16119 & n16123 ) ;
  assign n16723 = ( n16119 & n16721 ) | ( n16119 & n16722 ) | ( n16721 & n16722 ) ;
  assign n16724 = ( n16123 & ~n16722 ) | ( n16123 & n16721 ) | ( ~n16722 & n16721 ) ;
  assign n16725 = ( n16110 & ~n16723 ) | ( n16110 & n16724 ) | ( ~n16723 & n16724 ) ;
  assign n16714 = ( n16086 & ~n16088 ) | ( n16086 & 1'b0 ) | ( ~n16088 & 1'b0 ) ;
  assign n16715 = ( n16088 & ~n16714 ) | ( n16088 & n16098 ) | ( ~n16714 & n16098 ) ;
  assign n16717 = ( n16671 & n16714 ) | ( n16671 & n16715 ) | ( n16714 & n16715 ) ;
  assign n16716 = ( n16088 & ~n16715 ) | ( n16088 & n16671 ) | ( ~n16715 & n16671 ) ;
  assign n16718 = ( n16098 & ~n16717 ) | ( n16098 & n16716 ) | ( ~n16717 & n16716 ) ;
  assign n16698 = ~x22 & n16070 ;
  assign n16699 = ( x23 & ~n16698 ) | ( x23 & 1'b0 ) | ( ~n16698 & 1'b0 ) ;
  assign n16700 = n16089 | n16699 ;
  assign n16695 = ( n16070 & ~x22 ) | ( n16070 & n16081 ) | ( ~x22 & n16081 ) ;
  assign n16696 = x22 &  n16695 ;
  assign n16697 = ( n16076 & ~n16696 ) | ( n16076 & n16081 ) | ( ~n16696 & n16081 ) ;
  assign n16701 = ( n16671 & ~n16700 ) | ( n16671 & n16697 ) | ( ~n16700 & n16697 ) ;
  assign n16703 = ( n16671 & ~n16701 ) | ( n16671 & 1'b0 ) | ( ~n16701 & 1'b0 ) ;
  assign n16702 = ~n16697 & n16701 ;
  assign n16704 = ( n16700 & ~n16703 ) | ( n16700 & n16702 ) | ( ~n16703 & n16702 ) ;
  assign n16684 = ( n16070 & ~n16668 ) | ( n16070 & 1'b0 ) | ( ~n16668 & 1'b0 ) ;
  assign n16685 = ( n16659 & ~n16663 ) | ( n16659 & n16684 ) | ( ~n16663 & n16684 ) ;
  assign n16686 = ~n16659 & n16685 ;
  assign n16687 = n16651 &  n16686 ;
  assign n16683 = ~n16073 & n16671 ;
  assign n16688 = ( n16683 & ~n16687 ) | ( n16683 & 1'b0 ) | ( ~n16687 & 1'b0 ) ;
  assign n16689 = ( x22 & n16687 ) | ( x22 & n16688 ) | ( n16687 & n16688 ) ;
  assign n16690 = x22 | n16687 ;
  assign n16691 = n16683 | n16690 ;
  assign n16692 = ~n16689 & n16691 ;
  assign n16674 = ( x20 & ~n16671 ) | ( x20 & x21 ) | ( ~n16671 & x21 ) ;
  assign n16680 = ( x20 & ~x21 ) | ( x20 & 1'b0 ) | ( ~x21 & 1'b0 ) ;
  assign n16071 = x18 | x19 ;
  assign n16675 = ~x20 & n16071 ;
  assign n16676 = ( x20 & ~n16068 ) | ( x20 & n16675 ) | ( ~n16068 & n16675 ) ;
  assign n16677 = ( n16058 & ~n16050 ) | ( n16058 & n16676 ) | ( ~n16050 & n16676 ) ;
  assign n16678 = n16050 &  n16677 ;
  assign n16679 = ( n16671 & ~x21 ) | ( n16671 & n16678 ) | ( ~x21 & n16678 ) ;
  assign n16681 = ( n16674 & ~n16680 ) | ( n16674 & n16679 ) | ( ~n16680 & n16679 ) ;
  assign n16072 = x20 | n16071 ;
  assign n16672 = x20 &  n16671 ;
  assign n16673 = ( n16070 & ~n16072 ) | ( n16070 & n16672 ) | ( ~n16072 & n16672 ) ;
  assign n16705 = n15484 | n16673 ;
  assign n16706 = ( n16681 & ~n16705 ) | ( n16681 & 1'b0 ) | ( ~n16705 & 1'b0 ) ;
  assign n16707 = n16692 | n16706 ;
  assign n16708 = n16673 &  n16681 ;
  assign n16709 = ( n15484 & ~n16681 ) | ( n15484 & n16708 ) | ( ~n16681 & n16708 ) ;
  assign n16710 = n14905 | n16709 ;
  assign n16711 = ( n16707 & ~n16710 ) | ( n16707 & 1'b0 ) | ( ~n16710 & 1'b0 ) ;
  assign n16712 = n16704 | n16711 ;
  assign n16682 = ~n16673 & n16681 ;
  assign n16693 = ( n16682 & ~n15484 ) | ( n16682 & n16692 ) | ( ~n15484 & n16692 ) ;
  assign n16694 = ( n14905 & ~n16693 ) | ( n14905 & 1'b0 ) | ( ~n16693 & 1'b0 ) ;
  assign n16726 = n14341 | n16694 ;
  assign n16727 = ( n16712 & ~n16726 ) | ( n16712 & 1'b0 ) | ( ~n16726 & 1'b0 ) ;
  assign n16728 = n16718 | n16727 ;
  assign n16729 = ( n16707 & ~n16709 ) | ( n16707 & 1'b0 ) | ( ~n16709 & 1'b0 ) ;
  assign n16730 = ( n16704 & ~n14905 ) | ( n16704 & n16729 ) | ( ~n14905 & n16729 ) ;
  assign n16731 = ( n14341 & ~n16730 ) | ( n14341 & 1'b0 ) | ( ~n16730 & 1'b0 ) ;
  assign n16732 = n13784 | n16731 ;
  assign n16733 = ( n16728 & ~n16732 ) | ( n16728 & 1'b0 ) | ( ~n16732 & 1'b0 ) ;
  assign n16734 = n16725 | n16733 ;
  assign n16713 = ~n16694 & n16712 ;
  assign n16719 = ( n16713 & ~n14341 ) | ( n16713 & n16718 ) | ( ~n14341 & n16718 ) ;
  assign n16720 = ( n13784 & ~n16719 ) | ( n13784 & 1'b0 ) | ( ~n16719 & 1'b0 ) ;
  assign n16748 = n13242 | n16720 ;
  assign n16749 = ( n16734 & ~n16748 ) | ( n16734 & 1'b0 ) | ( ~n16748 & 1'b0 ) ;
  assign n16750 = n16740 | n16749 ;
  assign n16751 = ( n16728 & ~n16731 ) | ( n16728 & 1'b0 ) | ( ~n16731 & 1'b0 ) ;
  assign n16752 = ( n16725 & ~n13784 ) | ( n16725 & n16751 ) | ( ~n13784 & n16751 ) ;
  assign n16753 = ( n13242 & ~n16752 ) | ( n13242 & 1'b0 ) | ( ~n16752 & 1'b0 ) ;
  assign n16754 = n12707 | n16753 ;
  assign n16755 = ( n16750 & ~n16754 ) | ( n16750 & 1'b0 ) | ( ~n16754 & 1'b0 ) ;
  assign n16756 = n16747 | n16755 ;
  assign n16735 = ~n16720 & n16734 ;
  assign n16741 = ( n16735 & ~n13242 ) | ( n16735 & n16740 ) | ( ~n13242 & n16740 ) ;
  assign n16742 = ( n12707 & ~n16741 ) | ( n12707 & 1'b0 ) | ( ~n16741 & 1'b0 ) ;
  assign n16770 = n12187 | n16742 ;
  assign n16771 = ( n16756 & ~n16770 ) | ( n16756 & 1'b0 ) | ( ~n16770 & 1'b0 ) ;
  assign n16772 = n16762 | n16771 ;
  assign n16773 = ( n16750 & ~n16753 ) | ( n16750 & 1'b0 ) | ( ~n16753 & 1'b0 ) ;
  assign n16774 = ( n16747 & ~n12707 ) | ( n16747 & n16773 ) | ( ~n12707 & n16773 ) ;
  assign n16775 = ( n12187 & ~n16774 ) | ( n12187 & 1'b0 ) | ( ~n16774 & 1'b0 ) ;
  assign n16776 = n11674 | n16775 ;
  assign n16777 = ( n16772 & ~n16776 ) | ( n16772 & 1'b0 ) | ( ~n16776 & 1'b0 ) ;
  assign n16778 = n16769 | n16777 ;
  assign n16757 = ~n16742 & n16756 ;
  assign n16763 = ( n16757 & ~n12187 ) | ( n16757 & n16762 ) | ( ~n12187 & n16762 ) ;
  assign n16764 = ( n11674 & ~n16763 ) | ( n11674 & 1'b0 ) | ( ~n16763 & 1'b0 ) ;
  assign n16792 = n11176 | n16764 ;
  assign n16793 = ( n16778 & ~n16792 ) | ( n16778 & 1'b0 ) | ( ~n16792 & 1'b0 ) ;
  assign n16794 = n16784 | n16793 ;
  assign n16795 = ( n16772 & ~n16775 ) | ( n16772 & 1'b0 ) | ( ~n16775 & 1'b0 ) ;
  assign n16796 = ( n16769 & ~n11674 ) | ( n16769 & n16795 ) | ( ~n11674 & n16795 ) ;
  assign n16797 = ( n11176 & ~n16796 ) | ( n11176 & 1'b0 ) | ( ~n16796 & 1'b0 ) ;
  assign n16798 = n10685 | n16797 ;
  assign n16799 = ( n16794 & ~n16798 ) | ( n16794 & 1'b0 ) | ( ~n16798 & 1'b0 ) ;
  assign n16800 = n16791 | n16799 ;
  assign n16779 = ~n16764 & n16778 ;
  assign n16785 = ( n16779 & ~n11176 ) | ( n16779 & n16784 ) | ( ~n11176 & n16784 ) ;
  assign n16786 = ( n10685 & ~n16785 ) | ( n10685 & 1'b0 ) | ( ~n16785 & 1'b0 ) ;
  assign n16814 = n10209 | n16786 ;
  assign n16815 = ( n16800 & ~n16814 ) | ( n16800 & 1'b0 ) | ( ~n16814 & 1'b0 ) ;
  assign n16816 = n16806 | n16815 ;
  assign n16817 = ( n16794 & ~n16797 ) | ( n16794 & 1'b0 ) | ( ~n16797 & 1'b0 ) ;
  assign n16818 = ( n16791 & ~n10685 ) | ( n16791 & n16817 ) | ( ~n10685 & n16817 ) ;
  assign n16819 = ( n10209 & ~n16818 ) | ( n10209 & 1'b0 ) | ( ~n16818 & 1'b0 ) ;
  assign n16820 = ( n9740 & ~n16819 ) | ( n9740 & 1'b0 ) | ( ~n16819 & 1'b0 ) ;
  assign n16821 = n16816 &  n16820 ;
  assign n16822 = n16813 | n16821 ;
  assign n16801 = ~n16786 & n16800 ;
  assign n16807 = ( n16801 & ~n10209 ) | ( n16801 & n16806 ) | ( ~n10209 & n16806 ) ;
  assign n16808 = n9740 | n16807 ;
  assign n16836 = ~n9286 & n16808 ;
  assign n16837 = n16822 &  n16836 ;
  assign n16838 = n16828 | n16837 ;
  assign n16839 = ( n16816 & ~n16819 ) | ( n16816 & 1'b0 ) | ( ~n16819 & 1'b0 ) ;
  assign n16840 = ( n9740 & n16813 ) | ( n9740 & n16839 ) | ( n16813 & n16839 ) ;
  assign n16841 = ( n9286 & ~n16840 ) | ( n9286 & 1'b0 ) | ( ~n16840 & 1'b0 ) ;
  assign n16842 = n8839 | n16841 ;
  assign n16843 = ( n16838 & ~n16842 ) | ( n16838 & 1'b0 ) | ( ~n16842 & 1'b0 ) ;
  assign n16844 = n16835 | n16843 ;
  assign n16823 = n16808 &  n16822 ;
  assign n16829 = ( n16823 & ~n9286 ) | ( n16823 & n16828 ) | ( ~n9286 & n16828 ) ;
  assign n16830 = ( n8839 & ~n16829 ) | ( n8839 & 1'b0 ) | ( ~n16829 & 1'b0 ) ;
  assign n16858 = n8407 | n16830 ;
  assign n16859 = ( n16844 & ~n16858 ) | ( n16844 & 1'b0 ) | ( ~n16858 & 1'b0 ) ;
  assign n16860 = n16850 | n16859 ;
  assign n16861 = ( n16838 & ~n16841 ) | ( n16838 & 1'b0 ) | ( ~n16841 & 1'b0 ) ;
  assign n16862 = ( n16835 & ~n8839 ) | ( n16835 & n16861 ) | ( ~n8839 & n16861 ) ;
  assign n16863 = ( n8407 & ~n16862 ) | ( n8407 & 1'b0 ) | ( ~n16862 & 1'b0 ) ;
  assign n16864 = n7982 | n16863 ;
  assign n16865 = ( n16860 & ~n16864 ) | ( n16860 & 1'b0 ) | ( ~n16864 & 1'b0 ) ;
  assign n16866 = n16857 | n16865 ;
  assign n16845 = ~n16830 & n16844 ;
  assign n16851 = ( n16845 & ~n8407 ) | ( n16845 & n16850 ) | ( ~n8407 & n16850 ) ;
  assign n16852 = ( n7982 & ~n16851 ) | ( n7982 & 1'b0 ) | ( ~n16851 & 1'b0 ) ;
  assign n16880 = ( n7572 & ~n16852 ) | ( n7572 & 1'b0 ) | ( ~n16852 & 1'b0 ) ;
  assign n16881 = n16866 &  n16880 ;
  assign n16882 = n16872 | n16881 ;
  assign n16883 = ( n16860 & ~n16863 ) | ( n16860 & 1'b0 ) | ( ~n16863 & 1'b0 ) ;
  assign n16884 = ( n16857 & ~n7982 ) | ( n16857 & n16883 ) | ( ~n7982 & n16883 ) ;
  assign n16885 = n7572 | n16884 ;
  assign n16886 = n7169 &  n16885 ;
  assign n16887 = n16882 &  n16886 ;
  assign n16888 = n16879 | n16887 ;
  assign n16867 = ~n16852 & n16866 ;
  assign n16873 = ( n7572 & n16867 ) | ( n7572 & n16872 ) | ( n16867 & n16872 ) ;
  assign n16874 = n7169 | n16873 ;
  assign n16902 = ~n6781 & n16874 ;
  assign n16903 = n16888 &  n16902 ;
  assign n16904 = n16894 | n16903 ;
  assign n16905 = n16882 &  n16885 ;
  assign n16906 = ( n7169 & n16879 ) | ( n7169 & n16905 ) | ( n16879 & n16905 ) ;
  assign n16907 = ( n6781 & ~n16906 ) | ( n6781 & 1'b0 ) | ( ~n16906 & 1'b0 ) ;
  assign n16908 = ( n6399 & ~n16907 ) | ( n6399 & 1'b0 ) | ( ~n16907 & 1'b0 ) ;
  assign n16909 = n16904 &  n16908 ;
  assign n16910 = n16901 | n16909 ;
  assign n16889 = n16874 &  n16888 ;
  assign n16895 = ( n16889 & ~n6781 ) | ( n16889 & n16894 ) | ( ~n6781 & n16894 ) ;
  assign n16896 = n6399 | n16895 ;
  assign n16924 = ~n6032 & n16896 ;
  assign n16925 = n16910 &  n16924 ;
  assign n16926 = n16916 | n16925 ;
  assign n16927 = ( n16904 & ~n16907 ) | ( n16904 & 1'b0 ) | ( ~n16907 & 1'b0 ) ;
  assign n16928 = ( n6399 & n16901 ) | ( n6399 & n16927 ) | ( n16901 & n16927 ) ;
  assign n16929 = ( n6032 & ~n16928 ) | ( n6032 & 1'b0 ) | ( ~n16928 & 1'b0 ) ;
  assign n16930 = ( n5672 & ~n16929 ) | ( n5672 & 1'b0 ) | ( ~n16929 & 1'b0 ) ;
  assign n16931 = n16926 &  n16930 ;
  assign n16932 = n16923 | n16931 ;
  assign n16911 = n16896 &  n16910 ;
  assign n16917 = ( n16911 & ~n6032 ) | ( n16911 & n16916 ) | ( ~n6032 & n16916 ) ;
  assign n16918 = n5672 | n16917 ;
  assign n16946 = ~n5327 & n16918 ;
  assign n16947 = n16932 &  n16946 ;
  assign n16948 = n16938 | n16947 ;
  assign n16949 = ( n16926 & ~n16929 ) | ( n16926 & 1'b0 ) | ( ~n16929 & 1'b0 ) ;
  assign n16950 = ( n5672 & n16923 ) | ( n5672 & n16949 ) | ( n16923 & n16949 ) ;
  assign n16951 = ( n5327 & ~n16950 ) | ( n5327 & 1'b0 ) | ( ~n16950 & 1'b0 ) ;
  assign n16952 = n4990 | n16951 ;
  assign n16953 = ( n16948 & ~n16952 ) | ( n16948 & 1'b0 ) | ( ~n16952 & 1'b0 ) ;
  assign n16954 = n16945 | n16953 ;
  assign n16933 = n16918 &  n16932 ;
  assign n16939 = ( n16933 & ~n5327 ) | ( n16933 & n16938 ) | ( ~n5327 & n16938 ) ;
  assign n16940 = ( n4990 & ~n16939 ) | ( n4990 & 1'b0 ) | ( ~n16939 & 1'b0 ) ;
  assign n16968 = n4668 | n16940 ;
  assign n16969 = ( n16954 & ~n16968 ) | ( n16954 & 1'b0 ) | ( ~n16968 & 1'b0 ) ;
  assign n16970 = n16960 | n16969 ;
  assign n16971 = ( n16948 & ~n16951 ) | ( n16948 & 1'b0 ) | ( ~n16951 & 1'b0 ) ;
  assign n16972 = ( n16945 & ~n4990 ) | ( n16945 & n16971 ) | ( ~n4990 & n16971 ) ;
  assign n16973 = ( n4668 & ~n16972 ) | ( n4668 & 1'b0 ) | ( ~n16972 & 1'b0 ) ;
  assign n16974 = n4353 | n16973 ;
  assign n16975 = ( n16970 & ~n16974 ) | ( n16970 & 1'b0 ) | ( ~n16974 & 1'b0 ) ;
  assign n16976 = ( n16967 & ~n16975 ) | ( n16967 & 1'b0 ) | ( ~n16975 & 1'b0 ) ;
  assign n16955 = ~n16940 & n16954 ;
  assign n16961 = ( n16955 & ~n4668 ) | ( n16955 & n16960 ) | ( ~n4668 & n16960 ) ;
  assign n16962 = ( n4353 & ~n16961 ) | ( n4353 & 1'b0 ) | ( ~n16961 & 1'b0 ) ;
  assign n16990 = n4053 | n16962 ;
  assign n16991 = n16976 | n16990 ;
  assign n16992 = n16982 &  n16991 ;
  assign n16993 = ( n16970 & ~n16973 ) | ( n16970 & 1'b0 ) | ( ~n16973 & 1'b0 ) ;
  assign n16994 = ( n4353 & ~n16993 ) | ( n4353 & n16967 ) | ( ~n16993 & n16967 ) ;
  assign n16995 = n4053 &  n16994 ;
  assign n16996 = n3760 | n16995 ;
  assign n16997 = n16992 | n16996 ;
  assign n16998 = n16989 &  n16997 ;
  assign n16977 = n16962 | n16976 ;
  assign n16983 = ( n4053 & n16977 ) | ( n4053 & n16982 ) | ( n16977 & n16982 ) ;
  assign n16984 = n3760 &  n16983 ;
  assign n17012 = n3482 | n16984 ;
  assign n17013 = n16998 | n17012 ;
  assign n17014 = n17004 &  n17013 ;
  assign n17015 = n16992 | n16995 ;
  assign n17016 = ( n3760 & n16989 ) | ( n3760 & n17015 ) | ( n16989 & n17015 ) ;
  assign n17017 = n3482 &  n17016 ;
  assign n17018 = n3211 | n17017 ;
  assign n17019 = n17014 | n17018 ;
  assign n17020 = n17011 &  n17019 ;
  assign n16999 = n16984 | n16998 ;
  assign n17005 = ( n3482 & n16999 ) | ( n3482 & n17004 ) | ( n16999 & n17004 ) ;
  assign n17006 = n3211 &  n17005 ;
  assign n17034 = n2955 | n17006 ;
  assign n17035 = n17020 | n17034 ;
  assign n17036 = ~n17026 & n17035 ;
  assign n17037 = n17014 | n17017 ;
  assign n17038 = ( n3211 & n17011 ) | ( n3211 & n17037 ) | ( n17011 & n17037 ) ;
  assign n17039 = n2955 &  n17038 ;
  assign n17040 = n2706 | n17039 ;
  assign n17041 = n17036 | n17040 ;
  assign n17042 = ~n17033 & n17041 ;
  assign n17021 = n17006 | n17020 ;
  assign n17027 = ( n2955 & ~n17026 ) | ( n2955 & n17021 ) | ( ~n17026 & n17021 ) ;
  assign n17028 = n2706 &  n17027 ;
  assign n17056 = n2472 | n17028 ;
  assign n17057 = n17042 | n17056 ;
  assign n17058 = n17048 &  n17057 ;
  assign n17059 = n17036 | n17039 ;
  assign n17060 = ( n2706 & ~n17033 ) | ( n2706 & n17059 ) | ( ~n17033 & n17059 ) ;
  assign n17061 = n2472 &  n17060 ;
  assign n17062 = n2245 | n17061 ;
  assign n17063 = n17058 | n17062 ;
  assign n17064 = ~n17055 & n17063 ;
  assign n17043 = n17028 | n17042 ;
  assign n17049 = ( n2472 & n17043 ) | ( n2472 & n17048 ) | ( n17043 & n17048 ) ;
  assign n17050 = n2245 &  n17049 ;
  assign n17078 = ( n2033 & ~n17050 ) | ( n2033 & 1'b0 ) | ( ~n17050 & 1'b0 ) ;
  assign n17079 = ~n17064 & n17078 ;
  assign n17080 = ( n17070 & ~n17079 ) | ( n17070 & 1'b0 ) | ( ~n17079 & 1'b0 ) ;
  assign n17081 = n17058 | n17061 ;
  assign n17082 = ( n2245 & ~n17055 ) | ( n2245 & n17081 ) | ( ~n17055 & n17081 ) ;
  assign n17083 = ~n2033 & n17082 ;
  assign n17084 = n1827 | n17083 ;
  assign n17085 = n17080 | n17084 ;
  assign n17086 = n17077 &  n17085 ;
  assign n17065 = n17050 | n17064 ;
  assign n17071 = ( n17065 & ~n2033 ) | ( n17065 & n17070 ) | ( ~n2033 & n17070 ) ;
  assign n17072 = n1827 &  n17071 ;
  assign n17100 = ( n1636 & ~n17072 ) | ( n1636 & 1'b0 ) | ( ~n17072 & 1'b0 ) ;
  assign n17101 = ~n17086 & n17100 ;
  assign n17102 = n17092 | n17101 ;
  assign n17103 = n17080 | n17083 ;
  assign n17104 = ( n1827 & n17077 ) | ( n1827 & n17103 ) | ( n17077 & n17103 ) ;
  assign n17105 = ~n1636 & n17104 ;
  assign n17106 = ( n1452 & ~n17105 ) | ( n1452 & 1'b0 ) | ( ~n17105 & 1'b0 ) ;
  assign n17107 = n17102 &  n17106 ;
  assign n17108 = n17099 | n17107 ;
  assign n17087 = n17072 | n17086 ;
  assign n17093 = ( n1636 & ~n17087 ) | ( n1636 & n17092 ) | ( ~n17087 & n17092 ) ;
  assign n17094 = n1452 | n17093 ;
  assign n17122 = ~n1283 & n17094 ;
  assign n17123 = n17108 &  n17122 ;
  assign n17124 = n17114 | n17123 ;
  assign n17125 = ( n17102 & ~n17105 ) | ( n17102 & 1'b0 ) | ( ~n17105 & 1'b0 ) ;
  assign n17126 = ( n1452 & n17099 ) | ( n1452 & n17125 ) | ( n17099 & n17125 ) ;
  assign n17127 = ( n1283 & ~n17126 ) | ( n1283 & 1'b0 ) | ( ~n17126 & 1'b0 ) ;
  assign n17128 = ( n1122 & ~n17127 ) | ( n1122 & 1'b0 ) | ( ~n17127 & 1'b0 ) ;
  assign n17129 = n17124 &  n17128 ;
  assign n17130 = n17121 | n17129 ;
  assign n17109 = n17094 &  n17108 ;
  assign n17115 = ( n17109 & ~n1283 ) | ( n17109 & n17114 ) | ( ~n1283 & n17114 ) ;
  assign n17116 = n1122 | n17115 ;
  assign n17144 = n976 &  n17116 ;
  assign n17145 = n17130 &  n17144 ;
  assign n17146 = n17136 | n17145 ;
  assign n17147 = ( n17124 & ~n17127 ) | ( n17124 & 1'b0 ) | ( ~n17127 & 1'b0 ) ;
  assign n17148 = ( n1122 & n17121 ) | ( n1122 & n17147 ) | ( n17121 & n17147 ) ;
  assign n17149 = n976 | n17148 ;
  assign n17164 = n17146 &  n17149 ;
  assign n17139 = ( n16541 & ~n16671 ) | ( n16541 & 1'b0 ) | ( ~n16671 & 1'b0 ) ;
  assign n17140 = ( n16528 & n16537 ) | ( n16528 & n16541 ) | ( n16537 & n16541 ) ;
  assign n17141 = ( n17139 & ~n16537 ) | ( n17139 & n17140 ) | ( ~n16537 & n17140 ) ;
  assign n17142 = ( n16541 & ~n17140 ) | ( n16541 & n17139 ) | ( ~n17140 & n17139 ) ;
  assign n17143 = ( n16528 & ~n17141 ) | ( n16528 & n17142 ) | ( ~n17141 & n17142 ) ;
  assign n17165 = ( n837 & ~n17164 ) | ( n837 & n17143 ) | ( ~n17164 & n17143 ) ;
  assign n17166 = n713 &  n17165 ;
  assign n17247 = ( n16637 & ~n16656 ) | ( n16637 & 1'b0 ) | ( ~n16656 & 1'b0 ) ;
  assign n17248 = ( n16653 & n16671 ) | ( n16653 & n17247 ) | ( n16671 & n17247 ) ;
  assign n17249 = ~n16653 & n17248 ;
  assign n17250 = n16653 | n16656 ;
  assign n17251 = n16671 | n17250 ;
  assign n17252 = ( n16637 & ~n17250 ) | ( n16637 & n17251 ) | ( ~n17250 & n17251 ) ;
  assign n17253 = ~n17249 & n17252 ;
  assign n17254 = ~n16638 & n16645 ;
  assign n17255 = ~n16671 & n17254 ;
  assign n17256 = ( n16659 & ~n17255 ) | ( n16659 & n17254 ) | ( ~n17255 & n17254 ) ;
  assign n17257 = n17253 | n17256 ;
  assign n17241 = n16617 | n16671 ;
  assign n17242 = ( n16617 & ~n16630 ) | ( n16617 & n16622 ) | ( ~n16630 & n16622 ) ;
  assign n17243 = ( n16630 & n17241 ) | ( n16630 & n17242 ) | ( n17241 & n17242 ) ;
  assign n17244 = ( n16617 & ~n17242 ) | ( n16617 & n17241 ) | ( ~n17242 & n17241 ) ;
  assign n17245 = ( n16622 & ~n17243 ) | ( n16622 & n17244 ) | ( ~n17243 & n17244 ) ;
  assign n17219 = ~n16608 & n16671 ;
  assign n17220 = ( n16595 & ~n17219 ) | ( n16595 & n16671 ) | ( ~n17219 & n16671 ) ;
  assign n17221 = ( n16600 & ~n16595 ) | ( n16600 & n17220 ) | ( ~n16595 & n17220 ) ;
  assign n17222 = ( n16595 & ~n17220 ) | ( n16595 & n16600 ) | ( ~n17220 & n16600 ) ;
  assign n17223 = ( n17221 & ~n16600 ) | ( n17221 & n17222 ) | ( ~n16600 & n17222 ) ;
  assign n17131 = n17116 &  n17130 ;
  assign n17137 = ( n976 & n17131 ) | ( n976 & n17136 ) | ( n17131 & n17136 ) ;
  assign n17138 = ( n837 & ~n17137 ) | ( n837 & 1'b0 ) | ( ~n17137 & 1'b0 ) ;
  assign n17150 = ~n837 & n17149 ;
  assign n17151 = n17146 &  n17150 ;
  assign n17152 = ( n17143 & ~n17151 ) | ( n17143 & 1'b0 ) | ( ~n17151 & 1'b0 ) ;
  assign n17153 = n17138 | n17152 ;
  assign n17159 = ( n713 & ~n17158 ) | ( n713 & n17153 ) | ( ~n17158 & n17153 ) ;
  assign n17160 = n595 &  n17159 ;
  assign n17161 = n713 | n17138 ;
  assign n17162 = n17152 | n17161 ;
  assign n17163 = ~n17158 & n17162 ;
  assign n17167 = n595 | n17166 ;
  assign n17168 = n17163 | n17167 ;
  assign n17169 = ( n16549 & ~n16558 ) | ( n16549 & n16562 ) | ( ~n16558 & n16562 ) ;
  assign n17170 = ( n16558 & n16671 ) | ( n16558 & n17169 ) | ( n16671 & n17169 ) ;
  assign n17171 = ( n16562 & ~n17169 ) | ( n16562 & n16671 ) | ( ~n17169 & n16671 ) ;
  assign n17172 = ( n16549 & ~n17170 ) | ( n16549 & n17171 ) | ( ~n17170 & n17171 ) ;
  assign n17173 = ( n17168 & ~n17172 ) | ( n17168 & 1'b0 ) | ( ~n17172 & 1'b0 ) ;
  assign n17174 = n17160 | n17173 ;
  assign n17175 = n16564 &  n16671 ;
  assign n17176 = ( n16551 & ~n17175 ) | ( n16551 & n16671 ) | ( ~n17175 & n16671 ) ;
  assign n17177 = ( n16551 & ~n17176 ) | ( n16551 & n16556 ) | ( ~n17176 & n16556 ) ;
  assign n17178 = ( n16556 & ~n16551 ) | ( n16556 & n17176 ) | ( ~n16551 & n17176 ) ;
  assign n17179 = ( n17177 & ~n16556 ) | ( n17177 & n17178 ) | ( ~n16556 & n17178 ) ;
  assign n17180 = ( n492 & n17174 ) | ( n492 & n17179 ) | ( n17174 & n17179 ) ;
  assign n17181 = n396 &  n17180 ;
  assign n17183 = ( n16580 & ~n16571 ) | ( n16580 & n16584 ) | ( ~n16571 & n16584 ) ;
  assign n17182 = n16584 | n16671 ;
  assign n17185 = ( n16584 & ~n17183 ) | ( n16584 & n17182 ) | ( ~n17183 & n17182 ) ;
  assign n17184 = ( n17182 & ~n16580 ) | ( n17182 & n17183 ) | ( ~n16580 & n17183 ) ;
  assign n17186 = ( n16571 & ~n17185 ) | ( n16571 & n17184 ) | ( ~n17185 & n17184 ) ;
  assign n17187 = n492 | n17160 ;
  assign n17188 = n17173 | n17187 ;
  assign n17189 = n17179 &  n17188 ;
  assign n17190 = n17163 | n17166 ;
  assign n17191 = ( n595 & ~n17172 ) | ( n595 & n17190 ) | ( ~n17172 & n17190 ) ;
  assign n17192 = n492 &  n17191 ;
  assign n17193 = n396 | n17192 ;
  assign n17194 = n17189 | n17193 ;
  assign n17195 = ~n17186 & n17194 ;
  assign n17196 = n17181 | n17195 ;
  assign n17197 = ~n16586 & n16671 ;
  assign n17198 = ( n16573 & ~n17197 ) | ( n16573 & n16671 ) | ( ~n17197 & n16671 ) ;
  assign n17199 = ( n16573 & ~n17198 ) | ( n16573 & n16578 ) | ( ~n17198 & n16578 ) ;
  assign n17200 = ( n16578 & ~n16573 ) | ( n16578 & n17198 ) | ( ~n16573 & n17198 ) ;
  assign n17201 = ( n17199 & ~n16578 ) | ( n17199 & n17200 ) | ( ~n16578 & n17200 ) ;
  assign n17202 = ( n315 & n17196 ) | ( n315 & n17201 ) | ( n17196 & n17201 ) ;
  assign n17203 = n240 &  n17202 ;
  assign n17204 = n16606 | n16671 ;
  assign n17205 = ( n16593 & n16602 ) | ( n16593 & n16606 ) | ( n16602 & n16606 ) ;
  assign n17206 = ( n17204 & ~n16602 ) | ( n17204 & n17205 ) | ( ~n16602 & n17205 ) ;
  assign n17207 = ( n16606 & ~n17205 ) | ( n16606 & n17204 ) | ( ~n17205 & n17204 ) ;
  assign n17208 = ( n16593 & ~n17206 ) | ( n16593 & n17207 ) | ( ~n17206 & n17207 ) ;
  assign n17209 = n315 | n17181 ;
  assign n17210 = n17195 | n17209 ;
  assign n17211 = n17201 &  n17210 ;
  assign n17212 = n17189 | n17192 ;
  assign n17213 = ( n396 & ~n17186 ) | ( n396 & n17212 ) | ( ~n17186 & n17212 ) ;
  assign n17214 = n315 &  n17213 ;
  assign n17215 = n240 | n17214 ;
  assign n17216 = n17211 | n17215 ;
  assign n17217 = n17208 &  n17216 ;
  assign n17218 = n17203 | n17217 ;
  assign n17224 = ( n181 & ~n17223 ) | ( n181 & n17218 ) | ( ~n17223 & n17218 ) ;
  assign n17225 = ~n145 & n17224 ;
  assign n17227 = ( n16624 & ~n16615 ) | ( n16624 & n16628 ) | ( ~n16615 & n16628 ) ;
  assign n17226 = n16628 | n16671 ;
  assign n17229 = ( n16628 & ~n17227 ) | ( n16628 & n17226 ) | ( ~n17227 & n17226 ) ;
  assign n17228 = ( n17226 & ~n16624 ) | ( n17226 & n17227 ) | ( ~n16624 & n17227 ) ;
  assign n17230 = ( n16615 & ~n17229 ) | ( n16615 & n17228 ) | ( ~n17229 & n17228 ) ;
  assign n17231 = n181 | n17203 ;
  assign n17232 = n17217 | n17231 ;
  assign n17233 = ~n17223 & n17232 ;
  assign n17234 = n17211 | n17214 ;
  assign n17235 = ( n240 & n17208 ) | ( n240 & n17234 ) | ( n17208 & n17234 ) ;
  assign n17236 = n181 &  n17235 ;
  assign n17237 = ( n145 & ~n17236 ) | ( n145 & 1'b0 ) | ( ~n17236 & 1'b0 ) ;
  assign n17238 = ~n17233 & n17237 ;
  assign n17239 = ( n17230 & ~n17238 ) | ( n17230 & 1'b0 ) | ( ~n17238 & 1'b0 ) ;
  assign n17240 = n17225 | n17239 ;
  assign n17246 = ( n150 & ~n17245 ) | ( n150 & n17240 ) | ( ~n17245 & n17240 ) ;
  assign n17258 = n17246 | n17257 ;
  assign n17259 = ( n133 & ~n17257 ) | ( n133 & n17258 ) | ( ~n17257 & n17258 ) ;
  assign n17260 = n150 | n17225 ;
  assign n17261 = n17239 | n17260 ;
  assign n17266 = n17245 | n17261 ;
  assign n17262 = n17233 | n17236 ;
  assign n17263 = ( n17230 & ~n145 ) | ( n17230 & n17262 ) | ( ~n145 & n17262 ) ;
  assign n17264 = n150 &  n17263 ;
  assign n17265 = ( n17253 & ~n17264 ) | ( n17253 & 1'b0 ) | ( ~n17264 & 1'b0 ) ;
  assign n17267 = ( n17245 & ~n17266 ) | ( n17245 & n17265 ) | ( ~n17266 & n17265 ) ;
  assign n17269 = ( n133 & ~n16638 ) | ( n133 & n16645 ) | ( ~n16638 & n16645 ) ;
  assign n17268 = ( n16638 & ~n16645 ) | ( n16638 & n16671 ) | ( ~n16645 & n16671 ) ;
  assign n17270 = n16645 &  n17268 ;
  assign n17271 = ( n17269 & ~n16645 ) | ( n17269 & n17270 ) | ( ~n16645 & n17270 ) ;
  assign n17272 = n16641 | n16668 ;
  assign n17273 = ( n16663 & ~n16644 ) | ( n16663 & n17272 ) | ( ~n16644 & n17272 ) ;
  assign n17274 = n16644 | n17273 ;
  assign n17275 = ( n16651 & n16659 ) | ( n16651 & n17274 ) | ( n16659 & n17274 ) ;
  assign n17276 = ( n16651 & ~n17275 ) | ( n16651 & 1'b0 ) | ( ~n17275 & 1'b0 ) ;
  assign n17277 = n17271 | n17276 ;
  assign n17278 = n17267 | n17277 ;
  assign n17279 = ~n17259 |  n17278 ;
  assign n17784 = n17166 | n17279 ;
  assign n17785 = ( n17158 & n17162 ) | ( n17158 & n17166 ) | ( n17162 & n17166 ) ;
  assign n17786 = ( n17784 & ~n17162 ) | ( n17784 & n17785 ) | ( ~n17162 & n17785 ) ;
  assign n17787 = ( n17166 & ~n17785 ) | ( n17166 & n17784 ) | ( ~n17785 & n17784 ) ;
  assign n17788 = ( n17158 & ~n17786 ) | ( n17158 & n17787 ) | ( ~n17786 & n17787 ) ;
  assign n17668 = ( n17028 & ~n17033 ) | ( n17028 & n17041 ) | ( ~n17033 & n17041 ) ;
  assign n17667 = n17028 | n17279 ;
  assign n17670 = ( n17028 & ~n17668 ) | ( n17028 & n17667 ) | ( ~n17668 & n17667 ) ;
  assign n17669 = ( n17667 & ~n17041 ) | ( n17667 & n17668 ) | ( ~n17041 & n17668 ) ;
  assign n17671 = ( n17033 & ~n17670 ) | ( n17033 & n17669 ) | ( ~n17670 & n17669 ) ;
  assign n17286 = ( x18 & ~n17279 ) | ( x18 & x19 ) | ( ~n17279 & x19 ) ;
  assign n17292 = ( x18 & ~x19 ) | ( x18 & 1'b0 ) | ( ~x19 & 1'b0 ) ;
  assign n17282 = x16 | x17 ;
  assign n17287 = ~x18 & n17282 ;
  assign n17288 = ( x18 & ~n16669 ) | ( x18 & n17287 ) | ( ~n16669 & n17287 ) ;
  assign n17289 = ( n16651 & ~n17288 ) | ( n16651 & n16659 ) | ( ~n17288 & n16659 ) ;
  assign n17290 = ( n16651 & ~n17289 ) | ( n16651 & 1'b0 ) | ( ~n17289 & 1'b0 ) ;
  assign n17291 = ( n17279 & ~x19 ) | ( n17279 & n17290 ) | ( ~x19 & n17290 ) ;
  assign n17293 = ( n17286 & ~n17292 ) | ( n17286 & n17291 ) | ( ~n17292 & n17291 ) ;
  assign n17283 = x18 | n17282 ;
  assign n17284 = x18 &  n17279 ;
  assign n17285 = ( n16671 & ~n17283 ) | ( n16671 & n17284 ) | ( ~n17283 & n17284 ) ;
  assign n17294 = n17285 &  n17293 ;
  assign n17295 = ( n16070 & ~n17293 ) | ( n16070 & n17294 ) | ( ~n17293 & n17294 ) ;
  assign n17296 = n16070 | n17285 ;
  assign n17297 = ( n17293 & ~n17296 ) | ( n17293 & 1'b0 ) | ( ~n17296 & 1'b0 ) ;
  assign n17299 = ( n16671 & ~n17276 ) | ( n16671 & 1'b0 ) | ( ~n17276 & 1'b0 ) ;
  assign n17300 = ( n17267 & ~n17271 ) | ( n17267 & n17299 ) | ( ~n17271 & n17299 ) ;
  assign n17301 = ~n17267 & n17300 ;
  assign n17302 = n17259 &  n17301 ;
  assign n17298 = ~n16071 & n17279 ;
  assign n17303 = ( n17298 & ~n17302 ) | ( n17298 & 1'b0 ) | ( ~n17302 & 1'b0 ) ;
  assign n17304 = ( x20 & n17302 ) | ( x20 & n17303 ) | ( n17302 & n17303 ) ;
  assign n17305 = x20 | n17302 ;
  assign n17306 = n17298 | n17305 ;
  assign n17307 = ~n17304 & n17306 ;
  assign n17308 = n17297 | n17307 ;
  assign n17309 = ~n17295 & n17308 ;
  assign n17313 = ~x20 & n16671 ;
  assign n17314 = ( x21 & ~n17313 ) | ( x21 & 1'b0 ) | ( ~n17313 & 1'b0 ) ;
  assign n17315 = n16683 | n17314 ;
  assign n17310 = ( n16671 & ~x20 ) | ( n16671 & n16678 ) | ( ~x20 & n16678 ) ;
  assign n17311 = x20 &  n17310 ;
  assign n17312 = ( n16673 & ~n17311 ) | ( n16673 & n16678 ) | ( ~n17311 & n16678 ) ;
  assign n17316 = ( n17279 & ~n17315 ) | ( n17279 & n17312 ) | ( ~n17315 & n17312 ) ;
  assign n17318 = ( n17279 & ~n17316 ) | ( n17279 & 1'b0 ) | ( ~n17316 & 1'b0 ) ;
  assign n17317 = ~n17312 & n17316 ;
  assign n17319 = ( n17315 & ~n17318 ) | ( n17315 & n17317 ) | ( ~n17318 & n17317 ) ;
  assign n17320 = ( n17309 & ~n15484 ) | ( n17309 & n17319 ) | ( ~n15484 & n17319 ) ;
  assign n17321 = ( n14905 & ~n17320 ) | ( n14905 & 1'b0 ) | ( ~n17320 & 1'b0 ) ;
  assign n17322 = ~n16706 & n16709 ;
  assign n17323 = ( n16692 & ~n17322 ) | ( n16692 & n16706 ) | ( ~n17322 & n16706 ) ;
  assign n17324 = ( n17279 & n17322 ) | ( n17279 & n17323 ) | ( n17322 & n17323 ) ;
  assign n17325 = ( n16706 & ~n17323 ) | ( n16706 & n17279 ) | ( ~n17323 & n17279 ) ;
  assign n17326 = ( n16692 & ~n17324 ) | ( n16692 & n17325 ) | ( ~n17324 & n17325 ) ;
  assign n17327 = n15484 | n17295 ;
  assign n17328 = ( n17308 & ~n17327 ) | ( n17308 & 1'b0 ) | ( ~n17327 & 1'b0 ) ;
  assign n17329 = n17319 | n17328 ;
  assign n17330 = ~n17285 & n17293 ;
  assign n17331 = ( n17307 & ~n16070 ) | ( n17307 & n17330 ) | ( ~n16070 & n17330 ) ;
  assign n17332 = ( n15484 & ~n17331 ) | ( n15484 & 1'b0 ) | ( ~n17331 & 1'b0 ) ;
  assign n17333 = n14905 | n17332 ;
  assign n17334 = ( n17329 & ~n17333 ) | ( n17329 & 1'b0 ) | ( ~n17333 & 1'b0 ) ;
  assign n17335 = n17326 | n17334 ;
  assign n17336 = ~n17321 & n17335 ;
  assign n17337 = n16694 | n17279 ;
  assign n17338 = ( n16694 & ~n16711 ) | ( n16694 & n16704 ) | ( ~n16711 & n16704 ) ;
  assign n17339 = ( n16711 & n17337 ) | ( n16711 & n17338 ) | ( n17337 & n17338 ) ;
  assign n17340 = ( n16694 & ~n17338 ) | ( n16694 & n17337 ) | ( ~n17338 & n17337 ) ;
  assign n17341 = ( n16704 & ~n17339 ) | ( n16704 & n17340 ) | ( ~n17339 & n17340 ) ;
  assign n17342 = ( n17336 & ~n14341 ) | ( n17336 & n17341 ) | ( ~n14341 & n17341 ) ;
  assign n17343 = ( n13784 & ~n17342 ) | ( n13784 & 1'b0 ) | ( ~n17342 & 1'b0 ) ;
  assign n17344 = n16731 | n17279 ;
  assign n17345 = ( n16718 & ~n16731 ) | ( n16718 & n16727 ) | ( ~n16731 & n16727 ) ;
  assign n17347 = ( n16731 & n17344 ) | ( n16731 & n17345 ) | ( n17344 & n17345 ) ;
  assign n17346 = ( n16727 & ~n17345 ) | ( n16727 & n17344 ) | ( ~n17345 & n17344 ) ;
  assign n17348 = ( n16718 & ~n17347 ) | ( n16718 & n17346 ) | ( ~n17347 & n17346 ) ;
  assign n17349 = n14341 | n17321 ;
  assign n17350 = ( n17335 & ~n17349 ) | ( n17335 & 1'b0 ) | ( ~n17349 & 1'b0 ) ;
  assign n17351 = n17341 | n17350 ;
  assign n17352 = ( n17329 & ~n17332 ) | ( n17329 & 1'b0 ) | ( ~n17332 & 1'b0 ) ;
  assign n17353 = ( n17326 & ~n14905 ) | ( n17326 & n17352 ) | ( ~n14905 & n17352 ) ;
  assign n17354 = ( n14341 & ~n17353 ) | ( n14341 & 1'b0 ) | ( ~n17353 & 1'b0 ) ;
  assign n17355 = n13784 | n17354 ;
  assign n17356 = ( n17351 & ~n17355 ) | ( n17351 & 1'b0 ) | ( ~n17355 & 1'b0 ) ;
  assign n17357 = n17348 | n17356 ;
  assign n17358 = ~n17343 & n17357 ;
  assign n17360 = ( n16720 & ~n16725 ) | ( n16720 & n17279 ) | ( ~n16725 & n17279 ) ;
  assign n17359 = n16733 &  n17279 ;
  assign n17361 = ( n17279 & ~n17360 ) | ( n17279 & n17359 ) | ( ~n17360 & n17359 ) ;
  assign n17362 = ( n17359 & ~n16720 ) | ( n17359 & n17360 ) | ( ~n16720 & n17360 ) ;
  assign n17363 = ( n16725 & ~n17361 ) | ( n16725 & n17362 ) | ( ~n17361 & n17362 ) ;
  assign n17364 = ( n17358 & ~n13242 ) | ( n17358 & n17363 ) | ( ~n13242 & n17363 ) ;
  assign n17365 = ( n12707 & ~n17364 ) | ( n12707 & 1'b0 ) | ( ~n17364 & 1'b0 ) ;
  assign n17366 = n16753 | n17279 ;
  assign n17367 = ( n16740 & ~n16749 ) | ( n16740 & n16753 ) | ( ~n16749 & n16753 ) ;
  assign n17368 = ( n16749 & n17366 ) | ( n16749 & n17367 ) | ( n17366 & n17367 ) ;
  assign n17369 = ( n16753 & ~n17367 ) | ( n16753 & n17366 ) | ( ~n17367 & n17366 ) ;
  assign n17370 = ( n16740 & ~n17368 ) | ( n16740 & n17369 ) | ( ~n17368 & n17369 ) ;
  assign n17371 = n13242 | n17343 ;
  assign n17372 = ( n17357 & ~n17371 ) | ( n17357 & 1'b0 ) | ( ~n17371 & 1'b0 ) ;
  assign n17373 = n17363 | n17372 ;
  assign n17374 = ( n17351 & ~n17354 ) | ( n17351 & 1'b0 ) | ( ~n17354 & 1'b0 ) ;
  assign n17375 = ( n17348 & ~n13784 ) | ( n17348 & n17374 ) | ( ~n13784 & n17374 ) ;
  assign n17376 = ( n13242 & ~n17375 ) | ( n13242 & 1'b0 ) | ( ~n17375 & 1'b0 ) ;
  assign n17377 = n12707 | n17376 ;
  assign n17378 = ( n17373 & ~n17377 ) | ( n17373 & 1'b0 ) | ( ~n17377 & 1'b0 ) ;
  assign n17379 = n17370 | n17378 ;
  assign n17380 = ~n17365 & n17379 ;
  assign n17381 = n16742 | n17279 ;
  assign n17382 = ( n16747 & ~n16742 ) | ( n16747 & n16755 ) | ( ~n16742 & n16755 ) ;
  assign n17384 = ( n16742 & n17381 ) | ( n16742 & n17382 ) | ( n17381 & n17382 ) ;
  assign n17383 = ( n16755 & ~n17382 ) | ( n16755 & n17381 ) | ( ~n17382 & n17381 ) ;
  assign n17385 = ( n16747 & ~n17384 ) | ( n16747 & n17383 ) | ( ~n17384 & n17383 ) ;
  assign n17386 = ( n17380 & ~n12187 ) | ( n17380 & n17385 ) | ( ~n12187 & n17385 ) ;
  assign n17387 = ( n11674 & ~n17386 ) | ( n11674 & 1'b0 ) | ( ~n17386 & 1'b0 ) ;
  assign n17388 = n16775 | n17279 ;
  assign n17389 = ( n16762 & ~n16771 ) | ( n16762 & n16775 ) | ( ~n16771 & n16775 ) ;
  assign n17390 = ( n16771 & n17388 ) | ( n16771 & n17389 ) | ( n17388 & n17389 ) ;
  assign n17391 = ( n16775 & ~n17389 ) | ( n16775 & n17388 ) | ( ~n17389 & n17388 ) ;
  assign n17392 = ( n16762 & ~n17390 ) | ( n16762 & n17391 ) | ( ~n17390 & n17391 ) ;
  assign n17393 = n12187 | n17365 ;
  assign n17394 = ( n17379 & ~n17393 ) | ( n17379 & 1'b0 ) | ( ~n17393 & 1'b0 ) ;
  assign n17395 = n17385 | n17394 ;
  assign n17396 = ( n17373 & ~n17376 ) | ( n17373 & 1'b0 ) | ( ~n17376 & 1'b0 ) ;
  assign n17397 = ( n17370 & ~n12707 ) | ( n17370 & n17396 ) | ( ~n12707 & n17396 ) ;
  assign n17398 = ( n12187 & ~n17397 ) | ( n12187 & 1'b0 ) | ( ~n17397 & 1'b0 ) ;
  assign n17399 = n11674 | n17398 ;
  assign n17400 = ( n17395 & ~n17399 ) | ( n17395 & 1'b0 ) | ( ~n17399 & 1'b0 ) ;
  assign n17401 = n17392 | n17400 ;
  assign n17402 = ~n17387 & n17401 ;
  assign n17403 = n16764 | n17279 ;
  assign n17404 = ( n16764 & ~n16777 ) | ( n16764 & n16769 ) | ( ~n16777 & n16769 ) ;
  assign n17405 = ( n16777 & n17403 ) | ( n16777 & n17404 ) | ( n17403 & n17404 ) ;
  assign n17406 = ( n16764 & ~n17404 ) | ( n16764 & n17403 ) | ( ~n17404 & n17403 ) ;
  assign n17407 = ( n16769 & ~n17405 ) | ( n16769 & n17406 ) | ( ~n17405 & n17406 ) ;
  assign n17408 = ( n17402 & ~n11176 ) | ( n17402 & n17407 ) | ( ~n11176 & n17407 ) ;
  assign n17409 = ( n10685 & ~n17408 ) | ( n10685 & 1'b0 ) | ( ~n17408 & 1'b0 ) ;
  assign n17410 = n16797 | n17279 ;
  assign n17411 = ( n16784 & ~n16797 ) | ( n16784 & n16793 ) | ( ~n16797 & n16793 ) ;
  assign n17413 = ( n16797 & n17410 ) | ( n16797 & n17411 ) | ( n17410 & n17411 ) ;
  assign n17412 = ( n16793 & ~n17411 ) | ( n16793 & n17410 ) | ( ~n17411 & n17410 ) ;
  assign n17414 = ( n16784 & ~n17413 ) | ( n16784 & n17412 ) | ( ~n17413 & n17412 ) ;
  assign n17415 = n11176 | n17387 ;
  assign n17416 = ( n17401 & ~n17415 ) | ( n17401 & 1'b0 ) | ( ~n17415 & 1'b0 ) ;
  assign n17417 = n17407 | n17416 ;
  assign n17418 = ( n17395 & ~n17398 ) | ( n17395 & 1'b0 ) | ( ~n17398 & 1'b0 ) ;
  assign n17419 = ( n17392 & ~n11674 ) | ( n17392 & n17418 ) | ( ~n11674 & n17418 ) ;
  assign n17420 = ( n11176 & ~n17419 ) | ( n11176 & 1'b0 ) | ( ~n17419 & 1'b0 ) ;
  assign n17421 = n10685 | n17420 ;
  assign n17422 = ( n17417 & ~n17421 ) | ( n17417 & 1'b0 ) | ( ~n17421 & 1'b0 ) ;
  assign n17423 = n17414 | n17422 ;
  assign n17424 = ~n17409 & n17423 ;
  assign n17426 = ( n16786 & ~n16791 ) | ( n16786 & n17279 ) | ( ~n16791 & n17279 ) ;
  assign n17425 = n16799 &  n17279 ;
  assign n17427 = ( n17279 & ~n17426 ) | ( n17279 & n17425 ) | ( ~n17426 & n17425 ) ;
  assign n17428 = ( n17425 & ~n16786 ) | ( n17425 & n17426 ) | ( ~n16786 & n17426 ) ;
  assign n17429 = ( n16791 & ~n17427 ) | ( n16791 & n17428 ) | ( ~n17427 & n17428 ) ;
  assign n17430 = ( n17424 & ~n10209 ) | ( n17424 & n17429 ) | ( ~n10209 & n17429 ) ;
  assign n17431 = n9740 | n17430 ;
  assign n17432 = n16819 | n17279 ;
  assign n17433 = ( n16806 & ~n16815 ) | ( n16806 & n16819 ) | ( ~n16815 & n16819 ) ;
  assign n17434 = ( n16815 & n17432 ) | ( n16815 & n17433 ) | ( n17432 & n17433 ) ;
  assign n17435 = ( n16819 & ~n17433 ) | ( n16819 & n17432 ) | ( ~n17433 & n17432 ) ;
  assign n17436 = ( n16806 & ~n17434 ) | ( n16806 & n17435 ) | ( ~n17434 & n17435 ) ;
  assign n17437 = n10209 | n17409 ;
  assign n17438 = ( n17423 & ~n17437 ) | ( n17423 & 1'b0 ) | ( ~n17437 & 1'b0 ) ;
  assign n17439 = n17429 | n17438 ;
  assign n17440 = ( n17417 & ~n17420 ) | ( n17417 & 1'b0 ) | ( ~n17420 & 1'b0 ) ;
  assign n17441 = ( n17414 & ~n10685 ) | ( n17414 & n17440 ) | ( ~n10685 & n17440 ) ;
  assign n17442 = ( n10209 & ~n17441 ) | ( n10209 & 1'b0 ) | ( ~n17441 & 1'b0 ) ;
  assign n17443 = ( n9740 & ~n17442 ) | ( n9740 & 1'b0 ) | ( ~n17442 & 1'b0 ) ;
  assign n17444 = n17439 &  n17443 ;
  assign n17445 = n17436 | n17444 ;
  assign n17446 = n17431 &  n17445 ;
  assign n17447 = ( n16808 & ~n17279 ) | ( n16808 & 1'b0 ) | ( ~n17279 & 1'b0 ) ;
  assign n17448 = ( n16808 & n16813 ) | ( n16808 & n16821 ) | ( n16813 & n16821 ) ;
  assign n17449 = ( n17447 & ~n16821 ) | ( n17447 & n17448 ) | ( ~n16821 & n17448 ) ;
  assign n17450 = ( n16808 & ~n17448 ) | ( n16808 & n17447 ) | ( ~n17448 & n17447 ) ;
  assign n17451 = ( n16813 & ~n17449 ) | ( n16813 & n17450 ) | ( ~n17449 & n17450 ) ;
  assign n17452 = ( n17446 & ~n9286 ) | ( n17446 & n17451 ) | ( ~n9286 & n17451 ) ;
  assign n17453 = ( n8839 & ~n17452 ) | ( n8839 & 1'b0 ) | ( ~n17452 & 1'b0 ) ;
  assign n17454 = n16841 | n17279 ;
  assign n17455 = ( n16828 & ~n16837 ) | ( n16828 & n16841 ) | ( ~n16837 & n16841 ) ;
  assign n17456 = ( n16837 & n17454 ) | ( n16837 & n17455 ) | ( n17454 & n17455 ) ;
  assign n17457 = ( n16841 & ~n17455 ) | ( n16841 & n17454 ) | ( ~n17455 & n17454 ) ;
  assign n17458 = ( n16828 & ~n17456 ) | ( n16828 & n17457 ) | ( ~n17456 & n17457 ) ;
  assign n17459 = ~n9286 & n17431 ;
  assign n17460 = n17445 &  n17459 ;
  assign n17461 = n17451 | n17460 ;
  assign n17462 = ( n17439 & ~n17442 ) | ( n17439 & 1'b0 ) | ( ~n17442 & 1'b0 ) ;
  assign n17463 = ( n9740 & n17436 ) | ( n9740 & n17462 ) | ( n17436 & n17462 ) ;
  assign n17464 = ( n9286 & ~n17463 ) | ( n9286 & 1'b0 ) | ( ~n17463 & 1'b0 ) ;
  assign n17465 = n8839 | n17464 ;
  assign n17466 = ( n17461 & ~n17465 ) | ( n17461 & 1'b0 ) | ( ~n17465 & 1'b0 ) ;
  assign n17467 = n17458 | n17466 ;
  assign n17468 = ~n17453 & n17467 ;
  assign n17469 = n16830 | n17279 ;
  assign n17470 = ( n16830 & ~n16843 ) | ( n16830 & n16835 ) | ( ~n16843 & n16835 ) ;
  assign n17471 = ( n16843 & n17469 ) | ( n16843 & n17470 ) | ( n17469 & n17470 ) ;
  assign n17472 = ( n16830 & ~n17470 ) | ( n16830 & n17469 ) | ( ~n17470 & n17469 ) ;
  assign n17473 = ( n16835 & ~n17471 ) | ( n16835 & n17472 ) | ( ~n17471 & n17472 ) ;
  assign n17474 = ( n17468 & ~n8407 ) | ( n17468 & n17473 ) | ( ~n8407 & n17473 ) ;
  assign n17475 = ( n7982 & ~n17474 ) | ( n7982 & 1'b0 ) | ( ~n17474 & 1'b0 ) ;
  assign n17476 = n16863 | n17279 ;
  assign n17477 = ( n16850 & ~n16863 ) | ( n16850 & n16859 ) | ( ~n16863 & n16859 ) ;
  assign n17479 = ( n16863 & n17476 ) | ( n16863 & n17477 ) | ( n17476 & n17477 ) ;
  assign n17478 = ( n16859 & ~n17477 ) | ( n16859 & n17476 ) | ( ~n17477 & n17476 ) ;
  assign n17480 = ( n16850 & ~n17479 ) | ( n16850 & n17478 ) | ( ~n17479 & n17478 ) ;
  assign n17481 = n8407 | n17453 ;
  assign n17482 = ( n17467 & ~n17481 ) | ( n17467 & 1'b0 ) | ( ~n17481 & 1'b0 ) ;
  assign n17483 = n17473 | n17482 ;
  assign n17484 = ( n17461 & ~n17464 ) | ( n17461 & 1'b0 ) | ( ~n17464 & 1'b0 ) ;
  assign n17485 = ( n17458 & ~n8839 ) | ( n17458 & n17484 ) | ( ~n8839 & n17484 ) ;
  assign n17486 = ( n8407 & ~n17485 ) | ( n8407 & 1'b0 ) | ( ~n17485 & 1'b0 ) ;
  assign n17487 = n7982 | n17486 ;
  assign n17488 = ( n17483 & ~n17487 ) | ( n17483 & 1'b0 ) | ( ~n17487 & 1'b0 ) ;
  assign n17489 = n17480 | n17488 ;
  assign n17490 = ~n17475 & n17489 ;
  assign n17491 = n16852 | n17279 ;
  assign n17492 = ( n16857 & ~n16852 ) | ( n16857 & n16865 ) | ( ~n16852 & n16865 ) ;
  assign n17494 = ( n16852 & n17491 ) | ( n16852 & n17492 ) | ( n17491 & n17492 ) ;
  assign n17493 = ( n16865 & ~n17492 ) | ( n16865 & n17491 ) | ( ~n17492 & n17491 ) ;
  assign n17495 = ( n16857 & ~n17494 ) | ( n16857 & n17493 ) | ( ~n17494 & n17493 ) ;
  assign n17496 = ( n7572 & n17490 ) | ( n7572 & n17495 ) | ( n17490 & n17495 ) ;
  assign n17497 = n7169 | n17496 ;
  assign n17499 = ( n16881 & ~n16872 ) | ( n16881 & n16885 ) | ( ~n16872 & n16885 ) ;
  assign n17498 = ( n16885 & ~n17279 ) | ( n16885 & 1'b0 ) | ( ~n17279 & 1'b0 ) ;
  assign n17501 = ( n16885 & ~n17499 ) | ( n16885 & n17498 ) | ( ~n17499 & n17498 ) ;
  assign n17500 = ( n17498 & ~n16881 ) | ( n17498 & n17499 ) | ( ~n16881 & n17499 ) ;
  assign n17502 = ( n16872 & ~n17501 ) | ( n16872 & n17500 ) | ( ~n17501 & n17500 ) ;
  assign n17503 = ( n7572 & ~n17475 ) | ( n7572 & 1'b0 ) | ( ~n17475 & 1'b0 ) ;
  assign n17504 = n17489 &  n17503 ;
  assign n17505 = n17495 | n17504 ;
  assign n17506 = ( n17483 & ~n17486 ) | ( n17483 & 1'b0 ) | ( ~n17486 & 1'b0 ) ;
  assign n17507 = ( n17480 & ~n7982 ) | ( n17480 & n17506 ) | ( ~n7982 & n17506 ) ;
  assign n17508 = n7572 | n17507 ;
  assign n17509 = n7169 &  n17508 ;
  assign n17510 = n17505 &  n17509 ;
  assign n17511 = n17502 | n17510 ;
  assign n17512 = n17497 &  n17511 ;
  assign n17513 = ( n16874 & ~n17279 ) | ( n16874 & 1'b0 ) | ( ~n17279 & 1'b0 ) ;
  assign n17514 = ( n16874 & n16879 ) | ( n16874 & n16887 ) | ( n16879 & n16887 ) ;
  assign n17515 = ( n17513 & ~n16887 ) | ( n17513 & n17514 ) | ( ~n16887 & n17514 ) ;
  assign n17516 = ( n16874 & ~n17514 ) | ( n16874 & n17513 ) | ( ~n17514 & n17513 ) ;
  assign n17517 = ( n16879 & ~n17515 ) | ( n16879 & n17516 ) | ( ~n17515 & n17516 ) ;
  assign n17518 = ( n17512 & ~n6781 ) | ( n17512 & n17517 ) | ( ~n6781 & n17517 ) ;
  assign n17519 = n6399 | n17518 ;
  assign n17520 = n16907 | n17279 ;
  assign n17521 = ( n16894 & ~n16903 ) | ( n16894 & n16907 ) | ( ~n16903 & n16907 ) ;
  assign n17522 = ( n16903 & n17520 ) | ( n16903 & n17521 ) | ( n17520 & n17521 ) ;
  assign n17523 = ( n16907 & ~n17521 ) | ( n16907 & n17520 ) | ( ~n17521 & n17520 ) ;
  assign n17524 = ( n16894 & ~n17522 ) | ( n16894 & n17523 ) | ( ~n17522 & n17523 ) ;
  assign n17525 = ~n6781 & n17497 ;
  assign n17526 = n17511 &  n17525 ;
  assign n17527 = n17517 | n17526 ;
  assign n17528 = n17505 &  n17508 ;
  assign n17529 = ( n7169 & n17502 ) | ( n7169 & n17528 ) | ( n17502 & n17528 ) ;
  assign n17530 = ( n6781 & ~n17529 ) | ( n6781 & 1'b0 ) | ( ~n17529 & 1'b0 ) ;
  assign n17531 = ( n6399 & ~n17530 ) | ( n6399 & 1'b0 ) | ( ~n17530 & 1'b0 ) ;
  assign n17532 = n17527 &  n17531 ;
  assign n17533 = n17524 | n17532 ;
  assign n17534 = n17519 &  n17533 ;
  assign n17535 = ( n16896 & ~n17279 ) | ( n16896 & 1'b0 ) | ( ~n17279 & 1'b0 ) ;
  assign n17536 = ( n16896 & n16901 ) | ( n16896 & n16909 ) | ( n16901 & n16909 ) ;
  assign n17537 = ( n17535 & ~n16909 ) | ( n17535 & n17536 ) | ( ~n16909 & n17536 ) ;
  assign n17538 = ( n16896 & ~n17536 ) | ( n16896 & n17535 ) | ( ~n17536 & n17535 ) ;
  assign n17539 = ( n16901 & ~n17537 ) | ( n16901 & n17538 ) | ( ~n17537 & n17538 ) ;
  assign n17540 = ( n17534 & ~n6032 ) | ( n17534 & n17539 ) | ( ~n6032 & n17539 ) ;
  assign n17541 = n5672 | n17540 ;
  assign n17542 = n16929 | n17279 ;
  assign n17543 = ( n16916 & ~n16925 ) | ( n16916 & n16929 ) | ( ~n16925 & n16929 ) ;
  assign n17544 = ( n16925 & n17542 ) | ( n16925 & n17543 ) | ( n17542 & n17543 ) ;
  assign n17545 = ( n16929 & ~n17543 ) | ( n16929 & n17542 ) | ( ~n17543 & n17542 ) ;
  assign n17546 = ( n16916 & ~n17544 ) | ( n16916 & n17545 ) | ( ~n17544 & n17545 ) ;
  assign n17547 = ~n6032 & n17519 ;
  assign n17548 = n17533 &  n17547 ;
  assign n17549 = n17539 | n17548 ;
  assign n17550 = ( n17527 & ~n17530 ) | ( n17527 & 1'b0 ) | ( ~n17530 & 1'b0 ) ;
  assign n17551 = ( n6399 & n17524 ) | ( n6399 & n17550 ) | ( n17524 & n17550 ) ;
  assign n17552 = ( n6032 & ~n17551 ) | ( n6032 & 1'b0 ) | ( ~n17551 & 1'b0 ) ;
  assign n17553 = ( n5672 & ~n17552 ) | ( n5672 & 1'b0 ) | ( ~n17552 & 1'b0 ) ;
  assign n17554 = n17549 &  n17553 ;
  assign n17555 = n17546 | n17554 ;
  assign n17556 = n17541 &  n17555 ;
  assign n17557 = ( n16918 & ~n17279 ) | ( n16918 & 1'b0 ) | ( ~n17279 & 1'b0 ) ;
  assign n17558 = ( n16918 & n16923 ) | ( n16918 & n16931 ) | ( n16923 & n16931 ) ;
  assign n17559 = ( n17557 & ~n16931 ) | ( n17557 & n17558 ) | ( ~n16931 & n17558 ) ;
  assign n17560 = ( n16918 & ~n17558 ) | ( n16918 & n17557 ) | ( ~n17558 & n17557 ) ;
  assign n17561 = ( n16923 & ~n17559 ) | ( n16923 & n17560 ) | ( ~n17559 & n17560 ) ;
  assign n17562 = ( n17556 & ~n5327 ) | ( n17556 & n17561 ) | ( ~n5327 & n17561 ) ;
  assign n17563 = ( n4990 & ~n17562 ) | ( n4990 & 1'b0 ) | ( ~n17562 & 1'b0 ) ;
  assign n17564 = n16951 | n17279 ;
  assign n17565 = ( n16938 & ~n16947 ) | ( n16938 & n16951 ) | ( ~n16947 & n16951 ) ;
  assign n17566 = ( n16947 & n17564 ) | ( n16947 & n17565 ) | ( n17564 & n17565 ) ;
  assign n17567 = ( n16951 & ~n17565 ) | ( n16951 & n17564 ) | ( ~n17565 & n17564 ) ;
  assign n17568 = ( n16938 & ~n17566 ) | ( n16938 & n17567 ) | ( ~n17566 & n17567 ) ;
  assign n17569 = ~n5327 & n17541 ;
  assign n17570 = n17555 &  n17569 ;
  assign n17571 = n17561 | n17570 ;
  assign n17572 = ( n17549 & ~n17552 ) | ( n17549 & 1'b0 ) | ( ~n17552 & 1'b0 ) ;
  assign n17573 = ( n5672 & n17546 ) | ( n5672 & n17572 ) | ( n17546 & n17572 ) ;
  assign n17574 = ( n5327 & ~n17573 ) | ( n5327 & 1'b0 ) | ( ~n17573 & 1'b0 ) ;
  assign n17575 = n4990 | n17574 ;
  assign n17576 = ( n17571 & ~n17575 ) | ( n17571 & 1'b0 ) | ( ~n17575 & 1'b0 ) ;
  assign n17577 = n17568 | n17576 ;
  assign n17578 = ~n17563 & n17577 ;
  assign n17579 = n16940 | n17279 ;
  assign n17580 = ( n16945 & ~n16940 ) | ( n16945 & n16953 ) | ( ~n16940 & n16953 ) ;
  assign n17582 = ( n16940 & n17579 ) | ( n16940 & n17580 ) | ( n17579 & n17580 ) ;
  assign n17581 = ( n16953 & ~n17580 ) | ( n16953 & n17579 ) | ( ~n17580 & n17579 ) ;
  assign n17583 = ( n16945 & ~n17582 ) | ( n16945 & n17581 ) | ( ~n17582 & n17581 ) ;
  assign n17584 = ( n17578 & ~n4668 ) | ( n17578 & n17583 ) | ( ~n4668 & n17583 ) ;
  assign n17585 = ( n4353 & ~n17584 ) | ( n4353 & 1'b0 ) | ( ~n17584 & 1'b0 ) ;
  assign n17586 = n16973 | n17279 ;
  assign n17587 = ( n16960 & ~n16969 ) | ( n16960 & n16973 ) | ( ~n16969 & n16973 ) ;
  assign n17588 = ( n16969 & n17586 ) | ( n16969 & n17587 ) | ( n17586 & n17587 ) ;
  assign n17589 = ( n16973 & ~n17587 ) | ( n16973 & n17586 ) | ( ~n17587 & n17586 ) ;
  assign n17590 = ( n16960 & ~n17588 ) | ( n16960 & n17589 ) | ( ~n17588 & n17589 ) ;
  assign n17591 = n4668 | n17563 ;
  assign n17592 = ( n17577 & ~n17591 ) | ( n17577 & 1'b0 ) | ( ~n17591 & 1'b0 ) ;
  assign n17593 = n17583 | n17592 ;
  assign n17594 = ( n17571 & ~n17574 ) | ( n17571 & 1'b0 ) | ( ~n17574 & 1'b0 ) ;
  assign n17595 = ( n17568 & ~n4990 ) | ( n17568 & n17594 ) | ( ~n4990 & n17594 ) ;
  assign n17596 = ( n4668 & ~n17595 ) | ( n4668 & 1'b0 ) | ( ~n17595 & 1'b0 ) ;
  assign n17597 = n4353 | n17596 ;
  assign n17598 = ( n17593 & ~n17597 ) | ( n17593 & 1'b0 ) | ( ~n17597 & 1'b0 ) ;
  assign n17599 = n17590 | n17598 ;
  assign n17600 = ~n17585 & n17599 ;
  assign n17601 = n16962 | n17279 ;
  assign n17602 = ( n16962 & ~n16975 ) | ( n16962 & n16967 ) | ( ~n16975 & n16967 ) ;
  assign n17603 = ( n16975 & n17601 ) | ( n16975 & n17602 ) | ( n17601 & n17602 ) ;
  assign n17604 = ( n16962 & ~n17602 ) | ( n16962 & n17601 ) | ( ~n17602 & n17601 ) ;
  assign n17605 = ( n16967 & ~n17603 ) | ( n16967 & n17604 ) | ( ~n17603 & n17604 ) ;
  assign n17606 = ( n4053 & ~n17600 ) | ( n4053 & n17605 ) | ( ~n17600 & n17605 ) ;
  assign n17607 = n3760 &  n17606 ;
  assign n17609 = ( n16991 & ~n16982 ) | ( n16991 & n16995 ) | ( ~n16982 & n16995 ) ;
  assign n17608 = n16995 | n17279 ;
  assign n17611 = ( n16995 & ~n17609 ) | ( n16995 & n17608 ) | ( ~n17609 & n17608 ) ;
  assign n17610 = ( n17608 & ~n16991 ) | ( n17608 & n17609 ) | ( ~n16991 & n17609 ) ;
  assign n17612 = ( n16982 & ~n17611 ) | ( n16982 & n17610 ) | ( ~n17611 & n17610 ) ;
  assign n17613 = n4053 | n17585 ;
  assign n17614 = ( n17599 & ~n17613 ) | ( n17599 & 1'b0 ) | ( ~n17613 & 1'b0 ) ;
  assign n17615 = ( n17605 & ~n17614 ) | ( n17605 & 1'b0 ) | ( ~n17614 & 1'b0 ) ;
  assign n17616 = ( n17593 & ~n17596 ) | ( n17593 & 1'b0 ) | ( ~n17596 & 1'b0 ) ;
  assign n17617 = ( n17590 & ~n4353 ) | ( n17590 & n17616 ) | ( ~n4353 & n17616 ) ;
  assign n17618 = ( n4053 & ~n17617 ) | ( n4053 & 1'b0 ) | ( ~n17617 & 1'b0 ) ;
  assign n17619 = n3760 | n17618 ;
  assign n17620 = n17615 | n17619 ;
  assign n17621 = n17612 &  n17620 ;
  assign n17622 = n17607 | n17621 ;
  assign n17623 = n16984 | n17279 ;
  assign n17624 = ( n16984 & n16989 ) | ( n16984 & n16997 ) | ( n16989 & n16997 ) ;
  assign n17625 = ( n17623 & ~n16997 ) | ( n17623 & n17624 ) | ( ~n16997 & n17624 ) ;
  assign n17626 = ( n16984 & ~n17624 ) | ( n16984 & n17623 ) | ( ~n17624 & n17623 ) ;
  assign n17627 = ( n16989 & ~n17625 ) | ( n16989 & n17626 ) | ( ~n17625 & n17626 ) ;
  assign n17628 = ( n3482 & n17622 ) | ( n3482 & n17627 ) | ( n17622 & n17627 ) ;
  assign n17629 = n3211 &  n17628 ;
  assign n17631 = ( n17013 & ~n17004 ) | ( n17013 & n17017 ) | ( ~n17004 & n17017 ) ;
  assign n17630 = n17017 | n17279 ;
  assign n17633 = ( n17017 & ~n17631 ) | ( n17017 & n17630 ) | ( ~n17631 & n17630 ) ;
  assign n17632 = ( n17630 & ~n17013 ) | ( n17630 & n17631 ) | ( ~n17013 & n17631 ) ;
  assign n17634 = ( n17004 & ~n17633 ) | ( n17004 & n17632 ) | ( ~n17633 & n17632 ) ;
  assign n17635 = n3482 | n17607 ;
  assign n17636 = n17621 | n17635 ;
  assign n17637 = n17627 &  n17636 ;
  assign n17638 = n17615 | n17618 ;
  assign n17639 = ( n3760 & n17612 ) | ( n3760 & n17638 ) | ( n17612 & n17638 ) ;
  assign n17640 = n3482 &  n17639 ;
  assign n17641 = n3211 | n17640 ;
  assign n17642 = n17637 | n17641 ;
  assign n17643 = n17634 &  n17642 ;
  assign n17644 = n17629 | n17643 ;
  assign n17645 = n17006 | n17279 ;
  assign n17646 = ( n17006 & n17011 ) | ( n17006 & n17019 ) | ( n17011 & n17019 ) ;
  assign n17647 = ( n17645 & ~n17019 ) | ( n17645 & n17646 ) | ( ~n17019 & n17646 ) ;
  assign n17648 = ( n17006 & ~n17646 ) | ( n17006 & n17645 ) | ( ~n17646 & n17645 ) ;
  assign n17649 = ( n17011 & ~n17647 ) | ( n17011 & n17648 ) | ( ~n17647 & n17648 ) ;
  assign n17650 = ( n2955 & n17644 ) | ( n2955 & n17649 ) | ( n17644 & n17649 ) ;
  assign n17651 = n2706 &  n17650 ;
  assign n17652 = n17039 | n17279 ;
  assign n17653 = ( n17026 & n17035 ) | ( n17026 & n17039 ) | ( n17035 & n17039 ) ;
  assign n17654 = ( n17652 & ~n17035 ) | ( n17652 & n17653 ) | ( ~n17035 & n17653 ) ;
  assign n17655 = ( n17039 & ~n17653 ) | ( n17039 & n17652 ) | ( ~n17653 & n17652 ) ;
  assign n17656 = ( n17026 & ~n17654 ) | ( n17026 & n17655 ) | ( ~n17654 & n17655 ) ;
  assign n17657 = n2955 | n17629 ;
  assign n17658 = n17643 | n17657 ;
  assign n17659 = n17649 &  n17658 ;
  assign n17660 = n17637 | n17640 ;
  assign n17661 = ( n3211 & n17634 ) | ( n3211 & n17660 ) | ( n17634 & n17660 ) ;
  assign n17662 = n2955 &  n17661 ;
  assign n17663 = n2706 | n17662 ;
  assign n17664 = n17659 | n17663 ;
  assign n17665 = ~n17656 & n17664 ;
  assign n17666 = n17651 | n17665 ;
  assign n17672 = ( n2472 & ~n17671 ) | ( n2472 & n17666 ) | ( ~n17671 & n17666 ) ;
  assign n17673 = n2245 &  n17672 ;
  assign n17675 = ( n17057 & ~n17048 ) | ( n17057 & n17061 ) | ( ~n17048 & n17061 ) ;
  assign n17674 = n17061 | n17279 ;
  assign n17677 = ( n17061 & ~n17675 ) | ( n17061 & n17674 ) | ( ~n17675 & n17674 ) ;
  assign n17676 = ( n17674 & ~n17057 ) | ( n17674 & n17675 ) | ( ~n17057 & n17675 ) ;
  assign n17678 = ( n17048 & ~n17677 ) | ( n17048 & n17676 ) | ( ~n17677 & n17676 ) ;
  assign n17679 = n2472 | n17651 ;
  assign n17680 = n17665 | n17679 ;
  assign n17681 = ~n17671 & n17680 ;
  assign n17682 = n17659 | n17662 ;
  assign n17683 = ( n2706 & ~n17656 ) | ( n2706 & n17682 ) | ( ~n17656 & n17682 ) ;
  assign n17684 = n2472 &  n17683 ;
  assign n17685 = n2245 | n17684 ;
  assign n17686 = n17681 | n17685 ;
  assign n17687 = n17678 &  n17686 ;
  assign n17688 = n17673 | n17687 ;
  assign n17690 = ( n17050 & ~n17055 ) | ( n17050 & n17063 ) | ( ~n17055 & n17063 ) ;
  assign n17689 = n17050 | n17279 ;
  assign n17692 = ( n17050 & ~n17690 ) | ( n17050 & n17689 ) | ( ~n17690 & n17689 ) ;
  assign n17691 = ( n17689 & ~n17063 ) | ( n17689 & n17690 ) | ( ~n17063 & n17690 ) ;
  assign n17693 = ( n17055 & ~n17692 ) | ( n17055 & n17691 ) | ( ~n17692 & n17691 ) ;
  assign n17694 = ( n2033 & ~n17688 ) | ( n2033 & n17693 ) | ( ~n17688 & n17693 ) ;
  assign n17695 = ( n1827 & ~n17694 ) | ( n1827 & 1'b0 ) | ( ~n17694 & 1'b0 ) ;
  assign n17696 = n17083 | n17279 ;
  assign n17697 = ( n17070 & ~n17083 ) | ( n17070 & n17079 ) | ( ~n17083 & n17079 ) ;
  assign n17699 = ( n17083 & n17696 ) | ( n17083 & n17697 ) | ( n17696 & n17697 ) ;
  assign n17698 = ( n17079 & ~n17697 ) | ( n17079 & n17696 ) | ( ~n17697 & n17696 ) ;
  assign n17700 = ( n17070 & ~n17699 ) | ( n17070 & n17698 ) | ( ~n17699 & n17698 ) ;
  assign n17701 = ( n2033 & ~n17673 ) | ( n2033 & 1'b0 ) | ( ~n17673 & 1'b0 ) ;
  assign n17702 = ~n17687 & n17701 ;
  assign n17703 = n17693 | n17702 ;
  assign n17704 = n17681 | n17684 ;
  assign n17705 = ( n2245 & n17678 ) | ( n2245 & n17704 ) | ( n17678 & n17704 ) ;
  assign n17706 = ~n2033 & n17705 ;
  assign n17707 = n1827 | n17706 ;
  assign n17708 = ( n17703 & ~n17707 ) | ( n17703 & 1'b0 ) | ( ~n17707 & 1'b0 ) ;
  assign n17709 = ( n17700 & ~n17708 ) | ( n17700 & 1'b0 ) | ( ~n17708 & 1'b0 ) ;
  assign n17710 = n17695 | n17709 ;
  assign n17711 = n17072 | n17279 ;
  assign n17712 = ( n17072 & n17077 ) | ( n17072 & n17085 ) | ( n17077 & n17085 ) ;
  assign n17713 = ( n17711 & ~n17085 ) | ( n17711 & n17712 ) | ( ~n17085 & n17712 ) ;
  assign n17714 = ( n17072 & ~n17712 ) | ( n17072 & n17711 ) | ( ~n17712 & n17711 ) ;
  assign n17715 = ( n17077 & ~n17713 ) | ( n17077 & n17714 ) | ( ~n17713 & n17714 ) ;
  assign n17716 = ( n17710 & ~n1636 ) | ( n17710 & n17715 ) | ( ~n1636 & n17715 ) ;
  assign n17717 = ~n1452 & n17716 ;
  assign n17718 = n17105 | n17279 ;
  assign n17719 = ( n17092 & ~n17101 ) | ( n17092 & n17105 ) | ( ~n17101 & n17105 ) ;
  assign n17720 = ( n17101 & n17718 ) | ( n17101 & n17719 ) | ( n17718 & n17719 ) ;
  assign n17721 = ( n17105 & ~n17719 ) | ( n17105 & n17718 ) | ( ~n17719 & n17718 ) ;
  assign n17722 = ( n17092 & ~n17720 ) | ( n17092 & n17721 ) | ( ~n17720 & n17721 ) ;
  assign n17723 = ( n1636 & ~n17695 ) | ( n1636 & 1'b0 ) | ( ~n17695 & 1'b0 ) ;
  assign n17724 = ~n17709 & n17723 ;
  assign n17725 = ( n17715 & ~n17724 ) | ( n17715 & 1'b0 ) | ( ~n17724 & 1'b0 ) ;
  assign n17726 = ( n17703 & ~n17706 ) | ( n17703 & 1'b0 ) | ( ~n17706 & 1'b0 ) ;
  assign n17727 = ( n1827 & ~n17726 ) | ( n1827 & n17700 ) | ( ~n17726 & n17700 ) ;
  assign n17728 = ~n1636 & n17727 ;
  assign n17729 = ( n1452 & ~n17728 ) | ( n1452 & 1'b0 ) | ( ~n17728 & 1'b0 ) ;
  assign n17730 = ~n17725 & n17729 ;
  assign n17731 = n17722 | n17730 ;
  assign n17732 = ~n17717 & n17731 ;
  assign n17733 = ( n17094 & ~n17279 ) | ( n17094 & 1'b0 ) | ( ~n17279 & 1'b0 ) ;
  assign n17734 = ( n17094 & n17099 ) | ( n17094 & n17107 ) | ( n17099 & n17107 ) ;
  assign n17735 = ( n17733 & ~n17107 ) | ( n17733 & n17734 ) | ( ~n17107 & n17734 ) ;
  assign n17736 = ( n17094 & ~n17734 ) | ( n17094 & n17733 ) | ( ~n17734 & n17733 ) ;
  assign n17737 = ( n17099 & ~n17735 ) | ( n17099 & n17736 ) | ( ~n17735 & n17736 ) ;
  assign n17738 = ( n17732 & ~n1283 ) | ( n17732 & n17737 ) | ( ~n1283 & n17737 ) ;
  assign n17739 = n1122 | n17738 ;
  assign n17740 = n17127 | n17279 ;
  assign n17741 = ( n17114 & ~n17123 ) | ( n17114 & n17127 ) | ( ~n17123 & n17127 ) ;
  assign n17742 = ( n17123 & n17740 ) | ( n17123 & n17741 ) | ( n17740 & n17741 ) ;
  assign n17743 = ( n17127 & ~n17741 ) | ( n17127 & n17740 ) | ( ~n17741 & n17740 ) ;
  assign n17744 = ( n17114 & ~n17742 ) | ( n17114 & n17743 ) | ( ~n17742 & n17743 ) ;
  assign n17745 = n1283 | n17717 ;
  assign n17746 = ( n17731 & ~n17745 ) | ( n17731 & 1'b0 ) | ( ~n17745 & 1'b0 ) ;
  assign n17747 = n17737 | n17746 ;
  assign n17748 = n17725 | n17728 ;
  assign n17749 = ( n1452 & ~n17748 ) | ( n1452 & n17722 ) | ( ~n17748 & n17722 ) ;
  assign n17750 = ( n1283 & ~n17749 ) | ( n1283 & 1'b0 ) | ( ~n17749 & 1'b0 ) ;
  assign n17751 = ( n1122 & ~n17750 ) | ( n1122 & 1'b0 ) | ( ~n17750 & 1'b0 ) ;
  assign n17752 = n17747 &  n17751 ;
  assign n17753 = n17744 | n17752 ;
  assign n17754 = n17739 &  n17753 ;
  assign n17755 = ( n17116 & ~n17279 ) | ( n17116 & 1'b0 ) | ( ~n17279 & 1'b0 ) ;
  assign n17756 = ( n17116 & n17121 ) | ( n17116 & n17129 ) | ( n17121 & n17129 ) ;
  assign n17757 = ( n17755 & ~n17129 ) | ( n17755 & n17756 ) | ( ~n17129 & n17756 ) ;
  assign n17758 = ( n17116 & ~n17756 ) | ( n17116 & n17755 ) | ( ~n17756 & n17755 ) ;
  assign n17759 = ( n17121 & ~n17757 ) | ( n17121 & n17758 ) | ( ~n17757 & n17758 ) ;
  assign n17760 = ( n976 & n17754 ) | ( n976 & n17759 ) | ( n17754 & n17759 ) ;
  assign n17761 = ( n837 & ~n17760 ) | ( n837 & 1'b0 ) | ( ~n17760 & 1'b0 ) ;
  assign n17763 = ( n17145 & ~n17136 ) | ( n17145 & n17149 ) | ( ~n17136 & n17149 ) ;
  assign n17762 = ( n17149 & ~n17279 ) | ( n17149 & 1'b0 ) | ( ~n17279 & 1'b0 ) ;
  assign n17765 = ( n17149 & ~n17763 ) | ( n17149 & n17762 ) | ( ~n17763 & n17762 ) ;
  assign n17764 = ( n17762 & ~n17145 ) | ( n17762 & n17763 ) | ( ~n17145 & n17763 ) ;
  assign n17766 = ( n17136 & ~n17765 ) | ( n17136 & n17764 ) | ( ~n17765 & n17764 ) ;
  assign n17767 = n976 &  n17739 ;
  assign n17768 = n17753 &  n17767 ;
  assign n17769 = n17759 | n17768 ;
  assign n17770 = ( n17747 & ~n17750 ) | ( n17747 & 1'b0 ) | ( ~n17750 & 1'b0 ) ;
  assign n17771 = ( n1122 & n17744 ) | ( n1122 & n17770 ) | ( n17744 & n17770 ) ;
  assign n17772 = n976 | n17771 ;
  assign n17773 = ~n837 & n17772 ;
  assign n17774 = n17769 &  n17773 ;
  assign n17775 = n17766 | n17774 ;
  assign n17776 = ~n17761 & n17775 ;
  assign n17777 = n17138 | n17279 ;
  assign n17778 = ( n17138 & ~n17151 ) | ( n17138 & n17143 ) | ( ~n17151 & n17143 ) ;
  assign n17779 = ( n17151 & n17777 ) | ( n17151 & n17778 ) | ( n17777 & n17778 ) ;
  assign n17780 = ( n17138 & ~n17778 ) | ( n17138 & n17777 ) | ( ~n17778 & n17777 ) ;
  assign n17781 = ( n17143 & ~n17779 ) | ( n17143 & n17780 ) | ( ~n17779 & n17780 ) ;
  assign n17782 = ( n713 & ~n17776 ) | ( n713 & n17781 ) | ( ~n17776 & n17781 ) ;
  assign n17783 = n595 &  n17782 ;
  assign n17789 = n713 | n17761 ;
  assign n17790 = ( n17775 & ~n17789 ) | ( n17775 & 1'b0 ) | ( ~n17789 & 1'b0 ) ;
  assign n17791 = ( n17781 & ~n17790 ) | ( n17781 & 1'b0 ) | ( ~n17790 & 1'b0 ) ;
  assign n17792 = n17769 &  n17772 ;
  assign n17793 = ( n17766 & ~n837 ) | ( n17766 & n17792 ) | ( ~n837 & n17792 ) ;
  assign n17794 = ( n713 & ~n17793 ) | ( n713 & 1'b0 ) | ( ~n17793 & 1'b0 ) ;
  assign n17795 = n595 | n17794 ;
  assign n17796 = n17791 | n17795 ;
  assign n18430 = ( n17783 & ~n17788 ) | ( n17783 & n17796 ) | ( ~n17788 & n17796 ) ;
  assign n17870 = n17245 &  n17261 ;
  assign n17871 = ( n17264 & n17279 ) | ( n17264 & n17870 ) | ( n17279 & n17870 ) ;
  assign n17872 = ~n17264 & n17871 ;
  assign n17873 = ( n17261 & ~n17264 ) | ( n17261 & 1'b0 ) | ( ~n17264 & 1'b0 ) ;
  assign n17874 = ~n17279 & n17873 ;
  assign n17875 = ( n17245 & ~n17874 ) | ( n17245 & n17873 ) | ( ~n17874 & n17873 ) ;
  assign n17876 = ~n17872 & n17875 ;
  assign n17877 = ( n17246 & ~n17253 ) | ( n17246 & 1'b0 ) | ( ~n17253 & 1'b0 ) ;
  assign n17878 = ~n17279 & n17877 ;
  assign n17879 = ( n17267 & ~n17878 ) | ( n17267 & n17877 ) | ( ~n17878 & n17877 ) ;
  assign n17880 = n17876 | n17879 ;
  assign n17820 = ~n17194 & n17279 ;
  assign n17821 = ( n17181 & n17186 ) | ( n17181 & n17279 ) | ( n17186 & n17279 ) ;
  assign n17823 = ( n17820 & ~n17181 ) | ( n17820 & n17821 ) | ( ~n17181 & n17821 ) ;
  assign n17822 = ( n17279 & ~n17821 ) | ( n17279 & n17820 ) | ( ~n17821 & n17820 ) ;
  assign n17824 = ( n17186 & ~n17823 ) | ( n17186 & n17822 ) | ( ~n17823 & n17822 ) ;
  assign n17799 = ( n17160 & n17168 ) | ( n17160 & n17172 ) | ( n17168 & n17172 ) ;
  assign n17801 = ( n17279 & ~n17168 ) | ( n17279 & n17799 ) | ( ~n17168 & n17799 ) ;
  assign n17800 = ( n17160 & ~n17799 ) | ( n17160 & n17279 ) | ( ~n17799 & n17279 ) ;
  assign n17802 = ( n17172 & ~n17801 ) | ( n17172 & n17800 ) | ( ~n17801 & n17800 ) ;
  assign n17797 = ~n17788 & n17796 ;
  assign n17798 = n17783 | n17797 ;
  assign n17803 = ( n492 & ~n17802 ) | ( n492 & n17798 ) | ( ~n17802 & n17798 ) ;
  assign n17804 = n396 &  n17803 ;
  assign n17805 = n17192 | n17279 ;
  assign n17806 = ( n17179 & n17188 ) | ( n17179 & n17192 ) | ( n17188 & n17192 ) ;
  assign n17807 = ( n17805 & ~n17188 ) | ( n17805 & n17806 ) | ( ~n17188 & n17806 ) ;
  assign n17808 = ( n17192 & ~n17806 ) | ( n17192 & n17805 ) | ( ~n17806 & n17805 ) ;
  assign n17809 = ( n17179 & ~n17807 ) | ( n17179 & n17808 ) | ( ~n17807 & n17808 ) ;
  assign n17810 = n492 | n17783 ;
  assign n17811 = n17797 | n17810 ;
  assign n17812 = ~n17802 & n17811 ;
  assign n17813 = n17791 | n17794 ;
  assign n17814 = ( n595 & ~n17788 ) | ( n595 & n17813 ) | ( ~n17788 & n17813 ) ;
  assign n17815 = n492 &  n17814 ;
  assign n17816 = n396 | n17815 ;
  assign n17817 = n17812 | n17816 ;
  assign n17818 = n17809 &  n17817 ;
  assign n17819 = n17804 | n17818 ;
  assign n17825 = ( n315 & ~n17824 ) | ( n315 & n17819 ) | ( ~n17824 & n17819 ) ;
  assign n17826 = n240 &  n17825 ;
  assign n17827 = n17214 | n17279 ;
  assign n17828 = ( n17201 & n17210 ) | ( n17201 & n17214 ) | ( n17210 & n17214 ) ;
  assign n17829 = ( n17827 & ~n17210 ) | ( n17827 & n17828 ) | ( ~n17210 & n17828 ) ;
  assign n17830 = ( n17214 & ~n17828 ) | ( n17214 & n17827 ) | ( ~n17828 & n17827 ) ;
  assign n17831 = ( n17201 & ~n17829 ) | ( n17201 & n17830 ) | ( ~n17829 & n17830 ) ;
  assign n17832 = n315 | n17804 ;
  assign n17833 = n17818 | n17832 ;
  assign n17834 = ~n17824 & n17833 ;
  assign n17835 = n17812 | n17815 ;
  assign n17836 = ( n396 & n17809 ) | ( n396 & n17835 ) | ( n17809 & n17835 ) ;
  assign n17837 = n315 &  n17836 ;
  assign n17838 = n240 | n17837 ;
  assign n17839 = n17834 | n17838 ;
  assign n17840 = n17831 &  n17839 ;
  assign n17841 = n17826 | n17840 ;
  assign n17842 = ~n17216 & n17279 ;
  assign n17843 = ( n17203 & ~n17842 ) | ( n17203 & n17279 ) | ( ~n17842 & n17279 ) ;
  assign n17844 = ( n17203 & ~n17843 ) | ( n17203 & n17208 ) | ( ~n17843 & n17208 ) ;
  assign n17845 = ( n17208 & ~n17203 ) | ( n17208 & n17843 ) | ( ~n17203 & n17843 ) ;
  assign n17846 = ( n17844 & ~n17208 ) | ( n17844 & n17845 ) | ( ~n17208 & n17845 ) ;
  assign n17847 = ( n181 & n17841 ) | ( n181 & n17846 ) | ( n17841 & n17846 ) ;
  assign n17848 = ~n145 & n17847 ;
  assign n17849 = n17236 | n17279 ;
  assign n17850 = ( n17223 & n17232 ) | ( n17223 & n17236 ) | ( n17232 & n17236 ) ;
  assign n17851 = ( n17849 & ~n17232 ) | ( n17849 & n17850 ) | ( ~n17232 & n17850 ) ;
  assign n17852 = ( n17236 & ~n17850 ) | ( n17236 & n17849 ) | ( ~n17850 & n17849 ) ;
  assign n17853 = ( n17223 & ~n17851 ) | ( n17223 & n17852 ) | ( ~n17851 & n17852 ) ;
  assign n17854 = n181 | n17826 ;
  assign n17855 = n17840 | n17854 ;
  assign n17856 = n17846 &  n17855 ;
  assign n17857 = n17834 | n17837 ;
  assign n17858 = ( n240 & n17831 ) | ( n240 & n17857 ) | ( n17831 & n17857 ) ;
  assign n17859 = n181 &  n17858 ;
  assign n17860 = ( n145 & ~n17859 ) | ( n145 & 1'b0 ) | ( ~n17859 & 1'b0 ) ;
  assign n17861 = ~n17856 & n17860 ;
  assign n17862 = n17853 | n17861 ;
  assign n17863 = ~n17848 & n17862 ;
  assign n17864 = n17225 | n17279 ;
  assign n17865 = ( n17230 & ~n17225 ) | ( n17230 & n17238 ) | ( ~n17225 & n17238 ) ;
  assign n17867 = ( n17225 & n17864 ) | ( n17225 & n17865 ) | ( n17864 & n17865 ) ;
  assign n17866 = ( n17238 & ~n17865 ) | ( n17238 & n17864 ) | ( ~n17865 & n17864 ) ;
  assign n17868 = ( n17230 & ~n17867 ) | ( n17230 & n17866 ) | ( ~n17867 & n17866 ) ;
  assign n17869 = ( n150 & ~n17863 ) | ( n150 & n17868 ) | ( ~n17863 & n17868 ) ;
  assign n17881 = n17869 | n17880 ;
  assign n17882 = ( n133 & ~n17880 ) | ( n133 & n17881 ) | ( ~n17880 & n17881 ) ;
  assign n17885 = n17856 | n17859 ;
  assign n17886 = ( n145 & ~n17885 ) | ( n145 & n17853 ) | ( ~n17885 & n17853 ) ;
  assign n17887 = ( n150 & ~n17886 ) | ( n150 & 1'b0 ) | ( ~n17886 & 1'b0 ) ;
  assign n17888 = ( n17876 & ~n17887 ) | ( n17876 & 1'b0 ) | ( ~n17887 & 1'b0 ) ;
  assign n17883 = n150 | n17848 ;
  assign n17884 = ( n17862 & ~n17883 ) | ( n17862 & 1'b0 ) | ( ~n17883 & 1'b0 ) ;
  assign n17889 = n17868 &  n17884 ;
  assign n17890 = ( n17888 & ~n17868 ) | ( n17888 & n17889 ) | ( ~n17868 & n17889 ) ;
  assign n17892 = ( n133 & ~n17253 ) | ( n133 & n17246 ) | ( ~n17253 & n17246 ) ;
  assign n17891 = ( n17253 & ~n17246 ) | ( n17253 & n17279 ) | ( ~n17246 & n17279 ) ;
  assign n17893 = ~n17253 & n17891 ;
  assign n17894 = ( n17253 & n17892 ) | ( n17253 & n17893 ) | ( n17892 & n17893 ) ;
  assign n17895 = n17249 | n17276 ;
  assign n17896 = ( n17252 & n17271 ) | ( n17252 & n17895 ) | ( n17271 & n17895 ) ;
  assign n17897 = ( n17252 & ~n17896 ) | ( n17252 & 1'b0 ) | ( ~n17896 & 1'b0 ) ;
  assign n17898 = ( n17259 & ~n17897 ) | ( n17259 & n17267 ) | ( ~n17897 & n17267 ) ;
  assign n17899 = ( n17259 & ~n17898 ) | ( n17259 & 1'b0 ) | ( ~n17898 & 1'b0 ) ;
  assign n17900 = n17894 | n17899 ;
  assign n17901 = n17890 | n17900 ;
  assign n17902 = ~n17882 |  n17901 ;
  assign n18429 = n17783 | n17902 ;
  assign n18432 = ( n17783 & ~n18430 ) | ( n17783 & n18429 ) | ( ~n18430 & n18429 ) ;
  assign n18431 = ( n18429 & ~n17796 ) | ( n18429 & n18430 ) | ( ~n17796 & n18430 ) ;
  assign n18433 = ( n17788 & ~n18432 ) | ( n17788 & n18431 ) | ( ~n18432 & n18431 ) ;
  assign n18407 = n17761 | n17902 ;
  assign n18408 = ( n17766 & ~n17761 ) | ( n17766 & n17774 ) | ( ~n17761 & n17774 ) ;
  assign n18410 = ( n17761 & n18407 ) | ( n17761 & n18408 ) | ( n18407 & n18408 ) ;
  assign n18409 = ( n17774 & ~n18408 ) | ( n17774 & n18407 ) | ( ~n18408 & n18407 ) ;
  assign n18411 = ( n17766 & ~n18410 ) | ( n17766 & n18409 ) | ( ~n18410 & n18409 ) ;
  assign n18393 = ( n17768 & ~n17759 ) | ( n17768 & n17772 ) | ( ~n17759 & n17772 ) ;
  assign n18392 = ( n17772 & ~n17902 ) | ( n17772 & 1'b0 ) | ( ~n17902 & 1'b0 ) ;
  assign n18395 = ( n17772 & ~n18393 ) | ( n17772 & n18392 ) | ( ~n18393 & n18392 ) ;
  assign n18394 = ( n18392 & ~n17768 ) | ( n18392 & n18393 ) | ( ~n17768 & n18393 ) ;
  assign n18396 = ( n17759 & ~n18395 ) | ( n17759 & n18394 ) | ( ~n18395 & n18394 ) ;
  assign n18385 = ( n17739 & ~n17902 ) | ( n17739 & 1'b0 ) | ( ~n17902 & 1'b0 ) ;
  assign n18386 = ( n17739 & n17744 ) | ( n17739 & n17752 ) | ( n17744 & n17752 ) ;
  assign n18387 = ( n18385 & ~n17752 ) | ( n18385 & n18386 ) | ( ~n17752 & n18386 ) ;
  assign n18388 = ( n17739 & ~n18386 ) | ( n17739 & n18385 ) | ( ~n18386 & n18385 ) ;
  assign n18389 = ( n17744 & ~n18387 ) | ( n17744 & n18388 ) | ( ~n18387 & n18388 ) ;
  assign n18370 = n17750 | n17902 ;
  assign n18371 = ( n17737 & ~n17746 ) | ( n17737 & n17750 ) | ( ~n17746 & n17750 ) ;
  assign n18372 = ( n17746 & n18370 ) | ( n17746 & n18371 ) | ( n18370 & n18371 ) ;
  assign n18373 = ( n17750 & ~n18371 ) | ( n17750 & n18370 ) | ( ~n18371 & n18370 ) ;
  assign n18374 = ( n17737 & ~n18372 ) | ( n17737 & n18373 ) | ( ~n18372 & n18373 ) ;
  assign n18363 = n17717 | n17902 ;
  assign n18364 = ( n17722 & ~n17717 ) | ( n17722 & n17730 ) | ( ~n17717 & n17730 ) ;
  assign n18366 = ( n17717 & n18363 ) | ( n17717 & n18364 ) | ( n18363 & n18364 ) ;
  assign n18365 = ( n17730 & ~n18364 ) | ( n17730 & n18363 ) | ( ~n18364 & n18363 ) ;
  assign n18367 = ( n17722 & ~n18366 ) | ( n17722 & n18365 ) | ( ~n18366 & n18365 ) ;
  assign n18348 = n17728 | n17902 ;
  assign n18349 = ( n17715 & ~n17728 ) | ( n17715 & n17724 ) | ( ~n17728 & n17724 ) ;
  assign n18351 = ( n17728 & n18348 ) | ( n17728 & n18349 ) | ( n18348 & n18349 ) ;
  assign n18350 = ( n17724 & ~n18349 ) | ( n17724 & n18348 ) | ( ~n18349 & n18348 ) ;
  assign n18352 = ( n17715 & ~n18351 ) | ( n17715 & n18350 ) | ( ~n18351 & n18350 ) ;
  assign n18341 = n17695 | n17902 ;
  assign n18342 = ( n17695 & ~n17708 ) | ( n17695 & n17700 ) | ( ~n17708 & n17700 ) ;
  assign n18343 = ( n17708 & n18341 ) | ( n17708 & n18342 ) | ( n18341 & n18342 ) ;
  assign n18344 = ( n17695 & ~n18342 ) | ( n17695 & n18341 ) | ( ~n18342 & n18341 ) ;
  assign n18345 = ( n17700 & ~n18343 ) | ( n17700 & n18344 ) | ( ~n18343 & n18344 ) ;
  assign n18326 = n17706 | n17902 ;
  assign n18327 = ( n17693 & ~n17702 ) | ( n17693 & n17706 ) | ( ~n17702 & n17706 ) ;
  assign n18328 = ( n17702 & n18326 ) | ( n17702 & n18327 ) | ( n18326 & n18327 ) ;
  assign n18329 = ( n17706 & ~n18327 ) | ( n17706 & n18326 ) | ( ~n18327 & n18326 ) ;
  assign n18330 = ( n17693 & ~n18328 ) | ( n17693 & n18329 ) | ( ~n18328 & n18329 ) ;
  assign n18319 = n17673 | n17902 ;
  assign n18320 = ( n17673 & n17678 ) | ( n17673 & n17686 ) | ( n17678 & n17686 ) ;
  assign n18321 = ( n18319 & ~n17686 ) | ( n18319 & n18320 ) | ( ~n17686 & n18320 ) ;
  assign n18322 = ( n17673 & ~n18320 ) | ( n17673 & n18319 ) | ( ~n18320 & n18319 ) ;
  assign n18323 = ( n17678 & ~n18321 ) | ( n17678 & n18322 ) | ( ~n18321 & n18322 ) ;
  assign n18304 = n17684 | n17902 ;
  assign n18305 = ( n17671 & n17680 ) | ( n17671 & n17684 ) | ( n17680 & n17684 ) ;
  assign n18306 = ( n18304 & ~n17680 ) | ( n18304 & n18305 ) | ( ~n17680 & n18305 ) ;
  assign n18307 = ( n17684 & ~n18305 ) | ( n17684 & n18304 ) | ( ~n18305 & n18304 ) ;
  assign n18308 = ( n17671 & ~n18306 ) | ( n17671 & n18307 ) | ( ~n18306 & n18307 ) ;
  assign n18298 = ( n17651 & ~n17656 ) | ( n17651 & n17664 ) | ( ~n17656 & n17664 ) ;
  assign n18297 = n17651 | n17902 ;
  assign n18300 = ( n17651 & ~n18298 ) | ( n17651 & n18297 ) | ( ~n18298 & n18297 ) ;
  assign n18299 = ( n18297 & ~n17664 ) | ( n18297 & n18298 ) | ( ~n17664 & n18298 ) ;
  assign n18301 = ( n17656 & ~n18300 ) | ( n17656 & n18299 ) | ( ~n18300 & n18299 ) ;
  assign n18283 = ( n17658 & ~n17649 ) | ( n17658 & n17662 ) | ( ~n17649 & n17662 ) ;
  assign n18282 = n17662 | n17902 ;
  assign n18285 = ( n17662 & ~n18283 ) | ( n17662 & n18282 ) | ( ~n18283 & n18282 ) ;
  assign n18284 = ( n18282 & ~n17658 ) | ( n18282 & n18283 ) | ( ~n17658 & n18283 ) ;
  assign n18286 = ( n17649 & ~n18285 ) | ( n17649 & n18284 ) | ( ~n18285 & n18284 ) ;
  assign n18275 = n17629 | n17902 ;
  assign n18276 = ( n17629 & n17634 ) | ( n17629 & n17642 ) | ( n17634 & n17642 ) ;
  assign n18277 = ( n18275 & ~n17642 ) | ( n18275 & n18276 ) | ( ~n17642 & n18276 ) ;
  assign n18278 = ( n17629 & ~n18276 ) | ( n17629 & n18275 ) | ( ~n18276 & n18275 ) ;
  assign n18279 = ( n17634 & ~n18277 ) | ( n17634 & n18278 ) | ( ~n18277 & n18278 ) ;
  assign n18261 = ( n17636 & ~n17627 ) | ( n17636 & n17640 ) | ( ~n17627 & n17640 ) ;
  assign n18260 = n17640 | n17902 ;
  assign n18263 = ( n17640 & ~n18261 ) | ( n17640 & n18260 ) | ( ~n18261 & n18260 ) ;
  assign n18262 = ( n18260 & ~n17636 ) | ( n18260 & n18261 ) | ( ~n17636 & n18261 ) ;
  assign n18264 = ( n17627 & ~n18263 ) | ( n17627 & n18262 ) | ( ~n18263 & n18262 ) ;
  assign n18253 = n17607 | n17902 ;
  assign n18254 = ( n17607 & n17612 ) | ( n17607 & n17620 ) | ( n17612 & n17620 ) ;
  assign n18255 = ( n18253 & ~n17620 ) | ( n18253 & n18254 ) | ( ~n17620 & n18254 ) ;
  assign n18256 = ( n17607 & ~n18254 ) | ( n17607 & n18253 ) | ( ~n18254 & n18253 ) ;
  assign n18257 = ( n17612 & ~n18255 ) | ( n17612 & n18256 ) | ( ~n18255 & n18256 ) ;
  assign n18238 = n17618 | n17902 ;
  assign n18239 = ( n17605 & ~n17618 ) | ( n17605 & n17614 ) | ( ~n17618 & n17614 ) ;
  assign n18241 = ( n17618 & n18238 ) | ( n17618 & n18239 ) | ( n18238 & n18239 ) ;
  assign n18240 = ( n17614 & ~n18239 ) | ( n17614 & n18238 ) | ( ~n18239 & n18238 ) ;
  assign n18242 = ( n17605 & ~n18241 ) | ( n17605 & n18240 ) | ( ~n18241 & n18240 ) ;
  assign n18231 = n17585 | n17902 ;
  assign n18232 = ( n17590 & ~n17585 ) | ( n17590 & n17598 ) | ( ~n17585 & n17598 ) ;
  assign n18234 = ( n17585 & n18231 ) | ( n17585 & n18232 ) | ( n18231 & n18232 ) ;
  assign n18233 = ( n17598 & ~n18232 ) | ( n17598 & n18231 ) | ( ~n18232 & n18231 ) ;
  assign n18235 = ( n17590 & ~n18234 ) | ( n17590 & n18233 ) | ( ~n18234 & n18233 ) ;
  assign n18216 = n17596 | n17902 ;
  assign n18217 = ( n17583 & ~n17592 ) | ( n17583 & n17596 ) | ( ~n17592 & n17596 ) ;
  assign n18218 = ( n17592 & n18216 ) | ( n17592 & n18217 ) | ( n18216 & n18217 ) ;
  assign n18219 = ( n17596 & ~n18217 ) | ( n17596 & n18216 ) | ( ~n18217 & n18216 ) ;
  assign n18220 = ( n17583 & ~n18218 ) | ( n17583 & n18219 ) | ( ~n18218 & n18219 ) ;
  assign n18209 = n17563 | n17902 ;
  assign n18210 = ( n17568 & ~n17563 ) | ( n17568 & n17576 ) | ( ~n17563 & n17576 ) ;
  assign n18212 = ( n17563 & n18209 ) | ( n17563 & n18210 ) | ( n18209 & n18210 ) ;
  assign n18211 = ( n17576 & ~n18210 ) | ( n17576 & n18209 ) | ( ~n18210 & n18209 ) ;
  assign n18213 = ( n17568 & ~n18212 ) | ( n17568 & n18211 ) | ( ~n18212 & n18211 ) ;
  assign n18194 = n17574 | n17902 ;
  assign n18195 = ( n17561 & ~n17570 ) | ( n17561 & n17574 ) | ( ~n17570 & n17574 ) ;
  assign n18196 = ( n17570 & n18194 ) | ( n17570 & n18195 ) | ( n18194 & n18195 ) ;
  assign n18197 = ( n17574 & ~n18195 ) | ( n17574 & n18194 ) | ( ~n18195 & n18194 ) ;
  assign n18198 = ( n17561 & ~n18196 ) | ( n17561 & n18197 ) | ( ~n18196 & n18197 ) ;
  assign n18187 = ( n17541 & ~n17902 ) | ( n17541 & 1'b0 ) | ( ~n17902 & 1'b0 ) ;
  assign n18188 = ( n17541 & n17546 ) | ( n17541 & n17554 ) | ( n17546 & n17554 ) ;
  assign n18189 = ( n18187 & ~n17554 ) | ( n18187 & n18188 ) | ( ~n17554 & n18188 ) ;
  assign n18190 = ( n17541 & ~n18188 ) | ( n17541 & n18187 ) | ( ~n18188 & n18187 ) ;
  assign n18191 = ( n17546 & ~n18189 ) | ( n17546 & n18190 ) | ( ~n18189 & n18190 ) ;
  assign n18172 = n17552 | n17902 ;
  assign n18173 = ( n17539 & ~n17548 ) | ( n17539 & n17552 ) | ( ~n17548 & n17552 ) ;
  assign n18174 = ( n17548 & n18172 ) | ( n17548 & n18173 ) | ( n18172 & n18173 ) ;
  assign n18175 = ( n17552 & ~n18173 ) | ( n17552 & n18172 ) | ( ~n18173 & n18172 ) ;
  assign n18176 = ( n17539 & ~n18174 ) | ( n17539 & n18175 ) | ( ~n18174 & n18175 ) ;
  assign n18165 = ( n17519 & ~n17902 ) | ( n17519 & 1'b0 ) | ( ~n17902 & 1'b0 ) ;
  assign n18166 = ( n17519 & n17524 ) | ( n17519 & n17532 ) | ( n17524 & n17532 ) ;
  assign n18167 = ( n18165 & ~n17532 ) | ( n18165 & n18166 ) | ( ~n17532 & n18166 ) ;
  assign n18168 = ( n17519 & ~n18166 ) | ( n17519 & n18165 ) | ( ~n18166 & n18165 ) ;
  assign n18169 = ( n17524 & ~n18167 ) | ( n17524 & n18168 ) | ( ~n18167 & n18168 ) ;
  assign n18150 = n17530 | n17902 ;
  assign n18151 = ( n17517 & ~n17526 ) | ( n17517 & n17530 ) | ( ~n17526 & n17530 ) ;
  assign n18152 = ( n17526 & n18150 ) | ( n17526 & n18151 ) | ( n18150 & n18151 ) ;
  assign n18153 = ( n17530 & ~n18151 ) | ( n17530 & n18150 ) | ( ~n18151 & n18150 ) ;
  assign n18154 = ( n17517 & ~n18152 ) | ( n17517 & n18153 ) | ( ~n18152 & n18153 ) ;
  assign n18143 = ( n17497 & ~n17902 ) | ( n17497 & 1'b0 ) | ( ~n17902 & 1'b0 ) ;
  assign n18144 = ( n17497 & n17502 ) | ( n17497 & n17510 ) | ( n17502 & n17510 ) ;
  assign n18145 = ( n18143 & ~n17510 ) | ( n18143 & n18144 ) | ( ~n17510 & n18144 ) ;
  assign n18146 = ( n17497 & ~n18144 ) | ( n17497 & n18143 ) | ( ~n18144 & n18143 ) ;
  assign n18147 = ( n17502 & ~n18145 ) | ( n17502 & n18146 ) | ( ~n18145 & n18146 ) ;
  assign n18129 = ( n17504 & ~n17495 ) | ( n17504 & n17508 ) | ( ~n17495 & n17508 ) ;
  assign n18128 = ( n17508 & ~n17902 ) | ( n17508 & 1'b0 ) | ( ~n17902 & 1'b0 ) ;
  assign n18131 = ( n17508 & ~n18129 ) | ( n17508 & n18128 ) | ( ~n18129 & n18128 ) ;
  assign n18130 = ( n18128 & ~n17504 ) | ( n18128 & n18129 ) | ( ~n17504 & n18129 ) ;
  assign n18132 = ( n17495 & ~n18131 ) | ( n17495 & n18130 ) | ( ~n18131 & n18130 ) ;
  assign n18121 = n17475 | n17902 ;
  assign n18122 = ( n17480 & ~n17475 ) | ( n17480 & n17488 ) | ( ~n17475 & n17488 ) ;
  assign n18124 = ( n17475 & n18121 ) | ( n17475 & n18122 ) | ( n18121 & n18122 ) ;
  assign n18123 = ( n17488 & ~n18122 ) | ( n17488 & n18121 ) | ( ~n18122 & n18121 ) ;
  assign n18125 = ( n17480 & ~n18124 ) | ( n17480 & n18123 ) | ( ~n18124 & n18123 ) ;
  assign n18106 = n17486 | n17902 ;
  assign n18107 = ( n17473 & ~n17482 ) | ( n17473 & n17486 ) | ( ~n17482 & n17486 ) ;
  assign n18108 = ( n17482 & n18106 ) | ( n17482 & n18107 ) | ( n18106 & n18107 ) ;
  assign n18109 = ( n17486 & ~n18107 ) | ( n17486 & n18106 ) | ( ~n18107 & n18106 ) ;
  assign n18110 = ( n17473 & ~n18108 ) | ( n17473 & n18109 ) | ( ~n18108 & n18109 ) ;
  assign n18099 = n17453 | n17902 ;
  assign n18100 = ( n17458 & ~n17453 ) | ( n17458 & n17466 ) | ( ~n17453 & n17466 ) ;
  assign n18102 = ( n17453 & n18099 ) | ( n17453 & n18100 ) | ( n18099 & n18100 ) ;
  assign n18101 = ( n17466 & ~n18100 ) | ( n17466 & n18099 ) | ( ~n18100 & n18099 ) ;
  assign n18103 = ( n17458 & ~n18102 ) | ( n17458 & n18101 ) | ( ~n18102 & n18101 ) ;
  assign n18084 = n17464 | n17902 ;
  assign n18085 = ( n17451 & ~n17460 ) | ( n17451 & n17464 ) | ( ~n17460 & n17464 ) ;
  assign n18086 = ( n17460 & n18084 ) | ( n17460 & n18085 ) | ( n18084 & n18085 ) ;
  assign n18087 = ( n17464 & ~n18085 ) | ( n17464 & n18084 ) | ( ~n18085 & n18084 ) ;
  assign n18088 = ( n17451 & ~n18086 ) | ( n17451 & n18087 ) | ( ~n18086 & n18087 ) ;
  assign n18077 = n17444 &  n17902 ;
  assign n18078 = ( n17436 & ~n17431 ) | ( n17436 & n17902 ) | ( ~n17431 & n17902 ) ;
  assign n18080 = ( n18077 & n17431 ) | ( n18077 & n18078 ) | ( n17431 & n18078 ) ;
  assign n18079 = ( n17902 & ~n18078 ) | ( n17902 & n18077 ) | ( ~n18078 & n18077 ) ;
  assign n18081 = ( n17436 & ~n18080 ) | ( n17436 & n18079 ) | ( ~n18080 & n18079 ) ;
  assign n18062 = n17442 | n17902 ;
  assign n18063 = ( n17429 & ~n17442 ) | ( n17429 & n17438 ) | ( ~n17442 & n17438 ) ;
  assign n18065 = ( n17442 & n18062 ) | ( n17442 & n18063 ) | ( n18062 & n18063 ) ;
  assign n18064 = ( n17438 & ~n18063 ) | ( n17438 & n18062 ) | ( ~n18063 & n18062 ) ;
  assign n18066 = ( n17429 & ~n18065 ) | ( n17429 & n18064 ) | ( ~n18065 & n18064 ) ;
  assign n18055 = n17409 | n17902 ;
  assign n18056 = ( n17409 & ~n17422 ) | ( n17409 & n17414 ) | ( ~n17422 & n17414 ) ;
  assign n18057 = ( n17422 & n18055 ) | ( n17422 & n18056 ) | ( n18055 & n18056 ) ;
  assign n18058 = ( n17409 & ~n18056 ) | ( n17409 & n18055 ) | ( ~n18056 & n18055 ) ;
  assign n18059 = ( n17414 & ~n18057 ) | ( n17414 & n18058 ) | ( ~n18057 & n18058 ) ;
  assign n18040 = n17420 | n17902 ;
  assign n18041 = ( n17407 & ~n17416 ) | ( n17407 & n17420 ) | ( ~n17416 & n17420 ) ;
  assign n18042 = ( n17416 & n18040 ) | ( n17416 & n18041 ) | ( n18040 & n18041 ) ;
  assign n18043 = ( n17420 & ~n18041 ) | ( n17420 & n18040 ) | ( ~n18041 & n18040 ) ;
  assign n18044 = ( n17407 & ~n18042 ) | ( n17407 & n18043 ) | ( ~n18042 & n18043 ) ;
  assign n18033 = n17387 | n17902 ;
  assign n18034 = ( n17392 & ~n17387 ) | ( n17392 & n17400 ) | ( ~n17387 & n17400 ) ;
  assign n18036 = ( n17387 & n18033 ) | ( n17387 & n18034 ) | ( n18033 & n18034 ) ;
  assign n18035 = ( n17400 & ~n18034 ) | ( n17400 & n18033 ) | ( ~n18034 & n18033 ) ;
  assign n18037 = ( n17392 & ~n18036 ) | ( n17392 & n18035 ) | ( ~n18036 & n18035 ) ;
  assign n18018 = n17398 | n17902 ;
  assign n18019 = ( n17385 & ~n17394 ) | ( n17385 & n17398 ) | ( ~n17394 & n17398 ) ;
  assign n18020 = ( n17394 & n18018 ) | ( n17394 & n18019 ) | ( n18018 & n18019 ) ;
  assign n18021 = ( n17398 & ~n18019 ) | ( n17398 & n18018 ) | ( ~n18019 & n18018 ) ;
  assign n18022 = ( n17385 & ~n18020 ) | ( n17385 & n18021 ) | ( ~n18020 & n18021 ) ;
  assign n18011 = n17378 &  n17902 ;
  assign n18012 = ( n17365 & n17370 ) | ( n17365 & n17902 ) | ( n17370 & n17902 ) ;
  assign n18014 = ( n18011 & ~n17365 ) | ( n18011 & n18012 ) | ( ~n17365 & n18012 ) ;
  assign n18013 = ( n17902 & ~n18012 ) | ( n17902 & n18011 ) | ( ~n18012 & n18011 ) ;
  assign n18015 = ( n17370 & ~n18014 ) | ( n17370 & n18013 ) | ( ~n18014 & n18013 ) ;
  assign n17996 = n17376 | n17902 ;
  assign n17997 = ( n17363 & ~n17376 ) | ( n17363 & n17372 ) | ( ~n17376 & n17372 ) ;
  assign n17999 = ( n17376 & n17996 ) | ( n17376 & n17997 ) | ( n17996 & n17997 ) ;
  assign n17998 = ( n17372 & ~n17997 ) | ( n17372 & n17996 ) | ( ~n17997 & n17996 ) ;
  assign n18000 = ( n17363 & ~n17999 ) | ( n17363 & n17998 ) | ( ~n17999 & n17998 ) ;
  assign n17989 = n17343 | n17902 ;
  assign n17990 = ( n17343 & ~n17356 ) | ( n17343 & n17348 ) | ( ~n17356 & n17348 ) ;
  assign n17991 = ( n17356 & n17989 ) | ( n17356 & n17990 ) | ( n17989 & n17990 ) ;
  assign n17992 = ( n17343 & ~n17990 ) | ( n17343 & n17989 ) | ( ~n17990 & n17989 ) ;
  assign n17993 = ( n17348 & ~n17991 ) | ( n17348 & n17992 ) | ( ~n17991 & n17992 ) ;
  assign n17974 = n17354 | n17902 ;
  assign n17975 = ( n17341 & ~n17350 ) | ( n17341 & n17354 ) | ( ~n17350 & n17354 ) ;
  assign n17976 = ( n17350 & n17974 ) | ( n17350 & n17975 ) | ( n17974 & n17975 ) ;
  assign n17977 = ( n17354 & ~n17975 ) | ( n17354 & n17974 ) | ( ~n17975 & n17974 ) ;
  assign n17978 = ( n17341 & ~n17976 ) | ( n17341 & n17977 ) | ( ~n17976 & n17977 ) ;
  assign n17967 = n17321 | n17902 ;
  assign n17968 = ( n17326 & ~n17321 ) | ( n17326 & n17334 ) | ( ~n17321 & n17334 ) ;
  assign n17970 = ( n17321 & n17967 ) | ( n17321 & n17968 ) | ( n17967 & n17968 ) ;
  assign n17969 = ( n17334 & ~n17968 ) | ( n17334 & n17967 ) | ( ~n17968 & n17967 ) ;
  assign n17971 = ( n17326 & ~n17970 ) | ( n17326 & n17969 ) | ( ~n17970 & n17969 ) ;
  assign n17952 = n17332 | n17902 ;
  assign n17953 = ( n17319 & ~n17328 ) | ( n17319 & n17332 ) | ( ~n17328 & n17332 ) ;
  assign n17954 = ( n17328 & n17952 ) | ( n17328 & n17953 ) | ( n17952 & n17953 ) ;
  assign n17955 = ( n17332 & ~n17953 ) | ( n17332 & n17952 ) | ( ~n17953 & n17952 ) ;
  assign n17956 = ( n17319 & ~n17954 ) | ( n17319 & n17955 ) | ( ~n17954 & n17955 ) ;
  assign n17945 = ( n17295 & ~n17297 ) | ( n17295 & 1'b0 ) | ( ~n17297 & 1'b0 ) ;
  assign n17946 = ( n17297 & ~n17945 ) | ( n17297 & n17307 ) | ( ~n17945 & n17307 ) ;
  assign n17948 = ( n17902 & n17945 ) | ( n17902 & n17946 ) | ( n17945 & n17946 ) ;
  assign n17947 = ( n17297 & ~n17946 ) | ( n17297 & n17902 ) | ( ~n17946 & n17902 ) ;
  assign n17949 = ( n17307 & ~n17948 ) | ( n17307 & n17947 ) | ( ~n17948 & n17947 ) ;
  assign n17929 = ~x18 & n17279 ;
  assign n17930 = ( x19 & ~n17929 ) | ( x19 & 1'b0 ) | ( ~n17929 & 1'b0 ) ;
  assign n17931 = n17298 | n17930 ;
  assign n17926 = ( n17279 & ~x18 ) | ( n17279 & n17290 ) | ( ~x18 & n17290 ) ;
  assign n17927 = x18 &  n17926 ;
  assign n17928 = ( n17285 & ~n17927 ) | ( n17285 & n17290 ) | ( ~n17927 & n17290 ) ;
  assign n17932 = ( n17902 & ~n17931 ) | ( n17902 & n17928 ) | ( ~n17931 & n17928 ) ;
  assign n17934 = ( n17902 & ~n17932 ) | ( n17902 & 1'b0 ) | ( ~n17932 & 1'b0 ) ;
  assign n17933 = ~n17928 & n17932 ;
  assign n17935 = ( n17931 & ~n17934 ) | ( n17931 & n17933 ) | ( ~n17934 & n17933 ) ;
  assign n17915 = ( n17279 & ~n17899 ) | ( n17279 & 1'b0 ) | ( ~n17899 & 1'b0 ) ;
  assign n17916 = ( n17890 & ~n17894 ) | ( n17890 & n17915 ) | ( ~n17894 & n17915 ) ;
  assign n17917 = ~n17890 & n17916 ;
  assign n17918 = n17882 &  n17917 ;
  assign n17914 = ~n17282 & n17902 ;
  assign n17919 = ( n17914 & ~n17918 ) | ( n17914 & 1'b0 ) | ( ~n17918 & 1'b0 ) ;
  assign n17920 = ( x18 & n17918 ) | ( x18 & n17919 ) | ( n17918 & n17919 ) ;
  assign n17921 = x18 | n17918 ;
  assign n17922 = n17914 | n17921 ;
  assign n17923 = ~n17920 & n17922 ;
  assign n17905 = ( x16 & ~n17902 ) | ( x16 & x17 ) | ( ~n17902 & x17 ) ;
  assign n17911 = ( x16 & ~x17 ) | ( x16 & 1'b0 ) | ( ~x17 & 1'b0 ) ;
  assign n17280 = x14 | x15 ;
  assign n17906 = ~x16 & n17280 ;
  assign n17907 = ( x16 & ~n17277 ) | ( x16 & n17906 ) | ( ~n17277 & n17906 ) ;
  assign n17908 = ( n17259 & ~n17907 ) | ( n17259 & n17267 ) | ( ~n17907 & n17267 ) ;
  assign n17909 = ( n17259 & ~n17908 ) | ( n17259 & 1'b0 ) | ( ~n17908 & 1'b0 ) ;
  assign n17910 = ( n17902 & ~x17 ) | ( n17902 & n17909 ) | ( ~x17 & n17909 ) ;
  assign n17912 = ( n17905 & ~n17911 ) | ( n17905 & n17910 ) | ( ~n17911 & n17910 ) ;
  assign n17281 = x16 | n17280 ;
  assign n17903 = x16 &  n17902 ;
  assign n17904 = ( n17279 & ~n17281 ) | ( n17279 & n17903 ) | ( ~n17281 & n17903 ) ;
  assign n17936 = n16671 | n17904 ;
  assign n17937 = ( n17912 & ~n17936 ) | ( n17912 & 1'b0 ) | ( ~n17936 & 1'b0 ) ;
  assign n17938 = n17923 | n17937 ;
  assign n17939 = n17904 &  n17912 ;
  assign n17940 = ( n16671 & ~n17912 ) | ( n16671 & n17939 ) | ( ~n17912 & n17939 ) ;
  assign n17941 = n16070 | n17940 ;
  assign n17942 = ( n17938 & ~n17941 ) | ( n17938 & 1'b0 ) | ( ~n17941 & 1'b0 ) ;
  assign n17943 = n17935 | n17942 ;
  assign n17913 = ~n17904 & n17912 ;
  assign n17924 = ( n17913 & ~n16671 ) | ( n17913 & n17923 ) | ( ~n16671 & n17923 ) ;
  assign n17925 = ( n16070 & ~n17924 ) | ( n16070 & 1'b0 ) | ( ~n17924 & 1'b0 ) ;
  assign n17957 = n15484 | n17925 ;
  assign n17958 = ( n17943 & ~n17957 ) | ( n17943 & 1'b0 ) | ( ~n17957 & 1'b0 ) ;
  assign n17959 = n17949 | n17958 ;
  assign n17960 = ( n17938 & ~n17940 ) | ( n17938 & 1'b0 ) | ( ~n17940 & 1'b0 ) ;
  assign n17961 = ( n17935 & ~n16070 ) | ( n17935 & n17960 ) | ( ~n16070 & n17960 ) ;
  assign n17962 = ( n15484 & ~n17961 ) | ( n15484 & 1'b0 ) | ( ~n17961 & 1'b0 ) ;
  assign n17963 = n14905 | n17962 ;
  assign n17964 = ( n17959 & ~n17963 ) | ( n17959 & 1'b0 ) | ( ~n17963 & 1'b0 ) ;
  assign n17965 = n17956 | n17964 ;
  assign n17944 = ~n17925 & n17943 ;
  assign n17950 = ( n17944 & ~n15484 ) | ( n17944 & n17949 ) | ( ~n15484 & n17949 ) ;
  assign n17951 = ( n14905 & ~n17950 ) | ( n14905 & 1'b0 ) | ( ~n17950 & 1'b0 ) ;
  assign n17979 = n14341 | n17951 ;
  assign n17980 = ( n17965 & ~n17979 ) | ( n17965 & 1'b0 ) | ( ~n17979 & 1'b0 ) ;
  assign n17981 = n17971 | n17980 ;
  assign n17982 = ( n17959 & ~n17962 ) | ( n17959 & 1'b0 ) | ( ~n17962 & 1'b0 ) ;
  assign n17983 = ( n17956 & ~n14905 ) | ( n17956 & n17982 ) | ( ~n14905 & n17982 ) ;
  assign n17984 = ( n14341 & ~n17983 ) | ( n14341 & 1'b0 ) | ( ~n17983 & 1'b0 ) ;
  assign n17985 = n13784 | n17984 ;
  assign n17986 = ( n17981 & ~n17985 ) | ( n17981 & 1'b0 ) | ( ~n17985 & 1'b0 ) ;
  assign n17987 = n17978 | n17986 ;
  assign n17966 = ~n17951 & n17965 ;
  assign n17972 = ( n17966 & ~n14341 ) | ( n17966 & n17971 ) | ( ~n14341 & n17971 ) ;
  assign n17973 = ( n13784 & ~n17972 ) | ( n13784 & 1'b0 ) | ( ~n17972 & 1'b0 ) ;
  assign n18001 = n13242 | n17973 ;
  assign n18002 = ( n17987 & ~n18001 ) | ( n17987 & 1'b0 ) | ( ~n18001 & 1'b0 ) ;
  assign n18003 = n17993 | n18002 ;
  assign n18004 = ( n17981 & ~n17984 ) | ( n17981 & 1'b0 ) | ( ~n17984 & 1'b0 ) ;
  assign n18005 = ( n17978 & ~n13784 ) | ( n17978 & n18004 ) | ( ~n13784 & n18004 ) ;
  assign n18006 = ( n13242 & ~n18005 ) | ( n13242 & 1'b0 ) | ( ~n18005 & 1'b0 ) ;
  assign n18007 = n12707 | n18006 ;
  assign n18008 = ( n18003 & ~n18007 ) | ( n18003 & 1'b0 ) | ( ~n18007 & 1'b0 ) ;
  assign n18009 = n18000 | n18008 ;
  assign n17988 = ~n17973 & n17987 ;
  assign n17994 = ( n17988 & ~n13242 ) | ( n17988 & n17993 ) | ( ~n13242 & n17993 ) ;
  assign n17995 = ( n12707 & ~n17994 ) | ( n12707 & 1'b0 ) | ( ~n17994 & 1'b0 ) ;
  assign n18023 = n12187 | n17995 ;
  assign n18024 = ( n18009 & ~n18023 ) | ( n18009 & 1'b0 ) | ( ~n18023 & 1'b0 ) ;
  assign n18025 = n18015 | n18024 ;
  assign n18026 = ( n18003 & ~n18006 ) | ( n18003 & 1'b0 ) | ( ~n18006 & 1'b0 ) ;
  assign n18027 = ( n18000 & ~n12707 ) | ( n18000 & n18026 ) | ( ~n12707 & n18026 ) ;
  assign n18028 = ( n12187 & ~n18027 ) | ( n12187 & 1'b0 ) | ( ~n18027 & 1'b0 ) ;
  assign n18029 = n11674 | n18028 ;
  assign n18030 = ( n18025 & ~n18029 ) | ( n18025 & 1'b0 ) | ( ~n18029 & 1'b0 ) ;
  assign n18031 = n18022 | n18030 ;
  assign n18010 = ~n17995 & n18009 ;
  assign n18016 = ( n18010 & ~n12187 ) | ( n18010 & n18015 ) | ( ~n12187 & n18015 ) ;
  assign n18017 = ( n11674 & ~n18016 ) | ( n11674 & 1'b0 ) | ( ~n18016 & 1'b0 ) ;
  assign n18045 = n11176 | n18017 ;
  assign n18046 = ( n18031 & ~n18045 ) | ( n18031 & 1'b0 ) | ( ~n18045 & 1'b0 ) ;
  assign n18047 = n18037 | n18046 ;
  assign n18048 = ( n18025 & ~n18028 ) | ( n18025 & 1'b0 ) | ( ~n18028 & 1'b0 ) ;
  assign n18049 = ( n18022 & ~n11674 ) | ( n18022 & n18048 ) | ( ~n11674 & n18048 ) ;
  assign n18050 = ( n11176 & ~n18049 ) | ( n11176 & 1'b0 ) | ( ~n18049 & 1'b0 ) ;
  assign n18051 = n10685 | n18050 ;
  assign n18052 = ( n18047 & ~n18051 ) | ( n18047 & 1'b0 ) | ( ~n18051 & 1'b0 ) ;
  assign n18053 = n18044 | n18052 ;
  assign n18032 = ~n18017 & n18031 ;
  assign n18038 = ( n18032 & ~n11176 ) | ( n18032 & n18037 ) | ( ~n11176 & n18037 ) ;
  assign n18039 = ( n10685 & ~n18038 ) | ( n10685 & 1'b0 ) | ( ~n18038 & 1'b0 ) ;
  assign n18067 = n10209 | n18039 ;
  assign n18068 = ( n18053 & ~n18067 ) | ( n18053 & 1'b0 ) | ( ~n18067 & 1'b0 ) ;
  assign n18069 = n18059 | n18068 ;
  assign n18070 = ( n18047 & ~n18050 ) | ( n18047 & 1'b0 ) | ( ~n18050 & 1'b0 ) ;
  assign n18071 = ( n18044 & ~n10685 ) | ( n18044 & n18070 ) | ( ~n10685 & n18070 ) ;
  assign n18072 = ( n10209 & ~n18071 ) | ( n10209 & 1'b0 ) | ( ~n18071 & 1'b0 ) ;
  assign n18073 = ( n9740 & ~n18072 ) | ( n9740 & 1'b0 ) | ( ~n18072 & 1'b0 ) ;
  assign n18074 = n18069 &  n18073 ;
  assign n18075 = n18066 | n18074 ;
  assign n18054 = ~n18039 & n18053 ;
  assign n18060 = ( n18054 & ~n10209 ) | ( n18054 & n18059 ) | ( ~n10209 & n18059 ) ;
  assign n18061 = n9740 | n18060 ;
  assign n18089 = ~n9286 & n18061 ;
  assign n18090 = n18075 &  n18089 ;
  assign n18091 = n18081 | n18090 ;
  assign n18092 = ( n18069 & ~n18072 ) | ( n18069 & 1'b0 ) | ( ~n18072 & 1'b0 ) ;
  assign n18093 = ( n9740 & n18066 ) | ( n9740 & n18092 ) | ( n18066 & n18092 ) ;
  assign n18094 = ( n9286 & ~n18093 ) | ( n9286 & 1'b0 ) | ( ~n18093 & 1'b0 ) ;
  assign n18095 = n8839 | n18094 ;
  assign n18096 = ( n18091 & ~n18095 ) | ( n18091 & 1'b0 ) | ( ~n18095 & 1'b0 ) ;
  assign n18097 = n18088 | n18096 ;
  assign n18076 = n18061 &  n18075 ;
  assign n18082 = ( n18076 & ~n9286 ) | ( n18076 & n18081 ) | ( ~n9286 & n18081 ) ;
  assign n18083 = ( n8839 & ~n18082 ) | ( n8839 & 1'b0 ) | ( ~n18082 & 1'b0 ) ;
  assign n18111 = n8407 | n18083 ;
  assign n18112 = ( n18097 & ~n18111 ) | ( n18097 & 1'b0 ) | ( ~n18111 & 1'b0 ) ;
  assign n18113 = n18103 | n18112 ;
  assign n18114 = ( n18091 & ~n18094 ) | ( n18091 & 1'b0 ) | ( ~n18094 & 1'b0 ) ;
  assign n18115 = ( n18088 & ~n8839 ) | ( n18088 & n18114 ) | ( ~n8839 & n18114 ) ;
  assign n18116 = ( n8407 & ~n18115 ) | ( n8407 & 1'b0 ) | ( ~n18115 & 1'b0 ) ;
  assign n18117 = n7982 | n18116 ;
  assign n18118 = ( n18113 & ~n18117 ) | ( n18113 & 1'b0 ) | ( ~n18117 & 1'b0 ) ;
  assign n18119 = n18110 | n18118 ;
  assign n18098 = ~n18083 & n18097 ;
  assign n18104 = ( n18098 & ~n8407 ) | ( n18098 & n18103 ) | ( ~n8407 & n18103 ) ;
  assign n18105 = ( n7982 & ~n18104 ) | ( n7982 & 1'b0 ) | ( ~n18104 & 1'b0 ) ;
  assign n18133 = ( n7572 & ~n18105 ) | ( n7572 & 1'b0 ) | ( ~n18105 & 1'b0 ) ;
  assign n18134 = n18119 &  n18133 ;
  assign n18135 = n18125 | n18134 ;
  assign n18136 = ( n18113 & ~n18116 ) | ( n18113 & 1'b0 ) | ( ~n18116 & 1'b0 ) ;
  assign n18137 = ( n18110 & ~n7982 ) | ( n18110 & n18136 ) | ( ~n7982 & n18136 ) ;
  assign n18138 = n7572 | n18137 ;
  assign n18139 = n7169 &  n18138 ;
  assign n18140 = n18135 &  n18139 ;
  assign n18141 = n18132 | n18140 ;
  assign n18120 = ~n18105 & n18119 ;
  assign n18126 = ( n7572 & n18120 ) | ( n7572 & n18125 ) | ( n18120 & n18125 ) ;
  assign n18127 = n7169 | n18126 ;
  assign n18155 = ~n6781 & n18127 ;
  assign n18156 = n18141 &  n18155 ;
  assign n18157 = n18147 | n18156 ;
  assign n18158 = n18135 &  n18138 ;
  assign n18159 = ( n7169 & n18132 ) | ( n7169 & n18158 ) | ( n18132 & n18158 ) ;
  assign n18160 = ( n6781 & ~n18159 ) | ( n6781 & 1'b0 ) | ( ~n18159 & 1'b0 ) ;
  assign n18161 = ( n6399 & ~n18160 ) | ( n6399 & 1'b0 ) | ( ~n18160 & 1'b0 ) ;
  assign n18162 = n18157 &  n18161 ;
  assign n18163 = n18154 | n18162 ;
  assign n18142 = n18127 &  n18141 ;
  assign n18148 = ( n18142 & ~n6781 ) | ( n18142 & n18147 ) | ( ~n6781 & n18147 ) ;
  assign n18149 = n6399 | n18148 ;
  assign n18177 = ~n6032 & n18149 ;
  assign n18178 = n18163 &  n18177 ;
  assign n18179 = n18169 | n18178 ;
  assign n18180 = ( n18157 & ~n18160 ) | ( n18157 & 1'b0 ) | ( ~n18160 & 1'b0 ) ;
  assign n18181 = ( n6399 & n18154 ) | ( n6399 & n18180 ) | ( n18154 & n18180 ) ;
  assign n18182 = ( n6032 & ~n18181 ) | ( n6032 & 1'b0 ) | ( ~n18181 & 1'b0 ) ;
  assign n18183 = ( n5672 & ~n18182 ) | ( n5672 & 1'b0 ) | ( ~n18182 & 1'b0 ) ;
  assign n18184 = n18179 &  n18183 ;
  assign n18185 = n18176 | n18184 ;
  assign n18164 = n18149 &  n18163 ;
  assign n18170 = ( n18164 & ~n6032 ) | ( n18164 & n18169 ) | ( ~n6032 & n18169 ) ;
  assign n18171 = n5672 | n18170 ;
  assign n18199 = ~n5327 & n18171 ;
  assign n18200 = n18185 &  n18199 ;
  assign n18201 = n18191 | n18200 ;
  assign n18202 = ( n18179 & ~n18182 ) | ( n18179 & 1'b0 ) | ( ~n18182 & 1'b0 ) ;
  assign n18203 = ( n5672 & n18176 ) | ( n5672 & n18202 ) | ( n18176 & n18202 ) ;
  assign n18204 = ( n5327 & ~n18203 ) | ( n5327 & 1'b0 ) | ( ~n18203 & 1'b0 ) ;
  assign n18205 = n4990 | n18204 ;
  assign n18206 = ( n18201 & ~n18205 ) | ( n18201 & 1'b0 ) | ( ~n18205 & 1'b0 ) ;
  assign n18207 = n18198 | n18206 ;
  assign n18186 = n18171 &  n18185 ;
  assign n18192 = ( n18186 & ~n5327 ) | ( n18186 & n18191 ) | ( ~n5327 & n18191 ) ;
  assign n18193 = ( n4990 & ~n18192 ) | ( n4990 & 1'b0 ) | ( ~n18192 & 1'b0 ) ;
  assign n18221 = n4668 | n18193 ;
  assign n18222 = ( n18207 & ~n18221 ) | ( n18207 & 1'b0 ) | ( ~n18221 & 1'b0 ) ;
  assign n18223 = n18213 | n18222 ;
  assign n18224 = ( n18201 & ~n18204 ) | ( n18201 & 1'b0 ) | ( ~n18204 & 1'b0 ) ;
  assign n18225 = ( n18198 & ~n4990 ) | ( n18198 & n18224 ) | ( ~n4990 & n18224 ) ;
  assign n18226 = ( n4668 & ~n18225 ) | ( n4668 & 1'b0 ) | ( ~n18225 & 1'b0 ) ;
  assign n18227 = n4353 | n18226 ;
  assign n18228 = ( n18223 & ~n18227 ) | ( n18223 & 1'b0 ) | ( ~n18227 & 1'b0 ) ;
  assign n18229 = n18220 | n18228 ;
  assign n18208 = ~n18193 & n18207 ;
  assign n18214 = ( n18208 & ~n4668 ) | ( n18208 & n18213 ) | ( ~n4668 & n18213 ) ;
  assign n18215 = ( n4353 & ~n18214 ) | ( n4353 & 1'b0 ) | ( ~n18214 & 1'b0 ) ;
  assign n18243 = n4053 | n18215 ;
  assign n18244 = ( n18229 & ~n18243 ) | ( n18229 & 1'b0 ) | ( ~n18243 & 1'b0 ) ;
  assign n18245 = n18235 | n18244 ;
  assign n18246 = ( n18223 & ~n18226 ) | ( n18223 & 1'b0 ) | ( ~n18226 & 1'b0 ) ;
  assign n18247 = ( n18220 & ~n4353 ) | ( n18220 & n18246 ) | ( ~n4353 & n18246 ) ;
  assign n18248 = ( n4053 & ~n18247 ) | ( n4053 & 1'b0 ) | ( ~n18247 & 1'b0 ) ;
  assign n18249 = n3760 | n18248 ;
  assign n18250 = ( n18245 & ~n18249 ) | ( n18245 & 1'b0 ) | ( ~n18249 & 1'b0 ) ;
  assign n18251 = ( n18242 & ~n18250 ) | ( n18242 & 1'b0 ) | ( ~n18250 & 1'b0 ) ;
  assign n18230 = ~n18215 & n18229 ;
  assign n18236 = ( n18230 & ~n4053 ) | ( n18230 & n18235 ) | ( ~n4053 & n18235 ) ;
  assign n18237 = ( n3760 & ~n18236 ) | ( n3760 & 1'b0 ) | ( ~n18236 & 1'b0 ) ;
  assign n18265 = n3482 | n18237 ;
  assign n18266 = n18251 | n18265 ;
  assign n18267 = n18257 &  n18266 ;
  assign n18268 = ( n18245 & ~n18248 ) | ( n18245 & 1'b0 ) | ( ~n18248 & 1'b0 ) ;
  assign n18269 = ( n3760 & ~n18268 ) | ( n3760 & n18242 ) | ( ~n18268 & n18242 ) ;
  assign n18270 = n3482 &  n18269 ;
  assign n18271 = n3211 | n18270 ;
  assign n18272 = n18267 | n18271 ;
  assign n18273 = n18264 &  n18272 ;
  assign n18252 = n18237 | n18251 ;
  assign n18258 = ( n3482 & n18252 ) | ( n3482 & n18257 ) | ( n18252 & n18257 ) ;
  assign n18259 = n3211 &  n18258 ;
  assign n18287 = n2955 | n18259 ;
  assign n18288 = n18273 | n18287 ;
  assign n18289 = n18279 &  n18288 ;
  assign n18290 = n18267 | n18270 ;
  assign n18291 = ( n3211 & n18264 ) | ( n3211 & n18290 ) | ( n18264 & n18290 ) ;
  assign n18292 = n2955 &  n18291 ;
  assign n18293 = n2706 | n18292 ;
  assign n18294 = n18289 | n18293 ;
  assign n18295 = n18286 &  n18294 ;
  assign n18274 = n18259 | n18273 ;
  assign n18280 = ( n2955 & n18274 ) | ( n2955 & n18279 ) | ( n18274 & n18279 ) ;
  assign n18281 = n2706 &  n18280 ;
  assign n18309 = n2472 | n18281 ;
  assign n18310 = n18295 | n18309 ;
  assign n18311 = ~n18301 & n18310 ;
  assign n18312 = n18289 | n18292 ;
  assign n18313 = ( n2706 & n18286 ) | ( n2706 & n18312 ) | ( n18286 & n18312 ) ;
  assign n18314 = n2472 &  n18313 ;
  assign n18315 = n2245 | n18314 ;
  assign n18316 = n18311 | n18315 ;
  assign n18317 = ~n18308 & n18316 ;
  assign n18296 = n18281 | n18295 ;
  assign n18302 = ( n2472 & ~n18301 ) | ( n2472 & n18296 ) | ( ~n18301 & n18296 ) ;
  assign n18303 = n2245 &  n18302 ;
  assign n18331 = ( n2033 & ~n18303 ) | ( n2033 & 1'b0 ) | ( ~n18303 & 1'b0 ) ;
  assign n18332 = ~n18317 & n18331 ;
  assign n18333 = ( n18323 & ~n18332 ) | ( n18323 & 1'b0 ) | ( ~n18332 & 1'b0 ) ;
  assign n18334 = n18311 | n18314 ;
  assign n18335 = ( n2245 & ~n18308 ) | ( n2245 & n18334 ) | ( ~n18308 & n18334 ) ;
  assign n18336 = ~n2033 & n18335 ;
  assign n18337 = n1827 | n18336 ;
  assign n18338 = n18333 | n18337 ;
  assign n18339 = ~n18330 & n18338 ;
  assign n18318 = n18303 | n18317 ;
  assign n18324 = ( n18318 & ~n2033 ) | ( n18318 & n18323 ) | ( ~n2033 & n18323 ) ;
  assign n18325 = n1827 &  n18324 ;
  assign n18353 = ( n1636 & ~n18325 ) | ( n1636 & 1'b0 ) | ( ~n18325 & 1'b0 ) ;
  assign n18354 = ~n18339 & n18353 ;
  assign n18355 = ( n18345 & ~n18354 ) | ( n18345 & 1'b0 ) | ( ~n18354 & 1'b0 ) ;
  assign n18356 = n18333 | n18336 ;
  assign n18357 = ( n1827 & ~n18330 ) | ( n1827 & n18356 ) | ( ~n18330 & n18356 ) ;
  assign n18358 = ~n1636 & n18357 ;
  assign n18359 = ( n1452 & ~n18358 ) | ( n1452 & 1'b0 ) | ( ~n18358 & 1'b0 ) ;
  assign n18360 = ~n18355 & n18359 ;
  assign n18361 = ( n18352 & ~n18360 ) | ( n18352 & 1'b0 ) | ( ~n18360 & 1'b0 ) ;
  assign n18340 = n18325 | n18339 ;
  assign n18346 = ( n18340 & ~n1636 ) | ( n18340 & n18345 ) | ( ~n1636 & n18345 ) ;
  assign n18347 = ~n1452 & n18346 ;
  assign n18375 = n1283 | n18347 ;
  assign n18376 = n18361 | n18375 ;
  assign n18377 = ~n18367 & n18376 ;
  assign n18378 = n18355 | n18358 ;
  assign n18379 = ( n18352 & ~n1452 ) | ( n18352 & n18378 ) | ( ~n1452 & n18378 ) ;
  assign n18380 = n1283 &  n18379 ;
  assign n18381 = ( n1122 & ~n18380 ) | ( n1122 & 1'b0 ) | ( ~n18380 & 1'b0 ) ;
  assign n18382 = ~n18377 & n18381 ;
  assign n18383 = n18374 | n18382 ;
  assign n18362 = n18347 | n18361 ;
  assign n18368 = ( n1283 & ~n18367 ) | ( n1283 & n18362 ) | ( ~n18367 & n18362 ) ;
  assign n18369 = ~n1122 & n18368 ;
  assign n18397 = ( n976 & ~n18369 ) | ( n976 & 1'b0 ) | ( ~n18369 & 1'b0 ) ;
  assign n18398 = n18383 &  n18397 ;
  assign n18399 = n18389 | n18398 ;
  assign n18400 = n18377 | n18380 ;
  assign n18401 = ( n1122 & ~n18400 ) | ( n1122 & n18374 ) | ( ~n18400 & n18374 ) ;
  assign n18402 = n976 | n18401 ;
  assign n18403 = ~n837 & n18402 ;
  assign n18404 = n18399 &  n18403 ;
  assign n18405 = n18396 | n18404 ;
  assign n18384 = ~n18369 & n18383 ;
  assign n18390 = ( n976 & n18384 ) | ( n976 & n18389 ) | ( n18384 & n18389 ) ;
  assign n18391 = ( n837 & ~n18390 ) | ( n837 & 1'b0 ) | ( ~n18390 & 1'b0 ) ;
  assign n18419 = n713 | n18391 ;
  assign n18420 = ( n18405 & ~n18419 ) | ( n18405 & 1'b0 ) | ( ~n18419 & 1'b0 ) ;
  assign n18421 = n18411 | n18420 ;
  assign n18422 = n18399 &  n18402 ;
  assign n18423 = ( n18396 & ~n837 ) | ( n18396 & n18422 ) | ( ~n837 & n18422 ) ;
  assign n18424 = ( n713 & ~n18423 ) | ( n713 & 1'b0 ) | ( ~n18423 & 1'b0 ) ;
  assign n18439 = ( n18421 & ~n18424 ) | ( n18421 & 1'b0 ) | ( ~n18424 & 1'b0 ) ;
  assign n18414 = n17794 | n17902 ;
  assign n18415 = ( n17781 & ~n17794 ) | ( n17781 & n17790 ) | ( ~n17794 & n17790 ) ;
  assign n18417 = ( n17794 & n18414 ) | ( n17794 & n18415 ) | ( n18414 & n18415 ) ;
  assign n18416 = ( n17790 & ~n18415 ) | ( n17790 & n18414 ) | ( ~n18415 & n18414 ) ;
  assign n18418 = ( n17781 & ~n18417 ) | ( n17781 & n18416 ) | ( ~n18417 & n18416 ) ;
  assign n18440 = ( n595 & ~n18439 ) | ( n595 & n18418 ) | ( ~n18439 & n18418 ) ;
  assign n18441 = n492 &  n18440 ;
  assign n18494 = n17848 | n17902 ;
  assign n18495 = ( n17848 & ~n17861 ) | ( n17848 & n17853 ) | ( ~n17861 & n17853 ) ;
  assign n18496 = ( n17861 & n18494 ) | ( n17861 & n18495 ) | ( n18494 & n18495 ) ;
  assign n18497 = ( n17848 & ~n18495 ) | ( n17848 & n18494 ) | ( ~n18495 & n18494 ) ;
  assign n18498 = ( n17853 & ~n18496 ) | ( n17853 & n18497 ) | ( ~n18496 & n18497 ) ;
  assign n18406 = ~n18391 & n18405 ;
  assign n18412 = ( n18406 & ~n713 ) | ( n18406 & n18411 ) | ( ~n713 & n18411 ) ;
  assign n18413 = ( n595 & ~n18412 ) | ( n595 & 1'b0 ) | ( ~n18412 & 1'b0 ) ;
  assign n18425 = n595 | n18424 ;
  assign n18426 = ( n18421 & ~n18425 ) | ( n18421 & 1'b0 ) | ( ~n18425 & 1'b0 ) ;
  assign n18427 = ( n18418 & ~n18426 ) | ( n18418 & 1'b0 ) | ( ~n18426 & 1'b0 ) ;
  assign n18428 = n18413 | n18427 ;
  assign n18434 = ( n492 & ~n18433 ) | ( n492 & n18428 ) | ( ~n18433 & n18428 ) ;
  assign n18435 = n396 &  n18434 ;
  assign n18436 = n492 | n18413 ;
  assign n18437 = n18427 | n18436 ;
  assign n18438 = ~n18433 & n18437 ;
  assign n18442 = n396 | n18441 ;
  assign n18443 = n18438 | n18442 ;
  assign n18444 = ( n17802 & n17811 ) | ( n17802 & n17815 ) | ( n17811 & n17815 ) ;
  assign n18445 = ( n17902 & ~n17811 ) | ( n17902 & n18444 ) | ( ~n17811 & n18444 ) ;
  assign n18446 = ( n17815 & ~n18444 ) | ( n17815 & n17902 ) | ( ~n18444 & n17902 ) ;
  assign n18447 = ( n17802 & ~n18445 ) | ( n17802 & n18446 ) | ( ~n18445 & n18446 ) ;
  assign n18448 = ( n18443 & ~n18447 ) | ( n18443 & 1'b0 ) | ( ~n18447 & 1'b0 ) ;
  assign n18449 = n18435 | n18448 ;
  assign n18450 = ~n17817 & n17902 ;
  assign n18451 = ( n17804 & n17809 ) | ( n17804 & n17902 ) | ( n17809 & n17902 ) ;
  assign n18453 = ( n18450 & ~n17804 ) | ( n18450 & n18451 ) | ( ~n17804 & n18451 ) ;
  assign n18452 = ( n17902 & ~n18451 ) | ( n17902 & n18450 ) | ( ~n18451 & n18450 ) ;
  assign n18454 = ( n17809 & ~n18453 ) | ( n17809 & n18452 ) | ( ~n18453 & n18452 ) ;
  assign n18455 = ( n315 & n18449 ) | ( n315 & n18454 ) | ( n18449 & n18454 ) ;
  assign n18456 = n240 &  n18455 ;
  assign n18458 = ( n17833 & ~n17824 ) | ( n17833 & n17837 ) | ( ~n17824 & n17837 ) ;
  assign n18457 = n17837 | n17902 ;
  assign n18460 = ( n17837 & ~n18458 ) | ( n17837 & n18457 ) | ( ~n18458 & n18457 ) ;
  assign n18459 = ( n18457 & ~n17833 ) | ( n18457 & n18458 ) | ( ~n17833 & n18458 ) ;
  assign n18461 = ( n17824 & ~n18460 ) | ( n17824 & n18459 ) | ( ~n18460 & n18459 ) ;
  assign n18462 = n315 | n18435 ;
  assign n18463 = n18448 | n18462 ;
  assign n18464 = n18454 &  n18463 ;
  assign n18465 = n18438 | n18441 ;
  assign n18466 = ( n396 & ~n18447 ) | ( n396 & n18465 ) | ( ~n18447 & n18465 ) ;
  assign n18467 = n315 &  n18466 ;
  assign n18468 = n240 | n18467 ;
  assign n18469 = n18464 | n18468 ;
  assign n18470 = ~n18461 & n18469 ;
  assign n18471 = n18456 | n18470 ;
  assign n18472 = ~n17839 & n17902 ;
  assign n18473 = ( n17826 & n17831 ) | ( n17826 & n17902 ) | ( n17831 & n17902 ) ;
  assign n18475 = ( n18472 & ~n17826 ) | ( n18472 & n18473 ) | ( ~n17826 & n18473 ) ;
  assign n18474 = ( n17902 & ~n18473 ) | ( n17902 & n18472 ) | ( ~n18473 & n18472 ) ;
  assign n18476 = ( n17831 & ~n18475 ) | ( n17831 & n18474 ) | ( ~n18475 & n18474 ) ;
  assign n18477 = ( n181 & n18471 ) | ( n181 & n18476 ) | ( n18471 & n18476 ) ;
  assign n18478 = ~n145 & n18477 ;
  assign n18480 = ( n17855 & ~n17846 ) | ( n17855 & n17859 ) | ( ~n17846 & n17859 ) ;
  assign n18479 = n17859 | n17902 ;
  assign n18482 = ( n17859 & ~n18480 ) | ( n17859 & n18479 ) | ( ~n18480 & n18479 ) ;
  assign n18481 = ( n18479 & ~n17855 ) | ( n18479 & n18480 ) | ( ~n17855 & n18480 ) ;
  assign n18483 = ( n17846 & ~n18482 ) | ( n17846 & n18481 ) | ( ~n18482 & n18481 ) ;
  assign n18484 = n181 | n18456 ;
  assign n18485 = n18470 | n18484 ;
  assign n18486 = n18476 &  n18485 ;
  assign n18487 = n18464 | n18467 ;
  assign n18488 = ( n240 & ~n18461 ) | ( n240 & n18487 ) | ( ~n18461 & n18487 ) ;
  assign n18489 = n181 &  n18488 ;
  assign n18490 = ( n145 & ~n18489 ) | ( n145 & 1'b0 ) | ( ~n18489 & 1'b0 ) ;
  assign n18491 = ~n18486 & n18490 ;
  assign n18492 = ( n18483 & ~n18491 ) | ( n18483 & 1'b0 ) | ( ~n18491 & 1'b0 ) ;
  assign n18493 = n18478 | n18492 ;
  assign n18499 = ( n150 & ~n18498 ) | ( n150 & n18493 ) | ( ~n18498 & n18493 ) ;
  assign n18500 = n17868 | n17887 ;
  assign n18501 = ( n17884 & ~n18500 ) | ( n17884 & n17902 ) | ( ~n18500 & n17902 ) ;
  assign n18502 = ~n17884 & n18501 ;
  assign n18503 = n17884 | n17887 ;
  assign n18504 = n17902 | n18503 ;
  assign n18505 = ( n17868 & ~n18504 ) | ( n17868 & n18503 ) | ( ~n18504 & n18503 ) ;
  assign n18506 = n18502 | n18505 ;
  assign n18507 = ( n17869 & ~n17876 ) | ( n17869 & 1'b0 ) | ( ~n17876 & 1'b0 ) ;
  assign n18508 = ~n17902 & n18507 ;
  assign n18509 = ( n17890 & ~n18508 ) | ( n17890 & n18507 ) | ( ~n18508 & n18507 ) ;
  assign n18510 = ( n18506 & ~n18509 ) | ( n18506 & 1'b0 ) | ( ~n18509 & 1'b0 ) ;
  assign n18511 = ~n18499 & n18510 ;
  assign n18512 = ( n133 & ~n18511 ) | ( n133 & n18510 ) | ( ~n18511 & n18510 ) ;
  assign n18515 = n18486 | n18489 ;
  assign n18516 = ( n18483 & ~n145 ) | ( n18483 & n18515 ) | ( ~n145 & n18515 ) ;
  assign n18517 = n150 &  n18516 ;
  assign n18518 = n18506 | n18517 ;
  assign n18513 = n150 | n18478 ;
  assign n18514 = n18492 | n18513 ;
  assign n18519 = n18498 | n18514 ;
  assign n18520 = ( n18518 & ~n18498 ) | ( n18518 & n18519 ) | ( ~n18498 & n18519 ) ;
  assign n18522 = ( n133 & ~n17876 ) | ( n133 & n17869 ) | ( ~n17876 & n17869 ) ;
  assign n18521 = ( n17876 & ~n17869 ) | ( n17876 & n17902 ) | ( ~n17869 & n17902 ) ;
  assign n18523 = ~n17876 & n18521 ;
  assign n18524 = ( n17876 & n18522 ) | ( n17876 & n18523 ) | ( n18522 & n18523 ) ;
  assign n18525 = n17872 | n17899 ;
  assign n18526 = ( n17875 & n17894 ) | ( n17875 & n18525 ) | ( n17894 & n18525 ) ;
  assign n18527 = ( n17875 & ~n18526 ) | ( n17875 & 1'b0 ) | ( ~n18526 & 1'b0 ) ;
  assign n18528 = ( n17882 & ~n18527 ) | ( n17882 & n17890 ) | ( ~n18527 & n17890 ) ;
  assign n18529 = ( n17882 & ~n18528 ) | ( n17882 & 1'b0 ) | ( ~n18528 & 1'b0 ) ;
  assign n18530 = n18524 | n18529 ;
  assign n18531 = ( n18520 & ~n18530 ) | ( n18520 & 1'b0 ) | ( ~n18530 & 1'b0 ) ;
  assign n18532 = ~n18512 | ~n18531 ;
  assign n19081 = n18441 | n18532 ;
  assign n19082 = ( n18433 & n18437 ) | ( n18433 & n18441 ) | ( n18437 & n18441 ) ;
  assign n19083 = ( n19081 & ~n18437 ) | ( n19081 & n19082 ) | ( ~n18437 & n19082 ) ;
  assign n19084 = ( n18441 & ~n19082 ) | ( n18441 & n19081 ) | ( ~n19082 & n19081 ) ;
  assign n19085 = ( n18433 & ~n19083 ) | ( n18433 & n19084 ) | ( ~n19083 & n19084 ) ;
  assign n18539 = ( x14 & ~n18532 ) | ( x14 & x15 ) | ( ~n18532 & x15 ) ;
  assign n18545 = ( x14 & ~x15 ) | ( x14 & 1'b0 ) | ( ~x15 & 1'b0 ) ;
  assign n18535 = x12 | x13 ;
  assign n18540 = ~x14 & n18535 ;
  assign n18541 = ( x14 & ~n17900 ) | ( x14 & n18540 ) | ( ~n17900 & n18540 ) ;
  assign n18542 = ( n17882 & ~n18541 ) | ( n17882 & n17890 ) | ( ~n18541 & n17890 ) ;
  assign n18543 = ( n17882 & ~n18542 ) | ( n17882 & 1'b0 ) | ( ~n18542 & 1'b0 ) ;
  assign n18544 = ( n18532 & ~x15 ) | ( n18532 & n18543 ) | ( ~x15 & n18543 ) ;
  assign n18546 = ( n18539 & ~n18545 ) | ( n18539 & n18544 ) | ( ~n18545 & n18544 ) ;
  assign n18536 = x14 | n18535 ;
  assign n18537 = x14 &  n18532 ;
  assign n18538 = ( n17902 & ~n18536 ) | ( n17902 & n18537 ) | ( ~n18536 & n18537 ) ;
  assign n18547 = n18538 &  n18546 ;
  assign n18548 = ( n17279 & ~n18546 ) | ( n17279 & n18547 ) | ( ~n18546 & n18547 ) ;
  assign n18549 = n17279 | n18538 ;
  assign n18550 = ( n18546 & ~n18549 ) | ( n18546 & 1'b0 ) | ( ~n18549 & 1'b0 ) ;
  assign n18552 = ( n17902 & ~n18529 ) | ( n17902 & 1'b0 ) | ( ~n18529 & 1'b0 ) ;
  assign n18553 = ( n18520 & ~n18552 ) | ( n18520 & n18524 ) | ( ~n18552 & n18524 ) ;
  assign n18554 = ( n18520 & ~n18553 ) | ( n18520 & 1'b0 ) | ( ~n18553 & 1'b0 ) ;
  assign n18555 = n18512 &  n18554 ;
  assign n18551 = ~n17280 & n18532 ;
  assign n18556 = ( n18551 & ~n18555 ) | ( n18551 & 1'b0 ) | ( ~n18555 & 1'b0 ) ;
  assign n18557 = ( x16 & n18555 ) | ( x16 & n18556 ) | ( n18555 & n18556 ) ;
  assign n18558 = x16 | n18555 ;
  assign n18559 = n18551 | n18558 ;
  assign n18560 = ~n18557 & n18559 ;
  assign n18561 = n18550 | n18560 ;
  assign n18562 = ~n18548 & n18561 ;
  assign n18566 = ~x16 & n17902 ;
  assign n18567 = ( x17 & ~n18566 ) | ( x17 & 1'b0 ) | ( ~n18566 & 1'b0 ) ;
  assign n18568 = n17914 | n18567 ;
  assign n18563 = ( n17902 & ~x16 ) | ( n17902 & n17909 ) | ( ~x16 & n17909 ) ;
  assign n18564 = x16 &  n18563 ;
  assign n18565 = ( n17904 & ~n18564 ) | ( n17904 & n17909 ) | ( ~n18564 & n17909 ) ;
  assign n18569 = ( n18532 & ~n18568 ) | ( n18532 & n18565 ) | ( ~n18568 & n18565 ) ;
  assign n18571 = ( n18532 & ~n18569 ) | ( n18532 & 1'b0 ) | ( ~n18569 & 1'b0 ) ;
  assign n18570 = ~n18565 & n18569 ;
  assign n18572 = ( n18568 & ~n18571 ) | ( n18568 & n18570 ) | ( ~n18571 & n18570 ) ;
  assign n18573 = ( n18562 & ~n16671 ) | ( n18562 & n18572 ) | ( ~n16671 & n18572 ) ;
  assign n18574 = ( n16070 & ~n18573 ) | ( n16070 & 1'b0 ) | ( ~n18573 & 1'b0 ) ;
  assign n18575 = ~n17937 & n17940 ;
  assign n18576 = ( n17923 & ~n17937 ) | ( n17923 & n18575 ) | ( ~n17937 & n18575 ) ;
  assign n18578 = ( n18532 & n17937 ) | ( n18532 & n18576 ) | ( n17937 & n18576 ) ;
  assign n18577 = ( n18532 & ~n18576 ) | ( n18532 & n18575 ) | ( ~n18576 & n18575 ) ;
  assign n18579 = ( n17923 & ~n18578 ) | ( n17923 & n18577 ) | ( ~n18578 & n18577 ) ;
  assign n18580 = n16671 | n18548 ;
  assign n18581 = ( n18561 & ~n18580 ) | ( n18561 & 1'b0 ) | ( ~n18580 & 1'b0 ) ;
  assign n18582 = n18572 | n18581 ;
  assign n18583 = ~n18538 & n18546 ;
  assign n18584 = ( n18560 & ~n17279 ) | ( n18560 & n18583 ) | ( ~n17279 & n18583 ) ;
  assign n18585 = ( n16671 & ~n18584 ) | ( n16671 & 1'b0 ) | ( ~n18584 & 1'b0 ) ;
  assign n18586 = n16070 | n18585 ;
  assign n18587 = ( n18582 & ~n18586 ) | ( n18582 & 1'b0 ) | ( ~n18586 & 1'b0 ) ;
  assign n18588 = n18579 | n18587 ;
  assign n18589 = ~n18574 & n18588 ;
  assign n18590 = n17925 | n18532 ;
  assign n18591 = ( n17925 & ~n17942 ) | ( n17925 & n17935 ) | ( ~n17942 & n17935 ) ;
  assign n18592 = ( n17942 & n18590 ) | ( n17942 & n18591 ) | ( n18590 & n18591 ) ;
  assign n18593 = ( n17925 & ~n18591 ) | ( n17925 & n18590 ) | ( ~n18591 & n18590 ) ;
  assign n18594 = ( n17935 & ~n18592 ) | ( n17935 & n18593 ) | ( ~n18592 & n18593 ) ;
  assign n18595 = ( n18589 & ~n15484 ) | ( n18589 & n18594 ) | ( ~n15484 & n18594 ) ;
  assign n18596 = ( n14905 & ~n18595 ) | ( n14905 & 1'b0 ) | ( ~n18595 & 1'b0 ) ;
  assign n18597 = n17962 | n18532 ;
  assign n18598 = ( n17949 & ~n17962 ) | ( n17949 & n17958 ) | ( ~n17962 & n17958 ) ;
  assign n18600 = ( n17962 & n18597 ) | ( n17962 & n18598 ) | ( n18597 & n18598 ) ;
  assign n18599 = ( n17958 & ~n18598 ) | ( n17958 & n18597 ) | ( ~n18598 & n18597 ) ;
  assign n18601 = ( n17949 & ~n18600 ) | ( n17949 & n18599 ) | ( ~n18600 & n18599 ) ;
  assign n18602 = n15484 | n18574 ;
  assign n18603 = ( n18588 & ~n18602 ) | ( n18588 & 1'b0 ) | ( ~n18602 & 1'b0 ) ;
  assign n18604 = n18594 | n18603 ;
  assign n18605 = ( n18582 & ~n18585 ) | ( n18582 & 1'b0 ) | ( ~n18585 & 1'b0 ) ;
  assign n18606 = ( n18579 & ~n16070 ) | ( n18579 & n18605 ) | ( ~n16070 & n18605 ) ;
  assign n18607 = ( n15484 & ~n18606 ) | ( n15484 & 1'b0 ) | ( ~n18606 & 1'b0 ) ;
  assign n18608 = n14905 | n18607 ;
  assign n18609 = ( n18604 & ~n18608 ) | ( n18604 & 1'b0 ) | ( ~n18608 & 1'b0 ) ;
  assign n18610 = n18601 | n18609 ;
  assign n18611 = ~n18596 & n18610 ;
  assign n18612 = n17964 &  n18532 ;
  assign n18613 = ( n17951 & n17956 ) | ( n17951 & n18532 ) | ( n17956 & n18532 ) ;
  assign n18615 = ( n18612 & ~n17951 ) | ( n18612 & n18613 ) | ( ~n17951 & n18613 ) ;
  assign n18614 = ( n18532 & ~n18613 ) | ( n18532 & n18612 ) | ( ~n18613 & n18612 ) ;
  assign n18616 = ( n17956 & ~n18615 ) | ( n17956 & n18614 ) | ( ~n18615 & n18614 ) ;
  assign n18617 = ( n18611 & ~n14341 ) | ( n18611 & n18616 ) | ( ~n14341 & n18616 ) ;
  assign n18618 = ( n13784 & ~n18617 ) | ( n13784 & 1'b0 ) | ( ~n18617 & 1'b0 ) ;
  assign n18619 = n17984 | n18532 ;
  assign n18620 = ( n17971 & ~n17980 ) | ( n17971 & n17984 ) | ( ~n17980 & n17984 ) ;
  assign n18621 = ( n17980 & n18619 ) | ( n17980 & n18620 ) | ( n18619 & n18620 ) ;
  assign n18622 = ( n17984 & ~n18620 ) | ( n17984 & n18619 ) | ( ~n18620 & n18619 ) ;
  assign n18623 = ( n17971 & ~n18621 ) | ( n17971 & n18622 ) | ( ~n18621 & n18622 ) ;
  assign n18624 = n14341 | n18596 ;
  assign n18625 = ( n18610 & ~n18624 ) | ( n18610 & 1'b0 ) | ( ~n18624 & 1'b0 ) ;
  assign n18626 = n18616 | n18625 ;
  assign n18627 = ( n18604 & ~n18607 ) | ( n18604 & 1'b0 ) | ( ~n18607 & 1'b0 ) ;
  assign n18628 = ( n18601 & ~n14905 ) | ( n18601 & n18627 ) | ( ~n14905 & n18627 ) ;
  assign n18629 = ( n14341 & ~n18628 ) | ( n14341 & 1'b0 ) | ( ~n18628 & 1'b0 ) ;
  assign n18630 = n13784 | n18629 ;
  assign n18631 = ( n18626 & ~n18630 ) | ( n18626 & 1'b0 ) | ( ~n18630 & 1'b0 ) ;
  assign n18632 = n18623 | n18631 ;
  assign n18633 = ~n18618 & n18632 ;
  assign n18634 = n17973 | n18532 ;
  assign n18635 = ( n17978 & ~n17973 ) | ( n17978 & n17986 ) | ( ~n17973 & n17986 ) ;
  assign n18637 = ( n17973 & n18634 ) | ( n17973 & n18635 ) | ( n18634 & n18635 ) ;
  assign n18636 = ( n17986 & ~n18635 ) | ( n17986 & n18634 ) | ( ~n18635 & n18634 ) ;
  assign n18638 = ( n17978 & ~n18637 ) | ( n17978 & n18636 ) | ( ~n18637 & n18636 ) ;
  assign n18639 = ( n18633 & ~n13242 ) | ( n18633 & n18638 ) | ( ~n13242 & n18638 ) ;
  assign n18640 = ( n12707 & ~n18639 ) | ( n12707 & 1'b0 ) | ( ~n18639 & 1'b0 ) ;
  assign n18641 = n18006 | n18532 ;
  assign n18642 = ( n17993 & ~n18002 ) | ( n17993 & n18006 ) | ( ~n18002 & n18006 ) ;
  assign n18643 = ( n18002 & n18641 ) | ( n18002 & n18642 ) | ( n18641 & n18642 ) ;
  assign n18644 = ( n18006 & ~n18642 ) | ( n18006 & n18641 ) | ( ~n18642 & n18641 ) ;
  assign n18645 = ( n17993 & ~n18643 ) | ( n17993 & n18644 ) | ( ~n18643 & n18644 ) ;
  assign n18646 = n13242 | n18618 ;
  assign n18647 = ( n18632 & ~n18646 ) | ( n18632 & 1'b0 ) | ( ~n18646 & 1'b0 ) ;
  assign n18648 = n18638 | n18647 ;
  assign n18649 = ( n18626 & ~n18629 ) | ( n18626 & 1'b0 ) | ( ~n18629 & 1'b0 ) ;
  assign n18650 = ( n18623 & ~n13784 ) | ( n18623 & n18649 ) | ( ~n13784 & n18649 ) ;
  assign n18651 = ( n13242 & ~n18650 ) | ( n13242 & 1'b0 ) | ( ~n18650 & 1'b0 ) ;
  assign n18652 = n12707 | n18651 ;
  assign n18653 = ( n18648 & ~n18652 ) | ( n18648 & 1'b0 ) | ( ~n18652 & 1'b0 ) ;
  assign n18654 = n18645 | n18653 ;
  assign n18655 = ~n18640 & n18654 ;
  assign n18656 = n17995 | n18532 ;
  assign n18657 = ( n17995 & ~n18008 ) | ( n17995 & n18000 ) | ( ~n18008 & n18000 ) ;
  assign n18658 = ( n18008 & n18656 ) | ( n18008 & n18657 ) | ( n18656 & n18657 ) ;
  assign n18659 = ( n17995 & ~n18657 ) | ( n17995 & n18656 ) | ( ~n18657 & n18656 ) ;
  assign n18660 = ( n18000 & ~n18658 ) | ( n18000 & n18659 ) | ( ~n18658 & n18659 ) ;
  assign n18661 = ( n18655 & ~n12187 ) | ( n18655 & n18660 ) | ( ~n12187 & n18660 ) ;
  assign n18662 = ( n11674 & ~n18661 ) | ( n11674 & 1'b0 ) | ( ~n18661 & 1'b0 ) ;
  assign n18663 = n18028 | n18532 ;
  assign n18664 = ( n18015 & ~n18028 ) | ( n18015 & n18024 ) | ( ~n18028 & n18024 ) ;
  assign n18666 = ( n18028 & n18663 ) | ( n18028 & n18664 ) | ( n18663 & n18664 ) ;
  assign n18665 = ( n18024 & ~n18664 ) | ( n18024 & n18663 ) | ( ~n18664 & n18663 ) ;
  assign n18667 = ( n18015 & ~n18666 ) | ( n18015 & n18665 ) | ( ~n18666 & n18665 ) ;
  assign n18668 = n12187 | n18640 ;
  assign n18669 = ( n18654 & ~n18668 ) | ( n18654 & 1'b0 ) | ( ~n18668 & 1'b0 ) ;
  assign n18670 = n18660 | n18669 ;
  assign n18671 = ( n18648 & ~n18651 ) | ( n18648 & 1'b0 ) | ( ~n18651 & 1'b0 ) ;
  assign n18672 = ( n18645 & ~n12707 ) | ( n18645 & n18671 ) | ( ~n12707 & n18671 ) ;
  assign n18673 = ( n12187 & ~n18672 ) | ( n12187 & 1'b0 ) | ( ~n18672 & 1'b0 ) ;
  assign n18674 = n11674 | n18673 ;
  assign n18675 = ( n18670 & ~n18674 ) | ( n18670 & 1'b0 ) | ( ~n18674 & 1'b0 ) ;
  assign n18676 = n18667 | n18675 ;
  assign n18677 = ~n18662 & n18676 ;
  assign n18678 = n18030 &  n18532 ;
  assign n18679 = ( n18017 & n18022 ) | ( n18017 & n18532 ) | ( n18022 & n18532 ) ;
  assign n18681 = ( n18678 & ~n18017 ) | ( n18678 & n18679 ) | ( ~n18017 & n18679 ) ;
  assign n18680 = ( n18532 & ~n18679 ) | ( n18532 & n18678 ) | ( ~n18679 & n18678 ) ;
  assign n18682 = ( n18022 & ~n18681 ) | ( n18022 & n18680 ) | ( ~n18681 & n18680 ) ;
  assign n18683 = ( n18677 & ~n11176 ) | ( n18677 & n18682 ) | ( ~n11176 & n18682 ) ;
  assign n18684 = ( n10685 & ~n18683 ) | ( n10685 & 1'b0 ) | ( ~n18683 & 1'b0 ) ;
  assign n18685 = n18050 | n18532 ;
  assign n18686 = ( n18037 & ~n18046 ) | ( n18037 & n18050 ) | ( ~n18046 & n18050 ) ;
  assign n18687 = ( n18046 & n18685 ) | ( n18046 & n18686 ) | ( n18685 & n18686 ) ;
  assign n18688 = ( n18050 & ~n18686 ) | ( n18050 & n18685 ) | ( ~n18686 & n18685 ) ;
  assign n18689 = ( n18037 & ~n18687 ) | ( n18037 & n18688 ) | ( ~n18687 & n18688 ) ;
  assign n18690 = n11176 | n18662 ;
  assign n18691 = ( n18676 & ~n18690 ) | ( n18676 & 1'b0 ) | ( ~n18690 & 1'b0 ) ;
  assign n18692 = n18682 | n18691 ;
  assign n18693 = ( n18670 & ~n18673 ) | ( n18670 & 1'b0 ) | ( ~n18673 & 1'b0 ) ;
  assign n18694 = ( n18667 & ~n11674 ) | ( n18667 & n18693 ) | ( ~n11674 & n18693 ) ;
  assign n18695 = ( n11176 & ~n18694 ) | ( n11176 & 1'b0 ) | ( ~n18694 & 1'b0 ) ;
  assign n18696 = n10685 | n18695 ;
  assign n18697 = ( n18692 & ~n18696 ) | ( n18692 & 1'b0 ) | ( ~n18696 & 1'b0 ) ;
  assign n18698 = n18689 | n18697 ;
  assign n18699 = ~n18684 & n18698 ;
  assign n18700 = n18039 | n18532 ;
  assign n18701 = ( n18044 & ~n18039 ) | ( n18044 & n18052 ) | ( ~n18039 & n18052 ) ;
  assign n18703 = ( n18039 & n18700 ) | ( n18039 & n18701 ) | ( n18700 & n18701 ) ;
  assign n18702 = ( n18052 & ~n18701 ) | ( n18052 & n18700 ) | ( ~n18701 & n18700 ) ;
  assign n18704 = ( n18044 & ~n18703 ) | ( n18044 & n18702 ) | ( ~n18703 & n18702 ) ;
  assign n18705 = ( n18699 & ~n10209 ) | ( n18699 & n18704 ) | ( ~n10209 & n18704 ) ;
  assign n18706 = n9740 | n18705 ;
  assign n18707 = n18072 | n18532 ;
  assign n18708 = ( n18059 & ~n18068 ) | ( n18059 & n18072 ) | ( ~n18068 & n18072 ) ;
  assign n18709 = ( n18068 & n18707 ) | ( n18068 & n18708 ) | ( n18707 & n18708 ) ;
  assign n18710 = ( n18072 & ~n18708 ) | ( n18072 & n18707 ) | ( ~n18708 & n18707 ) ;
  assign n18711 = ( n18059 & ~n18709 ) | ( n18059 & n18710 ) | ( ~n18709 & n18710 ) ;
  assign n18712 = n10209 | n18684 ;
  assign n18713 = ( n18698 & ~n18712 ) | ( n18698 & 1'b0 ) | ( ~n18712 & 1'b0 ) ;
  assign n18714 = n18704 | n18713 ;
  assign n18715 = ( n18692 & ~n18695 ) | ( n18692 & 1'b0 ) | ( ~n18695 & 1'b0 ) ;
  assign n18716 = ( n18689 & ~n10685 ) | ( n18689 & n18715 ) | ( ~n10685 & n18715 ) ;
  assign n18717 = ( n10209 & ~n18716 ) | ( n10209 & 1'b0 ) | ( ~n18716 & 1'b0 ) ;
  assign n18718 = ( n9740 & ~n18717 ) | ( n9740 & 1'b0 ) | ( ~n18717 & 1'b0 ) ;
  assign n18719 = n18714 &  n18718 ;
  assign n18720 = n18711 | n18719 ;
  assign n18721 = n18706 &  n18720 ;
  assign n18723 = ( n18061 & ~n18066 ) | ( n18061 & n18074 ) | ( ~n18066 & n18074 ) ;
  assign n18722 = ( n18061 & ~n18532 ) | ( n18061 & 1'b0 ) | ( ~n18532 & 1'b0 ) ;
  assign n18725 = ( n18061 & ~n18723 ) | ( n18061 & n18722 ) | ( ~n18723 & n18722 ) ;
  assign n18724 = ( n18722 & ~n18074 ) | ( n18722 & n18723 ) | ( ~n18074 & n18723 ) ;
  assign n18726 = ( n18066 & ~n18725 ) | ( n18066 & n18724 ) | ( ~n18725 & n18724 ) ;
  assign n18727 = ( n18721 & ~n9286 ) | ( n18721 & n18726 ) | ( ~n9286 & n18726 ) ;
  assign n18728 = ( n8839 & ~n18727 ) | ( n8839 & 1'b0 ) | ( ~n18727 & 1'b0 ) ;
  assign n18729 = n18094 | n18532 ;
  assign n18730 = ( n18081 & ~n18094 ) | ( n18081 & n18090 ) | ( ~n18094 & n18090 ) ;
  assign n18732 = ( n18094 & n18729 ) | ( n18094 & n18730 ) | ( n18729 & n18730 ) ;
  assign n18731 = ( n18090 & ~n18730 ) | ( n18090 & n18729 ) | ( ~n18730 & n18729 ) ;
  assign n18733 = ( n18081 & ~n18732 ) | ( n18081 & n18731 ) | ( ~n18732 & n18731 ) ;
  assign n18734 = ~n9286 & n18706 ;
  assign n18735 = n18720 &  n18734 ;
  assign n18736 = n18726 | n18735 ;
  assign n18737 = ( n18714 & ~n18717 ) | ( n18714 & 1'b0 ) | ( ~n18717 & 1'b0 ) ;
  assign n18738 = ( n9740 & n18711 ) | ( n9740 & n18737 ) | ( n18711 & n18737 ) ;
  assign n18739 = ( n9286 & ~n18738 ) | ( n9286 & 1'b0 ) | ( ~n18738 & 1'b0 ) ;
  assign n18740 = n8839 | n18739 ;
  assign n18741 = ( n18736 & ~n18740 ) | ( n18736 & 1'b0 ) | ( ~n18740 & 1'b0 ) ;
  assign n18742 = n18733 | n18741 ;
  assign n18743 = ~n18728 & n18742 ;
  assign n18745 = ( n18083 & ~n18088 ) | ( n18083 & n18532 ) | ( ~n18088 & n18532 ) ;
  assign n18744 = n18096 &  n18532 ;
  assign n18746 = ( n18532 & ~n18745 ) | ( n18532 & n18744 ) | ( ~n18745 & n18744 ) ;
  assign n18747 = ( n18744 & ~n18083 ) | ( n18744 & n18745 ) | ( ~n18083 & n18745 ) ;
  assign n18748 = ( n18088 & ~n18746 ) | ( n18088 & n18747 ) | ( ~n18746 & n18747 ) ;
  assign n18749 = ( n18743 & ~n8407 ) | ( n18743 & n18748 ) | ( ~n8407 & n18748 ) ;
  assign n18750 = ( n7982 & ~n18749 ) | ( n7982 & 1'b0 ) | ( ~n18749 & 1'b0 ) ;
  assign n18751 = n18116 | n18532 ;
  assign n18752 = ( n18103 & ~n18112 ) | ( n18103 & n18116 ) | ( ~n18112 & n18116 ) ;
  assign n18753 = ( n18112 & n18751 ) | ( n18112 & n18752 ) | ( n18751 & n18752 ) ;
  assign n18754 = ( n18116 & ~n18752 ) | ( n18116 & n18751 ) | ( ~n18752 & n18751 ) ;
  assign n18755 = ( n18103 & ~n18753 ) | ( n18103 & n18754 ) | ( ~n18753 & n18754 ) ;
  assign n18756 = n8407 | n18728 ;
  assign n18757 = ( n18742 & ~n18756 ) | ( n18742 & 1'b0 ) | ( ~n18756 & 1'b0 ) ;
  assign n18758 = n18748 | n18757 ;
  assign n18759 = ( n18736 & ~n18739 ) | ( n18736 & 1'b0 ) | ( ~n18739 & 1'b0 ) ;
  assign n18760 = ( n18733 & ~n8839 ) | ( n18733 & n18759 ) | ( ~n8839 & n18759 ) ;
  assign n18761 = ( n8407 & ~n18760 ) | ( n8407 & 1'b0 ) | ( ~n18760 & 1'b0 ) ;
  assign n18762 = n7982 | n18761 ;
  assign n18763 = ( n18758 & ~n18762 ) | ( n18758 & 1'b0 ) | ( ~n18762 & 1'b0 ) ;
  assign n18764 = n18755 | n18763 ;
  assign n18765 = ~n18750 & n18764 ;
  assign n18766 = n18105 | n18532 ;
  assign n18767 = ( n18110 & ~n18105 ) | ( n18110 & n18118 ) | ( ~n18105 & n18118 ) ;
  assign n18769 = ( n18105 & n18766 ) | ( n18105 & n18767 ) | ( n18766 & n18767 ) ;
  assign n18768 = ( n18118 & ~n18767 ) | ( n18118 & n18766 ) | ( ~n18767 & n18766 ) ;
  assign n18770 = ( n18110 & ~n18769 ) | ( n18110 & n18768 ) | ( ~n18769 & n18768 ) ;
  assign n18771 = ( n7572 & n18765 ) | ( n7572 & n18770 ) | ( n18765 & n18770 ) ;
  assign n18772 = n7169 | n18771 ;
  assign n18774 = ( n18134 & ~n18125 ) | ( n18134 & n18138 ) | ( ~n18125 & n18138 ) ;
  assign n18773 = ( n18138 & ~n18532 ) | ( n18138 & 1'b0 ) | ( ~n18532 & 1'b0 ) ;
  assign n18776 = ( n18138 & ~n18774 ) | ( n18138 & n18773 ) | ( ~n18774 & n18773 ) ;
  assign n18775 = ( n18773 & ~n18134 ) | ( n18773 & n18774 ) | ( ~n18134 & n18774 ) ;
  assign n18777 = ( n18125 & ~n18776 ) | ( n18125 & n18775 ) | ( ~n18776 & n18775 ) ;
  assign n18778 = ( n7572 & ~n18750 ) | ( n7572 & 1'b0 ) | ( ~n18750 & 1'b0 ) ;
  assign n18779 = n18764 &  n18778 ;
  assign n18780 = n18770 | n18779 ;
  assign n18781 = ( n18758 & ~n18761 ) | ( n18758 & 1'b0 ) | ( ~n18761 & 1'b0 ) ;
  assign n18782 = ( n18755 & ~n7982 ) | ( n18755 & n18781 ) | ( ~n7982 & n18781 ) ;
  assign n18783 = n7572 | n18782 ;
  assign n18784 = n7169 &  n18783 ;
  assign n18785 = n18780 &  n18784 ;
  assign n18786 = n18777 | n18785 ;
  assign n18787 = n18772 &  n18786 ;
  assign n18788 = ( n18127 & ~n18532 ) | ( n18127 & 1'b0 ) | ( ~n18532 & 1'b0 ) ;
  assign n18789 = ( n18127 & n18132 ) | ( n18127 & n18140 ) | ( n18132 & n18140 ) ;
  assign n18790 = ( n18788 & ~n18140 ) | ( n18788 & n18789 ) | ( ~n18140 & n18789 ) ;
  assign n18791 = ( n18127 & ~n18789 ) | ( n18127 & n18788 ) | ( ~n18789 & n18788 ) ;
  assign n18792 = ( n18132 & ~n18790 ) | ( n18132 & n18791 ) | ( ~n18790 & n18791 ) ;
  assign n18793 = ( n18787 & ~n6781 ) | ( n18787 & n18792 ) | ( ~n6781 & n18792 ) ;
  assign n18794 = n6399 | n18793 ;
  assign n18795 = n18160 | n18532 ;
  assign n18796 = ( n18147 & ~n18156 ) | ( n18147 & n18160 ) | ( ~n18156 & n18160 ) ;
  assign n18797 = ( n18156 & n18795 ) | ( n18156 & n18796 ) | ( n18795 & n18796 ) ;
  assign n18798 = ( n18160 & ~n18796 ) | ( n18160 & n18795 ) | ( ~n18796 & n18795 ) ;
  assign n18799 = ( n18147 & ~n18797 ) | ( n18147 & n18798 ) | ( ~n18797 & n18798 ) ;
  assign n18800 = ~n6781 & n18772 ;
  assign n18801 = n18786 &  n18800 ;
  assign n18802 = n18792 | n18801 ;
  assign n18803 = n18780 &  n18783 ;
  assign n18804 = ( n7169 & n18777 ) | ( n7169 & n18803 ) | ( n18777 & n18803 ) ;
  assign n18805 = ( n6781 & ~n18804 ) | ( n6781 & 1'b0 ) | ( ~n18804 & 1'b0 ) ;
  assign n18806 = ( n6399 & ~n18805 ) | ( n6399 & 1'b0 ) | ( ~n18805 & 1'b0 ) ;
  assign n18807 = n18802 &  n18806 ;
  assign n18808 = n18799 | n18807 ;
  assign n18809 = n18794 &  n18808 ;
  assign n18810 = ( n18149 & ~n18532 ) | ( n18149 & 1'b0 ) | ( ~n18532 & 1'b0 ) ;
  assign n18811 = ( n18149 & n18154 ) | ( n18149 & n18162 ) | ( n18154 & n18162 ) ;
  assign n18812 = ( n18810 & ~n18162 ) | ( n18810 & n18811 ) | ( ~n18162 & n18811 ) ;
  assign n18813 = ( n18149 & ~n18811 ) | ( n18149 & n18810 ) | ( ~n18811 & n18810 ) ;
  assign n18814 = ( n18154 & ~n18812 ) | ( n18154 & n18813 ) | ( ~n18812 & n18813 ) ;
  assign n18815 = ( n18809 & ~n6032 ) | ( n18809 & n18814 ) | ( ~n6032 & n18814 ) ;
  assign n18816 = n5672 | n18815 ;
  assign n18817 = n18182 | n18532 ;
  assign n18818 = ( n18169 & ~n18178 ) | ( n18169 & n18182 ) | ( ~n18178 & n18182 ) ;
  assign n18819 = ( n18178 & n18817 ) | ( n18178 & n18818 ) | ( n18817 & n18818 ) ;
  assign n18820 = ( n18182 & ~n18818 ) | ( n18182 & n18817 ) | ( ~n18818 & n18817 ) ;
  assign n18821 = ( n18169 & ~n18819 ) | ( n18169 & n18820 ) | ( ~n18819 & n18820 ) ;
  assign n18822 = ~n6032 & n18794 ;
  assign n18823 = n18808 &  n18822 ;
  assign n18824 = n18814 | n18823 ;
  assign n18825 = ( n18802 & ~n18805 ) | ( n18802 & 1'b0 ) | ( ~n18805 & 1'b0 ) ;
  assign n18826 = ( n6399 & n18799 ) | ( n6399 & n18825 ) | ( n18799 & n18825 ) ;
  assign n18827 = ( n6032 & ~n18826 ) | ( n6032 & 1'b0 ) | ( ~n18826 & 1'b0 ) ;
  assign n18828 = ( n5672 & ~n18827 ) | ( n5672 & 1'b0 ) | ( ~n18827 & 1'b0 ) ;
  assign n18829 = n18824 &  n18828 ;
  assign n18830 = n18821 | n18829 ;
  assign n18831 = n18816 &  n18830 ;
  assign n18832 = ( n18171 & ~n18532 ) | ( n18171 & 1'b0 ) | ( ~n18532 & 1'b0 ) ;
  assign n18833 = ( n18171 & n18176 ) | ( n18171 & n18184 ) | ( n18176 & n18184 ) ;
  assign n18834 = ( n18832 & ~n18184 ) | ( n18832 & n18833 ) | ( ~n18184 & n18833 ) ;
  assign n18835 = ( n18171 & ~n18833 ) | ( n18171 & n18832 ) | ( ~n18833 & n18832 ) ;
  assign n18836 = ( n18176 & ~n18834 ) | ( n18176 & n18835 ) | ( ~n18834 & n18835 ) ;
  assign n18837 = ( n18831 & ~n5327 ) | ( n18831 & n18836 ) | ( ~n5327 & n18836 ) ;
  assign n18838 = ( n4990 & ~n18837 ) | ( n4990 & 1'b0 ) | ( ~n18837 & 1'b0 ) ;
  assign n18839 = n18204 | n18532 ;
  assign n18840 = ( n18191 & ~n18200 ) | ( n18191 & n18204 ) | ( ~n18200 & n18204 ) ;
  assign n18841 = ( n18200 & n18839 ) | ( n18200 & n18840 ) | ( n18839 & n18840 ) ;
  assign n18842 = ( n18204 & ~n18840 ) | ( n18204 & n18839 ) | ( ~n18840 & n18839 ) ;
  assign n18843 = ( n18191 & ~n18841 ) | ( n18191 & n18842 ) | ( ~n18841 & n18842 ) ;
  assign n18844 = ~n5327 & n18816 ;
  assign n18845 = n18830 &  n18844 ;
  assign n18846 = n18836 | n18845 ;
  assign n18847 = ( n18824 & ~n18827 ) | ( n18824 & 1'b0 ) | ( ~n18827 & 1'b0 ) ;
  assign n18848 = ( n5672 & n18821 ) | ( n5672 & n18847 ) | ( n18821 & n18847 ) ;
  assign n18849 = ( n5327 & ~n18848 ) | ( n5327 & 1'b0 ) | ( ~n18848 & 1'b0 ) ;
  assign n18850 = n4990 | n18849 ;
  assign n18851 = ( n18846 & ~n18850 ) | ( n18846 & 1'b0 ) | ( ~n18850 & 1'b0 ) ;
  assign n18852 = n18843 | n18851 ;
  assign n18853 = ~n18838 & n18852 ;
  assign n18854 = n18193 | n18532 ;
  assign n18855 = ( n18198 & ~n18193 ) | ( n18198 & n18206 ) | ( ~n18193 & n18206 ) ;
  assign n18857 = ( n18193 & n18854 ) | ( n18193 & n18855 ) | ( n18854 & n18855 ) ;
  assign n18856 = ( n18206 & ~n18855 ) | ( n18206 & n18854 ) | ( ~n18855 & n18854 ) ;
  assign n18858 = ( n18198 & ~n18857 ) | ( n18198 & n18856 ) | ( ~n18857 & n18856 ) ;
  assign n18859 = ( n18853 & ~n4668 ) | ( n18853 & n18858 ) | ( ~n4668 & n18858 ) ;
  assign n18860 = ( n4353 & ~n18859 ) | ( n4353 & 1'b0 ) | ( ~n18859 & 1'b0 ) ;
  assign n18861 = n18226 | n18532 ;
  assign n18862 = ( n18213 & ~n18222 ) | ( n18213 & n18226 ) | ( ~n18222 & n18226 ) ;
  assign n18863 = ( n18222 & n18861 ) | ( n18222 & n18862 ) | ( n18861 & n18862 ) ;
  assign n18864 = ( n18226 & ~n18862 ) | ( n18226 & n18861 ) | ( ~n18862 & n18861 ) ;
  assign n18865 = ( n18213 & ~n18863 ) | ( n18213 & n18864 ) | ( ~n18863 & n18864 ) ;
  assign n18866 = n4668 | n18838 ;
  assign n18867 = ( n18852 & ~n18866 ) | ( n18852 & 1'b0 ) | ( ~n18866 & 1'b0 ) ;
  assign n18868 = n18858 | n18867 ;
  assign n18869 = ( n18846 & ~n18849 ) | ( n18846 & 1'b0 ) | ( ~n18849 & 1'b0 ) ;
  assign n18870 = ( n18843 & ~n4990 ) | ( n18843 & n18869 ) | ( ~n4990 & n18869 ) ;
  assign n18871 = ( n4668 & ~n18870 ) | ( n4668 & 1'b0 ) | ( ~n18870 & 1'b0 ) ;
  assign n18872 = n4353 | n18871 ;
  assign n18873 = ( n18868 & ~n18872 ) | ( n18868 & 1'b0 ) | ( ~n18872 & 1'b0 ) ;
  assign n18874 = n18865 | n18873 ;
  assign n18875 = ~n18860 & n18874 ;
  assign n18876 = n18215 | n18532 ;
  assign n18877 = ( n18220 & ~n18215 ) | ( n18220 & n18228 ) | ( ~n18215 & n18228 ) ;
  assign n18879 = ( n18215 & n18876 ) | ( n18215 & n18877 ) | ( n18876 & n18877 ) ;
  assign n18878 = ( n18228 & ~n18877 ) | ( n18228 & n18876 ) | ( ~n18877 & n18876 ) ;
  assign n18880 = ( n18220 & ~n18879 ) | ( n18220 & n18878 ) | ( ~n18879 & n18878 ) ;
  assign n18881 = ( n18875 & ~n4053 ) | ( n18875 & n18880 ) | ( ~n4053 & n18880 ) ;
  assign n18882 = ( n3760 & ~n18881 ) | ( n3760 & 1'b0 ) | ( ~n18881 & 1'b0 ) ;
  assign n18883 = n18248 | n18532 ;
  assign n18884 = ( n18235 & ~n18244 ) | ( n18235 & n18248 ) | ( ~n18244 & n18248 ) ;
  assign n18885 = ( n18244 & n18883 ) | ( n18244 & n18884 ) | ( n18883 & n18884 ) ;
  assign n18886 = ( n18248 & ~n18884 ) | ( n18248 & n18883 ) | ( ~n18884 & n18883 ) ;
  assign n18887 = ( n18235 & ~n18885 ) | ( n18235 & n18886 ) | ( ~n18885 & n18886 ) ;
  assign n18888 = n4053 | n18860 ;
  assign n18889 = ( n18874 & ~n18888 ) | ( n18874 & 1'b0 ) | ( ~n18888 & 1'b0 ) ;
  assign n18890 = n18880 | n18889 ;
  assign n18891 = ( n18868 & ~n18871 ) | ( n18868 & 1'b0 ) | ( ~n18871 & 1'b0 ) ;
  assign n18892 = ( n18865 & ~n4353 ) | ( n18865 & n18891 ) | ( ~n4353 & n18891 ) ;
  assign n18893 = ( n4053 & ~n18892 ) | ( n4053 & 1'b0 ) | ( ~n18892 & 1'b0 ) ;
  assign n18894 = n3760 | n18893 ;
  assign n18895 = ( n18890 & ~n18894 ) | ( n18890 & 1'b0 ) | ( ~n18894 & 1'b0 ) ;
  assign n18896 = n18887 | n18895 ;
  assign n18897 = ~n18882 & n18896 ;
  assign n18898 = n18237 | n18532 ;
  assign n18899 = ( n18237 & ~n18250 ) | ( n18237 & n18242 ) | ( ~n18250 & n18242 ) ;
  assign n18900 = ( n18250 & n18898 ) | ( n18250 & n18899 ) | ( n18898 & n18899 ) ;
  assign n18901 = ( n18237 & ~n18899 ) | ( n18237 & n18898 ) | ( ~n18899 & n18898 ) ;
  assign n18902 = ( n18242 & ~n18900 ) | ( n18242 & n18901 ) | ( ~n18900 & n18901 ) ;
  assign n18903 = ( n3482 & ~n18897 ) | ( n3482 & n18902 ) | ( ~n18897 & n18902 ) ;
  assign n18904 = n3211 &  n18903 ;
  assign n18906 = ( n18266 & ~n18257 ) | ( n18266 & n18270 ) | ( ~n18257 & n18270 ) ;
  assign n18905 = n18270 | n18532 ;
  assign n18908 = ( n18270 & ~n18906 ) | ( n18270 & n18905 ) | ( ~n18906 & n18905 ) ;
  assign n18907 = ( n18905 & ~n18266 ) | ( n18905 & n18906 ) | ( ~n18266 & n18906 ) ;
  assign n18909 = ( n18257 & ~n18908 ) | ( n18257 & n18907 ) | ( ~n18908 & n18907 ) ;
  assign n18910 = n3482 | n18882 ;
  assign n18911 = ( n18896 & ~n18910 ) | ( n18896 & 1'b0 ) | ( ~n18910 & 1'b0 ) ;
  assign n18912 = ( n18902 & ~n18911 ) | ( n18902 & 1'b0 ) | ( ~n18911 & 1'b0 ) ;
  assign n18913 = ( n18890 & ~n18893 ) | ( n18890 & 1'b0 ) | ( ~n18893 & 1'b0 ) ;
  assign n18914 = ( n18887 & ~n3760 ) | ( n18887 & n18913 ) | ( ~n3760 & n18913 ) ;
  assign n18915 = ( n3482 & ~n18914 ) | ( n3482 & 1'b0 ) | ( ~n18914 & 1'b0 ) ;
  assign n18916 = n3211 | n18915 ;
  assign n18917 = n18912 | n18916 ;
  assign n18918 = n18909 &  n18917 ;
  assign n18919 = n18904 | n18918 ;
  assign n18920 = n18259 | n18532 ;
  assign n18921 = ( n18259 & n18264 ) | ( n18259 & n18272 ) | ( n18264 & n18272 ) ;
  assign n18922 = ( n18920 & ~n18272 ) | ( n18920 & n18921 ) | ( ~n18272 & n18921 ) ;
  assign n18923 = ( n18259 & ~n18921 ) | ( n18259 & n18920 ) | ( ~n18921 & n18920 ) ;
  assign n18924 = ( n18264 & ~n18922 ) | ( n18264 & n18923 ) | ( ~n18922 & n18923 ) ;
  assign n18925 = ( n2955 & n18919 ) | ( n2955 & n18924 ) | ( n18919 & n18924 ) ;
  assign n18926 = n2706 &  n18925 ;
  assign n18928 = ( n18288 & ~n18279 ) | ( n18288 & n18292 ) | ( ~n18279 & n18292 ) ;
  assign n18927 = n18292 | n18532 ;
  assign n18930 = ( n18292 & ~n18928 ) | ( n18292 & n18927 ) | ( ~n18928 & n18927 ) ;
  assign n18929 = ( n18927 & ~n18288 ) | ( n18927 & n18928 ) | ( ~n18288 & n18928 ) ;
  assign n18931 = ( n18279 & ~n18930 ) | ( n18279 & n18929 ) | ( ~n18930 & n18929 ) ;
  assign n18932 = n2955 | n18904 ;
  assign n18933 = n18918 | n18932 ;
  assign n18934 = n18924 &  n18933 ;
  assign n18935 = n18912 | n18915 ;
  assign n18936 = ( n3211 & n18909 ) | ( n3211 & n18935 ) | ( n18909 & n18935 ) ;
  assign n18937 = n2955 &  n18936 ;
  assign n18938 = n2706 | n18937 ;
  assign n18939 = n18934 | n18938 ;
  assign n18940 = n18931 &  n18939 ;
  assign n18941 = n18926 | n18940 ;
  assign n18942 = n18281 | n18532 ;
  assign n18943 = ( n18281 & n18286 ) | ( n18281 & n18294 ) | ( n18286 & n18294 ) ;
  assign n18944 = ( n18942 & ~n18294 ) | ( n18942 & n18943 ) | ( ~n18294 & n18943 ) ;
  assign n18945 = ( n18281 & ~n18943 ) | ( n18281 & n18942 ) | ( ~n18943 & n18942 ) ;
  assign n18946 = ( n18286 & ~n18944 ) | ( n18286 & n18945 ) | ( ~n18944 & n18945 ) ;
  assign n18947 = ( n2472 & n18941 ) | ( n2472 & n18946 ) | ( n18941 & n18946 ) ;
  assign n18948 = n2245 &  n18947 ;
  assign n18949 = n18314 | n18532 ;
  assign n18950 = ( n18301 & n18310 ) | ( n18301 & n18314 ) | ( n18310 & n18314 ) ;
  assign n18951 = ( n18949 & ~n18310 ) | ( n18949 & n18950 ) | ( ~n18310 & n18950 ) ;
  assign n18952 = ( n18314 & ~n18950 ) | ( n18314 & n18949 ) | ( ~n18950 & n18949 ) ;
  assign n18953 = ( n18301 & ~n18951 ) | ( n18301 & n18952 ) | ( ~n18951 & n18952 ) ;
  assign n18954 = n2472 | n18926 ;
  assign n18955 = n18940 | n18954 ;
  assign n18956 = n18946 &  n18955 ;
  assign n18957 = n18934 | n18937 ;
  assign n18958 = ( n2706 & n18931 ) | ( n2706 & n18957 ) | ( n18931 & n18957 ) ;
  assign n18959 = n2472 &  n18958 ;
  assign n18960 = n2245 | n18959 ;
  assign n18961 = n18956 | n18960 ;
  assign n18962 = ~n18953 & n18961 ;
  assign n18963 = n18948 | n18962 ;
  assign n18965 = ( n18303 & ~n18308 ) | ( n18303 & n18316 ) | ( ~n18308 & n18316 ) ;
  assign n18964 = n18303 | n18532 ;
  assign n18967 = ( n18303 & ~n18965 ) | ( n18303 & n18964 ) | ( ~n18965 & n18964 ) ;
  assign n18966 = ( n18964 & ~n18316 ) | ( n18964 & n18965 ) | ( ~n18316 & n18965 ) ;
  assign n18968 = ( n18308 & ~n18967 ) | ( n18308 & n18966 ) | ( ~n18967 & n18966 ) ;
  assign n18969 = ( n2033 & ~n18963 ) | ( n2033 & n18968 ) | ( ~n18963 & n18968 ) ;
  assign n18970 = ( n1827 & ~n18969 ) | ( n1827 & 1'b0 ) | ( ~n18969 & 1'b0 ) ;
  assign n18971 = n18336 | n18532 ;
  assign n18972 = ( n18323 & ~n18336 ) | ( n18323 & n18332 ) | ( ~n18336 & n18332 ) ;
  assign n18974 = ( n18336 & n18971 ) | ( n18336 & n18972 ) | ( n18971 & n18972 ) ;
  assign n18973 = ( n18332 & ~n18972 ) | ( n18332 & n18971 ) | ( ~n18972 & n18971 ) ;
  assign n18975 = ( n18323 & ~n18974 ) | ( n18323 & n18973 ) | ( ~n18974 & n18973 ) ;
  assign n18976 = ( n2033 & ~n18948 ) | ( n2033 & 1'b0 ) | ( ~n18948 & 1'b0 ) ;
  assign n18977 = ~n18962 & n18976 ;
  assign n18978 = n18968 | n18977 ;
  assign n18979 = n18956 | n18959 ;
  assign n18980 = ( n2245 & ~n18953 ) | ( n2245 & n18979 ) | ( ~n18953 & n18979 ) ;
  assign n18981 = ~n2033 & n18980 ;
  assign n18982 = n1827 | n18981 ;
  assign n18983 = ( n18978 & ~n18982 ) | ( n18978 & 1'b0 ) | ( ~n18982 & 1'b0 ) ;
  assign n18984 = ( n18975 & ~n18983 ) | ( n18975 & 1'b0 ) | ( ~n18983 & 1'b0 ) ;
  assign n18985 = n18970 | n18984 ;
  assign n18987 = ( n18325 & ~n18330 ) | ( n18325 & n18338 ) | ( ~n18330 & n18338 ) ;
  assign n18986 = n18325 | n18532 ;
  assign n18989 = ( n18325 & ~n18987 ) | ( n18325 & n18986 ) | ( ~n18987 & n18986 ) ;
  assign n18988 = ( n18986 & ~n18338 ) | ( n18986 & n18987 ) | ( ~n18338 & n18987 ) ;
  assign n18990 = ( n18330 & ~n18989 ) | ( n18330 & n18988 ) | ( ~n18989 & n18988 ) ;
  assign n18991 = ( n1636 & ~n18985 ) | ( n1636 & n18990 ) | ( ~n18985 & n18990 ) ;
  assign n18992 = n1452 | n18991 ;
  assign n18993 = n18358 | n18532 ;
  assign n18994 = ( n18345 & ~n18358 ) | ( n18345 & n18354 ) | ( ~n18358 & n18354 ) ;
  assign n18996 = ( n18358 & n18993 ) | ( n18358 & n18994 ) | ( n18993 & n18994 ) ;
  assign n18995 = ( n18354 & ~n18994 ) | ( n18354 & n18993 ) | ( ~n18994 & n18993 ) ;
  assign n18997 = ( n18345 & ~n18996 ) | ( n18345 & n18995 ) | ( ~n18996 & n18995 ) ;
  assign n18998 = ( n1636 & ~n18970 ) | ( n1636 & 1'b0 ) | ( ~n18970 & 1'b0 ) ;
  assign n18999 = ~n18984 & n18998 ;
  assign n19000 = n18990 | n18999 ;
  assign n19001 = ( n18978 & ~n18981 ) | ( n18978 & 1'b0 ) | ( ~n18981 & 1'b0 ) ;
  assign n19002 = ( n1827 & ~n19001 ) | ( n1827 & n18975 ) | ( ~n19001 & n18975 ) ;
  assign n19003 = ~n1636 & n19002 ;
  assign n19004 = ( n1452 & ~n19003 ) | ( n1452 & 1'b0 ) | ( ~n19003 & 1'b0 ) ;
  assign n19005 = n19000 &  n19004 ;
  assign n19006 = ( n18997 & ~n19005 ) | ( n18997 & 1'b0 ) | ( ~n19005 & 1'b0 ) ;
  assign n19007 = ( n18992 & ~n19006 ) | ( n18992 & 1'b0 ) | ( ~n19006 & 1'b0 ) ;
  assign n19008 = n18347 | n18532 ;
  assign n19009 = ( n18347 & ~n18360 ) | ( n18347 & n18352 ) | ( ~n18360 & n18352 ) ;
  assign n19010 = ( n18360 & n19008 ) | ( n18360 & n19009 ) | ( n19008 & n19009 ) ;
  assign n19011 = ( n18347 & ~n19009 ) | ( n18347 & n19008 ) | ( ~n19009 & n19008 ) ;
  assign n19012 = ( n18352 & ~n19010 ) | ( n18352 & n19011 ) | ( ~n19010 & n19011 ) ;
  assign n19013 = ( n1283 & ~n19007 ) | ( n1283 & n19012 ) | ( ~n19007 & n19012 ) ;
  assign n19014 = ~n1122 & n19013 ;
  assign n19015 = n18380 | n18532 ;
  assign n19016 = ( n18367 & n18376 ) | ( n18367 & n18380 ) | ( n18376 & n18380 ) ;
  assign n19017 = ( n19015 & ~n18376 ) | ( n19015 & n19016 ) | ( ~n18376 & n19016 ) ;
  assign n19018 = ( n18380 & ~n19016 ) | ( n18380 & n19015 ) | ( ~n19016 & n19015 ) ;
  assign n19019 = ( n18367 & ~n19017 ) | ( n18367 & n19018 ) | ( ~n19017 & n19018 ) ;
  assign n19020 = ~n1283 & n18992 ;
  assign n19021 = ~n19006 & n19020 ;
  assign n19022 = ( n19012 & ~n19021 ) | ( n19012 & 1'b0 ) | ( ~n19021 & 1'b0 ) ;
  assign n19023 = ( n19000 & ~n19003 ) | ( n19000 & 1'b0 ) | ( ~n19003 & 1'b0 ) ;
  assign n19024 = ( n1452 & ~n18997 ) | ( n1452 & n19023 ) | ( ~n18997 & n19023 ) ;
  assign n19025 = ( n1283 & ~n19024 ) | ( n1283 & 1'b0 ) | ( ~n19024 & 1'b0 ) ;
  assign n19026 = ( n1122 & ~n19025 ) | ( n1122 & 1'b0 ) | ( ~n19025 & 1'b0 ) ;
  assign n19027 = ~n19022 & n19026 ;
  assign n19028 = n19019 | n19027 ;
  assign n19029 = ~n19014 & n19028 ;
  assign n19030 = n18369 | n18532 ;
  assign n19031 = ( n18374 & ~n18369 ) | ( n18374 & n18382 ) | ( ~n18369 & n18382 ) ;
  assign n19033 = ( n18369 & n19030 ) | ( n18369 & n19031 ) | ( n19030 & n19031 ) ;
  assign n19032 = ( n18382 & ~n19031 ) | ( n18382 & n19030 ) | ( ~n19031 & n19030 ) ;
  assign n19034 = ( n18374 & ~n19033 ) | ( n18374 & n19032 ) | ( ~n19033 & n19032 ) ;
  assign n19035 = ( n976 & n19029 ) | ( n976 & n19034 ) | ( n19029 & n19034 ) ;
  assign n19036 = ( n837 & ~n19035 ) | ( n837 & 1'b0 ) | ( ~n19035 & 1'b0 ) ;
  assign n19038 = ( n18398 & ~n18389 ) | ( n18398 & n18402 ) | ( ~n18389 & n18402 ) ;
  assign n19037 = ( n18402 & ~n18532 ) | ( n18402 & 1'b0 ) | ( ~n18532 & 1'b0 ) ;
  assign n19040 = ( n18402 & ~n19038 ) | ( n18402 & n19037 ) | ( ~n19038 & n19037 ) ;
  assign n19039 = ( n19037 & ~n18398 ) | ( n19037 & n19038 ) | ( ~n18398 & n19038 ) ;
  assign n19041 = ( n18389 & ~n19040 ) | ( n18389 & n19039 ) | ( ~n19040 & n19039 ) ;
  assign n19042 = ( n976 & ~n19014 ) | ( n976 & 1'b0 ) | ( ~n19014 & 1'b0 ) ;
  assign n19043 = n19028 &  n19042 ;
  assign n19044 = n19034 | n19043 ;
  assign n19045 = n19022 | n19025 ;
  assign n19046 = ( n1122 & ~n19045 ) | ( n1122 & n19019 ) | ( ~n19045 & n19019 ) ;
  assign n19047 = n976 | n19046 ;
  assign n19048 = ~n837 & n19047 ;
  assign n19049 = n19044 &  n19048 ;
  assign n19050 = n19041 | n19049 ;
  assign n19051 = ~n19036 & n19050 ;
  assign n19052 = n18391 | n18532 ;
  assign n19053 = ( n18396 & ~n18391 ) | ( n18396 & n18404 ) | ( ~n18391 & n18404 ) ;
  assign n19055 = ( n18391 & n19052 ) | ( n18391 & n19053 ) | ( n19052 & n19053 ) ;
  assign n19054 = ( n18404 & ~n19053 ) | ( n18404 & n19052 ) | ( ~n19053 & n19052 ) ;
  assign n19056 = ( n18396 & ~n19055 ) | ( n18396 & n19054 ) | ( ~n19055 & n19054 ) ;
  assign n19057 = ( n19051 & ~n713 ) | ( n19051 & n19056 ) | ( ~n713 & n19056 ) ;
  assign n19058 = ( n595 & ~n19057 ) | ( n595 & 1'b0 ) | ( ~n19057 & 1'b0 ) ;
  assign n19059 = n18424 | n18532 ;
  assign n19060 = ( n18411 & ~n18420 ) | ( n18411 & n18424 ) | ( ~n18420 & n18424 ) ;
  assign n19061 = ( n18420 & n19059 ) | ( n18420 & n19060 ) | ( n19059 & n19060 ) ;
  assign n19062 = ( n18424 & ~n19060 ) | ( n18424 & n19059 ) | ( ~n19060 & n19059 ) ;
  assign n19063 = ( n18411 & ~n19061 ) | ( n18411 & n19062 ) | ( ~n19061 & n19062 ) ;
  assign n19064 = n713 | n19036 ;
  assign n19065 = ( n19050 & ~n19064 ) | ( n19050 & 1'b0 ) | ( ~n19064 & 1'b0 ) ;
  assign n19066 = n19056 | n19065 ;
  assign n19067 = n19044 &  n19047 ;
  assign n19068 = ( n19041 & ~n837 ) | ( n19041 & n19067 ) | ( ~n837 & n19067 ) ;
  assign n19069 = ( n713 & ~n19068 ) | ( n713 & 1'b0 ) | ( ~n19068 & 1'b0 ) ;
  assign n19070 = n595 | n19069 ;
  assign n19071 = ( n19066 & ~n19070 ) | ( n19066 & 1'b0 ) | ( ~n19070 & 1'b0 ) ;
  assign n19072 = n19063 | n19071 ;
  assign n19073 = ~n19058 & n19072 ;
  assign n19074 = n18413 | n18532 ;
  assign n19075 = ( n18413 & ~n18426 ) | ( n18413 & n18418 ) | ( ~n18426 & n18418 ) ;
  assign n19076 = ( n18426 & n19074 ) | ( n18426 & n19075 ) | ( n19074 & n19075 ) ;
  assign n19077 = ( n18413 & ~n19075 ) | ( n18413 & n19074 ) | ( ~n19075 & n19074 ) ;
  assign n19078 = ( n18418 & ~n19076 ) | ( n18418 & n19077 ) | ( ~n19076 & n19077 ) ;
  assign n19079 = ( n492 & ~n19073 ) | ( n492 & n19078 ) | ( ~n19073 & n19078 ) ;
  assign n19080 = n396 &  n19079 ;
  assign n19086 = n492 | n19058 ;
  assign n19087 = ( n19072 & ~n19086 ) | ( n19072 & 1'b0 ) | ( ~n19086 & 1'b0 ) ;
  assign n19088 = ( n19078 & ~n19087 ) | ( n19078 & 1'b0 ) | ( ~n19087 & 1'b0 ) ;
  assign n19089 = ( n19066 & ~n19069 ) | ( n19066 & 1'b0 ) | ( ~n19069 & 1'b0 ) ;
  assign n19090 = ( n19063 & ~n595 ) | ( n19063 & n19089 ) | ( ~n595 & n19089 ) ;
  assign n19091 = ( n492 & ~n19090 ) | ( n492 & 1'b0 ) | ( ~n19090 & 1'b0 ) ;
  assign n19092 = n396 | n19091 ;
  assign n19093 = n19088 | n19092 ;
  assign n19747 = ( n19080 & ~n19085 ) | ( n19080 & n19093 ) | ( ~n19085 & n19093 ) ;
  assign n19117 = ~n18469 & n18532 ;
  assign n19118 = ( n18456 & n18461 ) | ( n18456 & n18532 ) | ( n18461 & n18532 ) ;
  assign n19120 = ( n19117 & ~n18456 ) | ( n19117 & n19118 ) | ( ~n18456 & n19118 ) ;
  assign n19119 = ( n18532 & ~n19118 ) | ( n18532 & n19117 ) | ( ~n19118 & n19117 ) ;
  assign n19121 = ( n18461 & ~n19120 ) | ( n18461 & n19119 ) | ( ~n19120 & n19119 ) ;
  assign n19096 = ( n18435 & ~n18447 ) | ( n18435 & n18443 ) | ( ~n18447 & n18443 ) ;
  assign n19097 = ( n18435 & ~n19096 ) | ( n18435 & n18532 ) | ( ~n19096 & n18532 ) ;
  assign n19098 = ( n18532 & ~n18443 ) | ( n18532 & n19096 ) | ( ~n18443 & n19096 ) ;
  assign n19099 = ( n18447 & ~n19097 ) | ( n18447 & n19098 ) | ( ~n19097 & n19098 ) ;
  assign n19094 = ~n19085 & n19093 ;
  assign n19095 = n19080 | n19094 ;
  assign n19100 = ( n315 & ~n19099 ) | ( n315 & n19095 ) | ( ~n19099 & n19095 ) ;
  assign n19101 = n240 &  n19100 ;
  assign n19102 = n18467 | n18532 ;
  assign n19103 = ( n18454 & n18463 ) | ( n18454 & n18467 ) | ( n18463 & n18467 ) ;
  assign n19104 = ( n19102 & ~n18463 ) | ( n19102 & n19103 ) | ( ~n18463 & n19103 ) ;
  assign n19105 = ( n18467 & ~n19103 ) | ( n18467 & n19102 ) | ( ~n19103 & n19102 ) ;
  assign n19106 = ( n18454 & ~n19104 ) | ( n18454 & n19105 ) | ( ~n19104 & n19105 ) ;
  assign n19107 = n315 | n19080 ;
  assign n19108 = n19094 | n19107 ;
  assign n19109 = ~n19099 & n19108 ;
  assign n19110 = n19088 | n19091 ;
  assign n19111 = ( n396 & ~n19085 ) | ( n396 & n19110 ) | ( ~n19085 & n19110 ) ;
  assign n19112 = n315 &  n19111 ;
  assign n19113 = n240 | n19112 ;
  assign n19114 = n19109 | n19113 ;
  assign n19115 = n19106 &  n19114 ;
  assign n19116 = n19101 | n19115 ;
  assign n19122 = ( n181 & ~n19121 ) | ( n181 & n19116 ) | ( ~n19121 & n19116 ) ;
  assign n19123 = ~n145 & n19122 ;
  assign n19125 = ( n18485 & ~n18476 ) | ( n18485 & n18489 ) | ( ~n18476 & n18489 ) ;
  assign n19124 = n18489 | n18532 ;
  assign n19127 = ( n18489 & ~n19125 ) | ( n18489 & n19124 ) | ( ~n19125 & n19124 ) ;
  assign n19126 = ( n19124 & ~n18485 ) | ( n19124 & n19125 ) | ( ~n18485 & n19125 ) ;
  assign n19128 = ( n18476 & ~n19127 ) | ( n18476 & n19126 ) | ( ~n19127 & n19126 ) ;
  assign n19129 = n181 | n19101 ;
  assign n19130 = n19115 | n19129 ;
  assign n19131 = ~n19121 & n19130 ;
  assign n19132 = n19109 | n19112 ;
  assign n19133 = ( n240 & n19106 ) | ( n240 & n19132 ) | ( n19106 & n19132 ) ;
  assign n19134 = n181 &  n19133 ;
  assign n19135 = ( n145 & ~n19134 ) | ( n145 & 1'b0 ) | ( ~n19134 & 1'b0 ) ;
  assign n19136 = ~n19131 & n19135 ;
  assign n19137 = ( n19128 & ~n19136 ) | ( n19128 & 1'b0 ) | ( ~n19136 & 1'b0 ) ;
  assign n19138 = n19123 | n19137 ;
  assign n19139 = n18478 | n18532 ;
  assign n19140 = ( n18483 & ~n18478 ) | ( n18483 & n18491 ) | ( ~n18478 & n18491 ) ;
  assign n19142 = ( n18478 & n19139 ) | ( n18478 & n19140 ) | ( n19139 & n19140 ) ;
  assign n19141 = ( n18491 & ~n19140 ) | ( n18491 & n19139 ) | ( ~n19140 & n19139 ) ;
  assign n19143 = ( n18483 & ~n19142 ) | ( n18483 & n19141 ) | ( ~n19142 & n19141 ) ;
  assign n19144 = ( n150 & n19138 ) | ( n150 & n19143 ) | ( n19138 & n19143 ) ;
  assign n19146 = ( n18514 & ~n18498 ) | ( n18514 & n18517 ) | ( ~n18498 & n18517 ) ;
  assign n19145 = n18517 | n18532 ;
  assign n19148 = ( n18517 & ~n19146 ) | ( n18517 & n19145 ) | ( ~n19146 & n19145 ) ;
  assign n19147 = ( n19145 & ~n18514 ) | ( n19145 & n19146 ) | ( ~n18514 & n19146 ) ;
  assign n19149 = ( n18498 & ~n19148 ) | ( n18498 & n19147 ) | ( ~n19148 & n19147 ) ;
  assign n19150 = n18499 &  n18506 ;
  assign n19151 = ~n18532 & n19150 ;
  assign n19152 = ( n18520 & ~n19150 ) | ( n18520 & n19151 ) | ( ~n19150 & n19151 ) ;
  assign n19153 = ~n19149 & n19152 ;
  assign n19154 = ~n19144 & n19153 ;
  assign n19155 = ( n133 & ~n19154 ) | ( n133 & n19153 ) | ( ~n19154 & n19153 ) ;
  assign n19158 = n19131 | n19134 ;
  assign n19159 = ( n19128 & ~n145 ) | ( n19128 & n19158 ) | ( ~n145 & n19158 ) ;
  assign n19160 = n150 &  n19159 ;
  assign n19161 = ( n19149 & ~n19160 ) | ( n19149 & 1'b0 ) | ( ~n19160 & 1'b0 ) ;
  assign n19156 = n150 | n19123 ;
  assign n19157 = n19137 | n19156 ;
  assign n19162 = ( n19143 & ~n19157 ) | ( n19143 & 1'b0 ) | ( ~n19157 & 1'b0 ) ;
  assign n19163 = ( n19161 & ~n19143 ) | ( n19161 & n19162 ) | ( ~n19143 & n19162 ) ;
  assign n19165 = ( n133 & n18499 ) | ( n133 & n18506 ) | ( n18499 & n18506 ) ;
  assign n19164 = ( n18499 & ~n18532 ) | ( n18499 & n18506 ) | ( ~n18532 & n18506 ) ;
  assign n19166 = ( n18506 & ~n19164 ) | ( n18506 & 1'b0 ) | ( ~n19164 & 1'b0 ) ;
  assign n19167 = ( n19165 & ~n18506 ) | ( n19165 & n19166 ) | ( ~n18506 & n19166 ) ;
  assign n19168 = n18502 | n18529 ;
  assign n19169 = ( n18524 & ~n18505 ) | ( n18524 & n19168 ) | ( ~n18505 & n19168 ) ;
  assign n19170 = n18505 | n19169 ;
  assign n19171 = ( n18512 & ~n18520 ) | ( n18512 & n19170 ) | ( ~n18520 & n19170 ) ;
  assign n19172 = ( n18512 & ~n19171 ) | ( n18512 & 1'b0 ) | ( ~n19171 & 1'b0 ) ;
  assign n19173 = n19167 | n19172 ;
  assign n19174 = n19163 | n19173 ;
  assign n19175 = ~n19155 |  n19174 ;
  assign n19746 = n19080 | n19175 ;
  assign n19749 = ( n19080 & ~n19747 ) | ( n19080 & n19746 ) | ( ~n19747 & n19746 ) ;
  assign n19748 = ( n19746 & ~n19093 ) | ( n19746 & n19747 ) | ( ~n19093 & n19747 ) ;
  assign n19750 = ( n19085 & ~n19749 ) | ( n19085 & n19748 ) | ( ~n19749 & n19748 ) ;
  assign n19724 = n19058 | n19175 ;
  assign n19725 = ( n19063 & ~n19058 ) | ( n19063 & n19071 ) | ( ~n19058 & n19071 ) ;
  assign n19727 = ( n19058 & n19724 ) | ( n19058 & n19725 ) | ( n19724 & n19725 ) ;
  assign n19726 = ( n19071 & ~n19725 ) | ( n19071 & n19724 ) | ( ~n19725 & n19724 ) ;
  assign n19728 = ( n19063 & ~n19727 ) | ( n19063 & n19726 ) | ( ~n19727 & n19726 ) ;
  assign n19709 = n19069 | n19175 ;
  assign n19710 = ( n19056 & ~n19065 ) | ( n19056 & n19069 ) | ( ~n19065 & n19069 ) ;
  assign n19711 = ( n19065 & n19709 ) | ( n19065 & n19710 ) | ( n19709 & n19710 ) ;
  assign n19712 = ( n19069 & ~n19710 ) | ( n19069 & n19709 ) | ( ~n19710 & n19709 ) ;
  assign n19713 = ( n19056 & ~n19711 ) | ( n19056 & n19712 ) | ( ~n19711 & n19712 ) ;
  assign n19702 = n19036 | n19175 ;
  assign n19703 = ( n19041 & ~n19036 ) | ( n19041 & n19049 ) | ( ~n19036 & n19049 ) ;
  assign n19705 = ( n19036 & n19702 ) | ( n19036 & n19703 ) | ( n19702 & n19703 ) ;
  assign n19704 = ( n19049 & ~n19703 ) | ( n19049 & n19702 ) | ( ~n19703 & n19702 ) ;
  assign n19706 = ( n19041 & ~n19705 ) | ( n19041 & n19704 ) | ( ~n19705 & n19704 ) ;
  assign n19688 = ( n19043 & ~n19034 ) | ( n19043 & n19047 ) | ( ~n19034 & n19047 ) ;
  assign n19687 = ( n19047 & ~n19175 ) | ( n19047 & 1'b0 ) | ( ~n19175 & 1'b0 ) ;
  assign n19690 = ( n19047 & ~n19688 ) | ( n19047 & n19687 ) | ( ~n19688 & n19687 ) ;
  assign n19689 = ( n19687 & ~n19043 ) | ( n19687 & n19688 ) | ( ~n19043 & n19688 ) ;
  assign n19691 = ( n19034 & ~n19690 ) | ( n19034 & n19689 ) | ( ~n19690 & n19689 ) ;
  assign n19680 = n19014 | n19175 ;
  assign n19681 = ( n19019 & ~n19014 ) | ( n19019 & n19027 ) | ( ~n19014 & n19027 ) ;
  assign n19683 = ( n19014 & n19680 ) | ( n19014 & n19681 ) | ( n19680 & n19681 ) ;
  assign n19682 = ( n19027 & ~n19681 ) | ( n19027 & n19680 ) | ( ~n19681 & n19680 ) ;
  assign n19684 = ( n19019 & ~n19683 ) | ( n19019 & n19682 ) | ( ~n19683 & n19682 ) ;
  assign n19665 = n19025 | n19175 ;
  assign n19666 = ( n19012 & ~n19025 ) | ( n19012 & n19021 ) | ( ~n19025 & n19021 ) ;
  assign n19668 = ( n19025 & n19665 ) | ( n19025 & n19666 ) | ( n19665 & n19666 ) ;
  assign n19667 = ( n19021 & ~n19666 ) | ( n19021 & n19665 ) | ( ~n19666 & n19665 ) ;
  assign n19669 = ( n19012 & ~n19668 ) | ( n19012 & n19667 ) | ( ~n19668 & n19667 ) ;
  assign n19659 = ( n18992 & ~n18997 ) | ( n18992 & n19005 ) | ( ~n18997 & n19005 ) ;
  assign n19658 = ( n18992 & ~n19175 ) | ( n18992 & 1'b0 ) | ( ~n19175 & 1'b0 ) ;
  assign n19661 = ( n18992 & ~n19659 ) | ( n18992 & n19658 ) | ( ~n19659 & n19658 ) ;
  assign n19660 = ( n19658 & ~n19005 ) | ( n19658 & n19659 ) | ( ~n19005 & n19659 ) ;
  assign n19662 = ( n18997 & ~n19661 ) | ( n18997 & n19660 ) | ( ~n19661 & n19660 ) ;
  assign n19643 = n19003 | n19175 ;
  assign n19644 = ( n18990 & ~n18999 ) | ( n18990 & n19003 ) | ( ~n18999 & n19003 ) ;
  assign n19645 = ( n18999 & n19643 ) | ( n18999 & n19644 ) | ( n19643 & n19644 ) ;
  assign n19646 = ( n19003 & ~n19644 ) | ( n19003 & n19643 ) | ( ~n19644 & n19643 ) ;
  assign n19647 = ( n18990 & ~n19645 ) | ( n18990 & n19646 ) | ( ~n19645 & n19646 ) ;
  assign n19636 = n18970 | n19175 ;
  assign n19637 = ( n18970 & ~n18983 ) | ( n18970 & n18975 ) | ( ~n18983 & n18975 ) ;
  assign n19638 = ( n18983 & n19636 ) | ( n18983 & n19637 ) | ( n19636 & n19637 ) ;
  assign n19639 = ( n18970 & ~n19637 ) | ( n18970 & n19636 ) | ( ~n19637 & n19636 ) ;
  assign n19640 = ( n18975 & ~n19638 ) | ( n18975 & n19639 ) | ( ~n19638 & n19639 ) ;
  assign n19621 = n18981 | n19175 ;
  assign n19622 = ( n18968 & ~n18977 ) | ( n18968 & n18981 ) | ( ~n18977 & n18981 ) ;
  assign n19623 = ( n18977 & n19621 ) | ( n18977 & n19622 ) | ( n19621 & n19622 ) ;
  assign n19624 = ( n18981 & ~n19622 ) | ( n18981 & n19621 ) | ( ~n19622 & n19621 ) ;
  assign n19625 = ( n18968 & ~n19623 ) | ( n18968 & n19624 ) | ( ~n19623 & n19624 ) ;
  assign n19615 = ( n18948 & ~n18953 ) | ( n18948 & n18961 ) | ( ~n18953 & n18961 ) ;
  assign n19614 = n18948 | n19175 ;
  assign n19617 = ( n18948 & ~n19615 ) | ( n18948 & n19614 ) | ( ~n19615 & n19614 ) ;
  assign n19616 = ( n19614 & ~n18961 ) | ( n19614 & n19615 ) | ( ~n18961 & n19615 ) ;
  assign n19618 = ( n18953 & ~n19617 ) | ( n18953 & n19616 ) | ( ~n19617 & n19616 ) ;
  assign n19600 = ( n18955 & ~n18946 ) | ( n18955 & n18959 ) | ( ~n18946 & n18959 ) ;
  assign n19599 = n18959 | n19175 ;
  assign n19602 = ( n18959 & ~n19600 ) | ( n18959 & n19599 ) | ( ~n19600 & n19599 ) ;
  assign n19601 = ( n19599 & ~n18955 ) | ( n19599 & n19600 ) | ( ~n18955 & n19600 ) ;
  assign n19603 = ( n18946 & ~n19602 ) | ( n18946 & n19601 ) | ( ~n19602 & n19601 ) ;
  assign n19592 = n18926 | n19175 ;
  assign n19593 = ( n18926 & n18931 ) | ( n18926 & n18939 ) | ( n18931 & n18939 ) ;
  assign n19594 = ( n19592 & ~n18939 ) | ( n19592 & n19593 ) | ( ~n18939 & n19593 ) ;
  assign n19595 = ( n18926 & ~n19593 ) | ( n18926 & n19592 ) | ( ~n19593 & n19592 ) ;
  assign n19596 = ( n18931 & ~n19594 ) | ( n18931 & n19595 ) | ( ~n19594 & n19595 ) ;
  assign n19578 = ( n18933 & ~n18924 ) | ( n18933 & n18937 ) | ( ~n18924 & n18937 ) ;
  assign n19577 = n18937 | n19175 ;
  assign n19580 = ( n18937 & ~n19578 ) | ( n18937 & n19577 ) | ( ~n19578 & n19577 ) ;
  assign n19579 = ( n19577 & ~n18933 ) | ( n19577 & n19578 ) | ( ~n18933 & n19578 ) ;
  assign n19581 = ( n18924 & ~n19580 ) | ( n18924 & n19579 ) | ( ~n19580 & n19579 ) ;
  assign n19570 = n18904 | n19175 ;
  assign n19571 = ( n18904 & n18909 ) | ( n18904 & n18917 ) | ( n18909 & n18917 ) ;
  assign n19572 = ( n19570 & ~n18917 ) | ( n19570 & n19571 ) | ( ~n18917 & n19571 ) ;
  assign n19573 = ( n18904 & ~n19571 ) | ( n18904 & n19570 ) | ( ~n19571 & n19570 ) ;
  assign n19574 = ( n18909 & ~n19572 ) | ( n18909 & n19573 ) | ( ~n19572 & n19573 ) ;
  assign n19555 = n18915 | n19175 ;
  assign n19556 = ( n18902 & ~n18915 ) | ( n18902 & n18911 ) | ( ~n18915 & n18911 ) ;
  assign n19558 = ( n18915 & n19555 ) | ( n18915 & n19556 ) | ( n19555 & n19556 ) ;
  assign n19557 = ( n18911 & ~n19556 ) | ( n18911 & n19555 ) | ( ~n19556 & n19555 ) ;
  assign n19559 = ( n18902 & ~n19558 ) | ( n18902 & n19557 ) | ( ~n19558 & n19557 ) ;
  assign n19548 = n18882 | n19175 ;
  assign n19549 = ( n18887 & ~n18882 ) | ( n18887 & n18895 ) | ( ~n18882 & n18895 ) ;
  assign n19551 = ( n18882 & n19548 ) | ( n18882 & n19549 ) | ( n19548 & n19549 ) ;
  assign n19550 = ( n18895 & ~n19549 ) | ( n18895 & n19548 ) | ( ~n19549 & n19548 ) ;
  assign n19552 = ( n18887 & ~n19551 ) | ( n18887 & n19550 ) | ( ~n19551 & n19550 ) ;
  assign n19533 = n18893 | n19175 ;
  assign n19534 = ( n18880 & ~n18889 ) | ( n18880 & n18893 ) | ( ~n18889 & n18893 ) ;
  assign n19535 = ( n18889 & n19533 ) | ( n18889 & n19534 ) | ( n19533 & n19534 ) ;
  assign n19536 = ( n18893 & ~n19534 ) | ( n18893 & n19533 ) | ( ~n19534 & n19533 ) ;
  assign n19537 = ( n18880 & ~n19535 ) | ( n18880 & n19536 ) | ( ~n19535 & n19536 ) ;
  assign n19526 = n18860 | n19175 ;
  assign n19527 = ( n18865 & ~n18860 ) | ( n18865 & n18873 ) | ( ~n18860 & n18873 ) ;
  assign n19529 = ( n18860 & n19526 ) | ( n18860 & n19527 ) | ( n19526 & n19527 ) ;
  assign n19528 = ( n18873 & ~n19527 ) | ( n18873 & n19526 ) | ( ~n19527 & n19526 ) ;
  assign n19530 = ( n18865 & ~n19529 ) | ( n18865 & n19528 ) | ( ~n19529 & n19528 ) ;
  assign n19511 = n18871 | n19175 ;
  assign n19512 = ( n18858 & ~n18867 ) | ( n18858 & n18871 ) | ( ~n18867 & n18871 ) ;
  assign n19513 = ( n18867 & n19511 ) | ( n18867 & n19512 ) | ( n19511 & n19512 ) ;
  assign n19514 = ( n18871 & ~n19512 ) | ( n18871 & n19511 ) | ( ~n19512 & n19511 ) ;
  assign n19515 = ( n18858 & ~n19513 ) | ( n18858 & n19514 ) | ( ~n19513 & n19514 ) ;
  assign n19504 = n18838 | n19175 ;
  assign n19505 = ( n18843 & ~n18838 ) | ( n18843 & n18851 ) | ( ~n18838 & n18851 ) ;
  assign n19507 = ( n18838 & n19504 ) | ( n18838 & n19505 ) | ( n19504 & n19505 ) ;
  assign n19506 = ( n18851 & ~n19505 ) | ( n18851 & n19504 ) | ( ~n19505 & n19504 ) ;
  assign n19508 = ( n18843 & ~n19507 ) | ( n18843 & n19506 ) | ( ~n19507 & n19506 ) ;
  assign n19489 = n18849 | n19175 ;
  assign n19490 = ( n18836 & ~n18845 ) | ( n18836 & n18849 ) | ( ~n18845 & n18849 ) ;
  assign n19491 = ( n18845 & n19489 ) | ( n18845 & n19490 ) | ( n19489 & n19490 ) ;
  assign n19492 = ( n18849 & ~n19490 ) | ( n18849 & n19489 ) | ( ~n19490 & n19489 ) ;
  assign n19493 = ( n18836 & ~n19491 ) | ( n18836 & n19492 ) | ( ~n19491 & n19492 ) ;
  assign n19482 = ( n18816 & ~n19175 ) | ( n18816 & 1'b0 ) | ( ~n19175 & 1'b0 ) ;
  assign n19483 = ( n18816 & n18821 ) | ( n18816 & n18829 ) | ( n18821 & n18829 ) ;
  assign n19484 = ( n19482 & ~n18829 ) | ( n19482 & n19483 ) | ( ~n18829 & n19483 ) ;
  assign n19485 = ( n18816 & ~n19483 ) | ( n18816 & n19482 ) | ( ~n19483 & n19482 ) ;
  assign n19486 = ( n18821 & ~n19484 ) | ( n18821 & n19485 ) | ( ~n19484 & n19485 ) ;
  assign n19467 = n18827 | n19175 ;
  assign n19468 = ( n18814 & ~n18823 ) | ( n18814 & n18827 ) | ( ~n18823 & n18827 ) ;
  assign n19469 = ( n18823 & n19467 ) | ( n18823 & n19468 ) | ( n19467 & n19468 ) ;
  assign n19470 = ( n18827 & ~n19468 ) | ( n18827 & n19467 ) | ( ~n19468 & n19467 ) ;
  assign n19471 = ( n18814 & ~n19469 ) | ( n18814 & n19470 ) | ( ~n19469 & n19470 ) ;
  assign n19460 = ( n18794 & ~n19175 ) | ( n18794 & 1'b0 ) | ( ~n19175 & 1'b0 ) ;
  assign n19461 = ( n18794 & n18799 ) | ( n18794 & n18807 ) | ( n18799 & n18807 ) ;
  assign n19462 = ( n19460 & ~n18807 ) | ( n19460 & n19461 ) | ( ~n18807 & n19461 ) ;
  assign n19463 = ( n18794 & ~n19461 ) | ( n18794 & n19460 ) | ( ~n19461 & n19460 ) ;
  assign n19464 = ( n18799 & ~n19462 ) | ( n18799 & n19463 ) | ( ~n19462 & n19463 ) ;
  assign n19445 = n18805 | n19175 ;
  assign n19446 = ( n18792 & ~n18801 ) | ( n18792 & n18805 ) | ( ~n18801 & n18805 ) ;
  assign n19447 = ( n18801 & n19445 ) | ( n18801 & n19446 ) | ( n19445 & n19446 ) ;
  assign n19448 = ( n18805 & ~n19446 ) | ( n18805 & n19445 ) | ( ~n19446 & n19445 ) ;
  assign n19449 = ( n18792 & ~n19447 ) | ( n18792 & n19448 ) | ( ~n19447 & n19448 ) ;
  assign n19438 = ( n18772 & ~n19175 ) | ( n18772 & 1'b0 ) | ( ~n19175 & 1'b0 ) ;
  assign n19439 = ( n18772 & n18777 ) | ( n18772 & n18785 ) | ( n18777 & n18785 ) ;
  assign n19440 = ( n19438 & ~n18785 ) | ( n19438 & n19439 ) | ( ~n18785 & n19439 ) ;
  assign n19441 = ( n18772 & ~n19439 ) | ( n18772 & n19438 ) | ( ~n19439 & n19438 ) ;
  assign n19442 = ( n18777 & ~n19440 ) | ( n18777 & n19441 ) | ( ~n19440 & n19441 ) ;
  assign n19424 = ( n18779 & ~n18770 ) | ( n18779 & n18783 ) | ( ~n18770 & n18783 ) ;
  assign n19423 = ( n18783 & ~n19175 ) | ( n18783 & 1'b0 ) | ( ~n19175 & 1'b0 ) ;
  assign n19426 = ( n18783 & ~n19424 ) | ( n18783 & n19423 ) | ( ~n19424 & n19423 ) ;
  assign n19425 = ( n19423 & ~n18779 ) | ( n19423 & n19424 ) | ( ~n18779 & n19424 ) ;
  assign n19427 = ( n18770 & ~n19426 ) | ( n18770 & n19425 ) | ( ~n19426 & n19425 ) ;
  assign n19416 = n18750 | n19175 ;
  assign n19417 = ( n18755 & ~n18750 ) | ( n18755 & n18763 ) | ( ~n18750 & n18763 ) ;
  assign n19419 = ( n18750 & n19416 ) | ( n18750 & n19417 ) | ( n19416 & n19417 ) ;
  assign n19418 = ( n18763 & ~n19417 ) | ( n18763 & n19416 ) | ( ~n19417 & n19416 ) ;
  assign n19420 = ( n18755 & ~n19419 ) | ( n18755 & n19418 ) | ( ~n19419 & n19418 ) ;
  assign n19401 = n18761 | n19175 ;
  assign n19402 = ( n18748 & ~n18761 ) | ( n18748 & n18757 ) | ( ~n18761 & n18757 ) ;
  assign n19404 = ( n18761 & n19401 ) | ( n18761 & n19402 ) | ( n19401 & n19402 ) ;
  assign n19403 = ( n18757 & ~n19402 ) | ( n18757 & n19401 ) | ( ~n19402 & n19401 ) ;
  assign n19405 = ( n18748 & ~n19404 ) | ( n18748 & n19403 ) | ( ~n19404 & n19403 ) ;
  assign n19394 = n18728 | n19175 ;
  assign n19395 = ( n18728 & ~n18741 ) | ( n18728 & n18733 ) | ( ~n18741 & n18733 ) ;
  assign n19396 = ( n18741 & n19394 ) | ( n18741 & n19395 ) | ( n19394 & n19395 ) ;
  assign n19397 = ( n18728 & ~n19395 ) | ( n18728 & n19394 ) | ( ~n19395 & n19394 ) ;
  assign n19398 = ( n18733 & ~n19396 ) | ( n18733 & n19397 ) | ( ~n19396 & n19397 ) ;
  assign n19379 = n18739 | n19175 ;
  assign n19380 = ( n18726 & ~n18735 ) | ( n18726 & n18739 ) | ( ~n18735 & n18739 ) ;
  assign n19381 = ( n18735 & n19379 ) | ( n18735 & n19380 ) | ( n19379 & n19380 ) ;
  assign n19382 = ( n18739 & ~n19380 ) | ( n18739 & n19379 ) | ( ~n19380 & n19379 ) ;
  assign n19383 = ( n18726 & ~n19381 ) | ( n18726 & n19382 ) | ( ~n19381 & n19382 ) ;
  assign n19372 = ( n18706 & ~n19175 ) | ( n18706 & 1'b0 ) | ( ~n19175 & 1'b0 ) ;
  assign n19373 = ( n18706 & n18711 ) | ( n18706 & n18719 ) | ( n18711 & n18719 ) ;
  assign n19374 = ( n19372 & ~n18719 ) | ( n19372 & n19373 ) | ( ~n18719 & n19373 ) ;
  assign n19375 = ( n18706 & ~n19373 ) | ( n18706 & n19372 ) | ( ~n19373 & n19372 ) ;
  assign n19376 = ( n18711 & ~n19374 ) | ( n18711 & n19375 ) | ( ~n19374 & n19375 ) ;
  assign n19357 = n18717 | n19175 ;
  assign n19358 = ( n18704 & ~n18713 ) | ( n18704 & n18717 ) | ( ~n18713 & n18717 ) ;
  assign n19359 = ( n18713 & n19357 ) | ( n18713 & n19358 ) | ( n19357 & n19358 ) ;
  assign n19360 = ( n18717 & ~n19358 ) | ( n18717 & n19357 ) | ( ~n19358 & n19357 ) ;
  assign n19361 = ( n18704 & ~n19359 ) | ( n18704 & n19360 ) | ( ~n19359 & n19360 ) ;
  assign n19350 = n18697 &  n19175 ;
  assign n19351 = ( n18684 & n18689 ) | ( n18684 & n19175 ) | ( n18689 & n19175 ) ;
  assign n19353 = ( n19350 & ~n18684 ) | ( n19350 & n19351 ) | ( ~n18684 & n19351 ) ;
  assign n19352 = ( n19175 & ~n19351 ) | ( n19175 & n19350 ) | ( ~n19351 & n19350 ) ;
  assign n19354 = ( n18689 & ~n19353 ) | ( n18689 & n19352 ) | ( ~n19353 & n19352 ) ;
  assign n19335 = n18695 | n19175 ;
  assign n19336 = ( n18682 & ~n18695 ) | ( n18682 & n18691 ) | ( ~n18695 & n18691 ) ;
  assign n19338 = ( n18695 & n19335 ) | ( n18695 & n19336 ) | ( n19335 & n19336 ) ;
  assign n19337 = ( n18691 & ~n19336 ) | ( n18691 & n19335 ) | ( ~n19336 & n19335 ) ;
  assign n19339 = ( n18682 & ~n19338 ) | ( n18682 & n19337 ) | ( ~n19338 & n19337 ) ;
  assign n19328 = n18662 | n19175 ;
  assign n19329 = ( n18662 & ~n18675 ) | ( n18662 & n18667 ) | ( ~n18675 & n18667 ) ;
  assign n19330 = ( n18675 & n19328 ) | ( n18675 & n19329 ) | ( n19328 & n19329 ) ;
  assign n19331 = ( n18662 & ~n19329 ) | ( n18662 & n19328 ) | ( ~n19329 & n19328 ) ;
  assign n19332 = ( n18667 & ~n19330 ) | ( n18667 & n19331 ) | ( ~n19330 & n19331 ) ;
  assign n19313 = n18673 | n19175 ;
  assign n19314 = ( n18660 & ~n18669 ) | ( n18660 & n18673 ) | ( ~n18669 & n18673 ) ;
  assign n19315 = ( n18669 & n19313 ) | ( n18669 & n19314 ) | ( n19313 & n19314 ) ;
  assign n19316 = ( n18673 & ~n19314 ) | ( n18673 & n19313 ) | ( ~n19314 & n19313 ) ;
  assign n19317 = ( n18660 & ~n19315 ) | ( n18660 & n19316 ) | ( ~n19315 & n19316 ) ;
  assign n19306 = n18640 | n19175 ;
  assign n19307 = ( n18645 & ~n18640 ) | ( n18645 & n18653 ) | ( ~n18640 & n18653 ) ;
  assign n19309 = ( n18640 & n19306 ) | ( n18640 & n19307 ) | ( n19306 & n19307 ) ;
  assign n19308 = ( n18653 & ~n19307 ) | ( n18653 & n19306 ) | ( ~n19307 & n19306 ) ;
  assign n19310 = ( n18645 & ~n19309 ) | ( n18645 & n19308 ) | ( ~n19309 & n19308 ) ;
  assign n19291 = n18651 | n19175 ;
  assign n19292 = ( n18638 & ~n18647 ) | ( n18638 & n18651 ) | ( ~n18647 & n18651 ) ;
  assign n19293 = ( n18647 & n19291 ) | ( n18647 & n19292 ) | ( n19291 & n19292 ) ;
  assign n19294 = ( n18651 & ~n19292 ) | ( n18651 & n19291 ) | ( ~n19292 & n19291 ) ;
  assign n19295 = ( n18638 & ~n19293 ) | ( n18638 & n19294 ) | ( ~n19293 & n19294 ) ;
  assign n19284 = n18631 &  n19175 ;
  assign n19285 = ( n18618 & n18623 ) | ( n18618 & n19175 ) | ( n18623 & n19175 ) ;
  assign n19287 = ( n19284 & ~n18618 ) | ( n19284 & n19285 ) | ( ~n18618 & n19285 ) ;
  assign n19286 = ( n19175 & ~n19285 ) | ( n19175 & n19284 ) | ( ~n19285 & n19284 ) ;
  assign n19288 = ( n18623 & ~n19287 ) | ( n18623 & n19286 ) | ( ~n19287 & n19286 ) ;
  assign n19269 = n18629 | n19175 ;
  assign n19270 = ( n18616 & ~n18629 ) | ( n18616 & n18625 ) | ( ~n18629 & n18625 ) ;
  assign n19272 = ( n18629 & n19269 ) | ( n18629 & n19270 ) | ( n19269 & n19270 ) ;
  assign n19271 = ( n18625 & ~n19270 ) | ( n18625 & n19269 ) | ( ~n19270 & n19269 ) ;
  assign n19273 = ( n18616 & ~n19272 ) | ( n18616 & n19271 ) | ( ~n19272 & n19271 ) ;
  assign n19262 = n18596 | n19175 ;
  assign n19263 = ( n18596 & ~n18609 ) | ( n18596 & n18601 ) | ( ~n18609 & n18601 ) ;
  assign n19264 = ( n18609 & n19262 ) | ( n18609 & n19263 ) | ( n19262 & n19263 ) ;
  assign n19265 = ( n18596 & ~n19263 ) | ( n18596 & n19262 ) | ( ~n19263 & n19262 ) ;
  assign n19266 = ( n18601 & ~n19264 ) | ( n18601 & n19265 ) | ( ~n19264 & n19265 ) ;
  assign n19247 = n18607 | n19175 ;
  assign n19248 = ( n18594 & ~n18603 ) | ( n18594 & n18607 ) | ( ~n18603 & n18607 ) ;
  assign n19249 = ( n18603 & n19247 ) | ( n18603 & n19248 ) | ( n19247 & n19248 ) ;
  assign n19250 = ( n18607 & ~n19248 ) | ( n18607 & n19247 ) | ( ~n19248 & n19247 ) ;
  assign n19251 = ( n18594 & ~n19249 ) | ( n18594 & n19250 ) | ( ~n19249 & n19250 ) ;
  assign n19240 = n18574 | n19175 ;
  assign n19241 = ( n18579 & ~n18574 ) | ( n18579 & n18587 ) | ( ~n18574 & n18587 ) ;
  assign n19243 = ( n18574 & n19240 ) | ( n18574 & n19241 ) | ( n19240 & n19241 ) ;
  assign n19242 = ( n18587 & ~n19241 ) | ( n18587 & n19240 ) | ( ~n19241 & n19240 ) ;
  assign n19244 = ( n18579 & ~n19243 ) | ( n18579 & n19242 ) | ( ~n19243 & n19242 ) ;
  assign n19225 = n18585 | n19175 ;
  assign n19226 = ( n18572 & ~n18581 ) | ( n18572 & n18585 ) | ( ~n18581 & n18585 ) ;
  assign n19227 = ( n18581 & n19225 ) | ( n18581 & n19226 ) | ( n19225 & n19226 ) ;
  assign n19228 = ( n18585 & ~n19226 ) | ( n18585 & n19225 ) | ( ~n19226 & n19225 ) ;
  assign n19229 = ( n18572 & ~n19227 ) | ( n18572 & n19228 ) | ( ~n19227 & n19228 ) ;
  assign n19218 = ( n18548 & ~n18550 ) | ( n18548 & 1'b0 ) | ( ~n18550 & 1'b0 ) ;
  assign n19219 = ( n18550 & ~n19218 ) | ( n18550 & n18560 ) | ( ~n19218 & n18560 ) ;
  assign n19221 = ( n19175 & n19218 ) | ( n19175 & n19219 ) | ( n19218 & n19219 ) ;
  assign n19220 = ( n18550 & ~n19219 ) | ( n18550 & n19175 ) | ( ~n19219 & n19175 ) ;
  assign n19222 = ( n18560 & ~n19221 ) | ( n18560 & n19220 ) | ( ~n19221 & n19220 ) ;
  assign n19202 = ~x14 & n18532 ;
  assign n19203 = ( x15 & ~n19202 ) | ( x15 & 1'b0 ) | ( ~n19202 & 1'b0 ) ;
  assign n19204 = n18551 | n19203 ;
  assign n19199 = ( n18532 & ~x14 ) | ( n18532 & n18543 ) | ( ~x14 & n18543 ) ;
  assign n19200 = x14 &  n19199 ;
  assign n19201 = ( n18538 & ~n19200 ) | ( n18538 & n18543 ) | ( ~n19200 & n18543 ) ;
  assign n19205 = ( n19175 & ~n19204 ) | ( n19175 & n19201 ) | ( ~n19204 & n19201 ) ;
  assign n19207 = ( n19175 & ~n19205 ) | ( n19175 & 1'b0 ) | ( ~n19205 & 1'b0 ) ;
  assign n19206 = ~n19201 & n19205 ;
  assign n19208 = ( n19204 & ~n19207 ) | ( n19204 & n19206 ) | ( ~n19207 & n19206 ) ;
  assign n19188 = ( n18532 & ~n19172 ) | ( n18532 & 1'b0 ) | ( ~n19172 & 1'b0 ) ;
  assign n19189 = ( n19163 & ~n19167 ) | ( n19163 & n19188 ) | ( ~n19167 & n19188 ) ;
  assign n19190 = ~n19163 & n19189 ;
  assign n19191 = n19155 &  n19190 ;
  assign n19187 = ~n18535 & n19175 ;
  assign n19192 = ( n19187 & ~n19191 ) | ( n19187 & 1'b0 ) | ( ~n19191 & 1'b0 ) ;
  assign n19193 = ( x14 & n19191 ) | ( x14 & n19192 ) | ( n19191 & n19192 ) ;
  assign n19194 = x14 | n19191 ;
  assign n19195 = n19187 | n19194 ;
  assign n19196 = ~n19193 & n19195 ;
  assign n19178 = ( x12 & ~n19175 ) | ( x12 & x13 ) | ( ~n19175 & x13 ) ;
  assign n19184 = ( x12 & ~x13 ) | ( x12 & 1'b0 ) | ( ~x13 & 1'b0 ) ;
  assign n18533 = x10 | x11 ;
  assign n19179 = ~x12 & n18533 ;
  assign n19180 = ( x12 & ~n18530 ) | ( x12 & n19179 ) | ( ~n18530 & n19179 ) ;
  assign n19181 = ( n18520 & ~n18512 ) | ( n18520 & n19180 ) | ( ~n18512 & n19180 ) ;
  assign n19182 = n18512 &  n19181 ;
  assign n19183 = ( n19175 & ~x13 ) | ( n19175 & n19182 ) | ( ~x13 & n19182 ) ;
  assign n19185 = ( n19178 & ~n19184 ) | ( n19178 & n19183 ) | ( ~n19184 & n19183 ) ;
  assign n18534 = x12 | n18533 ;
  assign n19176 = x12 &  n19175 ;
  assign n19177 = ( n18532 & ~n18534 ) | ( n18532 & n19176 ) | ( ~n18534 & n19176 ) ;
  assign n19209 = n17902 | n19177 ;
  assign n19210 = ( n19185 & ~n19209 ) | ( n19185 & 1'b0 ) | ( ~n19209 & 1'b0 ) ;
  assign n19211 = n19196 | n19210 ;
  assign n19212 = n19177 &  n19185 ;
  assign n19213 = ( n17902 & ~n19185 ) | ( n17902 & n19212 ) | ( ~n19185 & n19212 ) ;
  assign n19214 = n17279 | n19213 ;
  assign n19215 = ( n19211 & ~n19214 ) | ( n19211 & 1'b0 ) | ( ~n19214 & 1'b0 ) ;
  assign n19216 = n19208 | n19215 ;
  assign n19186 = ~n19177 & n19185 ;
  assign n19197 = ( n19186 & ~n17902 ) | ( n19186 & n19196 ) | ( ~n17902 & n19196 ) ;
  assign n19198 = ( n17279 & ~n19197 ) | ( n17279 & 1'b0 ) | ( ~n19197 & 1'b0 ) ;
  assign n19230 = n16671 | n19198 ;
  assign n19231 = ( n19216 & ~n19230 ) | ( n19216 & 1'b0 ) | ( ~n19230 & 1'b0 ) ;
  assign n19232 = n19222 | n19231 ;
  assign n19233 = ( n19211 & ~n19213 ) | ( n19211 & 1'b0 ) | ( ~n19213 & 1'b0 ) ;
  assign n19234 = ( n19208 & ~n17279 ) | ( n19208 & n19233 ) | ( ~n17279 & n19233 ) ;
  assign n19235 = ( n16671 & ~n19234 ) | ( n16671 & 1'b0 ) | ( ~n19234 & 1'b0 ) ;
  assign n19236 = n16070 | n19235 ;
  assign n19237 = ( n19232 & ~n19236 ) | ( n19232 & 1'b0 ) | ( ~n19236 & 1'b0 ) ;
  assign n19238 = n19229 | n19237 ;
  assign n19217 = ~n19198 & n19216 ;
  assign n19223 = ( n19217 & ~n16671 ) | ( n19217 & n19222 ) | ( ~n16671 & n19222 ) ;
  assign n19224 = ( n16070 & ~n19223 ) | ( n16070 & 1'b0 ) | ( ~n19223 & 1'b0 ) ;
  assign n19252 = n15484 | n19224 ;
  assign n19253 = ( n19238 & ~n19252 ) | ( n19238 & 1'b0 ) | ( ~n19252 & 1'b0 ) ;
  assign n19254 = n19244 | n19253 ;
  assign n19255 = ( n19232 & ~n19235 ) | ( n19232 & 1'b0 ) | ( ~n19235 & 1'b0 ) ;
  assign n19256 = ( n19229 & ~n16070 ) | ( n19229 & n19255 ) | ( ~n16070 & n19255 ) ;
  assign n19257 = ( n15484 & ~n19256 ) | ( n15484 & 1'b0 ) | ( ~n19256 & 1'b0 ) ;
  assign n19258 = n14905 | n19257 ;
  assign n19259 = ( n19254 & ~n19258 ) | ( n19254 & 1'b0 ) | ( ~n19258 & 1'b0 ) ;
  assign n19260 = n19251 | n19259 ;
  assign n19239 = ~n19224 & n19238 ;
  assign n19245 = ( n19239 & ~n15484 ) | ( n19239 & n19244 ) | ( ~n15484 & n19244 ) ;
  assign n19246 = ( n14905 & ~n19245 ) | ( n14905 & 1'b0 ) | ( ~n19245 & 1'b0 ) ;
  assign n19274 = n14341 | n19246 ;
  assign n19275 = ( n19260 & ~n19274 ) | ( n19260 & 1'b0 ) | ( ~n19274 & 1'b0 ) ;
  assign n19276 = n19266 | n19275 ;
  assign n19277 = ( n19254 & ~n19257 ) | ( n19254 & 1'b0 ) | ( ~n19257 & 1'b0 ) ;
  assign n19278 = ( n19251 & ~n14905 ) | ( n19251 & n19277 ) | ( ~n14905 & n19277 ) ;
  assign n19279 = ( n14341 & ~n19278 ) | ( n14341 & 1'b0 ) | ( ~n19278 & 1'b0 ) ;
  assign n19280 = n13784 | n19279 ;
  assign n19281 = ( n19276 & ~n19280 ) | ( n19276 & 1'b0 ) | ( ~n19280 & 1'b0 ) ;
  assign n19282 = n19273 | n19281 ;
  assign n19261 = ~n19246 & n19260 ;
  assign n19267 = ( n19261 & ~n14341 ) | ( n19261 & n19266 ) | ( ~n14341 & n19266 ) ;
  assign n19268 = ( n13784 & ~n19267 ) | ( n13784 & 1'b0 ) | ( ~n19267 & 1'b0 ) ;
  assign n19296 = n13242 | n19268 ;
  assign n19297 = ( n19282 & ~n19296 ) | ( n19282 & 1'b0 ) | ( ~n19296 & 1'b0 ) ;
  assign n19298 = n19288 | n19297 ;
  assign n19299 = ( n19276 & ~n19279 ) | ( n19276 & 1'b0 ) | ( ~n19279 & 1'b0 ) ;
  assign n19300 = ( n19273 & ~n13784 ) | ( n19273 & n19299 ) | ( ~n13784 & n19299 ) ;
  assign n19301 = ( n13242 & ~n19300 ) | ( n13242 & 1'b0 ) | ( ~n19300 & 1'b0 ) ;
  assign n19302 = n12707 | n19301 ;
  assign n19303 = ( n19298 & ~n19302 ) | ( n19298 & 1'b0 ) | ( ~n19302 & 1'b0 ) ;
  assign n19304 = n19295 | n19303 ;
  assign n19283 = ~n19268 & n19282 ;
  assign n19289 = ( n19283 & ~n13242 ) | ( n19283 & n19288 ) | ( ~n13242 & n19288 ) ;
  assign n19290 = ( n12707 & ~n19289 ) | ( n12707 & 1'b0 ) | ( ~n19289 & 1'b0 ) ;
  assign n19318 = n12187 | n19290 ;
  assign n19319 = ( n19304 & ~n19318 ) | ( n19304 & 1'b0 ) | ( ~n19318 & 1'b0 ) ;
  assign n19320 = n19310 | n19319 ;
  assign n19321 = ( n19298 & ~n19301 ) | ( n19298 & 1'b0 ) | ( ~n19301 & 1'b0 ) ;
  assign n19322 = ( n19295 & ~n12707 ) | ( n19295 & n19321 ) | ( ~n12707 & n19321 ) ;
  assign n19323 = ( n12187 & ~n19322 ) | ( n12187 & 1'b0 ) | ( ~n19322 & 1'b0 ) ;
  assign n19324 = n11674 | n19323 ;
  assign n19325 = ( n19320 & ~n19324 ) | ( n19320 & 1'b0 ) | ( ~n19324 & 1'b0 ) ;
  assign n19326 = n19317 | n19325 ;
  assign n19305 = ~n19290 & n19304 ;
  assign n19311 = ( n19305 & ~n12187 ) | ( n19305 & n19310 ) | ( ~n12187 & n19310 ) ;
  assign n19312 = ( n11674 & ~n19311 ) | ( n11674 & 1'b0 ) | ( ~n19311 & 1'b0 ) ;
  assign n19340 = n11176 | n19312 ;
  assign n19341 = ( n19326 & ~n19340 ) | ( n19326 & 1'b0 ) | ( ~n19340 & 1'b0 ) ;
  assign n19342 = n19332 | n19341 ;
  assign n19343 = ( n19320 & ~n19323 ) | ( n19320 & 1'b0 ) | ( ~n19323 & 1'b0 ) ;
  assign n19344 = ( n19317 & ~n11674 ) | ( n19317 & n19343 ) | ( ~n11674 & n19343 ) ;
  assign n19345 = ( n11176 & ~n19344 ) | ( n11176 & 1'b0 ) | ( ~n19344 & 1'b0 ) ;
  assign n19346 = n10685 | n19345 ;
  assign n19347 = ( n19342 & ~n19346 ) | ( n19342 & 1'b0 ) | ( ~n19346 & 1'b0 ) ;
  assign n19348 = n19339 | n19347 ;
  assign n19327 = ~n19312 & n19326 ;
  assign n19333 = ( n19327 & ~n11176 ) | ( n19327 & n19332 ) | ( ~n11176 & n19332 ) ;
  assign n19334 = ( n10685 & ~n19333 ) | ( n10685 & 1'b0 ) | ( ~n19333 & 1'b0 ) ;
  assign n19362 = n10209 | n19334 ;
  assign n19363 = ( n19348 & ~n19362 ) | ( n19348 & 1'b0 ) | ( ~n19362 & 1'b0 ) ;
  assign n19364 = n19354 | n19363 ;
  assign n19365 = ( n19342 & ~n19345 ) | ( n19342 & 1'b0 ) | ( ~n19345 & 1'b0 ) ;
  assign n19366 = ( n19339 & ~n10685 ) | ( n19339 & n19365 ) | ( ~n10685 & n19365 ) ;
  assign n19367 = ( n10209 & ~n19366 ) | ( n10209 & 1'b0 ) | ( ~n19366 & 1'b0 ) ;
  assign n19368 = ( n9740 & ~n19367 ) | ( n9740 & 1'b0 ) | ( ~n19367 & 1'b0 ) ;
  assign n19369 = n19364 &  n19368 ;
  assign n19370 = n19361 | n19369 ;
  assign n19349 = ~n19334 & n19348 ;
  assign n19355 = ( n19349 & ~n10209 ) | ( n19349 & n19354 ) | ( ~n10209 & n19354 ) ;
  assign n19356 = n9740 | n19355 ;
  assign n19384 = ~n9286 & n19356 ;
  assign n19385 = n19370 &  n19384 ;
  assign n19386 = n19376 | n19385 ;
  assign n19387 = ( n19364 & ~n19367 ) | ( n19364 & 1'b0 ) | ( ~n19367 & 1'b0 ) ;
  assign n19388 = ( n9740 & n19361 ) | ( n9740 & n19387 ) | ( n19361 & n19387 ) ;
  assign n19389 = ( n9286 & ~n19388 ) | ( n9286 & 1'b0 ) | ( ~n19388 & 1'b0 ) ;
  assign n19390 = n8839 | n19389 ;
  assign n19391 = ( n19386 & ~n19390 ) | ( n19386 & 1'b0 ) | ( ~n19390 & 1'b0 ) ;
  assign n19392 = n19383 | n19391 ;
  assign n19371 = n19356 &  n19370 ;
  assign n19377 = ( n19371 & ~n9286 ) | ( n19371 & n19376 ) | ( ~n9286 & n19376 ) ;
  assign n19378 = ( n8839 & ~n19377 ) | ( n8839 & 1'b0 ) | ( ~n19377 & 1'b0 ) ;
  assign n19406 = n8407 | n19378 ;
  assign n19407 = ( n19392 & ~n19406 ) | ( n19392 & 1'b0 ) | ( ~n19406 & 1'b0 ) ;
  assign n19408 = n19398 | n19407 ;
  assign n19409 = ( n19386 & ~n19389 ) | ( n19386 & 1'b0 ) | ( ~n19389 & 1'b0 ) ;
  assign n19410 = ( n19383 & ~n8839 ) | ( n19383 & n19409 ) | ( ~n8839 & n19409 ) ;
  assign n19411 = ( n8407 & ~n19410 ) | ( n8407 & 1'b0 ) | ( ~n19410 & 1'b0 ) ;
  assign n19412 = n7982 | n19411 ;
  assign n19413 = ( n19408 & ~n19412 ) | ( n19408 & 1'b0 ) | ( ~n19412 & 1'b0 ) ;
  assign n19414 = n19405 | n19413 ;
  assign n19393 = ~n19378 & n19392 ;
  assign n19399 = ( n19393 & ~n8407 ) | ( n19393 & n19398 ) | ( ~n8407 & n19398 ) ;
  assign n19400 = ( n7982 & ~n19399 ) | ( n7982 & 1'b0 ) | ( ~n19399 & 1'b0 ) ;
  assign n19428 = ( n7572 & ~n19400 ) | ( n7572 & 1'b0 ) | ( ~n19400 & 1'b0 ) ;
  assign n19429 = n19414 &  n19428 ;
  assign n19430 = n19420 | n19429 ;
  assign n19431 = ( n19408 & ~n19411 ) | ( n19408 & 1'b0 ) | ( ~n19411 & 1'b0 ) ;
  assign n19432 = ( n19405 & ~n7982 ) | ( n19405 & n19431 ) | ( ~n7982 & n19431 ) ;
  assign n19433 = n7572 | n19432 ;
  assign n19434 = n7169 &  n19433 ;
  assign n19435 = n19430 &  n19434 ;
  assign n19436 = n19427 | n19435 ;
  assign n19415 = ~n19400 & n19414 ;
  assign n19421 = ( n7572 & n19415 ) | ( n7572 & n19420 ) | ( n19415 & n19420 ) ;
  assign n19422 = n7169 | n19421 ;
  assign n19450 = ~n6781 & n19422 ;
  assign n19451 = n19436 &  n19450 ;
  assign n19452 = n19442 | n19451 ;
  assign n19453 = n19430 &  n19433 ;
  assign n19454 = ( n7169 & n19427 ) | ( n7169 & n19453 ) | ( n19427 & n19453 ) ;
  assign n19455 = ( n6781 & ~n19454 ) | ( n6781 & 1'b0 ) | ( ~n19454 & 1'b0 ) ;
  assign n19456 = ( n6399 & ~n19455 ) | ( n6399 & 1'b0 ) | ( ~n19455 & 1'b0 ) ;
  assign n19457 = n19452 &  n19456 ;
  assign n19458 = n19449 | n19457 ;
  assign n19437 = n19422 &  n19436 ;
  assign n19443 = ( n19437 & ~n6781 ) | ( n19437 & n19442 ) | ( ~n6781 & n19442 ) ;
  assign n19444 = n6399 | n19443 ;
  assign n19472 = ~n6032 & n19444 ;
  assign n19473 = n19458 &  n19472 ;
  assign n19474 = n19464 | n19473 ;
  assign n19475 = ( n19452 & ~n19455 ) | ( n19452 & 1'b0 ) | ( ~n19455 & 1'b0 ) ;
  assign n19476 = ( n6399 & n19449 ) | ( n6399 & n19475 ) | ( n19449 & n19475 ) ;
  assign n19477 = ( n6032 & ~n19476 ) | ( n6032 & 1'b0 ) | ( ~n19476 & 1'b0 ) ;
  assign n19478 = ( n5672 & ~n19477 ) | ( n5672 & 1'b0 ) | ( ~n19477 & 1'b0 ) ;
  assign n19479 = n19474 &  n19478 ;
  assign n19480 = n19471 | n19479 ;
  assign n19459 = n19444 &  n19458 ;
  assign n19465 = ( n19459 & ~n6032 ) | ( n19459 & n19464 ) | ( ~n6032 & n19464 ) ;
  assign n19466 = n5672 | n19465 ;
  assign n19494 = ~n5327 & n19466 ;
  assign n19495 = n19480 &  n19494 ;
  assign n19496 = n19486 | n19495 ;
  assign n19497 = ( n19474 & ~n19477 ) | ( n19474 & 1'b0 ) | ( ~n19477 & 1'b0 ) ;
  assign n19498 = ( n5672 & n19471 ) | ( n5672 & n19497 ) | ( n19471 & n19497 ) ;
  assign n19499 = ( n5327 & ~n19498 ) | ( n5327 & 1'b0 ) | ( ~n19498 & 1'b0 ) ;
  assign n19500 = n4990 | n19499 ;
  assign n19501 = ( n19496 & ~n19500 ) | ( n19496 & 1'b0 ) | ( ~n19500 & 1'b0 ) ;
  assign n19502 = n19493 | n19501 ;
  assign n19481 = n19466 &  n19480 ;
  assign n19487 = ( n19481 & ~n5327 ) | ( n19481 & n19486 ) | ( ~n5327 & n19486 ) ;
  assign n19488 = ( n4990 & ~n19487 ) | ( n4990 & 1'b0 ) | ( ~n19487 & 1'b0 ) ;
  assign n19516 = n4668 | n19488 ;
  assign n19517 = ( n19502 & ~n19516 ) | ( n19502 & 1'b0 ) | ( ~n19516 & 1'b0 ) ;
  assign n19518 = n19508 | n19517 ;
  assign n19519 = ( n19496 & ~n19499 ) | ( n19496 & 1'b0 ) | ( ~n19499 & 1'b0 ) ;
  assign n19520 = ( n19493 & ~n4990 ) | ( n19493 & n19519 ) | ( ~n4990 & n19519 ) ;
  assign n19521 = ( n4668 & ~n19520 ) | ( n4668 & 1'b0 ) | ( ~n19520 & 1'b0 ) ;
  assign n19522 = n4353 | n19521 ;
  assign n19523 = ( n19518 & ~n19522 ) | ( n19518 & 1'b0 ) | ( ~n19522 & 1'b0 ) ;
  assign n19524 = n19515 | n19523 ;
  assign n19503 = ~n19488 & n19502 ;
  assign n19509 = ( n19503 & ~n4668 ) | ( n19503 & n19508 ) | ( ~n4668 & n19508 ) ;
  assign n19510 = ( n4353 & ~n19509 ) | ( n4353 & 1'b0 ) | ( ~n19509 & 1'b0 ) ;
  assign n19538 = n4053 | n19510 ;
  assign n19539 = ( n19524 & ~n19538 ) | ( n19524 & 1'b0 ) | ( ~n19538 & 1'b0 ) ;
  assign n19540 = n19530 | n19539 ;
  assign n19541 = ( n19518 & ~n19521 ) | ( n19518 & 1'b0 ) | ( ~n19521 & 1'b0 ) ;
  assign n19542 = ( n19515 & ~n4353 ) | ( n19515 & n19541 ) | ( ~n4353 & n19541 ) ;
  assign n19543 = ( n4053 & ~n19542 ) | ( n4053 & 1'b0 ) | ( ~n19542 & 1'b0 ) ;
  assign n19544 = n3760 | n19543 ;
  assign n19545 = ( n19540 & ~n19544 ) | ( n19540 & 1'b0 ) | ( ~n19544 & 1'b0 ) ;
  assign n19546 = n19537 | n19545 ;
  assign n19525 = ~n19510 & n19524 ;
  assign n19531 = ( n19525 & ~n4053 ) | ( n19525 & n19530 ) | ( ~n4053 & n19530 ) ;
  assign n19532 = ( n3760 & ~n19531 ) | ( n3760 & 1'b0 ) | ( ~n19531 & 1'b0 ) ;
  assign n19560 = n3482 | n19532 ;
  assign n19561 = ( n19546 & ~n19560 ) | ( n19546 & 1'b0 ) | ( ~n19560 & 1'b0 ) ;
  assign n19562 = n19552 | n19561 ;
  assign n19563 = ( n19540 & ~n19543 ) | ( n19540 & 1'b0 ) | ( ~n19543 & 1'b0 ) ;
  assign n19564 = ( n19537 & ~n3760 ) | ( n19537 & n19563 ) | ( ~n3760 & n19563 ) ;
  assign n19565 = ( n3482 & ~n19564 ) | ( n3482 & 1'b0 ) | ( ~n19564 & 1'b0 ) ;
  assign n19566 = n3211 | n19565 ;
  assign n19567 = ( n19562 & ~n19566 ) | ( n19562 & 1'b0 ) | ( ~n19566 & 1'b0 ) ;
  assign n19568 = ( n19559 & ~n19567 ) | ( n19559 & 1'b0 ) | ( ~n19567 & 1'b0 ) ;
  assign n19547 = ~n19532 & n19546 ;
  assign n19553 = ( n19547 & ~n3482 ) | ( n19547 & n19552 ) | ( ~n3482 & n19552 ) ;
  assign n19554 = ( n3211 & ~n19553 ) | ( n3211 & 1'b0 ) | ( ~n19553 & 1'b0 ) ;
  assign n19582 = n2955 | n19554 ;
  assign n19583 = n19568 | n19582 ;
  assign n19584 = n19574 &  n19583 ;
  assign n19585 = ( n19562 & ~n19565 ) | ( n19562 & 1'b0 ) | ( ~n19565 & 1'b0 ) ;
  assign n19586 = ( n3211 & ~n19585 ) | ( n3211 & n19559 ) | ( ~n19585 & n19559 ) ;
  assign n19587 = n2955 &  n19586 ;
  assign n19588 = n2706 | n19587 ;
  assign n19589 = n19584 | n19588 ;
  assign n19590 = n19581 &  n19589 ;
  assign n19569 = n19554 | n19568 ;
  assign n19575 = ( n2955 & n19569 ) | ( n2955 & n19574 ) | ( n19569 & n19574 ) ;
  assign n19576 = n2706 &  n19575 ;
  assign n19604 = n2472 | n19576 ;
  assign n19605 = n19590 | n19604 ;
  assign n19606 = n19596 &  n19605 ;
  assign n19607 = n19584 | n19587 ;
  assign n19608 = ( n2706 & n19581 ) | ( n2706 & n19607 ) | ( n19581 & n19607 ) ;
  assign n19609 = n2472 &  n19608 ;
  assign n19610 = n2245 | n19609 ;
  assign n19611 = n19606 | n19610 ;
  assign n19612 = n19603 &  n19611 ;
  assign n19591 = n19576 | n19590 ;
  assign n19597 = ( n2472 & n19591 ) | ( n2472 & n19596 ) | ( n19591 & n19596 ) ;
  assign n19598 = n2245 &  n19597 ;
  assign n19626 = ( n2033 & ~n19598 ) | ( n2033 & 1'b0 ) | ( ~n19598 & 1'b0 ) ;
  assign n19627 = ~n19612 & n19626 ;
  assign n19628 = n19618 | n19627 ;
  assign n19629 = n19606 | n19609 ;
  assign n19630 = ( n2245 & n19603 ) | ( n2245 & n19629 ) | ( n19603 & n19629 ) ;
  assign n19631 = ~n2033 & n19630 ;
  assign n19632 = n1827 | n19631 ;
  assign n19633 = ( n19628 & ~n19632 ) | ( n19628 & 1'b0 ) | ( ~n19632 & 1'b0 ) ;
  assign n19634 = n19625 | n19633 ;
  assign n19613 = n19598 | n19612 ;
  assign n19619 = ( n2033 & ~n19613 ) | ( n2033 & n19618 ) | ( ~n19613 & n19618 ) ;
  assign n19620 = ( n1827 & ~n19619 ) | ( n1827 & 1'b0 ) | ( ~n19619 & 1'b0 ) ;
  assign n19648 = ( n1636 & ~n19620 ) | ( n1636 & 1'b0 ) | ( ~n19620 & 1'b0 ) ;
  assign n19649 = n19634 &  n19648 ;
  assign n19650 = ( n19640 & ~n19649 ) | ( n19640 & 1'b0 ) | ( ~n19649 & 1'b0 ) ;
  assign n19651 = ( n19628 & ~n19631 ) | ( n19628 & 1'b0 ) | ( ~n19631 & 1'b0 ) ;
  assign n19652 = ( n19625 & ~n1827 ) | ( n19625 & n19651 ) | ( ~n1827 & n19651 ) ;
  assign n19653 = n1636 | n19652 ;
  assign n19654 = n1452 &  n19653 ;
  assign n19655 = ~n19650 & n19654 ;
  assign n19656 = n19647 | n19655 ;
  assign n19635 = ~n19620 & n19634 ;
  assign n19641 = ( n1636 & ~n19640 ) | ( n1636 & n19635 ) | ( ~n19640 & n19635 ) ;
  assign n19642 = n1452 | n19641 ;
  assign n19670 = ~n1283 & n19642 ;
  assign n19671 = n19656 &  n19670 ;
  assign n19672 = ( n19662 & ~n19671 ) | ( n19662 & 1'b0 ) | ( ~n19671 & 1'b0 ) ;
  assign n19673 = ~n19650 & n19653 ;
  assign n19674 = ( n1452 & n19647 ) | ( n1452 & n19673 ) | ( n19647 & n19673 ) ;
  assign n19675 = ( n1283 & ~n19674 ) | ( n1283 & 1'b0 ) | ( ~n19674 & 1'b0 ) ;
  assign n19676 = ( n1122 & ~n19675 ) | ( n1122 & 1'b0 ) | ( ~n19675 & 1'b0 ) ;
  assign n19677 = ~n19672 & n19676 ;
  assign n19678 = ( n19669 & ~n19677 ) | ( n19669 & 1'b0 ) | ( ~n19677 & 1'b0 ) ;
  assign n19657 = n19642 &  n19656 ;
  assign n19663 = ( n1283 & ~n19657 ) | ( n1283 & n19662 ) | ( ~n19657 & n19662 ) ;
  assign n19664 = ~n1122 & n19663 ;
  assign n19692 = ( n976 & ~n19664 ) | ( n976 & 1'b0 ) | ( ~n19664 & 1'b0 ) ;
  assign n19693 = ~n19678 & n19692 ;
  assign n19694 = n19684 | n19693 ;
  assign n19695 = n19672 | n19675 ;
  assign n19696 = ( n19669 & ~n1122 ) | ( n19669 & n19695 ) | ( ~n1122 & n19695 ) ;
  assign n19697 = ~n976 & n19696 ;
  assign n19698 = n837 | n19697 ;
  assign n19699 = ( n19694 & ~n19698 ) | ( n19694 & 1'b0 ) | ( ~n19698 & 1'b0 ) ;
  assign n19700 = n19691 | n19699 ;
  assign n19679 = n19664 | n19678 ;
  assign n19685 = ( n976 & ~n19679 ) | ( n976 & n19684 ) | ( ~n19679 & n19684 ) ;
  assign n19686 = ( n837 & ~n19685 ) | ( n837 & 1'b0 ) | ( ~n19685 & 1'b0 ) ;
  assign n19714 = n713 | n19686 ;
  assign n19715 = ( n19700 & ~n19714 ) | ( n19700 & 1'b0 ) | ( ~n19714 & 1'b0 ) ;
  assign n19716 = n19706 | n19715 ;
  assign n19717 = ( n19694 & ~n19697 ) | ( n19694 & 1'b0 ) | ( ~n19697 & 1'b0 ) ;
  assign n19718 = ( n19691 & ~n837 ) | ( n19691 & n19717 ) | ( ~n837 & n19717 ) ;
  assign n19719 = ( n713 & ~n19718 ) | ( n713 & 1'b0 ) | ( ~n19718 & 1'b0 ) ;
  assign n19720 = n595 | n19719 ;
  assign n19721 = ( n19716 & ~n19720 ) | ( n19716 & 1'b0 ) | ( ~n19720 & 1'b0 ) ;
  assign n19722 = n19713 | n19721 ;
  assign n19701 = ~n19686 & n19700 ;
  assign n19707 = ( n19701 & ~n713 ) | ( n19701 & n19706 ) | ( ~n713 & n19706 ) ;
  assign n19708 = ( n595 & ~n19707 ) | ( n595 & 1'b0 ) | ( ~n19707 & 1'b0 ) ;
  assign n19736 = n492 | n19708 ;
  assign n19737 = ( n19722 & ~n19736 ) | ( n19722 & 1'b0 ) | ( ~n19736 & 1'b0 ) ;
  assign n19738 = n19728 | n19737 ;
  assign n19739 = ( n19716 & ~n19719 ) | ( n19716 & 1'b0 ) | ( ~n19719 & 1'b0 ) ;
  assign n19740 = ( n19713 & ~n595 ) | ( n19713 & n19739 ) | ( ~n595 & n19739 ) ;
  assign n19741 = ( n492 & ~n19740 ) | ( n492 & 1'b0 ) | ( ~n19740 & 1'b0 ) ;
  assign n19756 = ( n19738 & ~n19741 ) | ( n19738 & 1'b0 ) | ( ~n19741 & 1'b0 ) ;
  assign n19731 = n19091 | n19175 ;
  assign n19732 = ( n19078 & ~n19091 ) | ( n19078 & n19087 ) | ( ~n19091 & n19087 ) ;
  assign n19734 = ( n19091 & n19731 ) | ( n19091 & n19732 ) | ( n19731 & n19732 ) ;
  assign n19733 = ( n19087 & ~n19732 ) | ( n19087 & n19731 ) | ( ~n19732 & n19731 ) ;
  assign n19735 = ( n19078 & ~n19734 ) | ( n19078 & n19733 ) | ( ~n19734 & n19733 ) ;
  assign n19757 = ( n396 & ~n19756 ) | ( n396 & n19735 ) | ( ~n19756 & n19735 ) ;
  assign n19758 = n315 &  n19757 ;
  assign n19723 = ~n19708 & n19722 ;
  assign n19729 = ( n19723 & ~n492 ) | ( n19723 & n19728 ) | ( ~n492 & n19728 ) ;
  assign n19730 = ( n396 & ~n19729 ) | ( n396 & 1'b0 ) | ( ~n19729 & 1'b0 ) ;
  assign n19742 = n396 | n19741 ;
  assign n19743 = ( n19738 & ~n19742 ) | ( n19738 & 1'b0 ) | ( ~n19742 & 1'b0 ) ;
  assign n19744 = ( n19735 & ~n19743 ) | ( n19735 & 1'b0 ) | ( ~n19743 & 1'b0 ) ;
  assign n19745 = n19730 | n19744 ;
  assign n19751 = ( n315 & ~n19750 ) | ( n315 & n19745 ) | ( ~n19750 & n19745 ) ;
  assign n19752 = n240 &  n19751 ;
  assign n19753 = n315 | n19730 ;
  assign n19754 = n19744 | n19753 ;
  assign n19755 = ~n19750 & n19754 ;
  assign n19759 = n240 | n19758 ;
  assign n19760 = n19755 | n19759 ;
  assign n19761 = ( n19099 & n19108 ) | ( n19099 & n19112 ) | ( n19108 & n19112 ) ;
  assign n19762 = ( n19175 & ~n19108 ) | ( n19175 & n19761 ) | ( ~n19108 & n19761 ) ;
  assign n19763 = ( n19112 & ~n19761 ) | ( n19112 & n19175 ) | ( ~n19761 & n19175 ) ;
  assign n19764 = ( n19099 & ~n19762 ) | ( n19099 & n19763 ) | ( ~n19762 & n19763 ) ;
  assign n19765 = ( n19760 & ~n19764 ) | ( n19760 & 1'b0 ) | ( ~n19764 & 1'b0 ) ;
  assign n19766 = n19752 | n19765 ;
  assign n19768 = ( n19101 & ~n19106 ) | ( n19101 & n19175 ) | ( ~n19106 & n19175 ) ;
  assign n19767 = ~n19114 & n19175 ;
  assign n19769 = ( n19175 & ~n19768 ) | ( n19175 & n19767 ) | ( ~n19768 & n19767 ) ;
  assign n19770 = ( n19767 & ~n19101 ) | ( n19767 & n19768 ) | ( ~n19101 & n19768 ) ;
  assign n19771 = ( n19106 & ~n19769 ) | ( n19106 & n19770 ) | ( ~n19769 & n19770 ) ;
  assign n19772 = ( n181 & n19766 ) | ( n181 & n19771 ) | ( n19766 & n19771 ) ;
  assign n19773 = ~n145 & n19772 ;
  assign n19774 = n19134 | n19175 ;
  assign n19775 = ( n19121 & n19130 ) | ( n19121 & n19134 ) | ( n19130 & n19134 ) ;
  assign n19776 = ( n19774 & ~n19130 ) | ( n19774 & n19775 ) | ( ~n19130 & n19775 ) ;
  assign n19777 = ( n19134 & ~n19775 ) | ( n19134 & n19774 ) | ( ~n19775 & n19774 ) ;
  assign n19778 = ( n19121 & ~n19776 ) | ( n19121 & n19777 ) | ( ~n19776 & n19777 ) ;
  assign n19779 = n181 | n19752 ;
  assign n19780 = n19765 | n19779 ;
  assign n19781 = n19771 &  n19780 ;
  assign n19782 = n19755 | n19758 ;
  assign n19783 = ( n240 & ~n19764 ) | ( n240 & n19782 ) | ( ~n19764 & n19782 ) ;
  assign n19784 = n181 &  n19783 ;
  assign n19785 = ( n145 & ~n19784 ) | ( n145 & 1'b0 ) | ( ~n19784 & 1'b0 ) ;
  assign n19786 = ~n19781 & n19785 ;
  assign n19787 = n19778 | n19786 ;
  assign n19788 = ~n19773 & n19787 ;
  assign n19789 = n19123 | n19175 ;
  assign n19790 = ( n19128 & ~n19123 ) | ( n19128 & n19136 ) | ( ~n19123 & n19136 ) ;
  assign n19792 = ( n19123 & n19789 ) | ( n19123 & n19790 ) | ( n19789 & n19790 ) ;
  assign n19791 = ( n19136 & ~n19790 ) | ( n19136 & n19789 ) | ( ~n19790 & n19789 ) ;
  assign n19793 = ( n19128 & ~n19792 ) | ( n19128 & n19791 ) | ( ~n19792 & n19791 ) ;
  assign n19794 = ( n150 & ~n19788 ) | ( n150 & n19793 ) | ( ~n19788 & n19793 ) ;
  assign n19795 = n19160 | n19175 ;
  assign n19796 = ( n19143 & n19157 ) | ( n19143 & n19160 ) | ( n19157 & n19160 ) ;
  assign n19797 = ( n19795 & ~n19157 ) | ( n19795 & n19796 ) | ( ~n19157 & n19796 ) ;
  assign n19798 = ( n19160 & ~n19796 ) | ( n19160 & n19795 ) | ( ~n19796 & n19795 ) ;
  assign n19799 = ( n19143 & ~n19797 ) | ( n19143 & n19798 ) | ( ~n19797 & n19798 ) ;
  assign n19800 = ( n19144 & ~n19149 ) | ( n19144 & 1'b0 ) | ( ~n19149 & 1'b0 ) ;
  assign n19801 = ~n19175 & n19800 ;
  assign n19802 = ( n19163 & ~n19801 ) | ( n19163 & n19800 ) | ( ~n19801 & n19800 ) ;
  assign n19803 = ( n19799 & ~n19802 ) | ( n19799 & 1'b0 ) | ( ~n19802 & 1'b0 ) ;
  assign n19804 = ~n19794 & n19803 ;
  assign n19805 = ( n133 & ~n19804 ) | ( n133 & n19803 ) | ( ~n19804 & n19803 ) ;
  assign n19806 = n150 | n19773 ;
  assign n19807 = ( n19787 & ~n19806 ) | ( n19787 & 1'b0 ) | ( ~n19806 & 1'b0 ) ;
  assign n19812 = n19807 &  n19793 ;
  assign n19808 = n19781 | n19784 ;
  assign n19809 = ( n145 & ~n19808 ) | ( n145 & n19778 ) | ( ~n19808 & n19778 ) ;
  assign n19810 = ( n150 & ~n19809 ) | ( n150 & 1'b0 ) | ( ~n19809 & 1'b0 ) ;
  assign n19811 = n19799 | n19810 ;
  assign n19813 = ( n19793 & ~n19812 ) | ( n19793 & n19811 ) | ( ~n19812 & n19811 ) ;
  assign n19815 = ( n133 & ~n19149 ) | ( n133 & n19144 ) | ( ~n19149 & n19144 ) ;
  assign n19814 = ( n19149 & ~n19144 ) | ( n19149 & n19175 ) | ( ~n19144 & n19175 ) ;
  assign n19816 = ~n19149 & n19814 ;
  assign n19817 = ( n19149 & n19815 ) | ( n19149 & n19816 ) | ( n19815 & n19816 ) ;
  assign n19818 = ( n19813 & ~n19817 ) | ( n19813 & 1'b0 ) | ( ~n19817 & 1'b0 ) ;
  assign n19819 = ~n19805 | ~n19818 ;
  assign n20409 = n19758 | n19819 ;
  assign n20410 = ( n19750 & n19754 ) | ( n19750 & n19758 ) | ( n19754 & n19758 ) ;
  assign n20411 = ( n20409 & ~n19754 ) | ( n20409 & n20410 ) | ( ~n19754 & n20410 ) ;
  assign n20412 = ( n19758 & ~n20410 ) | ( n19758 & n20409 ) | ( ~n20410 & n20409 ) ;
  assign n20413 = ( n19750 & ~n20411 ) | ( n19750 & n20412 ) | ( ~n20411 & n20412 ) ;
  assign n20336 = n19664 | n19819 ;
  assign n20337 = ( n19664 & ~n19677 ) | ( n19664 & n19669 ) | ( ~n19677 & n19669 ) ;
  assign n20338 = ( n19677 & n20336 ) | ( n19677 & n20337 ) | ( n20336 & n20337 ) ;
  assign n20339 = ( n19664 & ~n20337 ) | ( n19664 & n20336 ) | ( ~n20337 & n20336 ) ;
  assign n20340 = ( n19669 & ~n20338 ) | ( n19669 & n20339 ) | ( ~n20338 & n20339 ) ;
  assign n19824 = ( x10 & ~n19819 ) | ( x10 & x11 ) | ( ~n19819 & x11 ) ;
  assign n19830 = ( x10 & ~x11 ) | ( x10 & 1'b0 ) | ( ~x11 & 1'b0 ) ;
  assign n19820 = x8 | x9 ;
  assign n19825 = ~x10 & n19820 ;
  assign n19826 = ( x10 & ~n19173 ) | ( x10 & n19825 ) | ( ~n19173 & n19825 ) ;
  assign n19827 = ( n19155 & ~n19826 ) | ( n19155 & n19163 ) | ( ~n19826 & n19163 ) ;
  assign n19828 = ( n19155 & ~n19827 ) | ( n19155 & 1'b0 ) | ( ~n19827 & 1'b0 ) ;
  assign n19829 = ( n19819 & ~x11 ) | ( n19819 & n19828 ) | ( ~x11 & n19828 ) ;
  assign n19831 = ( n19824 & ~n19830 ) | ( n19824 & n19829 ) | ( ~n19830 & n19829 ) ;
  assign n19821 = x10 | n19820 ;
  assign n19822 = x10 &  n19819 ;
  assign n19823 = ( n19175 & ~n19821 ) | ( n19175 & n19822 ) | ( ~n19821 & n19822 ) ;
  assign n19832 = n19823 &  n19831 ;
  assign n19833 = ( n18532 & ~n19831 ) | ( n18532 & n19832 ) | ( ~n19831 & n19832 ) ;
  assign n19834 = n18532 | n19823 ;
  assign n19835 = ( n19831 & ~n19834 ) | ( n19831 & 1'b0 ) | ( ~n19834 & 1'b0 ) ;
  assign n19837 = ( n19175 & ~n19817 ) | ( n19175 & 1'b0 ) | ( ~n19817 & 1'b0 ) ;
  assign n19838 = ( n19813 & ~n19805 ) | ( n19813 & n19837 ) | ( ~n19805 & n19837 ) ;
  assign n19839 = n19805 &  n19838 ;
  assign n19836 = ~n18533 & n19819 ;
  assign n19840 = ~n19839 & n19836 ;
  assign n19841 = ( x12 & n19840 ) | ( x12 & n19839 ) | ( n19840 & n19839 ) ;
  assign n19842 = x12 | n19839 ;
  assign n19843 = n19836 | n19842 ;
  assign n19844 = ~n19841 & n19843 ;
  assign n19845 = n19835 | n19844 ;
  assign n19846 = ~n19833 & n19845 ;
  assign n19850 = ~x12 & n19175 ;
  assign n19851 = ( x13 & ~n19850 ) | ( x13 & 1'b0 ) | ( ~n19850 & 1'b0 ) ;
  assign n19852 = n19187 | n19851 ;
  assign n19847 = ( n19175 & ~x12 ) | ( n19175 & n19182 ) | ( ~x12 & n19182 ) ;
  assign n19848 = x12 &  n19847 ;
  assign n19849 = ( n19177 & ~n19848 ) | ( n19177 & n19182 ) | ( ~n19848 & n19182 ) ;
  assign n19853 = ( n19819 & ~n19852 ) | ( n19819 & n19849 ) | ( ~n19852 & n19849 ) ;
  assign n19855 = ( n19819 & ~n19853 ) | ( n19819 & 1'b0 ) | ( ~n19853 & 1'b0 ) ;
  assign n19854 = ~n19849 & n19853 ;
  assign n19856 = ( n19852 & ~n19855 ) | ( n19852 & n19854 ) | ( ~n19855 & n19854 ) ;
  assign n19857 = ( n19846 & ~n17902 ) | ( n19846 & n19856 ) | ( ~n17902 & n19856 ) ;
  assign n19858 = ( n17279 & ~n19857 ) | ( n17279 & 1'b0 ) | ( ~n19857 & 1'b0 ) ;
  assign n19859 = ~n19210 & n19213 ;
  assign n19860 = ( n19196 & ~n19210 ) | ( n19196 & n19859 ) | ( ~n19210 & n19859 ) ;
  assign n19862 = ( n19819 & n19210 ) | ( n19819 & n19860 ) | ( n19210 & n19860 ) ;
  assign n19861 = ( n19819 & ~n19860 ) | ( n19819 & n19859 ) | ( ~n19860 & n19859 ) ;
  assign n19863 = ( n19196 & ~n19862 ) | ( n19196 & n19861 ) | ( ~n19862 & n19861 ) ;
  assign n19864 = n17902 | n19833 ;
  assign n19865 = ( n19845 & ~n19864 ) | ( n19845 & 1'b0 ) | ( ~n19864 & 1'b0 ) ;
  assign n19866 = n19856 | n19865 ;
  assign n19867 = ~n19823 & n19831 ;
  assign n19868 = ( n19844 & ~n18532 ) | ( n19844 & n19867 ) | ( ~n18532 & n19867 ) ;
  assign n19869 = ( n17902 & ~n19868 ) | ( n17902 & 1'b0 ) | ( ~n19868 & 1'b0 ) ;
  assign n19870 = n17279 | n19869 ;
  assign n19871 = ( n19866 & ~n19870 ) | ( n19866 & 1'b0 ) | ( ~n19870 & 1'b0 ) ;
  assign n19872 = n19863 | n19871 ;
  assign n19873 = ~n19858 & n19872 ;
  assign n19875 = ( n19198 & ~n19208 ) | ( n19198 & n19819 ) | ( ~n19208 & n19819 ) ;
  assign n19874 = n19215 &  n19819 ;
  assign n19876 = ( n19819 & ~n19875 ) | ( n19819 & n19874 ) | ( ~n19875 & n19874 ) ;
  assign n19877 = ( n19874 & ~n19198 ) | ( n19874 & n19875 ) | ( ~n19198 & n19875 ) ;
  assign n19878 = ( n19208 & ~n19876 ) | ( n19208 & n19877 ) | ( ~n19876 & n19877 ) ;
  assign n19879 = ( n19873 & ~n16671 ) | ( n19873 & n19878 ) | ( ~n16671 & n19878 ) ;
  assign n19880 = ( n16070 & ~n19879 ) | ( n16070 & 1'b0 ) | ( ~n19879 & 1'b0 ) ;
  assign n19881 = n19235 | n19819 ;
  assign n19882 = ( n19222 & ~n19235 ) | ( n19222 & n19231 ) | ( ~n19235 & n19231 ) ;
  assign n19884 = ( n19235 & n19881 ) | ( n19235 & n19882 ) | ( n19881 & n19882 ) ;
  assign n19883 = ( n19231 & ~n19882 ) | ( n19231 & n19881 ) | ( ~n19882 & n19881 ) ;
  assign n19885 = ( n19222 & ~n19884 ) | ( n19222 & n19883 ) | ( ~n19884 & n19883 ) ;
  assign n19886 = n16671 | n19858 ;
  assign n19887 = ( n19872 & ~n19886 ) | ( n19872 & 1'b0 ) | ( ~n19886 & 1'b0 ) ;
  assign n19888 = n19878 | n19887 ;
  assign n19889 = ( n19866 & ~n19869 ) | ( n19866 & 1'b0 ) | ( ~n19869 & 1'b0 ) ;
  assign n19890 = ( n19863 & ~n17279 ) | ( n19863 & n19889 ) | ( ~n17279 & n19889 ) ;
  assign n19891 = ( n16671 & ~n19890 ) | ( n16671 & 1'b0 ) | ( ~n19890 & 1'b0 ) ;
  assign n19892 = n16070 | n19891 ;
  assign n19893 = ( n19888 & ~n19892 ) | ( n19888 & 1'b0 ) | ( ~n19892 & 1'b0 ) ;
  assign n19894 = n19885 | n19893 ;
  assign n19895 = ~n19880 & n19894 ;
  assign n19896 = n19237 &  n19819 ;
  assign n19897 = ( n19224 & n19229 ) | ( n19224 & n19819 ) | ( n19229 & n19819 ) ;
  assign n19899 = ( n19896 & ~n19224 ) | ( n19896 & n19897 ) | ( ~n19224 & n19897 ) ;
  assign n19898 = ( n19819 & ~n19897 ) | ( n19819 & n19896 ) | ( ~n19897 & n19896 ) ;
  assign n19900 = ( n19229 & ~n19899 ) | ( n19229 & n19898 ) | ( ~n19899 & n19898 ) ;
  assign n19901 = ( n19895 & ~n15484 ) | ( n19895 & n19900 ) | ( ~n15484 & n19900 ) ;
  assign n19902 = ( n14905 & ~n19901 ) | ( n14905 & 1'b0 ) | ( ~n19901 & 1'b0 ) ;
  assign n19903 = n19257 | n19819 ;
  assign n19904 = ( n19244 & ~n19253 ) | ( n19244 & n19257 ) | ( ~n19253 & n19257 ) ;
  assign n19905 = ( n19253 & n19903 ) | ( n19253 & n19904 ) | ( n19903 & n19904 ) ;
  assign n19906 = ( n19257 & ~n19904 ) | ( n19257 & n19903 ) | ( ~n19904 & n19903 ) ;
  assign n19907 = ( n19244 & ~n19905 ) | ( n19244 & n19906 ) | ( ~n19905 & n19906 ) ;
  assign n19908 = n15484 | n19880 ;
  assign n19909 = ( n19894 & ~n19908 ) | ( n19894 & 1'b0 ) | ( ~n19908 & 1'b0 ) ;
  assign n19910 = n19900 | n19909 ;
  assign n19911 = ( n19888 & ~n19891 ) | ( n19888 & 1'b0 ) | ( ~n19891 & 1'b0 ) ;
  assign n19912 = ( n19885 & ~n16070 ) | ( n19885 & n19911 ) | ( ~n16070 & n19911 ) ;
  assign n19913 = ( n15484 & ~n19912 ) | ( n15484 & 1'b0 ) | ( ~n19912 & 1'b0 ) ;
  assign n19914 = n14905 | n19913 ;
  assign n19915 = ( n19910 & ~n19914 ) | ( n19910 & 1'b0 ) | ( ~n19914 & 1'b0 ) ;
  assign n19916 = n19907 | n19915 ;
  assign n19917 = ~n19902 & n19916 ;
  assign n19918 = n19246 | n19819 ;
  assign n19919 = ( n19251 & ~n19246 ) | ( n19251 & n19259 ) | ( ~n19246 & n19259 ) ;
  assign n19921 = ( n19246 & n19918 ) | ( n19246 & n19919 ) | ( n19918 & n19919 ) ;
  assign n19920 = ( n19259 & ~n19919 ) | ( n19259 & n19918 ) | ( ~n19919 & n19918 ) ;
  assign n19922 = ( n19251 & ~n19921 ) | ( n19251 & n19920 ) | ( ~n19921 & n19920 ) ;
  assign n19923 = ( n19917 & ~n14341 ) | ( n19917 & n19922 ) | ( ~n14341 & n19922 ) ;
  assign n19924 = ( n13784 & ~n19923 ) | ( n13784 & 1'b0 ) | ( ~n19923 & 1'b0 ) ;
  assign n19925 = n19279 | n19819 ;
  assign n19926 = ( n19266 & ~n19275 ) | ( n19266 & n19279 ) | ( ~n19275 & n19279 ) ;
  assign n19927 = ( n19275 & n19925 ) | ( n19275 & n19926 ) | ( n19925 & n19926 ) ;
  assign n19928 = ( n19279 & ~n19926 ) | ( n19279 & n19925 ) | ( ~n19926 & n19925 ) ;
  assign n19929 = ( n19266 & ~n19927 ) | ( n19266 & n19928 ) | ( ~n19927 & n19928 ) ;
  assign n19930 = n14341 | n19902 ;
  assign n19931 = ( n19916 & ~n19930 ) | ( n19916 & 1'b0 ) | ( ~n19930 & 1'b0 ) ;
  assign n19932 = n19922 | n19931 ;
  assign n19933 = ( n19910 & ~n19913 ) | ( n19910 & 1'b0 ) | ( ~n19913 & 1'b0 ) ;
  assign n19934 = ( n19907 & ~n14905 ) | ( n19907 & n19933 ) | ( ~n14905 & n19933 ) ;
  assign n19935 = ( n14341 & ~n19934 ) | ( n14341 & 1'b0 ) | ( ~n19934 & 1'b0 ) ;
  assign n19936 = n13784 | n19935 ;
  assign n19937 = ( n19932 & ~n19936 ) | ( n19932 & 1'b0 ) | ( ~n19936 & 1'b0 ) ;
  assign n19938 = n19929 | n19937 ;
  assign n19939 = ~n19924 & n19938 ;
  assign n19940 = n19268 | n19819 ;
  assign n19941 = ( n19268 & ~n19281 ) | ( n19268 & n19273 ) | ( ~n19281 & n19273 ) ;
  assign n19942 = ( n19281 & n19940 ) | ( n19281 & n19941 ) | ( n19940 & n19941 ) ;
  assign n19943 = ( n19268 & ~n19941 ) | ( n19268 & n19940 ) | ( ~n19941 & n19940 ) ;
  assign n19944 = ( n19273 & ~n19942 ) | ( n19273 & n19943 ) | ( ~n19942 & n19943 ) ;
  assign n19945 = ( n19939 & ~n13242 ) | ( n19939 & n19944 ) | ( ~n13242 & n19944 ) ;
  assign n19946 = ( n12707 & ~n19945 ) | ( n12707 & 1'b0 ) | ( ~n19945 & 1'b0 ) ;
  assign n19947 = n19301 | n19819 ;
  assign n19948 = ( n19288 & ~n19301 ) | ( n19288 & n19297 ) | ( ~n19301 & n19297 ) ;
  assign n19950 = ( n19301 & n19947 ) | ( n19301 & n19948 ) | ( n19947 & n19948 ) ;
  assign n19949 = ( n19297 & ~n19948 ) | ( n19297 & n19947 ) | ( ~n19948 & n19947 ) ;
  assign n19951 = ( n19288 & ~n19950 ) | ( n19288 & n19949 ) | ( ~n19950 & n19949 ) ;
  assign n19952 = n13242 | n19924 ;
  assign n19953 = ( n19938 & ~n19952 ) | ( n19938 & 1'b0 ) | ( ~n19952 & 1'b0 ) ;
  assign n19954 = n19944 | n19953 ;
  assign n19955 = ( n19932 & ~n19935 ) | ( n19932 & 1'b0 ) | ( ~n19935 & 1'b0 ) ;
  assign n19956 = ( n19929 & ~n13784 ) | ( n19929 & n19955 ) | ( ~n13784 & n19955 ) ;
  assign n19957 = ( n13242 & ~n19956 ) | ( n13242 & 1'b0 ) | ( ~n19956 & 1'b0 ) ;
  assign n19958 = n12707 | n19957 ;
  assign n19959 = ( n19954 & ~n19958 ) | ( n19954 & 1'b0 ) | ( ~n19958 & 1'b0 ) ;
  assign n19960 = n19951 | n19959 ;
  assign n19961 = ~n19946 & n19960 ;
  assign n19962 = n19303 &  n19819 ;
  assign n19963 = ( n19290 & n19295 ) | ( n19290 & n19819 ) | ( n19295 & n19819 ) ;
  assign n19965 = ( n19962 & ~n19290 ) | ( n19962 & n19963 ) | ( ~n19290 & n19963 ) ;
  assign n19964 = ( n19819 & ~n19963 ) | ( n19819 & n19962 ) | ( ~n19963 & n19962 ) ;
  assign n19966 = ( n19295 & ~n19965 ) | ( n19295 & n19964 ) | ( ~n19965 & n19964 ) ;
  assign n19967 = ( n19961 & ~n12187 ) | ( n19961 & n19966 ) | ( ~n12187 & n19966 ) ;
  assign n19968 = ( n11674 & ~n19967 ) | ( n11674 & 1'b0 ) | ( ~n19967 & 1'b0 ) ;
  assign n19969 = n19323 | n19819 ;
  assign n19970 = ( n19310 & ~n19319 ) | ( n19310 & n19323 ) | ( ~n19319 & n19323 ) ;
  assign n19971 = ( n19319 & n19969 ) | ( n19319 & n19970 ) | ( n19969 & n19970 ) ;
  assign n19972 = ( n19323 & ~n19970 ) | ( n19323 & n19969 ) | ( ~n19970 & n19969 ) ;
  assign n19973 = ( n19310 & ~n19971 ) | ( n19310 & n19972 ) | ( ~n19971 & n19972 ) ;
  assign n19974 = n12187 | n19946 ;
  assign n19975 = ( n19960 & ~n19974 ) | ( n19960 & 1'b0 ) | ( ~n19974 & 1'b0 ) ;
  assign n19976 = n19966 | n19975 ;
  assign n19977 = ( n19954 & ~n19957 ) | ( n19954 & 1'b0 ) | ( ~n19957 & 1'b0 ) ;
  assign n19978 = ( n19951 & ~n12707 ) | ( n19951 & n19977 ) | ( ~n12707 & n19977 ) ;
  assign n19979 = ( n12187 & ~n19978 ) | ( n12187 & 1'b0 ) | ( ~n19978 & 1'b0 ) ;
  assign n19980 = n11674 | n19979 ;
  assign n19981 = ( n19976 & ~n19980 ) | ( n19976 & 1'b0 ) | ( ~n19980 & 1'b0 ) ;
  assign n19982 = n19973 | n19981 ;
  assign n19983 = ~n19968 & n19982 ;
  assign n19984 = n19312 | n19819 ;
  assign n19985 = ( n19317 & ~n19312 ) | ( n19317 & n19325 ) | ( ~n19312 & n19325 ) ;
  assign n19987 = ( n19312 & n19984 ) | ( n19312 & n19985 ) | ( n19984 & n19985 ) ;
  assign n19986 = ( n19325 & ~n19985 ) | ( n19325 & n19984 ) | ( ~n19985 & n19984 ) ;
  assign n19988 = ( n19317 & ~n19987 ) | ( n19317 & n19986 ) | ( ~n19987 & n19986 ) ;
  assign n19989 = ( n19983 & ~n11176 ) | ( n19983 & n19988 ) | ( ~n11176 & n19988 ) ;
  assign n19990 = ( n10685 & ~n19989 ) | ( n10685 & 1'b0 ) | ( ~n19989 & 1'b0 ) ;
  assign n19991 = n19345 | n19819 ;
  assign n19992 = ( n19332 & ~n19341 ) | ( n19332 & n19345 ) | ( ~n19341 & n19345 ) ;
  assign n19993 = ( n19341 & n19991 ) | ( n19341 & n19992 ) | ( n19991 & n19992 ) ;
  assign n19994 = ( n19345 & ~n19992 ) | ( n19345 & n19991 ) | ( ~n19992 & n19991 ) ;
  assign n19995 = ( n19332 & ~n19993 ) | ( n19332 & n19994 ) | ( ~n19993 & n19994 ) ;
  assign n19996 = n11176 | n19968 ;
  assign n19997 = ( n19982 & ~n19996 ) | ( n19982 & 1'b0 ) | ( ~n19996 & 1'b0 ) ;
  assign n19998 = n19988 | n19997 ;
  assign n19999 = ( n19976 & ~n19979 ) | ( n19976 & 1'b0 ) | ( ~n19979 & 1'b0 ) ;
  assign n20000 = ( n19973 & ~n11674 ) | ( n19973 & n19999 ) | ( ~n11674 & n19999 ) ;
  assign n20001 = ( n11176 & ~n20000 ) | ( n11176 & 1'b0 ) | ( ~n20000 & 1'b0 ) ;
  assign n20002 = n10685 | n20001 ;
  assign n20003 = ( n19998 & ~n20002 ) | ( n19998 & 1'b0 ) | ( ~n20002 & 1'b0 ) ;
  assign n20004 = n19995 | n20003 ;
  assign n20005 = ~n19990 & n20004 ;
  assign n20006 = n19334 | n19819 ;
  assign n20007 = ( n19334 & ~n19347 ) | ( n19334 & n19339 ) | ( ~n19347 & n19339 ) ;
  assign n20008 = ( n19347 & n20006 ) | ( n19347 & n20007 ) | ( n20006 & n20007 ) ;
  assign n20009 = ( n19334 & ~n20007 ) | ( n19334 & n20006 ) | ( ~n20007 & n20006 ) ;
  assign n20010 = ( n19339 & ~n20008 ) | ( n19339 & n20009 ) | ( ~n20008 & n20009 ) ;
  assign n20011 = ( n20005 & ~n10209 ) | ( n20005 & n20010 ) | ( ~n10209 & n20010 ) ;
  assign n20012 = n9740 | n20011 ;
  assign n20013 = n19367 | n19819 ;
  assign n20014 = ( n19354 & ~n19367 ) | ( n19354 & n19363 ) | ( ~n19367 & n19363 ) ;
  assign n20016 = ( n19367 & n20013 ) | ( n19367 & n20014 ) | ( n20013 & n20014 ) ;
  assign n20015 = ( n19363 & ~n20014 ) | ( n19363 & n20013 ) | ( ~n20014 & n20013 ) ;
  assign n20017 = ( n19354 & ~n20016 ) | ( n19354 & n20015 ) | ( ~n20016 & n20015 ) ;
  assign n20018 = n10209 | n19990 ;
  assign n20019 = ( n20004 & ~n20018 ) | ( n20004 & 1'b0 ) | ( ~n20018 & 1'b0 ) ;
  assign n20020 = n20010 | n20019 ;
  assign n20021 = ( n19998 & ~n20001 ) | ( n19998 & 1'b0 ) | ( ~n20001 & 1'b0 ) ;
  assign n20022 = ( n19995 & ~n10685 ) | ( n19995 & n20021 ) | ( ~n10685 & n20021 ) ;
  assign n20023 = ( n10209 & ~n20022 ) | ( n10209 & 1'b0 ) | ( ~n20022 & 1'b0 ) ;
  assign n20024 = ( n9740 & ~n20023 ) | ( n9740 & 1'b0 ) | ( ~n20023 & 1'b0 ) ;
  assign n20025 = n20020 &  n20024 ;
  assign n20026 = n20017 | n20025 ;
  assign n20027 = n20012 &  n20026 ;
  assign n20028 = n19369 &  n19819 ;
  assign n20029 = ( n19361 & ~n19356 ) | ( n19361 & n19819 ) | ( ~n19356 & n19819 ) ;
  assign n20031 = ( n20028 & n19356 ) | ( n20028 & n20029 ) | ( n19356 & n20029 ) ;
  assign n20030 = ( n19819 & ~n20029 ) | ( n19819 & n20028 ) | ( ~n20029 & n20028 ) ;
  assign n20032 = ( n19361 & ~n20031 ) | ( n19361 & n20030 ) | ( ~n20031 & n20030 ) ;
  assign n20033 = ( n20027 & ~n9286 ) | ( n20027 & n20032 ) | ( ~n9286 & n20032 ) ;
  assign n20034 = ( n8839 & ~n20033 ) | ( n8839 & 1'b0 ) | ( ~n20033 & 1'b0 ) ;
  assign n20035 = n19389 | n19819 ;
  assign n20036 = ( n19376 & ~n19385 ) | ( n19376 & n19389 ) | ( ~n19385 & n19389 ) ;
  assign n20037 = ( n19385 & n20035 ) | ( n19385 & n20036 ) | ( n20035 & n20036 ) ;
  assign n20038 = ( n19389 & ~n20036 ) | ( n19389 & n20035 ) | ( ~n20036 & n20035 ) ;
  assign n20039 = ( n19376 & ~n20037 ) | ( n19376 & n20038 ) | ( ~n20037 & n20038 ) ;
  assign n20040 = ~n9286 & n20012 ;
  assign n20041 = n20026 &  n20040 ;
  assign n20042 = n20032 | n20041 ;
  assign n20043 = ( n20020 & ~n20023 ) | ( n20020 & 1'b0 ) | ( ~n20023 & 1'b0 ) ;
  assign n20044 = ( n9740 & n20017 ) | ( n9740 & n20043 ) | ( n20017 & n20043 ) ;
  assign n20045 = ( n9286 & ~n20044 ) | ( n9286 & 1'b0 ) | ( ~n20044 & 1'b0 ) ;
  assign n20046 = n8839 | n20045 ;
  assign n20047 = ( n20042 & ~n20046 ) | ( n20042 & 1'b0 ) | ( ~n20046 & 1'b0 ) ;
  assign n20048 = n20039 | n20047 ;
  assign n20049 = ~n20034 & n20048 ;
  assign n20050 = n19378 | n19819 ;
  assign n20051 = ( n19383 & ~n19378 ) | ( n19383 & n19391 ) | ( ~n19378 & n19391 ) ;
  assign n20053 = ( n19378 & n20050 ) | ( n19378 & n20051 ) | ( n20050 & n20051 ) ;
  assign n20052 = ( n19391 & ~n20051 ) | ( n19391 & n20050 ) | ( ~n20051 & n20050 ) ;
  assign n20054 = ( n19383 & ~n20053 ) | ( n19383 & n20052 ) | ( ~n20053 & n20052 ) ;
  assign n20055 = ( n20049 & ~n8407 ) | ( n20049 & n20054 ) | ( ~n8407 & n20054 ) ;
  assign n20056 = ( n7982 & ~n20055 ) | ( n7982 & 1'b0 ) | ( ~n20055 & 1'b0 ) ;
  assign n20057 = n19411 | n19819 ;
  assign n20058 = ( n19398 & ~n19407 ) | ( n19398 & n19411 ) | ( ~n19407 & n19411 ) ;
  assign n20059 = ( n19407 & n20057 ) | ( n19407 & n20058 ) | ( n20057 & n20058 ) ;
  assign n20060 = ( n19411 & ~n20058 ) | ( n19411 & n20057 ) | ( ~n20058 & n20057 ) ;
  assign n20061 = ( n19398 & ~n20059 ) | ( n19398 & n20060 ) | ( ~n20059 & n20060 ) ;
  assign n20062 = n8407 | n20034 ;
  assign n20063 = ( n20048 & ~n20062 ) | ( n20048 & 1'b0 ) | ( ~n20062 & 1'b0 ) ;
  assign n20064 = n20054 | n20063 ;
  assign n20065 = ( n20042 & ~n20045 ) | ( n20042 & 1'b0 ) | ( ~n20045 & 1'b0 ) ;
  assign n20066 = ( n20039 & ~n8839 ) | ( n20039 & n20065 ) | ( ~n8839 & n20065 ) ;
  assign n20067 = ( n8407 & ~n20066 ) | ( n8407 & 1'b0 ) | ( ~n20066 & 1'b0 ) ;
  assign n20068 = n7982 | n20067 ;
  assign n20069 = ( n20064 & ~n20068 ) | ( n20064 & 1'b0 ) | ( ~n20068 & 1'b0 ) ;
  assign n20070 = n20061 | n20069 ;
  assign n20071 = ~n20056 & n20070 ;
  assign n20072 = n19400 | n19819 ;
  assign n20073 = ( n19405 & ~n19400 ) | ( n19405 & n19413 ) | ( ~n19400 & n19413 ) ;
  assign n20075 = ( n19400 & n20072 ) | ( n19400 & n20073 ) | ( n20072 & n20073 ) ;
  assign n20074 = ( n19413 & ~n20073 ) | ( n19413 & n20072 ) | ( ~n20073 & n20072 ) ;
  assign n20076 = ( n19405 & ~n20075 ) | ( n19405 & n20074 ) | ( ~n20075 & n20074 ) ;
  assign n20077 = ( n7572 & n20071 ) | ( n7572 & n20076 ) | ( n20071 & n20076 ) ;
  assign n20078 = n7169 | n20077 ;
  assign n20080 = ( n19429 & ~n19420 ) | ( n19429 & n19433 ) | ( ~n19420 & n19433 ) ;
  assign n20079 = ( n19433 & ~n19819 ) | ( n19433 & 1'b0 ) | ( ~n19819 & 1'b0 ) ;
  assign n20082 = ( n19433 & ~n20080 ) | ( n19433 & n20079 ) | ( ~n20080 & n20079 ) ;
  assign n20081 = ( n20079 & ~n19429 ) | ( n20079 & n20080 ) | ( ~n19429 & n20080 ) ;
  assign n20083 = ( n19420 & ~n20082 ) | ( n19420 & n20081 ) | ( ~n20082 & n20081 ) ;
  assign n20084 = ( n7572 & ~n20056 ) | ( n7572 & 1'b0 ) | ( ~n20056 & 1'b0 ) ;
  assign n20085 = n20070 &  n20084 ;
  assign n20086 = n20076 | n20085 ;
  assign n20087 = ( n20064 & ~n20067 ) | ( n20064 & 1'b0 ) | ( ~n20067 & 1'b0 ) ;
  assign n20088 = ( n20061 & ~n7982 ) | ( n20061 & n20087 ) | ( ~n7982 & n20087 ) ;
  assign n20089 = n7572 | n20088 ;
  assign n20090 = n7169 &  n20089 ;
  assign n20091 = n20086 &  n20090 ;
  assign n20092 = n20083 | n20091 ;
  assign n20093 = n20078 &  n20092 ;
  assign n20094 = ( n19422 & ~n19819 ) | ( n19422 & 1'b0 ) | ( ~n19819 & 1'b0 ) ;
  assign n20095 = ( n19422 & n19427 ) | ( n19422 & n19435 ) | ( n19427 & n19435 ) ;
  assign n20096 = ( n20094 & ~n19435 ) | ( n20094 & n20095 ) | ( ~n19435 & n20095 ) ;
  assign n20097 = ( n19422 & ~n20095 ) | ( n19422 & n20094 ) | ( ~n20095 & n20094 ) ;
  assign n20098 = ( n19427 & ~n20096 ) | ( n19427 & n20097 ) | ( ~n20096 & n20097 ) ;
  assign n20099 = ( n20093 & ~n6781 ) | ( n20093 & n20098 ) | ( ~n6781 & n20098 ) ;
  assign n20100 = n6399 | n20099 ;
  assign n20101 = n19455 | n19819 ;
  assign n20102 = ( n19442 & ~n19451 ) | ( n19442 & n19455 ) | ( ~n19451 & n19455 ) ;
  assign n20103 = ( n19451 & n20101 ) | ( n19451 & n20102 ) | ( n20101 & n20102 ) ;
  assign n20104 = ( n19455 & ~n20102 ) | ( n19455 & n20101 ) | ( ~n20102 & n20101 ) ;
  assign n20105 = ( n19442 & ~n20103 ) | ( n19442 & n20104 ) | ( ~n20103 & n20104 ) ;
  assign n20106 = ~n6781 & n20078 ;
  assign n20107 = n20092 &  n20106 ;
  assign n20108 = n20098 | n20107 ;
  assign n20109 = n20086 &  n20089 ;
  assign n20110 = ( n7169 & n20083 ) | ( n7169 & n20109 ) | ( n20083 & n20109 ) ;
  assign n20111 = ( n6781 & ~n20110 ) | ( n6781 & 1'b0 ) | ( ~n20110 & 1'b0 ) ;
  assign n20112 = ( n6399 & ~n20111 ) | ( n6399 & 1'b0 ) | ( ~n20111 & 1'b0 ) ;
  assign n20113 = n20108 &  n20112 ;
  assign n20114 = n20105 | n20113 ;
  assign n20115 = n20100 &  n20114 ;
  assign n20116 = ( n19444 & ~n19819 ) | ( n19444 & 1'b0 ) | ( ~n19819 & 1'b0 ) ;
  assign n20117 = ( n19444 & n19449 ) | ( n19444 & n19457 ) | ( n19449 & n19457 ) ;
  assign n20118 = ( n20116 & ~n19457 ) | ( n20116 & n20117 ) | ( ~n19457 & n20117 ) ;
  assign n20119 = ( n19444 & ~n20117 ) | ( n19444 & n20116 ) | ( ~n20117 & n20116 ) ;
  assign n20120 = ( n19449 & ~n20118 ) | ( n19449 & n20119 ) | ( ~n20118 & n20119 ) ;
  assign n20121 = ( n20115 & ~n6032 ) | ( n20115 & n20120 ) | ( ~n6032 & n20120 ) ;
  assign n20122 = n5672 | n20121 ;
  assign n20123 = n19477 | n19819 ;
  assign n20124 = ( n19464 & ~n19473 ) | ( n19464 & n19477 ) | ( ~n19473 & n19477 ) ;
  assign n20125 = ( n19473 & n20123 ) | ( n19473 & n20124 ) | ( n20123 & n20124 ) ;
  assign n20126 = ( n19477 & ~n20124 ) | ( n19477 & n20123 ) | ( ~n20124 & n20123 ) ;
  assign n20127 = ( n19464 & ~n20125 ) | ( n19464 & n20126 ) | ( ~n20125 & n20126 ) ;
  assign n20128 = ~n6032 & n20100 ;
  assign n20129 = n20114 &  n20128 ;
  assign n20130 = n20120 | n20129 ;
  assign n20131 = ( n20108 & ~n20111 ) | ( n20108 & 1'b0 ) | ( ~n20111 & 1'b0 ) ;
  assign n20132 = ( n6399 & n20105 ) | ( n6399 & n20131 ) | ( n20105 & n20131 ) ;
  assign n20133 = ( n6032 & ~n20132 ) | ( n6032 & 1'b0 ) | ( ~n20132 & 1'b0 ) ;
  assign n20134 = ( n5672 & ~n20133 ) | ( n5672 & 1'b0 ) | ( ~n20133 & 1'b0 ) ;
  assign n20135 = n20130 &  n20134 ;
  assign n20136 = n20127 | n20135 ;
  assign n20137 = n20122 &  n20136 ;
  assign n20138 = ( n19466 & ~n19819 ) | ( n19466 & 1'b0 ) | ( ~n19819 & 1'b0 ) ;
  assign n20139 = ( n19466 & n19471 ) | ( n19466 & n19479 ) | ( n19471 & n19479 ) ;
  assign n20140 = ( n20138 & ~n19479 ) | ( n20138 & n20139 ) | ( ~n19479 & n20139 ) ;
  assign n20141 = ( n19466 & ~n20139 ) | ( n19466 & n20138 ) | ( ~n20139 & n20138 ) ;
  assign n20142 = ( n19471 & ~n20140 ) | ( n19471 & n20141 ) | ( ~n20140 & n20141 ) ;
  assign n20143 = ( n20137 & ~n5327 ) | ( n20137 & n20142 ) | ( ~n5327 & n20142 ) ;
  assign n20144 = ( n4990 & ~n20143 ) | ( n4990 & 1'b0 ) | ( ~n20143 & 1'b0 ) ;
  assign n20145 = n19499 | n19819 ;
  assign n20146 = ( n19486 & ~n19495 ) | ( n19486 & n19499 ) | ( ~n19495 & n19499 ) ;
  assign n20147 = ( n19495 & n20145 ) | ( n19495 & n20146 ) | ( n20145 & n20146 ) ;
  assign n20148 = ( n19499 & ~n20146 ) | ( n19499 & n20145 ) | ( ~n20146 & n20145 ) ;
  assign n20149 = ( n19486 & ~n20147 ) | ( n19486 & n20148 ) | ( ~n20147 & n20148 ) ;
  assign n20150 = ~n5327 & n20122 ;
  assign n20151 = n20136 &  n20150 ;
  assign n20152 = n20142 | n20151 ;
  assign n20153 = ( n20130 & ~n20133 ) | ( n20130 & 1'b0 ) | ( ~n20133 & 1'b0 ) ;
  assign n20154 = ( n5672 & n20127 ) | ( n5672 & n20153 ) | ( n20127 & n20153 ) ;
  assign n20155 = ( n5327 & ~n20154 ) | ( n5327 & 1'b0 ) | ( ~n20154 & 1'b0 ) ;
  assign n20156 = n4990 | n20155 ;
  assign n20157 = ( n20152 & ~n20156 ) | ( n20152 & 1'b0 ) | ( ~n20156 & 1'b0 ) ;
  assign n20158 = n20149 | n20157 ;
  assign n20159 = ~n20144 & n20158 ;
  assign n20160 = n19488 | n19819 ;
  assign n20161 = ( n19493 & ~n19488 ) | ( n19493 & n19501 ) | ( ~n19488 & n19501 ) ;
  assign n20163 = ( n19488 & n20160 ) | ( n19488 & n20161 ) | ( n20160 & n20161 ) ;
  assign n20162 = ( n19501 & ~n20161 ) | ( n19501 & n20160 ) | ( ~n20161 & n20160 ) ;
  assign n20164 = ( n19493 & ~n20163 ) | ( n19493 & n20162 ) | ( ~n20163 & n20162 ) ;
  assign n20165 = ( n20159 & ~n4668 ) | ( n20159 & n20164 ) | ( ~n4668 & n20164 ) ;
  assign n20166 = ( n4353 & ~n20165 ) | ( n4353 & 1'b0 ) | ( ~n20165 & 1'b0 ) ;
  assign n20167 = n19521 | n19819 ;
  assign n20168 = ( n19508 & ~n19517 ) | ( n19508 & n19521 ) | ( ~n19517 & n19521 ) ;
  assign n20169 = ( n19517 & n20167 ) | ( n19517 & n20168 ) | ( n20167 & n20168 ) ;
  assign n20170 = ( n19521 & ~n20168 ) | ( n19521 & n20167 ) | ( ~n20168 & n20167 ) ;
  assign n20171 = ( n19508 & ~n20169 ) | ( n19508 & n20170 ) | ( ~n20169 & n20170 ) ;
  assign n20172 = n4668 | n20144 ;
  assign n20173 = ( n20158 & ~n20172 ) | ( n20158 & 1'b0 ) | ( ~n20172 & 1'b0 ) ;
  assign n20174 = n20164 | n20173 ;
  assign n20175 = ( n20152 & ~n20155 ) | ( n20152 & 1'b0 ) | ( ~n20155 & 1'b0 ) ;
  assign n20176 = ( n20149 & ~n4990 ) | ( n20149 & n20175 ) | ( ~n4990 & n20175 ) ;
  assign n20177 = ( n4668 & ~n20176 ) | ( n4668 & 1'b0 ) | ( ~n20176 & 1'b0 ) ;
  assign n20178 = n4353 | n20177 ;
  assign n20179 = ( n20174 & ~n20178 ) | ( n20174 & 1'b0 ) | ( ~n20178 & 1'b0 ) ;
  assign n20180 = n20171 | n20179 ;
  assign n20181 = ~n20166 & n20180 ;
  assign n20182 = n19510 | n19819 ;
  assign n20183 = ( n19515 & ~n19510 ) | ( n19515 & n19523 ) | ( ~n19510 & n19523 ) ;
  assign n20185 = ( n19510 & n20182 ) | ( n19510 & n20183 ) | ( n20182 & n20183 ) ;
  assign n20184 = ( n19523 & ~n20183 ) | ( n19523 & n20182 ) | ( ~n20183 & n20182 ) ;
  assign n20186 = ( n19515 & ~n20185 ) | ( n19515 & n20184 ) | ( ~n20185 & n20184 ) ;
  assign n20187 = ( n20181 & ~n4053 ) | ( n20181 & n20186 ) | ( ~n4053 & n20186 ) ;
  assign n20188 = ( n3760 & ~n20187 ) | ( n3760 & 1'b0 ) | ( ~n20187 & 1'b0 ) ;
  assign n20189 = n19543 | n19819 ;
  assign n20190 = ( n19530 & ~n19539 ) | ( n19530 & n19543 ) | ( ~n19539 & n19543 ) ;
  assign n20191 = ( n19539 & n20189 ) | ( n19539 & n20190 ) | ( n20189 & n20190 ) ;
  assign n20192 = ( n19543 & ~n20190 ) | ( n19543 & n20189 ) | ( ~n20190 & n20189 ) ;
  assign n20193 = ( n19530 & ~n20191 ) | ( n19530 & n20192 ) | ( ~n20191 & n20192 ) ;
  assign n20194 = n4053 | n20166 ;
  assign n20195 = ( n20180 & ~n20194 ) | ( n20180 & 1'b0 ) | ( ~n20194 & 1'b0 ) ;
  assign n20196 = n20186 | n20195 ;
  assign n20197 = ( n20174 & ~n20177 ) | ( n20174 & 1'b0 ) | ( ~n20177 & 1'b0 ) ;
  assign n20198 = ( n20171 & ~n4353 ) | ( n20171 & n20197 ) | ( ~n4353 & n20197 ) ;
  assign n20199 = ( n4053 & ~n20198 ) | ( n4053 & 1'b0 ) | ( ~n20198 & 1'b0 ) ;
  assign n20200 = n3760 | n20199 ;
  assign n20201 = ( n20196 & ~n20200 ) | ( n20196 & 1'b0 ) | ( ~n20200 & 1'b0 ) ;
  assign n20202 = n20193 | n20201 ;
  assign n20203 = ~n20188 & n20202 ;
  assign n20204 = n19532 | n19819 ;
  assign n20205 = ( n19537 & ~n19532 ) | ( n19537 & n19545 ) | ( ~n19532 & n19545 ) ;
  assign n20207 = ( n19532 & n20204 ) | ( n19532 & n20205 ) | ( n20204 & n20205 ) ;
  assign n20206 = ( n19545 & ~n20205 ) | ( n19545 & n20204 ) | ( ~n20205 & n20204 ) ;
  assign n20208 = ( n19537 & ~n20207 ) | ( n19537 & n20206 ) | ( ~n20207 & n20206 ) ;
  assign n20209 = ( n20203 & ~n3482 ) | ( n20203 & n20208 ) | ( ~n3482 & n20208 ) ;
  assign n20210 = ( n3211 & ~n20209 ) | ( n3211 & 1'b0 ) | ( ~n20209 & 1'b0 ) ;
  assign n20211 = n19565 | n19819 ;
  assign n20212 = ( n19552 & ~n19561 ) | ( n19552 & n19565 ) | ( ~n19561 & n19565 ) ;
  assign n20213 = ( n19561 & n20211 ) | ( n19561 & n20212 ) | ( n20211 & n20212 ) ;
  assign n20214 = ( n19565 & ~n20212 ) | ( n19565 & n20211 ) | ( ~n20212 & n20211 ) ;
  assign n20215 = ( n19552 & ~n20213 ) | ( n19552 & n20214 ) | ( ~n20213 & n20214 ) ;
  assign n20216 = n3482 | n20188 ;
  assign n20217 = ( n20202 & ~n20216 ) | ( n20202 & 1'b0 ) | ( ~n20216 & 1'b0 ) ;
  assign n20218 = n20208 | n20217 ;
  assign n20219 = ( n20196 & ~n20199 ) | ( n20196 & 1'b0 ) | ( ~n20199 & 1'b0 ) ;
  assign n20220 = ( n20193 & ~n3760 ) | ( n20193 & n20219 ) | ( ~n3760 & n20219 ) ;
  assign n20221 = ( n3482 & ~n20220 ) | ( n3482 & 1'b0 ) | ( ~n20220 & 1'b0 ) ;
  assign n20222 = n3211 | n20221 ;
  assign n20223 = ( n20218 & ~n20222 ) | ( n20218 & 1'b0 ) | ( ~n20222 & 1'b0 ) ;
  assign n20224 = n20215 | n20223 ;
  assign n20225 = ~n20210 & n20224 ;
  assign n20226 = n19554 | n19819 ;
  assign n20227 = ( n19554 & ~n19567 ) | ( n19554 & n19559 ) | ( ~n19567 & n19559 ) ;
  assign n20228 = ( n19567 & n20226 ) | ( n19567 & n20227 ) | ( n20226 & n20227 ) ;
  assign n20229 = ( n19554 & ~n20227 ) | ( n19554 & n20226 ) | ( ~n20227 & n20226 ) ;
  assign n20230 = ( n19559 & ~n20228 ) | ( n19559 & n20229 ) | ( ~n20228 & n20229 ) ;
  assign n20231 = ( n2955 & ~n20225 ) | ( n2955 & n20230 ) | ( ~n20225 & n20230 ) ;
  assign n20232 = n2706 &  n20231 ;
  assign n20234 = ( n19583 & ~n19574 ) | ( n19583 & n19587 ) | ( ~n19574 & n19587 ) ;
  assign n20233 = n19587 | n19819 ;
  assign n20236 = ( n19587 & ~n20234 ) | ( n19587 & n20233 ) | ( ~n20234 & n20233 ) ;
  assign n20235 = ( n20233 & ~n19583 ) | ( n20233 & n20234 ) | ( ~n19583 & n20234 ) ;
  assign n20237 = ( n19574 & ~n20236 ) | ( n19574 & n20235 ) | ( ~n20236 & n20235 ) ;
  assign n20238 = n2955 | n20210 ;
  assign n20239 = ( n20224 & ~n20238 ) | ( n20224 & 1'b0 ) | ( ~n20238 & 1'b0 ) ;
  assign n20240 = ( n20230 & ~n20239 ) | ( n20230 & 1'b0 ) | ( ~n20239 & 1'b0 ) ;
  assign n20241 = ( n20218 & ~n20221 ) | ( n20218 & 1'b0 ) | ( ~n20221 & 1'b0 ) ;
  assign n20242 = ( n20215 & ~n3211 ) | ( n20215 & n20241 ) | ( ~n3211 & n20241 ) ;
  assign n20243 = ( n2955 & ~n20242 ) | ( n2955 & 1'b0 ) | ( ~n20242 & 1'b0 ) ;
  assign n20244 = n2706 | n20243 ;
  assign n20245 = n20240 | n20244 ;
  assign n20246 = n20237 &  n20245 ;
  assign n20247 = n20232 | n20246 ;
  assign n20248 = n19576 | n19819 ;
  assign n20249 = ( n19576 & n19581 ) | ( n19576 & n19589 ) | ( n19581 & n19589 ) ;
  assign n20250 = ( n20248 & ~n19589 ) | ( n20248 & n20249 ) | ( ~n19589 & n20249 ) ;
  assign n20251 = ( n19576 & ~n20249 ) | ( n19576 & n20248 ) | ( ~n20249 & n20248 ) ;
  assign n20252 = ( n19581 & ~n20250 ) | ( n19581 & n20251 ) | ( ~n20250 & n20251 ) ;
  assign n20253 = ( n2472 & n20247 ) | ( n2472 & n20252 ) | ( n20247 & n20252 ) ;
  assign n20254 = n2245 &  n20253 ;
  assign n20256 = ( n19605 & ~n19596 ) | ( n19605 & n19609 ) | ( ~n19596 & n19609 ) ;
  assign n20255 = n19609 | n19819 ;
  assign n20258 = ( n19609 & ~n20256 ) | ( n19609 & n20255 ) | ( ~n20256 & n20255 ) ;
  assign n20257 = ( n20255 & ~n19605 ) | ( n20255 & n20256 ) | ( ~n19605 & n20256 ) ;
  assign n20259 = ( n19596 & ~n20258 ) | ( n19596 & n20257 ) | ( ~n20258 & n20257 ) ;
  assign n20260 = n2472 | n20232 ;
  assign n20261 = n20246 | n20260 ;
  assign n20262 = n20252 &  n20261 ;
  assign n20263 = n20240 | n20243 ;
  assign n20264 = ( n2706 & n20237 ) | ( n2706 & n20263 ) | ( n20237 & n20263 ) ;
  assign n20265 = n2472 &  n20264 ;
  assign n20266 = n2245 | n20265 ;
  assign n20267 = n20262 | n20266 ;
  assign n20268 = n20259 &  n20267 ;
  assign n20269 = n20254 | n20268 ;
  assign n20270 = n19598 | n19819 ;
  assign n20271 = ( n19598 & n19603 ) | ( n19598 & n19611 ) | ( n19603 & n19611 ) ;
  assign n20272 = ( n20270 & ~n19611 ) | ( n20270 & n20271 ) | ( ~n19611 & n20271 ) ;
  assign n20273 = ( n19598 & ~n20271 ) | ( n19598 & n20270 ) | ( ~n20271 & n20270 ) ;
  assign n20274 = ( n19603 & ~n20272 ) | ( n19603 & n20273 ) | ( ~n20272 & n20273 ) ;
  assign n20275 = ( n20269 & ~n2033 ) | ( n20269 & n20274 ) | ( ~n2033 & n20274 ) ;
  assign n20276 = n1827 &  n20275 ;
  assign n20277 = n19631 | n19819 ;
  assign n20278 = ( n19618 & ~n19627 ) | ( n19618 & n19631 ) | ( ~n19627 & n19631 ) ;
  assign n20279 = ( n19627 & n20277 ) | ( n19627 & n20278 ) | ( n20277 & n20278 ) ;
  assign n20280 = ( n19631 & ~n20278 ) | ( n19631 & n20277 ) | ( ~n20278 & n20277 ) ;
  assign n20281 = ( n19618 & ~n20279 ) | ( n19618 & n20280 ) | ( ~n20279 & n20280 ) ;
  assign n20282 = ( n2033 & ~n20254 ) | ( n2033 & 1'b0 ) | ( ~n20254 & 1'b0 ) ;
  assign n20283 = ~n20268 & n20282 ;
  assign n20284 = ( n20274 & ~n20283 ) | ( n20274 & 1'b0 ) | ( ~n20283 & 1'b0 ) ;
  assign n20285 = n20262 | n20265 ;
  assign n20286 = ( n2245 & n20259 ) | ( n2245 & n20285 ) | ( n20259 & n20285 ) ;
  assign n20287 = ~n2033 & n20286 ;
  assign n20288 = n1827 | n20287 ;
  assign n20289 = n20284 | n20288 ;
  assign n20290 = ~n20281 & n20289 ;
  assign n20291 = n20276 | n20290 ;
  assign n20292 = n19620 | n19819 ;
  assign n20293 = ( n19625 & ~n19620 ) | ( n19625 & n19633 ) | ( ~n19620 & n19633 ) ;
  assign n20295 = ( n19620 & n20292 ) | ( n19620 & n20293 ) | ( n20292 & n20293 ) ;
  assign n20294 = ( n19633 & ~n20293 ) | ( n19633 & n20292 ) | ( ~n20293 & n20292 ) ;
  assign n20296 = ( n19625 & ~n20295 ) | ( n19625 & n20294 ) | ( ~n20295 & n20294 ) ;
  assign n20297 = ( n1636 & ~n20291 ) | ( n1636 & n20296 ) | ( ~n20291 & n20296 ) ;
  assign n20298 = n1452 | n20297 ;
  assign n20299 = ( n19653 & ~n19819 ) | ( n19653 & 1'b0 ) | ( ~n19819 & 1'b0 ) ;
  assign n20300 = ( n19640 & n19649 ) | ( n19640 & n19653 ) | ( n19649 & n19653 ) ;
  assign n20301 = ( n20299 & ~n19649 ) | ( n20299 & n20300 ) | ( ~n19649 & n20300 ) ;
  assign n20302 = ( n19653 & ~n20300 ) | ( n19653 & n20299 ) | ( ~n20300 & n20299 ) ;
  assign n20303 = ( n19640 & ~n20301 ) | ( n19640 & n20302 ) | ( ~n20301 & n20302 ) ;
  assign n20304 = ( n1636 & ~n20276 ) | ( n1636 & 1'b0 ) | ( ~n20276 & 1'b0 ) ;
  assign n20305 = ~n20290 & n20304 ;
  assign n20306 = n20296 | n20305 ;
  assign n20307 = n20284 | n20287 ;
  assign n20308 = ( n1827 & ~n20281 ) | ( n1827 & n20307 ) | ( ~n20281 & n20307 ) ;
  assign n20309 = ~n1636 & n20308 ;
  assign n20310 = ( n1452 & ~n20309 ) | ( n1452 & 1'b0 ) | ( ~n20309 & 1'b0 ) ;
  assign n20311 = n20306 &  n20310 ;
  assign n20312 = ( n20303 & ~n20311 ) | ( n20303 & 1'b0 ) | ( ~n20311 & 1'b0 ) ;
  assign n20313 = ( n20298 & ~n20312 ) | ( n20298 & 1'b0 ) | ( ~n20312 & 1'b0 ) ;
  assign n20314 = ( n19642 & ~n19819 ) | ( n19642 & 1'b0 ) | ( ~n19819 & 1'b0 ) ;
  assign n20315 = ( n19642 & n19647 ) | ( n19642 & n19655 ) | ( n19647 & n19655 ) ;
  assign n20316 = ( n20314 & ~n19655 ) | ( n20314 & n20315 ) | ( ~n19655 & n20315 ) ;
  assign n20317 = ( n19642 & ~n20315 ) | ( n19642 & n20314 ) | ( ~n20315 & n20314 ) ;
  assign n20318 = ( n19647 & ~n20316 ) | ( n19647 & n20317 ) | ( ~n20316 & n20317 ) ;
  assign n20319 = ( n20313 & ~n1283 ) | ( n20313 & n20318 ) | ( ~n1283 & n20318 ) ;
  assign n20320 = n1122 | n20319 ;
  assign n20321 = n19675 | n19819 ;
  assign n20322 = ( n19662 & ~n19675 ) | ( n19662 & n19671 ) | ( ~n19675 & n19671 ) ;
  assign n20324 = ( n19675 & n20321 ) | ( n19675 & n20322 ) | ( n20321 & n20322 ) ;
  assign n20323 = ( n19671 & ~n20322 ) | ( n19671 & n20321 ) | ( ~n20322 & n20321 ) ;
  assign n20325 = ( n19662 & ~n20324 ) | ( n19662 & n20323 ) | ( ~n20324 & n20323 ) ;
  assign n20326 = ~n1283 & n20298 ;
  assign n20327 = ~n20312 & n20326 ;
  assign n20328 = n20318 | n20327 ;
  assign n20329 = ( n20306 & ~n20309 ) | ( n20306 & 1'b0 ) | ( ~n20309 & 1'b0 ) ;
  assign n20330 = ( n1452 & ~n20303 ) | ( n1452 & n20329 ) | ( ~n20303 & n20329 ) ;
  assign n20331 = ( n1283 & ~n20330 ) | ( n1283 & 1'b0 ) | ( ~n20330 & 1'b0 ) ;
  assign n20332 = ( n1122 & ~n20331 ) | ( n1122 & 1'b0 ) | ( ~n20331 & 1'b0 ) ;
  assign n20333 = n20328 &  n20332 ;
  assign n20334 = ( n20325 & ~n20333 ) | ( n20325 & 1'b0 ) | ( ~n20333 & 1'b0 ) ;
  assign n20335 = ( n20320 & ~n20334 ) | ( n20320 & 1'b0 ) | ( ~n20334 & 1'b0 ) ;
  assign n20341 = ( n976 & ~n20340 ) | ( n976 & n20335 ) | ( ~n20340 & n20335 ) ;
  assign n20342 = ( n837 & ~n20341 ) | ( n837 & 1'b0 ) | ( ~n20341 & 1'b0 ) ;
  assign n20343 = n19697 | n19819 ;
  assign n20344 = ( n19684 & ~n19693 ) | ( n19684 & n19697 ) | ( ~n19693 & n19697 ) ;
  assign n20345 = ( n19693 & n20343 ) | ( n19693 & n20344 ) | ( n20343 & n20344 ) ;
  assign n20346 = ( n19697 & ~n20344 ) | ( n19697 & n20343 ) | ( ~n20344 & n20343 ) ;
  assign n20347 = ( n19684 & ~n20345 ) | ( n19684 & n20346 ) | ( ~n20345 & n20346 ) ;
  assign n20348 = n976 &  n20320 ;
  assign n20349 = ~n20334 & n20348 ;
  assign n20350 = ( n20340 & ~n20349 ) | ( n20340 & 1'b0 ) | ( ~n20349 & 1'b0 ) ;
  assign n20351 = ( n20328 & ~n20331 ) | ( n20328 & 1'b0 ) | ( ~n20331 & 1'b0 ) ;
  assign n20352 = ( n1122 & ~n20325 ) | ( n1122 & n20351 ) | ( ~n20325 & n20351 ) ;
  assign n20353 = n976 | n20352 ;
  assign n20354 = ~n837 & n20353 ;
  assign n20355 = ~n20350 & n20354 ;
  assign n20356 = n20347 | n20355 ;
  assign n20357 = ~n20342 & n20356 ;
  assign n20358 = n19686 | n19819 ;
  assign n20359 = ( n19691 & ~n19686 ) | ( n19691 & n19699 ) | ( ~n19686 & n19699 ) ;
  assign n20361 = ( n19686 & n20358 ) | ( n19686 & n20359 ) | ( n20358 & n20359 ) ;
  assign n20360 = ( n19699 & ~n20359 ) | ( n19699 & n20358 ) | ( ~n20359 & n20358 ) ;
  assign n20362 = ( n19691 & ~n20361 ) | ( n19691 & n20360 ) | ( ~n20361 & n20360 ) ;
  assign n20363 = ( n20357 & ~n713 ) | ( n20357 & n20362 ) | ( ~n713 & n20362 ) ;
  assign n20364 = ( n595 & ~n20363 ) | ( n595 & 1'b0 ) | ( ~n20363 & 1'b0 ) ;
  assign n20365 = n19719 | n19819 ;
  assign n20366 = ( n19706 & ~n19715 ) | ( n19706 & n19719 ) | ( ~n19715 & n19719 ) ;
  assign n20367 = ( n19715 & n20365 ) | ( n19715 & n20366 ) | ( n20365 & n20366 ) ;
  assign n20368 = ( n19719 & ~n20366 ) | ( n19719 & n20365 ) | ( ~n20366 & n20365 ) ;
  assign n20369 = ( n19706 & ~n20367 ) | ( n19706 & n20368 ) | ( ~n20367 & n20368 ) ;
  assign n20370 = n713 | n20342 ;
  assign n20371 = ( n20356 & ~n20370 ) | ( n20356 & 1'b0 ) | ( ~n20370 & 1'b0 ) ;
  assign n20372 = n20362 | n20371 ;
  assign n20373 = ~n20350 & n20353 ;
  assign n20374 = ( n20347 & ~n837 ) | ( n20347 & n20373 ) | ( ~n837 & n20373 ) ;
  assign n20375 = ( n713 & ~n20374 ) | ( n713 & 1'b0 ) | ( ~n20374 & 1'b0 ) ;
  assign n20376 = n595 | n20375 ;
  assign n20377 = ( n20372 & ~n20376 ) | ( n20372 & 1'b0 ) | ( ~n20376 & 1'b0 ) ;
  assign n20378 = n20369 | n20377 ;
  assign n20379 = ~n20364 & n20378 ;
  assign n20380 = n19708 | n19819 ;
  assign n20381 = ( n19713 & ~n19708 ) | ( n19713 & n19721 ) | ( ~n19708 & n19721 ) ;
  assign n20383 = ( n19708 & n20380 ) | ( n19708 & n20381 ) | ( n20380 & n20381 ) ;
  assign n20382 = ( n19721 & ~n20381 ) | ( n19721 & n20380 ) | ( ~n20381 & n20380 ) ;
  assign n20384 = ( n19713 & ~n20383 ) | ( n19713 & n20382 ) | ( ~n20383 & n20382 ) ;
  assign n20385 = ( n20379 & ~n492 ) | ( n20379 & n20384 ) | ( ~n492 & n20384 ) ;
  assign n20386 = ( n396 & ~n20385 ) | ( n396 & 1'b0 ) | ( ~n20385 & 1'b0 ) ;
  assign n20387 = n19741 | n19819 ;
  assign n20388 = ( n19728 & ~n19737 ) | ( n19728 & n19741 ) | ( ~n19737 & n19741 ) ;
  assign n20389 = ( n19737 & n20387 ) | ( n19737 & n20388 ) | ( n20387 & n20388 ) ;
  assign n20390 = ( n19741 & ~n20388 ) | ( n19741 & n20387 ) | ( ~n20388 & n20387 ) ;
  assign n20391 = ( n19728 & ~n20389 ) | ( n19728 & n20390 ) | ( ~n20389 & n20390 ) ;
  assign n20392 = n492 | n20364 ;
  assign n20393 = ( n20378 & ~n20392 ) | ( n20378 & 1'b0 ) | ( ~n20392 & 1'b0 ) ;
  assign n20394 = n20384 | n20393 ;
  assign n20395 = ( n20372 & ~n20375 ) | ( n20372 & 1'b0 ) | ( ~n20375 & 1'b0 ) ;
  assign n20396 = ( n20369 & ~n595 ) | ( n20369 & n20395 ) | ( ~n595 & n20395 ) ;
  assign n20397 = ( n492 & ~n20396 ) | ( n492 & 1'b0 ) | ( ~n20396 & 1'b0 ) ;
  assign n20398 = n396 | n20397 ;
  assign n20399 = ( n20394 & ~n20398 ) | ( n20394 & 1'b0 ) | ( ~n20398 & 1'b0 ) ;
  assign n20400 = n20391 | n20399 ;
  assign n20401 = ~n20386 & n20400 ;
  assign n20402 = n19730 | n19819 ;
  assign n20403 = ( n19730 & ~n19743 ) | ( n19730 & n19735 ) | ( ~n19743 & n19735 ) ;
  assign n20404 = ( n19743 & n20402 ) | ( n19743 & n20403 ) | ( n20402 & n20403 ) ;
  assign n20405 = ( n19730 & ~n20403 ) | ( n19730 & n20402 ) | ( ~n20403 & n20402 ) ;
  assign n20406 = ( n19735 & ~n20404 ) | ( n19735 & n20405 ) | ( ~n20404 & n20405 ) ;
  assign n20407 = ( n315 & ~n20401 ) | ( n315 & n20406 ) | ( ~n20401 & n20406 ) ;
  assign n20408 = n240 &  n20407 ;
  assign n20414 = n315 | n20386 ;
  assign n20415 = ( n20400 & ~n20414 ) | ( n20400 & 1'b0 ) | ( ~n20414 & 1'b0 ) ;
  assign n20416 = ( n20406 & ~n20415 ) | ( n20406 & 1'b0 ) | ( ~n20415 & 1'b0 ) ;
  assign n20417 = ( n20394 & ~n20397 ) | ( n20394 & 1'b0 ) | ( ~n20397 & 1'b0 ) ;
  assign n20418 = ( n20391 & ~n396 ) | ( n20391 & n20417 ) | ( ~n396 & n20417 ) ;
  assign n20419 = ( n315 & ~n20418 ) | ( n315 & 1'b0 ) | ( ~n20418 & 1'b0 ) ;
  assign n20420 = n240 | n20419 ;
  assign n20421 = n20416 | n20420 ;
  assign n21093 = ( n20408 & ~n20413 ) | ( n20408 & n20421 ) | ( ~n20413 & n20421 ) ;
  assign n20445 = n19773 | n19819 ;
  assign n20446 = ( n19773 & ~n19786 ) | ( n19773 & n19778 ) | ( ~n19786 & n19778 ) ;
  assign n20447 = ( n19786 & n20445 ) | ( n19786 & n20446 ) | ( n20445 & n20446 ) ;
  assign n20448 = ( n19773 & ~n20446 ) | ( n19773 & n20445 ) | ( ~n20446 & n20445 ) ;
  assign n20449 = ( n19778 & ~n20447 ) | ( n19778 & n20448 ) | ( ~n20447 & n20448 ) ;
  assign n20424 = ( n19752 & ~n19764 ) | ( n19752 & n19760 ) | ( ~n19764 & n19760 ) ;
  assign n20425 = ( n19752 & ~n20424 ) | ( n19752 & n19819 ) | ( ~n20424 & n19819 ) ;
  assign n20426 = ( n19819 & ~n19760 ) | ( n19819 & n20424 ) | ( ~n19760 & n20424 ) ;
  assign n20427 = ( n19764 & ~n20425 ) | ( n19764 & n20426 ) | ( ~n20425 & n20426 ) ;
  assign n20422 = ~n20413 & n20421 ;
  assign n20423 = n20408 | n20422 ;
  assign n20428 = ( n181 & ~n20427 ) | ( n181 & n20423 ) | ( ~n20427 & n20423 ) ;
  assign n20429 = ~n145 & n20428 ;
  assign n20430 = n19784 | n19819 ;
  assign n20431 = ( n19771 & n19780 ) | ( n19771 & n19784 ) | ( n19780 & n19784 ) ;
  assign n20432 = ( n20430 & ~n19780 ) | ( n20430 & n20431 ) | ( ~n19780 & n20431 ) ;
  assign n20433 = ( n19784 & ~n20431 ) | ( n19784 & n20430 ) | ( ~n20431 & n20430 ) ;
  assign n20434 = ( n19771 & ~n20432 ) | ( n19771 & n20433 ) | ( ~n20432 & n20433 ) ;
  assign n20435 = n181 | n20408 ;
  assign n20436 = n20422 | n20435 ;
  assign n20437 = ~n20427 & n20436 ;
  assign n20438 = n20416 | n20419 ;
  assign n20439 = ( n240 & ~n20413 ) | ( n240 & n20438 ) | ( ~n20413 & n20438 ) ;
  assign n20440 = n181 &  n20439 ;
  assign n20441 = ( n145 & ~n20440 ) | ( n145 & 1'b0 ) | ( ~n20440 & 1'b0 ) ;
  assign n20442 = ~n20437 & n20441 ;
  assign n20443 = ( n20434 & ~n20442 ) | ( n20434 & 1'b0 ) | ( ~n20442 & 1'b0 ) ;
  assign n20444 = n20429 | n20443 ;
  assign n20450 = ( n150 & ~n20449 ) | ( n150 & n20444 ) | ( ~n20449 & n20444 ) ;
  assign n20451 = n19810 | n19819 ;
  assign n20452 = ( n19793 & ~n19807 ) | ( n19793 & n19810 ) | ( ~n19807 & n19810 ) ;
  assign n20453 = ( n19807 & n20451 ) | ( n19807 & n20452 ) | ( n20451 & n20452 ) ;
  assign n20454 = ( n19810 & ~n20452 ) | ( n19810 & n20451 ) | ( ~n20452 & n20451 ) ;
  assign n20455 = ( n19793 & ~n20453 ) | ( n19793 & n20454 ) | ( ~n20453 & n20454 ) ;
  assign n20456 = n19794 &  n19799 ;
  assign n20457 = ~n19819 & n20456 ;
  assign n20458 = ( n19813 & ~n20456 ) | ( n19813 & n20457 ) | ( ~n20456 & n20457 ) ;
  assign n20459 = n20455 &  n20458 ;
  assign n20460 = ~n20450 & n20459 ;
  assign n20461 = ( n133 & ~n20460 ) | ( n133 & n20459 ) | ( ~n20460 & n20459 ) ;
  assign n20464 = n20437 | n20440 ;
  assign n20465 = ( n20434 & ~n145 ) | ( n20434 & n20464 ) | ( ~n145 & n20464 ) ;
  assign n20466 = n150 &  n20465 ;
  assign n20467 = n20455 | n20466 ;
  assign n20462 = n150 | n20429 ;
  assign n20463 = n20443 | n20462 ;
  assign n20468 = n20449 | n20463 ;
  assign n20469 = ( n20467 & ~n20449 ) | ( n20467 & n20468 ) | ( ~n20449 & n20468 ) ;
  assign n20471 = ( n133 & n19794 ) | ( n133 & n19799 ) | ( n19794 & n19799 ) ;
  assign n20470 = ( n19794 & ~n19819 ) | ( n19794 & n19799 ) | ( ~n19819 & n19799 ) ;
  assign n20472 = ( n19799 & ~n20470 ) | ( n19799 & 1'b0 ) | ( ~n20470 & 1'b0 ) ;
  assign n20473 = ( n20471 & ~n19799 ) | ( n20471 & n20472 ) | ( ~n19799 & n20472 ) ;
  assign n20474 = ( n20469 & ~n20473 ) | ( n20469 & 1'b0 ) | ( ~n20473 & 1'b0 ) ;
  assign n20475 = ~n20461 | ~n20474 ;
  assign n21092 = n20408 | n20475 ;
  assign n21095 = ( n20408 & ~n21093 ) | ( n20408 & n21092 ) | ( ~n21093 & n21092 ) ;
  assign n21094 = ( n21092 & ~n20421 ) | ( n21092 & n21093 ) | ( ~n20421 & n21093 ) ;
  assign n21096 = ( n20413 & ~n21095 ) | ( n20413 & n21094 ) | ( ~n21095 & n21094 ) ;
  assign n21077 = n20419 | n20475 ;
  assign n21078 = ( n20406 & ~n20419 ) | ( n20406 & n20415 ) | ( ~n20419 & n20415 ) ;
  assign n21080 = ( n20419 & n21077 ) | ( n20419 & n21078 ) | ( n21077 & n21078 ) ;
  assign n21079 = ( n20415 & ~n21078 ) | ( n20415 & n21077 ) | ( ~n21078 & n21077 ) ;
  assign n21081 = ( n20406 & ~n21080 ) | ( n20406 & n21079 ) | ( ~n21080 & n21079 ) ;
  assign n21070 = n20386 | n20475 ;
  assign n21071 = ( n20391 & ~n20386 ) | ( n20391 & n20399 ) | ( ~n20386 & n20399 ) ;
  assign n21073 = ( n20386 & n21070 ) | ( n20386 & n21071 ) | ( n21070 & n21071 ) ;
  assign n21072 = ( n20399 & ~n21071 ) | ( n20399 & n21070 ) | ( ~n21071 & n21070 ) ;
  assign n21074 = ( n20391 & ~n21073 ) | ( n20391 & n21072 ) | ( ~n21073 & n21072 ) ;
  assign n21055 = n20397 | n20475 ;
  assign n21056 = ( n20384 & ~n20393 ) | ( n20384 & n20397 ) | ( ~n20393 & n20397 ) ;
  assign n21057 = ( n20393 & n21055 ) | ( n20393 & n21056 ) | ( n21055 & n21056 ) ;
  assign n21058 = ( n20397 & ~n21056 ) | ( n20397 & n21055 ) | ( ~n21056 & n21055 ) ;
  assign n21059 = ( n20384 & ~n21057 ) | ( n20384 & n21058 ) | ( ~n21057 & n21058 ) ;
  assign n21048 = n20364 | n20475 ;
  assign n21049 = ( n20369 & ~n20364 ) | ( n20369 & n20377 ) | ( ~n20364 & n20377 ) ;
  assign n21051 = ( n20364 & n21048 ) | ( n20364 & n21049 ) | ( n21048 & n21049 ) ;
  assign n21050 = ( n20377 & ~n21049 ) | ( n20377 & n21048 ) | ( ~n21049 & n21048 ) ;
  assign n21052 = ( n20369 & ~n21051 ) | ( n20369 & n21050 ) | ( ~n21051 & n21050 ) ;
  assign n21033 = n20375 | n20475 ;
  assign n21034 = ( n20362 & ~n20371 ) | ( n20362 & n20375 ) | ( ~n20371 & n20375 ) ;
  assign n21035 = ( n20371 & n21033 ) | ( n20371 & n21034 ) | ( n21033 & n21034 ) ;
  assign n21036 = ( n20375 & ~n21034 ) | ( n20375 & n21033 ) | ( ~n21034 & n21033 ) ;
  assign n21037 = ( n20362 & ~n21035 ) | ( n20362 & n21036 ) | ( ~n21035 & n21036 ) ;
  assign n21026 = n20342 | n20475 ;
  assign n21027 = ( n20347 & ~n20342 ) | ( n20347 & n20355 ) | ( ~n20342 & n20355 ) ;
  assign n21029 = ( n20342 & n21026 ) | ( n20342 & n21027 ) | ( n21026 & n21027 ) ;
  assign n21028 = ( n20355 & ~n21027 ) | ( n20355 & n21026 ) | ( ~n21027 & n21026 ) ;
  assign n21030 = ( n20347 & ~n21029 ) | ( n20347 & n21028 ) | ( ~n21029 & n21028 ) ;
  assign n21011 = ( n20353 & ~n20475 ) | ( n20353 & 1'b0 ) | ( ~n20475 & 1'b0 ) ;
  assign n21012 = ( n20340 & n20349 ) | ( n20340 & n20353 ) | ( n20349 & n20353 ) ;
  assign n21013 = ( n21011 & ~n20349 ) | ( n21011 & n21012 ) | ( ~n20349 & n21012 ) ;
  assign n21014 = ( n20353 & ~n21012 ) | ( n20353 & n21011 ) | ( ~n21012 & n21011 ) ;
  assign n21015 = ( n20340 & ~n21013 ) | ( n20340 & n21014 ) | ( ~n21013 & n21014 ) ;
  assign n21005 = ( n20320 & ~n20325 ) | ( n20320 & n20333 ) | ( ~n20325 & n20333 ) ;
  assign n21004 = ( n20320 & ~n20475 ) | ( n20320 & 1'b0 ) | ( ~n20475 & 1'b0 ) ;
  assign n21007 = ( n20320 & ~n21005 ) | ( n20320 & n21004 ) | ( ~n21005 & n21004 ) ;
  assign n21006 = ( n21004 & ~n20333 ) | ( n21004 & n21005 ) | ( ~n20333 & n21005 ) ;
  assign n21008 = ( n20325 & ~n21007 ) | ( n20325 & n21006 ) | ( ~n21007 & n21006 ) ;
  assign n20989 = n20331 | n20475 ;
  assign n20990 = ( n20318 & ~n20327 ) | ( n20318 & n20331 ) | ( ~n20327 & n20331 ) ;
  assign n20991 = ( n20327 & n20989 ) | ( n20327 & n20990 ) | ( n20989 & n20990 ) ;
  assign n20992 = ( n20331 & ~n20990 ) | ( n20331 & n20989 ) | ( ~n20990 & n20989 ) ;
  assign n20993 = ( n20318 & ~n20991 ) | ( n20318 & n20992 ) | ( ~n20991 & n20992 ) ;
  assign n20983 = ( n20298 & ~n20303 ) | ( n20298 & n20311 ) | ( ~n20303 & n20311 ) ;
  assign n20982 = ( n20298 & ~n20475 ) | ( n20298 & 1'b0 ) | ( ~n20475 & 1'b0 ) ;
  assign n20985 = ( n20298 & ~n20983 ) | ( n20298 & n20982 ) | ( ~n20983 & n20982 ) ;
  assign n20984 = ( n20982 & ~n20311 ) | ( n20982 & n20983 ) | ( ~n20311 & n20983 ) ;
  assign n20986 = ( n20303 & ~n20985 ) | ( n20303 & n20984 ) | ( ~n20985 & n20984 ) ;
  assign n20967 = n20309 | n20475 ;
  assign n20968 = ( n20296 & ~n20305 ) | ( n20296 & n20309 ) | ( ~n20305 & n20309 ) ;
  assign n20969 = ( n20305 & n20967 ) | ( n20305 & n20968 ) | ( n20967 & n20968 ) ;
  assign n20970 = ( n20309 & ~n20968 ) | ( n20309 & n20967 ) | ( ~n20968 & n20967 ) ;
  assign n20971 = ( n20296 & ~n20969 ) | ( n20296 & n20970 ) | ( ~n20969 & n20970 ) ;
  assign n20961 = ( n20276 & ~n20281 ) | ( n20276 & n20289 ) | ( ~n20281 & n20289 ) ;
  assign n20960 = n20276 | n20475 ;
  assign n20963 = ( n20276 & ~n20961 ) | ( n20276 & n20960 ) | ( ~n20961 & n20960 ) ;
  assign n20962 = ( n20960 & ~n20289 ) | ( n20960 & n20961 ) | ( ~n20289 & n20961 ) ;
  assign n20964 = ( n20281 & ~n20963 ) | ( n20281 & n20962 ) | ( ~n20963 & n20962 ) ;
  assign n20945 = n20287 | n20475 ;
  assign n20946 = ( n20274 & ~n20287 ) | ( n20274 & n20283 ) | ( ~n20287 & n20283 ) ;
  assign n20948 = ( n20287 & n20945 ) | ( n20287 & n20946 ) | ( n20945 & n20946 ) ;
  assign n20947 = ( n20283 & ~n20946 ) | ( n20283 & n20945 ) | ( ~n20946 & n20945 ) ;
  assign n20949 = ( n20274 & ~n20948 ) | ( n20274 & n20947 ) | ( ~n20948 & n20947 ) ;
  assign n20938 = n20254 | n20475 ;
  assign n20939 = ( n20254 & n20259 ) | ( n20254 & n20267 ) | ( n20259 & n20267 ) ;
  assign n20940 = ( n20938 & ~n20267 ) | ( n20938 & n20939 ) | ( ~n20267 & n20939 ) ;
  assign n20941 = ( n20254 & ~n20939 ) | ( n20254 & n20938 ) | ( ~n20939 & n20938 ) ;
  assign n20942 = ( n20259 & ~n20940 ) | ( n20259 & n20941 ) | ( ~n20940 & n20941 ) ;
  assign n20924 = ( n20261 & ~n20252 ) | ( n20261 & n20265 ) | ( ~n20252 & n20265 ) ;
  assign n20923 = n20265 | n20475 ;
  assign n20926 = ( n20265 & ~n20924 ) | ( n20265 & n20923 ) | ( ~n20924 & n20923 ) ;
  assign n20925 = ( n20923 & ~n20261 ) | ( n20923 & n20924 ) | ( ~n20261 & n20924 ) ;
  assign n20927 = ( n20252 & ~n20926 ) | ( n20252 & n20925 ) | ( ~n20926 & n20925 ) ;
  assign n20916 = n20232 | n20475 ;
  assign n20917 = ( n20232 & n20237 ) | ( n20232 & n20245 ) | ( n20237 & n20245 ) ;
  assign n20918 = ( n20916 & ~n20245 ) | ( n20916 & n20917 ) | ( ~n20245 & n20917 ) ;
  assign n20919 = ( n20232 & ~n20917 ) | ( n20232 & n20916 ) | ( ~n20917 & n20916 ) ;
  assign n20920 = ( n20237 & ~n20918 ) | ( n20237 & n20919 ) | ( ~n20918 & n20919 ) ;
  assign n20901 = n20243 | n20475 ;
  assign n20902 = ( n20230 & ~n20243 ) | ( n20230 & n20239 ) | ( ~n20243 & n20239 ) ;
  assign n20904 = ( n20243 & n20901 ) | ( n20243 & n20902 ) | ( n20901 & n20902 ) ;
  assign n20903 = ( n20239 & ~n20902 ) | ( n20239 & n20901 ) | ( ~n20902 & n20901 ) ;
  assign n20905 = ( n20230 & ~n20904 ) | ( n20230 & n20903 ) | ( ~n20904 & n20903 ) ;
  assign n20894 = n20210 | n20475 ;
  assign n20895 = ( n20215 & ~n20210 ) | ( n20215 & n20223 ) | ( ~n20210 & n20223 ) ;
  assign n20897 = ( n20210 & n20894 ) | ( n20210 & n20895 ) | ( n20894 & n20895 ) ;
  assign n20896 = ( n20223 & ~n20895 ) | ( n20223 & n20894 ) | ( ~n20895 & n20894 ) ;
  assign n20898 = ( n20215 & ~n20897 ) | ( n20215 & n20896 ) | ( ~n20897 & n20896 ) ;
  assign n20879 = n20221 | n20475 ;
  assign n20880 = ( n20208 & ~n20217 ) | ( n20208 & n20221 ) | ( ~n20217 & n20221 ) ;
  assign n20881 = ( n20217 & n20879 ) | ( n20217 & n20880 ) | ( n20879 & n20880 ) ;
  assign n20882 = ( n20221 & ~n20880 ) | ( n20221 & n20879 ) | ( ~n20880 & n20879 ) ;
  assign n20883 = ( n20208 & ~n20881 ) | ( n20208 & n20882 ) | ( ~n20881 & n20882 ) ;
  assign n20872 = n20188 | n20475 ;
  assign n20873 = ( n20193 & ~n20188 ) | ( n20193 & n20201 ) | ( ~n20188 & n20201 ) ;
  assign n20875 = ( n20188 & n20872 ) | ( n20188 & n20873 ) | ( n20872 & n20873 ) ;
  assign n20874 = ( n20201 & ~n20873 ) | ( n20201 & n20872 ) | ( ~n20873 & n20872 ) ;
  assign n20876 = ( n20193 & ~n20875 ) | ( n20193 & n20874 ) | ( ~n20875 & n20874 ) ;
  assign n20857 = n20199 | n20475 ;
  assign n20858 = ( n20186 & ~n20195 ) | ( n20186 & n20199 ) | ( ~n20195 & n20199 ) ;
  assign n20859 = ( n20195 & n20857 ) | ( n20195 & n20858 ) | ( n20857 & n20858 ) ;
  assign n20860 = ( n20199 & ~n20858 ) | ( n20199 & n20857 ) | ( ~n20858 & n20857 ) ;
  assign n20861 = ( n20186 & ~n20859 ) | ( n20186 & n20860 ) | ( ~n20859 & n20860 ) ;
  assign n20850 = n20166 | n20475 ;
  assign n20851 = ( n20171 & ~n20166 ) | ( n20171 & n20179 ) | ( ~n20166 & n20179 ) ;
  assign n20853 = ( n20166 & n20850 ) | ( n20166 & n20851 ) | ( n20850 & n20851 ) ;
  assign n20852 = ( n20179 & ~n20851 ) | ( n20179 & n20850 ) | ( ~n20851 & n20850 ) ;
  assign n20854 = ( n20171 & ~n20853 ) | ( n20171 & n20852 ) | ( ~n20853 & n20852 ) ;
  assign n20835 = n20177 | n20475 ;
  assign n20836 = ( n20164 & ~n20173 ) | ( n20164 & n20177 ) | ( ~n20173 & n20177 ) ;
  assign n20837 = ( n20173 & n20835 ) | ( n20173 & n20836 ) | ( n20835 & n20836 ) ;
  assign n20838 = ( n20177 & ~n20836 ) | ( n20177 & n20835 ) | ( ~n20836 & n20835 ) ;
  assign n20839 = ( n20164 & ~n20837 ) | ( n20164 & n20838 ) | ( ~n20837 & n20838 ) ;
  assign n20828 = n20144 | n20475 ;
  assign n20829 = ( n20149 & ~n20144 ) | ( n20149 & n20157 ) | ( ~n20144 & n20157 ) ;
  assign n20831 = ( n20144 & n20828 ) | ( n20144 & n20829 ) | ( n20828 & n20829 ) ;
  assign n20830 = ( n20157 & ~n20829 ) | ( n20157 & n20828 ) | ( ~n20829 & n20828 ) ;
  assign n20832 = ( n20149 & ~n20831 ) | ( n20149 & n20830 ) | ( ~n20831 & n20830 ) ;
  assign n20813 = n20155 | n20475 ;
  assign n20814 = ( n20142 & ~n20151 ) | ( n20142 & n20155 ) | ( ~n20151 & n20155 ) ;
  assign n20815 = ( n20151 & n20813 ) | ( n20151 & n20814 ) | ( n20813 & n20814 ) ;
  assign n20816 = ( n20155 & ~n20814 ) | ( n20155 & n20813 ) | ( ~n20814 & n20813 ) ;
  assign n20817 = ( n20142 & ~n20815 ) | ( n20142 & n20816 ) | ( ~n20815 & n20816 ) ;
  assign n20806 = ( n20122 & ~n20475 ) | ( n20122 & 1'b0 ) | ( ~n20475 & 1'b0 ) ;
  assign n20807 = ( n20122 & n20127 ) | ( n20122 & n20135 ) | ( n20127 & n20135 ) ;
  assign n20808 = ( n20806 & ~n20135 ) | ( n20806 & n20807 ) | ( ~n20135 & n20807 ) ;
  assign n20809 = ( n20122 & ~n20807 ) | ( n20122 & n20806 ) | ( ~n20807 & n20806 ) ;
  assign n20810 = ( n20127 & ~n20808 ) | ( n20127 & n20809 ) | ( ~n20808 & n20809 ) ;
  assign n20791 = n20133 | n20475 ;
  assign n20792 = ( n20120 & ~n20129 ) | ( n20120 & n20133 ) | ( ~n20129 & n20133 ) ;
  assign n20793 = ( n20129 & n20791 ) | ( n20129 & n20792 ) | ( n20791 & n20792 ) ;
  assign n20794 = ( n20133 & ~n20792 ) | ( n20133 & n20791 ) | ( ~n20792 & n20791 ) ;
  assign n20795 = ( n20120 & ~n20793 ) | ( n20120 & n20794 ) | ( ~n20793 & n20794 ) ;
  assign n20784 = ( n20100 & ~n20475 ) | ( n20100 & 1'b0 ) | ( ~n20475 & 1'b0 ) ;
  assign n20785 = ( n20100 & n20105 ) | ( n20100 & n20113 ) | ( n20105 & n20113 ) ;
  assign n20786 = ( n20784 & ~n20113 ) | ( n20784 & n20785 ) | ( ~n20113 & n20785 ) ;
  assign n20787 = ( n20100 & ~n20785 ) | ( n20100 & n20784 ) | ( ~n20785 & n20784 ) ;
  assign n20788 = ( n20105 & ~n20786 ) | ( n20105 & n20787 ) | ( ~n20786 & n20787 ) ;
  assign n20769 = n20111 | n20475 ;
  assign n20770 = ( n20098 & ~n20107 ) | ( n20098 & n20111 ) | ( ~n20107 & n20111 ) ;
  assign n20771 = ( n20107 & n20769 ) | ( n20107 & n20770 ) | ( n20769 & n20770 ) ;
  assign n20772 = ( n20111 & ~n20770 ) | ( n20111 & n20769 ) | ( ~n20770 & n20769 ) ;
  assign n20773 = ( n20098 & ~n20771 ) | ( n20098 & n20772 ) | ( ~n20771 & n20772 ) ;
  assign n20762 = ( n20078 & ~n20475 ) | ( n20078 & 1'b0 ) | ( ~n20475 & 1'b0 ) ;
  assign n20763 = ( n20078 & n20083 ) | ( n20078 & n20091 ) | ( n20083 & n20091 ) ;
  assign n20764 = ( n20762 & ~n20091 ) | ( n20762 & n20763 ) | ( ~n20091 & n20763 ) ;
  assign n20765 = ( n20078 & ~n20763 ) | ( n20078 & n20762 ) | ( ~n20763 & n20762 ) ;
  assign n20766 = ( n20083 & ~n20764 ) | ( n20083 & n20765 ) | ( ~n20764 & n20765 ) ;
  assign n20748 = ( n20085 & ~n20076 ) | ( n20085 & n20089 ) | ( ~n20076 & n20089 ) ;
  assign n20747 = ( n20089 & ~n20475 ) | ( n20089 & 1'b0 ) | ( ~n20475 & 1'b0 ) ;
  assign n20750 = ( n20089 & ~n20748 ) | ( n20089 & n20747 ) | ( ~n20748 & n20747 ) ;
  assign n20749 = ( n20747 & ~n20085 ) | ( n20747 & n20748 ) | ( ~n20085 & n20748 ) ;
  assign n20751 = ( n20076 & ~n20750 ) | ( n20076 & n20749 ) | ( ~n20750 & n20749 ) ;
  assign n20740 = n20056 | n20475 ;
  assign n20741 = ( n20061 & ~n20056 ) | ( n20061 & n20069 ) | ( ~n20056 & n20069 ) ;
  assign n20743 = ( n20056 & n20740 ) | ( n20056 & n20741 ) | ( n20740 & n20741 ) ;
  assign n20742 = ( n20069 & ~n20741 ) | ( n20069 & n20740 ) | ( ~n20741 & n20740 ) ;
  assign n20744 = ( n20061 & ~n20743 ) | ( n20061 & n20742 ) | ( ~n20743 & n20742 ) ;
  assign n20725 = n20067 | n20475 ;
  assign n20726 = ( n20054 & ~n20063 ) | ( n20054 & n20067 ) | ( ~n20063 & n20067 ) ;
  assign n20727 = ( n20063 & n20725 ) | ( n20063 & n20726 ) | ( n20725 & n20726 ) ;
  assign n20728 = ( n20067 & ~n20726 ) | ( n20067 & n20725 ) | ( ~n20726 & n20725 ) ;
  assign n20729 = ( n20054 & ~n20727 ) | ( n20054 & n20728 ) | ( ~n20727 & n20728 ) ;
  assign n20718 = n20047 &  n20475 ;
  assign n20719 = ( n20034 & n20039 ) | ( n20034 & n20475 ) | ( n20039 & n20475 ) ;
  assign n20721 = ( n20718 & ~n20034 ) | ( n20718 & n20719 ) | ( ~n20034 & n20719 ) ;
  assign n20720 = ( n20475 & ~n20719 ) | ( n20475 & n20718 ) | ( ~n20719 & n20718 ) ;
  assign n20722 = ( n20039 & ~n20721 ) | ( n20039 & n20720 ) | ( ~n20721 & n20720 ) ;
  assign n20703 = n20045 | n20475 ;
  assign n20704 = ( n20032 & ~n20045 ) | ( n20032 & n20041 ) | ( ~n20045 & n20041 ) ;
  assign n20706 = ( n20045 & n20703 ) | ( n20045 & n20704 ) | ( n20703 & n20704 ) ;
  assign n20705 = ( n20041 & ~n20704 ) | ( n20041 & n20703 ) | ( ~n20704 & n20703 ) ;
  assign n20707 = ( n20032 & ~n20706 ) | ( n20032 & n20705 ) | ( ~n20706 & n20705 ) ;
  assign n20697 = ( n20012 & ~n20017 ) | ( n20012 & n20025 ) | ( ~n20017 & n20025 ) ;
  assign n20696 = ( n20012 & ~n20475 ) | ( n20012 & 1'b0 ) | ( ~n20475 & 1'b0 ) ;
  assign n20699 = ( n20012 & ~n20697 ) | ( n20012 & n20696 ) | ( ~n20697 & n20696 ) ;
  assign n20698 = ( n20696 & ~n20025 ) | ( n20696 & n20697 ) | ( ~n20025 & n20697 ) ;
  assign n20700 = ( n20017 & ~n20699 ) | ( n20017 & n20698 ) | ( ~n20699 & n20698 ) ;
  assign n20681 = n20023 | n20475 ;
  assign n20682 = ( n20010 & ~n20019 ) | ( n20010 & n20023 ) | ( ~n20019 & n20023 ) ;
  assign n20683 = ( n20019 & n20681 ) | ( n20019 & n20682 ) | ( n20681 & n20682 ) ;
  assign n20684 = ( n20023 & ~n20682 ) | ( n20023 & n20681 ) | ( ~n20682 & n20681 ) ;
  assign n20685 = ( n20010 & ~n20683 ) | ( n20010 & n20684 ) | ( ~n20683 & n20684 ) ;
  assign n20674 = n19990 | n20475 ;
  assign n20675 = ( n19995 & ~n19990 ) | ( n19995 & n20003 ) | ( ~n19990 & n20003 ) ;
  assign n20677 = ( n19990 & n20674 ) | ( n19990 & n20675 ) | ( n20674 & n20675 ) ;
  assign n20676 = ( n20003 & ~n20675 ) | ( n20003 & n20674 ) | ( ~n20675 & n20674 ) ;
  assign n20678 = ( n19995 & ~n20677 ) | ( n19995 & n20676 ) | ( ~n20677 & n20676 ) ;
  assign n20659 = n20001 | n20475 ;
  assign n20660 = ( n19988 & ~n19997 ) | ( n19988 & n20001 ) | ( ~n19997 & n20001 ) ;
  assign n20661 = ( n19997 & n20659 ) | ( n19997 & n20660 ) | ( n20659 & n20660 ) ;
  assign n20662 = ( n20001 & ~n20660 ) | ( n20001 & n20659 ) | ( ~n20660 & n20659 ) ;
  assign n20663 = ( n19988 & ~n20661 ) | ( n19988 & n20662 ) | ( ~n20661 & n20662 ) ;
  assign n20652 = n19981 &  n20475 ;
  assign n20653 = ( n19968 & n19973 ) | ( n19968 & n20475 ) | ( n19973 & n20475 ) ;
  assign n20655 = ( n20652 & ~n19968 ) | ( n20652 & n20653 ) | ( ~n19968 & n20653 ) ;
  assign n20654 = ( n20475 & ~n20653 ) | ( n20475 & n20652 ) | ( ~n20653 & n20652 ) ;
  assign n20656 = ( n19973 & ~n20655 ) | ( n19973 & n20654 ) | ( ~n20655 & n20654 ) ;
  assign n20637 = n19979 | n20475 ;
  assign n20638 = ( n19966 & ~n19979 ) | ( n19966 & n19975 ) | ( ~n19979 & n19975 ) ;
  assign n20640 = ( n19979 & n20637 ) | ( n19979 & n20638 ) | ( n20637 & n20638 ) ;
  assign n20639 = ( n19975 & ~n20638 ) | ( n19975 & n20637 ) | ( ~n20638 & n20637 ) ;
  assign n20641 = ( n19966 & ~n20640 ) | ( n19966 & n20639 ) | ( ~n20640 & n20639 ) ;
  assign n20631 = ( n19946 & ~n19951 ) | ( n19946 & n20475 ) | ( ~n19951 & n20475 ) ;
  assign n20630 = n19959 &  n20475 ;
  assign n20632 = ( n20475 & ~n20631 ) | ( n20475 & n20630 ) | ( ~n20631 & n20630 ) ;
  assign n20633 = ( n20630 & ~n19946 ) | ( n20630 & n20631 ) | ( ~n19946 & n20631 ) ;
  assign n20634 = ( n19951 & ~n20632 ) | ( n19951 & n20633 ) | ( ~n20632 & n20633 ) ;
  assign n20615 = n19957 | n20475 ;
  assign n20616 = ( n19944 & ~n19953 ) | ( n19944 & n19957 ) | ( ~n19953 & n19957 ) ;
  assign n20617 = ( n19953 & n20615 ) | ( n19953 & n20616 ) | ( n20615 & n20616 ) ;
  assign n20618 = ( n19957 & ~n20616 ) | ( n19957 & n20615 ) | ( ~n20616 & n20615 ) ;
  assign n20619 = ( n19944 & ~n20617 ) | ( n19944 & n20618 ) | ( ~n20617 & n20618 ) ;
  assign n20609 = ( n19924 & ~n19929 ) | ( n19924 & n20475 ) | ( ~n19929 & n20475 ) ;
  assign n20608 = n19937 &  n20475 ;
  assign n20610 = ( n20475 & ~n20609 ) | ( n20475 & n20608 ) | ( ~n20609 & n20608 ) ;
  assign n20611 = ( n20608 & ~n19924 ) | ( n20608 & n20609 ) | ( ~n19924 & n20609 ) ;
  assign n20612 = ( n19929 & ~n20610 ) | ( n19929 & n20611 ) | ( ~n20610 & n20611 ) ;
  assign n20593 = n19935 | n20475 ;
  assign n20594 = ( n19922 & ~n19931 ) | ( n19922 & n19935 ) | ( ~n19931 & n19935 ) ;
  assign n20595 = ( n19931 & n20593 ) | ( n19931 & n20594 ) | ( n20593 & n20594 ) ;
  assign n20596 = ( n19935 & ~n20594 ) | ( n19935 & n20593 ) | ( ~n20594 & n20593 ) ;
  assign n20597 = ( n19922 & ~n20595 ) | ( n19922 & n20596 ) | ( ~n20595 & n20596 ) ;
  assign n20586 = n19915 &  n20475 ;
  assign n20587 = ( n19902 & n19907 ) | ( n19902 & n20475 ) | ( n19907 & n20475 ) ;
  assign n20589 = ( n20586 & ~n19902 ) | ( n20586 & n20587 ) | ( ~n19902 & n20587 ) ;
  assign n20588 = ( n20475 & ~n20587 ) | ( n20475 & n20586 ) | ( ~n20587 & n20586 ) ;
  assign n20590 = ( n19907 & ~n20589 ) | ( n19907 & n20588 ) | ( ~n20589 & n20588 ) ;
  assign n20571 = n19913 | n20475 ;
  assign n20572 = ( n19900 & ~n19913 ) | ( n19900 & n19909 ) | ( ~n19913 & n19909 ) ;
  assign n20574 = ( n19913 & n20571 ) | ( n19913 & n20572 ) | ( n20571 & n20572 ) ;
  assign n20573 = ( n19909 & ~n20572 ) | ( n19909 & n20571 ) | ( ~n20572 & n20571 ) ;
  assign n20575 = ( n19900 & ~n20574 ) | ( n19900 & n20573 ) | ( ~n20574 & n20573 ) ;
  assign n20565 = ( n19880 & ~n19885 ) | ( n19880 & n20475 ) | ( ~n19885 & n20475 ) ;
  assign n20564 = n19893 &  n20475 ;
  assign n20566 = ( n20475 & ~n20565 ) | ( n20475 & n20564 ) | ( ~n20565 & n20564 ) ;
  assign n20567 = ( n20564 & ~n19880 ) | ( n20564 & n20565 ) | ( ~n19880 & n20565 ) ;
  assign n20568 = ( n19885 & ~n20566 ) | ( n19885 & n20567 ) | ( ~n20566 & n20567 ) ;
  assign n20549 = n19891 | n20475 ;
  assign n20550 = ( n19878 & ~n19891 ) | ( n19878 & n19887 ) | ( ~n19891 & n19887 ) ;
  assign n20552 = ( n19891 & n20549 ) | ( n19891 & n20550 ) | ( n20549 & n20550 ) ;
  assign n20551 = ( n19887 & ~n20550 ) | ( n19887 & n20549 ) | ( ~n20550 & n20549 ) ;
  assign n20553 = ( n19878 & ~n20552 ) | ( n19878 & n20551 ) | ( ~n20552 & n20551 ) ;
  assign n20542 = n19858 | n20475 ;
  assign n20543 = ( n19863 & ~n19858 ) | ( n19863 & n19871 ) | ( ~n19858 & n19871 ) ;
  assign n20545 = ( n19858 & n20542 ) | ( n19858 & n20543 ) | ( n20542 & n20543 ) ;
  assign n20544 = ( n19871 & ~n20543 ) | ( n19871 & n20542 ) | ( ~n20543 & n20542 ) ;
  assign n20546 = ( n19863 & ~n20545 ) | ( n19863 & n20544 ) | ( ~n20545 & n20544 ) ;
  assign n20527 = n19869 | n20475 ;
  assign n20528 = ( n19856 & ~n19865 ) | ( n19856 & n19869 ) | ( ~n19865 & n19869 ) ;
  assign n20529 = ( n19865 & n20527 ) | ( n19865 & n20528 ) | ( n20527 & n20528 ) ;
  assign n20530 = ( n19869 & ~n20528 ) | ( n19869 & n20527 ) | ( ~n20528 & n20527 ) ;
  assign n20531 = ( n19856 & ~n20529 ) | ( n19856 & n20530 ) | ( ~n20529 & n20530 ) ;
  assign n20520 = ( n19833 & ~n19835 ) | ( n19833 & 1'b0 ) | ( ~n19835 & 1'b0 ) ;
  assign n20521 = ( n19835 & ~n20520 ) | ( n19835 & n19844 ) | ( ~n20520 & n19844 ) ;
  assign n20523 = ( n20475 & n20520 ) | ( n20475 & n20521 ) | ( n20520 & n20521 ) ;
  assign n20522 = ( n19835 & ~n20521 ) | ( n19835 & n20475 ) | ( ~n20521 & n20475 ) ;
  assign n20524 = ( n19844 & ~n20523 ) | ( n19844 & n20522 ) | ( ~n20523 & n20522 ) ;
  assign n20504 = ~x10 & n19819 ;
  assign n20505 = ( x11 & ~n20504 ) | ( x11 & 1'b0 ) | ( ~n20504 & 1'b0 ) ;
  assign n20506 = n19836 | n20505 ;
  assign n20501 = ( n19819 & ~x10 ) | ( n19819 & n19828 ) | ( ~x10 & n19828 ) ;
  assign n20502 = x10 &  n20501 ;
  assign n20503 = ( n19823 & ~n20502 ) | ( n19823 & n19828 ) | ( ~n20502 & n19828 ) ;
  assign n20507 = ( n20475 & ~n20506 ) | ( n20475 & n20503 ) | ( ~n20506 & n20503 ) ;
  assign n20509 = ( n20475 & ~n20507 ) | ( n20475 & 1'b0 ) | ( ~n20507 & 1'b0 ) ;
  assign n20508 = ~n20503 & n20507 ;
  assign n20510 = ( n20506 & ~n20509 ) | ( n20506 & n20508 ) | ( ~n20509 & n20508 ) ;
  assign n20491 = ( n19819 & ~n20473 ) | ( n19819 & 1'b0 ) | ( ~n20473 & 1'b0 ) ;
  assign n20492 = ( n20469 & ~n20461 ) | ( n20469 & n20491 ) | ( ~n20461 & n20491 ) ;
  assign n20493 = n20461 &  n20492 ;
  assign n20490 = ~n19820 & n20475 ;
  assign n20494 = ~n20493 & n20490 ;
  assign n20495 = ( x10 & n20494 ) | ( x10 & n20493 ) | ( n20494 & n20493 ) ;
  assign n20496 = x10 | n20493 ;
  assign n20497 = n20490 | n20496 ;
  assign n20498 = ~n20495 & n20497 ;
  assign n20482 = ( x8 & ~n20475 ) | ( x8 & x9 ) | ( ~n20475 & x9 ) ;
  assign n20487 = ( x8 & ~x9 ) | ( x8 & 1'b0 ) | ( ~x9 & 1'b0 ) ;
  assign n20478 = x6 | x7 ;
  assign n20483 = ~x8 & n20478 ;
  assign n20484 = ( x8 & n20483 ) | ( x8 & n19818 ) | ( n20483 & n19818 ) ;
  assign n20485 = n19805 &  n20484 ;
  assign n20486 = ( n20475 & ~x9 ) | ( n20475 & n20485 ) | ( ~x9 & n20485 ) ;
  assign n20488 = ( n20482 & ~n20487 ) | ( n20482 & n20486 ) | ( ~n20487 & n20486 ) ;
  assign n20479 = x8 | n20478 ;
  assign n20480 = x8 &  n20475 ;
  assign n20481 = ( n19819 & ~n20479 ) | ( n19819 & n20480 ) | ( ~n20479 & n20480 ) ;
  assign n20511 = n19175 | n20481 ;
  assign n20512 = ( n20488 & ~n20511 ) | ( n20488 & 1'b0 ) | ( ~n20511 & 1'b0 ) ;
  assign n20513 = n20498 | n20512 ;
  assign n20514 = n20481 &  n20488 ;
  assign n20515 = ( n19175 & ~n20488 ) | ( n19175 & n20514 ) | ( ~n20488 & n20514 ) ;
  assign n20516 = n18532 | n20515 ;
  assign n20517 = ( n20513 & ~n20516 ) | ( n20513 & 1'b0 ) | ( ~n20516 & 1'b0 ) ;
  assign n20518 = n20510 | n20517 ;
  assign n20489 = ~n20481 & n20488 ;
  assign n20499 = ( n20489 & ~n19175 ) | ( n20489 & n20498 ) | ( ~n19175 & n20498 ) ;
  assign n20500 = ( n18532 & ~n20499 ) | ( n18532 & 1'b0 ) | ( ~n20499 & 1'b0 ) ;
  assign n20532 = n17902 | n20500 ;
  assign n20533 = ( n20518 & ~n20532 ) | ( n20518 & 1'b0 ) | ( ~n20532 & 1'b0 ) ;
  assign n20534 = n20524 | n20533 ;
  assign n20535 = ( n20513 & ~n20515 ) | ( n20513 & 1'b0 ) | ( ~n20515 & 1'b0 ) ;
  assign n20536 = ( n20510 & ~n18532 ) | ( n20510 & n20535 ) | ( ~n18532 & n20535 ) ;
  assign n20537 = ( n17902 & ~n20536 ) | ( n17902 & 1'b0 ) | ( ~n20536 & 1'b0 ) ;
  assign n20538 = n17279 | n20537 ;
  assign n20539 = ( n20534 & ~n20538 ) | ( n20534 & 1'b0 ) | ( ~n20538 & 1'b0 ) ;
  assign n20540 = n20531 | n20539 ;
  assign n20519 = ~n20500 & n20518 ;
  assign n20525 = ( n20519 & ~n17902 ) | ( n20519 & n20524 ) | ( ~n17902 & n20524 ) ;
  assign n20526 = ( n17279 & ~n20525 ) | ( n17279 & 1'b0 ) | ( ~n20525 & 1'b0 ) ;
  assign n20554 = n16671 | n20526 ;
  assign n20555 = ( n20540 & ~n20554 ) | ( n20540 & 1'b0 ) | ( ~n20554 & 1'b0 ) ;
  assign n20556 = n20546 | n20555 ;
  assign n20557 = ( n20534 & ~n20537 ) | ( n20534 & 1'b0 ) | ( ~n20537 & 1'b0 ) ;
  assign n20558 = ( n20531 & ~n17279 ) | ( n20531 & n20557 ) | ( ~n17279 & n20557 ) ;
  assign n20559 = ( n16671 & ~n20558 ) | ( n16671 & 1'b0 ) | ( ~n20558 & 1'b0 ) ;
  assign n20560 = n16070 | n20559 ;
  assign n20561 = ( n20556 & ~n20560 ) | ( n20556 & 1'b0 ) | ( ~n20560 & 1'b0 ) ;
  assign n20562 = n20553 | n20561 ;
  assign n20541 = ~n20526 & n20540 ;
  assign n20547 = ( n20541 & ~n16671 ) | ( n20541 & n20546 ) | ( ~n16671 & n20546 ) ;
  assign n20548 = ( n16070 & ~n20547 ) | ( n16070 & 1'b0 ) | ( ~n20547 & 1'b0 ) ;
  assign n20576 = n15484 | n20548 ;
  assign n20577 = ( n20562 & ~n20576 ) | ( n20562 & 1'b0 ) | ( ~n20576 & 1'b0 ) ;
  assign n20578 = n20568 | n20577 ;
  assign n20579 = ( n20556 & ~n20559 ) | ( n20556 & 1'b0 ) | ( ~n20559 & 1'b0 ) ;
  assign n20580 = ( n20553 & ~n16070 ) | ( n20553 & n20579 ) | ( ~n16070 & n20579 ) ;
  assign n20581 = ( n15484 & ~n20580 ) | ( n15484 & 1'b0 ) | ( ~n20580 & 1'b0 ) ;
  assign n20582 = n14905 | n20581 ;
  assign n20583 = ( n20578 & ~n20582 ) | ( n20578 & 1'b0 ) | ( ~n20582 & 1'b0 ) ;
  assign n20584 = n20575 | n20583 ;
  assign n20563 = ~n20548 & n20562 ;
  assign n20569 = ( n20563 & ~n15484 ) | ( n20563 & n20568 ) | ( ~n15484 & n20568 ) ;
  assign n20570 = ( n14905 & ~n20569 ) | ( n14905 & 1'b0 ) | ( ~n20569 & 1'b0 ) ;
  assign n20598 = n14341 | n20570 ;
  assign n20599 = ( n20584 & ~n20598 ) | ( n20584 & 1'b0 ) | ( ~n20598 & 1'b0 ) ;
  assign n20600 = n20590 | n20599 ;
  assign n20601 = ( n20578 & ~n20581 ) | ( n20578 & 1'b0 ) | ( ~n20581 & 1'b0 ) ;
  assign n20602 = ( n20575 & ~n14905 ) | ( n20575 & n20601 ) | ( ~n14905 & n20601 ) ;
  assign n20603 = ( n14341 & ~n20602 ) | ( n14341 & 1'b0 ) | ( ~n20602 & 1'b0 ) ;
  assign n20604 = n13784 | n20603 ;
  assign n20605 = ( n20600 & ~n20604 ) | ( n20600 & 1'b0 ) | ( ~n20604 & 1'b0 ) ;
  assign n20606 = n20597 | n20605 ;
  assign n20585 = ~n20570 & n20584 ;
  assign n20591 = ( n20585 & ~n14341 ) | ( n20585 & n20590 ) | ( ~n14341 & n20590 ) ;
  assign n20592 = ( n13784 & ~n20591 ) | ( n13784 & 1'b0 ) | ( ~n20591 & 1'b0 ) ;
  assign n20620 = n13242 | n20592 ;
  assign n20621 = ( n20606 & ~n20620 ) | ( n20606 & 1'b0 ) | ( ~n20620 & 1'b0 ) ;
  assign n20622 = n20612 | n20621 ;
  assign n20623 = ( n20600 & ~n20603 ) | ( n20600 & 1'b0 ) | ( ~n20603 & 1'b0 ) ;
  assign n20624 = ( n20597 & ~n13784 ) | ( n20597 & n20623 ) | ( ~n13784 & n20623 ) ;
  assign n20625 = ( n13242 & ~n20624 ) | ( n13242 & 1'b0 ) | ( ~n20624 & 1'b0 ) ;
  assign n20626 = n12707 | n20625 ;
  assign n20627 = ( n20622 & ~n20626 ) | ( n20622 & 1'b0 ) | ( ~n20626 & 1'b0 ) ;
  assign n20628 = n20619 | n20627 ;
  assign n20607 = ~n20592 & n20606 ;
  assign n20613 = ( n20607 & ~n13242 ) | ( n20607 & n20612 ) | ( ~n13242 & n20612 ) ;
  assign n20614 = ( n12707 & ~n20613 ) | ( n12707 & 1'b0 ) | ( ~n20613 & 1'b0 ) ;
  assign n20642 = n12187 | n20614 ;
  assign n20643 = ( n20628 & ~n20642 ) | ( n20628 & 1'b0 ) | ( ~n20642 & 1'b0 ) ;
  assign n20644 = n20634 | n20643 ;
  assign n20645 = ( n20622 & ~n20625 ) | ( n20622 & 1'b0 ) | ( ~n20625 & 1'b0 ) ;
  assign n20646 = ( n20619 & ~n12707 ) | ( n20619 & n20645 ) | ( ~n12707 & n20645 ) ;
  assign n20647 = ( n12187 & ~n20646 ) | ( n12187 & 1'b0 ) | ( ~n20646 & 1'b0 ) ;
  assign n20648 = n11674 | n20647 ;
  assign n20649 = ( n20644 & ~n20648 ) | ( n20644 & 1'b0 ) | ( ~n20648 & 1'b0 ) ;
  assign n20650 = n20641 | n20649 ;
  assign n20629 = ~n20614 & n20628 ;
  assign n20635 = ( n20629 & ~n12187 ) | ( n20629 & n20634 ) | ( ~n12187 & n20634 ) ;
  assign n20636 = ( n11674 & ~n20635 ) | ( n11674 & 1'b0 ) | ( ~n20635 & 1'b0 ) ;
  assign n20664 = n11176 | n20636 ;
  assign n20665 = ( n20650 & ~n20664 ) | ( n20650 & 1'b0 ) | ( ~n20664 & 1'b0 ) ;
  assign n20666 = n20656 | n20665 ;
  assign n20667 = ( n20644 & ~n20647 ) | ( n20644 & 1'b0 ) | ( ~n20647 & 1'b0 ) ;
  assign n20668 = ( n20641 & ~n11674 ) | ( n20641 & n20667 ) | ( ~n11674 & n20667 ) ;
  assign n20669 = ( n11176 & ~n20668 ) | ( n11176 & 1'b0 ) | ( ~n20668 & 1'b0 ) ;
  assign n20670 = n10685 | n20669 ;
  assign n20671 = ( n20666 & ~n20670 ) | ( n20666 & 1'b0 ) | ( ~n20670 & 1'b0 ) ;
  assign n20672 = n20663 | n20671 ;
  assign n20651 = ~n20636 & n20650 ;
  assign n20657 = ( n20651 & ~n11176 ) | ( n20651 & n20656 ) | ( ~n11176 & n20656 ) ;
  assign n20658 = ( n10685 & ~n20657 ) | ( n10685 & 1'b0 ) | ( ~n20657 & 1'b0 ) ;
  assign n20686 = n10209 | n20658 ;
  assign n20687 = ( n20672 & ~n20686 ) | ( n20672 & 1'b0 ) | ( ~n20686 & 1'b0 ) ;
  assign n20688 = n20678 | n20687 ;
  assign n20689 = ( n20666 & ~n20669 ) | ( n20666 & 1'b0 ) | ( ~n20669 & 1'b0 ) ;
  assign n20690 = ( n20663 & ~n10685 ) | ( n20663 & n20689 ) | ( ~n10685 & n20689 ) ;
  assign n20691 = ( n10209 & ~n20690 ) | ( n10209 & 1'b0 ) | ( ~n20690 & 1'b0 ) ;
  assign n20692 = ( n9740 & ~n20691 ) | ( n9740 & 1'b0 ) | ( ~n20691 & 1'b0 ) ;
  assign n20693 = n20688 &  n20692 ;
  assign n20694 = n20685 | n20693 ;
  assign n20673 = ~n20658 & n20672 ;
  assign n20679 = ( n20673 & ~n10209 ) | ( n20673 & n20678 ) | ( ~n10209 & n20678 ) ;
  assign n20680 = n9740 | n20679 ;
  assign n20708 = ~n9286 & n20680 ;
  assign n20709 = n20694 &  n20708 ;
  assign n20710 = n20700 | n20709 ;
  assign n20711 = ( n20688 & ~n20691 ) | ( n20688 & 1'b0 ) | ( ~n20691 & 1'b0 ) ;
  assign n20712 = ( n9740 & n20685 ) | ( n9740 & n20711 ) | ( n20685 & n20711 ) ;
  assign n20713 = ( n9286 & ~n20712 ) | ( n9286 & 1'b0 ) | ( ~n20712 & 1'b0 ) ;
  assign n20714 = n8839 | n20713 ;
  assign n20715 = ( n20710 & ~n20714 ) | ( n20710 & 1'b0 ) | ( ~n20714 & 1'b0 ) ;
  assign n20716 = n20707 | n20715 ;
  assign n20695 = n20680 &  n20694 ;
  assign n20701 = ( n20695 & ~n9286 ) | ( n20695 & n20700 ) | ( ~n9286 & n20700 ) ;
  assign n20702 = ( n8839 & ~n20701 ) | ( n8839 & 1'b0 ) | ( ~n20701 & 1'b0 ) ;
  assign n20730 = n8407 | n20702 ;
  assign n20731 = ( n20716 & ~n20730 ) | ( n20716 & 1'b0 ) | ( ~n20730 & 1'b0 ) ;
  assign n20732 = n20722 | n20731 ;
  assign n20733 = ( n20710 & ~n20713 ) | ( n20710 & 1'b0 ) | ( ~n20713 & 1'b0 ) ;
  assign n20734 = ( n20707 & ~n8839 ) | ( n20707 & n20733 ) | ( ~n8839 & n20733 ) ;
  assign n20735 = ( n8407 & ~n20734 ) | ( n8407 & 1'b0 ) | ( ~n20734 & 1'b0 ) ;
  assign n20736 = n7982 | n20735 ;
  assign n20737 = ( n20732 & ~n20736 ) | ( n20732 & 1'b0 ) | ( ~n20736 & 1'b0 ) ;
  assign n20738 = n20729 | n20737 ;
  assign n20717 = ~n20702 & n20716 ;
  assign n20723 = ( n20717 & ~n8407 ) | ( n20717 & n20722 ) | ( ~n8407 & n20722 ) ;
  assign n20724 = ( n7982 & ~n20723 ) | ( n7982 & 1'b0 ) | ( ~n20723 & 1'b0 ) ;
  assign n20752 = ( n7572 & ~n20724 ) | ( n7572 & 1'b0 ) | ( ~n20724 & 1'b0 ) ;
  assign n20753 = n20738 &  n20752 ;
  assign n20754 = n20744 | n20753 ;
  assign n20755 = ( n20732 & ~n20735 ) | ( n20732 & 1'b0 ) | ( ~n20735 & 1'b0 ) ;
  assign n20756 = ( n20729 & ~n7982 ) | ( n20729 & n20755 ) | ( ~n7982 & n20755 ) ;
  assign n20757 = n7572 | n20756 ;
  assign n20758 = n7169 &  n20757 ;
  assign n20759 = n20754 &  n20758 ;
  assign n20760 = n20751 | n20759 ;
  assign n20739 = ~n20724 & n20738 ;
  assign n20745 = ( n7572 & n20739 ) | ( n7572 & n20744 ) | ( n20739 & n20744 ) ;
  assign n20746 = n7169 | n20745 ;
  assign n20774 = ~n6781 & n20746 ;
  assign n20775 = n20760 &  n20774 ;
  assign n20776 = n20766 | n20775 ;
  assign n20777 = n20754 &  n20757 ;
  assign n20778 = ( n7169 & n20751 ) | ( n7169 & n20777 ) | ( n20751 & n20777 ) ;
  assign n20779 = ( n6781 & ~n20778 ) | ( n6781 & 1'b0 ) | ( ~n20778 & 1'b0 ) ;
  assign n20780 = ( n6399 & ~n20779 ) | ( n6399 & 1'b0 ) | ( ~n20779 & 1'b0 ) ;
  assign n20781 = n20776 &  n20780 ;
  assign n20782 = n20773 | n20781 ;
  assign n20761 = n20746 &  n20760 ;
  assign n20767 = ( n20761 & ~n6781 ) | ( n20761 & n20766 ) | ( ~n6781 & n20766 ) ;
  assign n20768 = n6399 | n20767 ;
  assign n20796 = ~n6032 & n20768 ;
  assign n20797 = n20782 &  n20796 ;
  assign n20798 = n20788 | n20797 ;
  assign n20799 = ( n20776 & ~n20779 ) | ( n20776 & 1'b0 ) | ( ~n20779 & 1'b0 ) ;
  assign n20800 = ( n6399 & n20773 ) | ( n6399 & n20799 ) | ( n20773 & n20799 ) ;
  assign n20801 = ( n6032 & ~n20800 ) | ( n6032 & 1'b0 ) | ( ~n20800 & 1'b0 ) ;
  assign n20802 = ( n5672 & ~n20801 ) | ( n5672 & 1'b0 ) | ( ~n20801 & 1'b0 ) ;
  assign n20803 = n20798 &  n20802 ;
  assign n20804 = n20795 | n20803 ;
  assign n20783 = n20768 &  n20782 ;
  assign n20789 = ( n20783 & ~n6032 ) | ( n20783 & n20788 ) | ( ~n6032 & n20788 ) ;
  assign n20790 = n5672 | n20789 ;
  assign n20818 = ~n5327 & n20790 ;
  assign n20819 = n20804 &  n20818 ;
  assign n20820 = n20810 | n20819 ;
  assign n20821 = ( n20798 & ~n20801 ) | ( n20798 & 1'b0 ) | ( ~n20801 & 1'b0 ) ;
  assign n20822 = ( n5672 & n20795 ) | ( n5672 & n20821 ) | ( n20795 & n20821 ) ;
  assign n20823 = ( n5327 & ~n20822 ) | ( n5327 & 1'b0 ) | ( ~n20822 & 1'b0 ) ;
  assign n20824 = n4990 | n20823 ;
  assign n20825 = ( n20820 & ~n20824 ) | ( n20820 & 1'b0 ) | ( ~n20824 & 1'b0 ) ;
  assign n20826 = n20817 | n20825 ;
  assign n20805 = n20790 &  n20804 ;
  assign n20811 = ( n20805 & ~n5327 ) | ( n20805 & n20810 ) | ( ~n5327 & n20810 ) ;
  assign n20812 = ( n4990 & ~n20811 ) | ( n4990 & 1'b0 ) | ( ~n20811 & 1'b0 ) ;
  assign n20840 = n4668 | n20812 ;
  assign n20841 = ( n20826 & ~n20840 ) | ( n20826 & 1'b0 ) | ( ~n20840 & 1'b0 ) ;
  assign n20842 = n20832 | n20841 ;
  assign n20843 = ( n20820 & ~n20823 ) | ( n20820 & 1'b0 ) | ( ~n20823 & 1'b0 ) ;
  assign n20844 = ( n20817 & ~n4990 ) | ( n20817 & n20843 ) | ( ~n4990 & n20843 ) ;
  assign n20845 = ( n4668 & ~n20844 ) | ( n4668 & 1'b0 ) | ( ~n20844 & 1'b0 ) ;
  assign n20846 = n4353 | n20845 ;
  assign n20847 = ( n20842 & ~n20846 ) | ( n20842 & 1'b0 ) | ( ~n20846 & 1'b0 ) ;
  assign n20848 = n20839 | n20847 ;
  assign n20827 = ~n20812 & n20826 ;
  assign n20833 = ( n20827 & ~n4668 ) | ( n20827 & n20832 ) | ( ~n4668 & n20832 ) ;
  assign n20834 = ( n4353 & ~n20833 ) | ( n4353 & 1'b0 ) | ( ~n20833 & 1'b0 ) ;
  assign n20862 = n4053 | n20834 ;
  assign n20863 = ( n20848 & ~n20862 ) | ( n20848 & 1'b0 ) | ( ~n20862 & 1'b0 ) ;
  assign n20864 = n20854 | n20863 ;
  assign n20865 = ( n20842 & ~n20845 ) | ( n20842 & 1'b0 ) | ( ~n20845 & 1'b0 ) ;
  assign n20866 = ( n20839 & ~n4353 ) | ( n20839 & n20865 ) | ( ~n4353 & n20865 ) ;
  assign n20867 = ( n4053 & ~n20866 ) | ( n4053 & 1'b0 ) | ( ~n20866 & 1'b0 ) ;
  assign n20868 = n3760 | n20867 ;
  assign n20869 = ( n20864 & ~n20868 ) | ( n20864 & 1'b0 ) | ( ~n20868 & 1'b0 ) ;
  assign n20870 = n20861 | n20869 ;
  assign n20849 = ~n20834 & n20848 ;
  assign n20855 = ( n20849 & ~n4053 ) | ( n20849 & n20854 ) | ( ~n4053 & n20854 ) ;
  assign n20856 = ( n3760 & ~n20855 ) | ( n3760 & 1'b0 ) | ( ~n20855 & 1'b0 ) ;
  assign n20884 = n3482 | n20856 ;
  assign n20885 = ( n20870 & ~n20884 ) | ( n20870 & 1'b0 ) | ( ~n20884 & 1'b0 ) ;
  assign n20886 = n20876 | n20885 ;
  assign n20887 = ( n20864 & ~n20867 ) | ( n20864 & 1'b0 ) | ( ~n20867 & 1'b0 ) ;
  assign n20888 = ( n20861 & ~n3760 ) | ( n20861 & n20887 ) | ( ~n3760 & n20887 ) ;
  assign n20889 = ( n3482 & ~n20888 ) | ( n3482 & 1'b0 ) | ( ~n20888 & 1'b0 ) ;
  assign n20890 = n3211 | n20889 ;
  assign n20891 = ( n20886 & ~n20890 ) | ( n20886 & 1'b0 ) | ( ~n20890 & 1'b0 ) ;
  assign n20892 = n20883 | n20891 ;
  assign n20871 = ~n20856 & n20870 ;
  assign n20877 = ( n20871 & ~n3482 ) | ( n20871 & n20876 ) | ( ~n3482 & n20876 ) ;
  assign n20878 = ( n3211 & ~n20877 ) | ( n3211 & 1'b0 ) | ( ~n20877 & 1'b0 ) ;
  assign n20906 = n2955 | n20878 ;
  assign n20907 = ( n20892 & ~n20906 ) | ( n20892 & 1'b0 ) | ( ~n20906 & 1'b0 ) ;
  assign n20908 = n20898 | n20907 ;
  assign n20909 = ( n20886 & ~n20889 ) | ( n20886 & 1'b0 ) | ( ~n20889 & 1'b0 ) ;
  assign n20910 = ( n20883 & ~n3211 ) | ( n20883 & n20909 ) | ( ~n3211 & n20909 ) ;
  assign n20911 = ( n2955 & ~n20910 ) | ( n2955 & 1'b0 ) | ( ~n20910 & 1'b0 ) ;
  assign n20912 = n2706 | n20911 ;
  assign n20913 = ( n20908 & ~n20912 ) | ( n20908 & 1'b0 ) | ( ~n20912 & 1'b0 ) ;
  assign n20914 = ( n20905 & ~n20913 ) | ( n20905 & 1'b0 ) | ( ~n20913 & 1'b0 ) ;
  assign n20893 = ~n20878 & n20892 ;
  assign n20899 = ( n20893 & ~n2955 ) | ( n20893 & n20898 ) | ( ~n2955 & n20898 ) ;
  assign n20900 = ( n2706 & ~n20899 ) | ( n2706 & 1'b0 ) | ( ~n20899 & 1'b0 ) ;
  assign n20928 = n2472 | n20900 ;
  assign n20929 = n20914 | n20928 ;
  assign n20930 = n20920 &  n20929 ;
  assign n20931 = ( n20908 & ~n20911 ) | ( n20908 & 1'b0 ) | ( ~n20911 & 1'b0 ) ;
  assign n20932 = ( n2706 & ~n20931 ) | ( n2706 & n20905 ) | ( ~n20931 & n20905 ) ;
  assign n20933 = n2472 &  n20932 ;
  assign n20934 = n2245 | n20933 ;
  assign n20935 = n20930 | n20934 ;
  assign n20936 = n20927 &  n20935 ;
  assign n20915 = n20900 | n20914 ;
  assign n20921 = ( n2472 & n20915 ) | ( n2472 & n20920 ) | ( n20915 & n20920 ) ;
  assign n20922 = n2245 &  n20921 ;
  assign n20950 = ( n2033 & ~n20922 ) | ( n2033 & 1'b0 ) | ( ~n20922 & 1'b0 ) ;
  assign n20951 = ~n20936 & n20950 ;
  assign n20952 = ( n20942 & ~n20951 ) | ( n20942 & 1'b0 ) | ( ~n20951 & 1'b0 ) ;
  assign n20953 = n20930 | n20933 ;
  assign n20954 = ( n2245 & n20927 ) | ( n2245 & n20953 ) | ( n20927 & n20953 ) ;
  assign n20955 = ~n2033 & n20954 ;
  assign n20956 = n1827 | n20955 ;
  assign n20957 = n20952 | n20956 ;
  assign n20958 = n20949 &  n20957 ;
  assign n20937 = n20922 | n20936 ;
  assign n20943 = ( n20937 & ~n2033 ) | ( n20937 & n20942 ) | ( ~n2033 & n20942 ) ;
  assign n20944 = n1827 &  n20943 ;
  assign n20972 = ( n1636 & ~n20944 ) | ( n1636 & 1'b0 ) | ( ~n20944 & 1'b0 ) ;
  assign n20973 = ~n20958 & n20972 ;
  assign n20974 = n20964 | n20973 ;
  assign n20975 = n20952 | n20955 ;
  assign n20976 = ( n1827 & n20949 ) | ( n1827 & n20975 ) | ( n20949 & n20975 ) ;
  assign n20977 = ~n1636 & n20976 ;
  assign n20978 = ( n1452 & ~n20977 ) | ( n1452 & 1'b0 ) | ( ~n20977 & 1'b0 ) ;
  assign n20979 = n20974 &  n20978 ;
  assign n20980 = n20971 | n20979 ;
  assign n20959 = n20944 | n20958 ;
  assign n20965 = ( n1636 & ~n20959 ) | ( n1636 & n20964 ) | ( ~n20959 & n20964 ) ;
  assign n20966 = n1452 | n20965 ;
  assign n20994 = ~n1283 & n20966 ;
  assign n20995 = n20980 &  n20994 ;
  assign n20996 = ( n20986 & ~n20995 ) | ( n20986 & 1'b0 ) | ( ~n20995 & 1'b0 ) ;
  assign n20997 = ( n20974 & ~n20977 ) | ( n20974 & 1'b0 ) | ( ~n20977 & 1'b0 ) ;
  assign n20998 = ( n1452 & n20971 ) | ( n1452 & n20997 ) | ( n20971 & n20997 ) ;
  assign n20999 = ( n1283 & ~n20998 ) | ( n1283 & 1'b0 ) | ( ~n20998 & 1'b0 ) ;
  assign n21000 = ( n1122 & ~n20999 ) | ( n1122 & 1'b0 ) | ( ~n20999 & 1'b0 ) ;
  assign n21001 = ~n20996 & n21000 ;
  assign n21002 = n20993 | n21001 ;
  assign n20981 = n20966 &  n20980 ;
  assign n20987 = ( n1283 & ~n20981 ) | ( n1283 & n20986 ) | ( ~n20981 & n20986 ) ;
  assign n20988 = ~n1122 & n20987 ;
  assign n21016 = ( n976 & ~n20988 ) | ( n976 & 1'b0 ) | ( ~n20988 & 1'b0 ) ;
  assign n21017 = n21002 &  n21016 ;
  assign n21018 = ( n21008 & ~n21017 ) | ( n21008 & 1'b0 ) | ( ~n21017 & 1'b0 ) ;
  assign n21019 = n20996 | n20999 ;
  assign n21020 = ( n1122 & ~n21019 ) | ( n1122 & n20993 ) | ( ~n21019 & n20993 ) ;
  assign n21021 = n976 | n21020 ;
  assign n21022 = ~n837 & n21021 ;
  assign n21023 = ~n21018 & n21022 ;
  assign n21024 = ( n21015 & ~n21023 ) | ( n21015 & 1'b0 ) | ( ~n21023 & 1'b0 ) ;
  assign n21003 = ~n20988 & n21002 ;
  assign n21009 = ( n976 & ~n21008 ) | ( n976 & n21003 ) | ( ~n21008 & n21003 ) ;
  assign n21010 = ( n837 & ~n21009 ) | ( n837 & 1'b0 ) | ( ~n21009 & 1'b0 ) ;
  assign n21038 = n713 | n21010 ;
  assign n21039 = n21024 | n21038 ;
  assign n21040 = ~n21030 & n21039 ;
  assign n21041 = ~n21018 & n21021 ;
  assign n21042 = ( n837 & ~n21041 ) | ( n837 & n21015 ) | ( ~n21041 & n21015 ) ;
  assign n21043 = n713 &  n21042 ;
  assign n21044 = n595 | n21043 ;
  assign n21045 = n21040 | n21044 ;
  assign n21046 = ~n21037 & n21045 ;
  assign n21025 = n21010 | n21024 ;
  assign n21031 = ( n713 & ~n21030 ) | ( n713 & n21025 ) | ( ~n21030 & n21025 ) ;
  assign n21032 = n595 &  n21031 ;
  assign n21060 = n492 | n21032 ;
  assign n21061 = n21046 | n21060 ;
  assign n21062 = ~n21052 & n21061 ;
  assign n21063 = n21040 | n21043 ;
  assign n21064 = ( n595 & ~n21037 ) | ( n595 & n21063 ) | ( ~n21037 & n21063 ) ;
  assign n21065 = n492 &  n21064 ;
  assign n21066 = n396 | n21065 ;
  assign n21067 = n21062 | n21066 ;
  assign n21068 = ~n21059 & n21067 ;
  assign n21047 = n21032 | n21046 ;
  assign n21053 = ( n492 & ~n21052 ) | ( n492 & n21047 ) | ( ~n21052 & n21047 ) ;
  assign n21054 = n396 &  n21053 ;
  assign n21082 = n315 | n21054 ;
  assign n21083 = n21068 | n21082 ;
  assign n21084 = ~n21074 & n21083 ;
  assign n21085 = n21062 | n21065 ;
  assign n21086 = ( n396 & ~n21059 ) | ( n396 & n21085 ) | ( ~n21059 & n21085 ) ;
  assign n21087 = n315 &  n21086 ;
  assign n21102 = n21084 | n21087 ;
  assign n21103 = ( n240 & n21081 ) | ( n240 & n21102 ) | ( n21081 & n21102 ) ;
  assign n21104 = n181 &  n21103 ;
  assign n21069 = n21054 | n21068 ;
  assign n21075 = ( n315 & ~n21074 ) | ( n315 & n21069 ) | ( ~n21074 & n21069 ) ;
  assign n21076 = n240 &  n21075 ;
  assign n21088 = n240 | n21087 ;
  assign n21089 = n21084 | n21088 ;
  assign n21090 = n21081 &  n21089 ;
  assign n21091 = n21076 | n21090 ;
  assign n21097 = ( n181 & ~n21096 ) | ( n181 & n21091 ) | ( ~n21096 & n21091 ) ;
  assign n21098 = ~n145 & n21097 ;
  assign n21099 = n181 | n21076 ;
  assign n21100 = n21090 | n21099 ;
  assign n21101 = ~n21096 & n21100 ;
  assign n21105 = ( n145 & ~n21104 ) | ( n145 & 1'b0 ) | ( ~n21104 & 1'b0 ) ;
  assign n21106 = ~n21101 & n21105 ;
  assign n21107 = ( n20436 & ~n20427 ) | ( n20436 & n20440 ) | ( ~n20427 & n20440 ) ;
  assign n21109 = ( n20440 & ~n21107 ) | ( n20440 & n20475 ) | ( ~n21107 & n20475 ) ;
  assign n21108 = ( n20475 & ~n20436 ) | ( n20475 & n21107 ) | ( ~n20436 & n21107 ) ;
  assign n21110 = ( n20427 & ~n21109 ) | ( n20427 & n21108 ) | ( ~n21109 & n21108 ) ;
  assign n21111 = n21106 | n21110 ;
  assign n21112 = ~n21098 & n21111 ;
  assign n21113 = n20429 | n20475 ;
  assign n21114 = ( n20434 & ~n20429 ) | ( n20434 & n20442 ) | ( ~n20429 & n20442 ) ;
  assign n21116 = ( n20429 & n21113 ) | ( n20429 & n21114 ) | ( n21113 & n21114 ) ;
  assign n21115 = ( n20442 & ~n21114 ) | ( n20442 & n21113 ) | ( ~n21114 & n21113 ) ;
  assign n21117 = ( n20434 & ~n21116 ) | ( n20434 & n21115 ) | ( ~n21116 & n21115 ) ;
  assign n21118 = ( n150 & ~n21112 ) | ( n150 & n21117 ) | ( ~n21112 & n21117 ) ;
  assign n21120 = ( n20463 & ~n20449 ) | ( n20463 & n20466 ) | ( ~n20449 & n20466 ) ;
  assign n21119 = n20466 | n20475 ;
  assign n21122 = ( n20466 & ~n21120 ) | ( n20466 & n21119 ) | ( ~n21120 & n21119 ) ;
  assign n21121 = ( n21119 & ~n20463 ) | ( n21119 & n21120 ) | ( ~n20463 & n21120 ) ;
  assign n21123 = ( n20449 & ~n21122 ) | ( n20449 & n21121 ) | ( ~n21122 & n21121 ) ;
  assign n21124 = n20450 &  n20455 ;
  assign n21125 = ~n20475 & n21124 ;
  assign n21126 = ( n20469 & ~n21124 ) | ( n20469 & n21125 ) | ( ~n21124 & n21125 ) ;
  assign n21127 = ~n21123 & n21126 ;
  assign n21128 = ~n21118 & n21127 ;
  assign n21129 = ( n133 & ~n21128 ) | ( n133 & n21127 ) | ( ~n21128 & n21127 ) ;
  assign n21132 = n21101 | n21104 ;
  assign n21133 = ( n145 & ~n21132 ) | ( n145 & n21110 ) | ( ~n21132 & n21110 ) ;
  assign n21134 = ( n150 & ~n21133 ) | ( n150 & 1'b0 ) | ( ~n21133 & 1'b0 ) ;
  assign n21135 = ( n21123 & ~n21134 ) | ( n21123 & 1'b0 ) | ( ~n21134 & 1'b0 ) ;
  assign n21130 = n150 | n21098 ;
  assign n21131 = ( n21111 & ~n21130 ) | ( n21111 & 1'b0 ) | ( ~n21130 & 1'b0 ) ;
  assign n21136 = n21117 &  n21131 ;
  assign n21137 = ( n21135 & ~n21117 ) | ( n21135 & n21136 ) | ( ~n21117 & n21136 ) ;
  assign n21139 = ( n133 & n20450 ) | ( n133 & n20455 ) | ( n20450 & n20455 ) ;
  assign n21138 = ( n20450 & ~n20475 ) | ( n20450 & n20455 ) | ( ~n20475 & n20455 ) ;
  assign n21140 = ( n20455 & ~n21138 ) | ( n20455 & 1'b0 ) | ( ~n21138 & 1'b0 ) ;
  assign n21141 = ( n21139 & ~n20455 ) | ( n21139 & n21140 ) | ( ~n20455 & n21140 ) ;
  assign n21142 = n21137 | n21141 ;
  assign n21143 = ~n21129 |  n21142 ;
  assign n21774 = n21104 | n21143 ;
  assign n21775 = ( n21096 & n21100 ) | ( n21096 & n21104 ) | ( n21100 & n21104 ) ;
  assign n21776 = ( n21774 & ~n21100 ) | ( n21774 & n21775 ) | ( ~n21100 & n21775 ) ;
  assign n21777 = ( n21104 & ~n21775 ) | ( n21104 & n21774 ) | ( ~n21775 & n21774 ) ;
  assign n21778 = ( n21096 & ~n21776 ) | ( n21096 & n21777 ) | ( ~n21776 & n21777 ) ;
  assign n21746 = ( n21054 & ~n21059 ) | ( n21054 & n21067 ) | ( ~n21059 & n21067 ) ;
  assign n21745 = n21054 | n21143 ;
  assign n21748 = ( n21054 & ~n21746 ) | ( n21054 & n21745 ) | ( ~n21746 & n21745 ) ;
  assign n21747 = ( n21745 & ~n21067 ) | ( n21745 & n21746 ) | ( ~n21067 & n21746 ) ;
  assign n21749 = ( n21059 & ~n21748 ) | ( n21059 & n21747 ) | ( ~n21748 & n21747 ) ;
  assign n21724 = ( n21032 & ~n21037 ) | ( n21032 & n21045 ) | ( ~n21037 & n21045 ) ;
  assign n21723 = n21032 | n21143 ;
  assign n21726 = ( n21032 & ~n21724 ) | ( n21032 & n21723 ) | ( ~n21724 & n21723 ) ;
  assign n21725 = ( n21723 & ~n21045 ) | ( n21723 & n21724 ) | ( ~n21045 & n21724 ) ;
  assign n21727 = ( n21037 & ~n21726 ) | ( n21037 & n21725 ) | ( ~n21726 & n21725 ) ;
  assign n21146 = ( x6 & ~n21143 ) | ( x6 & x7 ) | ( ~n21143 & x7 ) ;
  assign n21151 = ( x6 & ~x7 ) | ( x6 & 1'b0 ) | ( ~x7 & 1'b0 ) ;
  assign n20476 = x4 | x5 ;
  assign n21147 = ~x6 & n20476 ;
  assign n21148 = ( x6 & n21147 ) | ( x6 & n20474 ) | ( n21147 & n20474 ) ;
  assign n21149 = n20461 &  n21148 ;
  assign n21150 = ( n21143 & ~x7 ) | ( n21143 & n21149 ) | ( ~x7 & n21149 ) ;
  assign n21152 = ( n21146 & ~n21151 ) | ( n21146 & n21150 ) | ( ~n21151 & n21150 ) ;
  assign n20477 = x6 | n20476 ;
  assign n21144 = x6 &  n21143 ;
  assign n21145 = ( n20475 & ~n20477 ) | ( n20475 & n21144 ) | ( ~n20477 & n21144 ) ;
  assign n21153 = n21145 &  n21152 ;
  assign n21154 = ( n19819 & ~n21152 ) | ( n19819 & n21153 ) | ( ~n21152 & n21153 ) ;
  assign n21155 = n19819 | n21145 ;
  assign n21156 = ( n21152 & ~n21155 ) | ( n21152 & 1'b0 ) | ( ~n21155 & 1'b0 ) ;
  assign n21158 = ( n20475 & ~n21141 ) | ( n20475 & 1'b0 ) | ( ~n21141 & 1'b0 ) ;
  assign n21159 = ( n21129 & ~n21158 ) | ( n21129 & n21137 ) | ( ~n21158 & n21137 ) ;
  assign n21160 = ( n21129 & ~n21159 ) | ( n21129 & 1'b0 ) | ( ~n21159 & 1'b0 ) ;
  assign n21157 = ~n20478 & n21143 ;
  assign n21161 = ~n21160 & n21157 ;
  assign n21162 = ( x8 & n21161 ) | ( x8 & n21160 ) | ( n21161 & n21160 ) ;
  assign n21163 = x8 | n21160 ;
  assign n21164 = n21157 | n21163 ;
  assign n21165 = ~n21162 & n21164 ;
  assign n21166 = n21156 | n21165 ;
  assign n21167 = ~n21154 & n21166 ;
  assign n21171 = ~x8 & n20475 ;
  assign n21172 = ( x9 & ~n21171 ) | ( x9 & 1'b0 ) | ( ~n21171 & 1'b0 ) ;
  assign n21173 = n20490 | n21172 ;
  assign n21168 = ( n20475 & ~x8 ) | ( n20475 & n20485 ) | ( ~x8 & n20485 ) ;
  assign n21169 = x8 &  n21168 ;
  assign n21170 = ( n20481 & ~n21169 ) | ( n20481 & n20485 ) | ( ~n21169 & n20485 ) ;
  assign n21174 = ( n21143 & ~n21173 ) | ( n21143 & n21170 ) | ( ~n21173 & n21170 ) ;
  assign n21176 = ( n21143 & ~n21174 ) | ( n21143 & 1'b0 ) | ( ~n21174 & 1'b0 ) ;
  assign n21175 = ~n21170 & n21174 ;
  assign n21177 = ( n21173 & ~n21176 ) | ( n21173 & n21175 ) | ( ~n21176 & n21175 ) ;
  assign n21178 = ( n21167 & ~n19175 ) | ( n21167 & n21177 ) | ( ~n19175 & n21177 ) ;
  assign n21179 = ( n18532 & ~n21178 ) | ( n18532 & 1'b0 ) | ( ~n21178 & 1'b0 ) ;
  assign n21180 = ~n20512 & n20515 ;
  assign n21181 = ( n20498 & ~n21180 ) | ( n20498 & n20512 ) | ( ~n21180 & n20512 ) ;
  assign n21182 = ( n21143 & n21180 ) | ( n21143 & n21181 ) | ( n21180 & n21181 ) ;
  assign n21183 = ( n20512 & ~n21181 ) | ( n20512 & n21143 ) | ( ~n21181 & n21143 ) ;
  assign n21184 = ( n20498 & ~n21182 ) | ( n20498 & n21183 ) | ( ~n21182 & n21183 ) ;
  assign n21185 = n19175 | n21154 ;
  assign n21186 = ( n21166 & ~n21185 ) | ( n21166 & 1'b0 ) | ( ~n21185 & 1'b0 ) ;
  assign n21187 = n21177 | n21186 ;
  assign n21188 = ~n21145 & n21152 ;
  assign n21189 = ( n21165 & ~n19819 ) | ( n21165 & n21188 ) | ( ~n19819 & n21188 ) ;
  assign n21190 = ( n19175 & ~n21189 ) | ( n19175 & 1'b0 ) | ( ~n21189 & 1'b0 ) ;
  assign n21191 = n18532 | n21190 ;
  assign n21192 = ( n21187 & ~n21191 ) | ( n21187 & 1'b0 ) | ( ~n21191 & 1'b0 ) ;
  assign n21193 = n21184 | n21192 ;
  assign n21194 = ~n21179 & n21193 ;
  assign n21195 = n20517 &  n21143 ;
  assign n21196 = ( n20500 & n20510 ) | ( n20500 & n21143 ) | ( n20510 & n21143 ) ;
  assign n21198 = ( n21195 & ~n20500 ) | ( n21195 & n21196 ) | ( ~n20500 & n21196 ) ;
  assign n21197 = ( n21143 & ~n21196 ) | ( n21143 & n21195 ) | ( ~n21196 & n21195 ) ;
  assign n21199 = ( n20510 & ~n21198 ) | ( n20510 & n21197 ) | ( ~n21198 & n21197 ) ;
  assign n21200 = ( n21194 & ~n17902 ) | ( n21194 & n21199 ) | ( ~n17902 & n21199 ) ;
  assign n21201 = ( n17279 & ~n21200 ) | ( n17279 & 1'b0 ) | ( ~n21200 & 1'b0 ) ;
  assign n21202 = n20537 | n21143 ;
  assign n21203 = ( n20524 & ~n20537 ) | ( n20524 & n20533 ) | ( ~n20537 & n20533 ) ;
  assign n21205 = ( n20537 & n21202 ) | ( n20537 & n21203 ) | ( n21202 & n21203 ) ;
  assign n21204 = ( n20533 & ~n21203 ) | ( n20533 & n21202 ) | ( ~n21203 & n21202 ) ;
  assign n21206 = ( n20524 & ~n21205 ) | ( n20524 & n21204 ) | ( ~n21205 & n21204 ) ;
  assign n21207 = n17902 | n21179 ;
  assign n21208 = ( n21193 & ~n21207 ) | ( n21193 & 1'b0 ) | ( ~n21207 & 1'b0 ) ;
  assign n21209 = n21199 | n21208 ;
  assign n21210 = ( n21187 & ~n21190 ) | ( n21187 & 1'b0 ) | ( ~n21190 & 1'b0 ) ;
  assign n21211 = ( n21184 & ~n18532 ) | ( n21184 & n21210 ) | ( ~n18532 & n21210 ) ;
  assign n21212 = ( n17902 & ~n21211 ) | ( n17902 & 1'b0 ) | ( ~n21211 & 1'b0 ) ;
  assign n21213 = n17279 | n21212 ;
  assign n21214 = ( n21209 & ~n21213 ) | ( n21209 & 1'b0 ) | ( ~n21213 & 1'b0 ) ;
  assign n21215 = n21206 | n21214 ;
  assign n21216 = ~n21201 & n21215 ;
  assign n21217 = n20539 &  n21143 ;
  assign n21218 = ( n20526 & n20531 ) | ( n20526 & n21143 ) | ( n20531 & n21143 ) ;
  assign n21220 = ( n21217 & ~n20526 ) | ( n21217 & n21218 ) | ( ~n20526 & n21218 ) ;
  assign n21219 = ( n21143 & ~n21218 ) | ( n21143 & n21217 ) | ( ~n21218 & n21217 ) ;
  assign n21221 = ( n20531 & ~n21220 ) | ( n20531 & n21219 ) | ( ~n21220 & n21219 ) ;
  assign n21222 = ( n21216 & ~n16671 ) | ( n21216 & n21221 ) | ( ~n16671 & n21221 ) ;
  assign n21223 = ( n16070 & ~n21222 ) | ( n16070 & 1'b0 ) | ( ~n21222 & 1'b0 ) ;
  assign n21224 = n20559 | n21143 ;
  assign n21225 = ( n20546 & ~n20555 ) | ( n20546 & n20559 ) | ( ~n20555 & n20559 ) ;
  assign n21226 = ( n20555 & n21224 ) | ( n20555 & n21225 ) | ( n21224 & n21225 ) ;
  assign n21227 = ( n20559 & ~n21225 ) | ( n20559 & n21224 ) | ( ~n21225 & n21224 ) ;
  assign n21228 = ( n20546 & ~n21226 ) | ( n20546 & n21227 ) | ( ~n21226 & n21227 ) ;
  assign n21229 = n16671 | n21201 ;
  assign n21230 = ( n21215 & ~n21229 ) | ( n21215 & 1'b0 ) | ( ~n21229 & 1'b0 ) ;
  assign n21231 = n21221 | n21230 ;
  assign n21232 = ( n21209 & ~n21212 ) | ( n21209 & 1'b0 ) | ( ~n21212 & 1'b0 ) ;
  assign n21233 = ( n21206 & ~n17279 ) | ( n21206 & n21232 ) | ( ~n17279 & n21232 ) ;
  assign n21234 = ( n16671 & ~n21233 ) | ( n16671 & 1'b0 ) | ( ~n21233 & 1'b0 ) ;
  assign n21235 = n16070 | n21234 ;
  assign n21236 = ( n21231 & ~n21235 ) | ( n21231 & 1'b0 ) | ( ~n21235 & 1'b0 ) ;
  assign n21237 = n21228 | n21236 ;
  assign n21238 = ~n21223 & n21237 ;
  assign n21240 = ( n20548 & ~n20553 ) | ( n20548 & n21143 ) | ( ~n20553 & n21143 ) ;
  assign n21239 = n20561 &  n21143 ;
  assign n21241 = ( n21143 & ~n21240 ) | ( n21143 & n21239 ) | ( ~n21240 & n21239 ) ;
  assign n21242 = ( n21239 & ~n20548 ) | ( n21239 & n21240 ) | ( ~n20548 & n21240 ) ;
  assign n21243 = ( n20553 & ~n21241 ) | ( n20553 & n21242 ) | ( ~n21241 & n21242 ) ;
  assign n21244 = ( n21238 & ~n15484 ) | ( n21238 & n21243 ) | ( ~n15484 & n21243 ) ;
  assign n21245 = ( n14905 & ~n21244 ) | ( n14905 & 1'b0 ) | ( ~n21244 & 1'b0 ) ;
  assign n21246 = n20581 | n21143 ;
  assign n21247 = ( n20568 & ~n20581 ) | ( n20568 & n20577 ) | ( ~n20581 & n20577 ) ;
  assign n21249 = ( n20581 & n21246 ) | ( n20581 & n21247 ) | ( n21246 & n21247 ) ;
  assign n21248 = ( n20577 & ~n21247 ) | ( n20577 & n21246 ) | ( ~n21247 & n21246 ) ;
  assign n21250 = ( n20568 & ~n21249 ) | ( n20568 & n21248 ) | ( ~n21249 & n21248 ) ;
  assign n21251 = n15484 | n21223 ;
  assign n21252 = ( n21237 & ~n21251 ) | ( n21237 & 1'b0 ) | ( ~n21251 & 1'b0 ) ;
  assign n21253 = n21243 | n21252 ;
  assign n21254 = ( n21231 & ~n21234 ) | ( n21231 & 1'b0 ) | ( ~n21234 & 1'b0 ) ;
  assign n21255 = ( n21228 & ~n16070 ) | ( n21228 & n21254 ) | ( ~n16070 & n21254 ) ;
  assign n21256 = ( n15484 & ~n21255 ) | ( n15484 & 1'b0 ) | ( ~n21255 & 1'b0 ) ;
  assign n21257 = n14905 | n21256 ;
  assign n21258 = ( n21253 & ~n21257 ) | ( n21253 & 1'b0 ) | ( ~n21257 & 1'b0 ) ;
  assign n21259 = n21250 | n21258 ;
  assign n21260 = ~n21245 & n21259 ;
  assign n21262 = ( n20570 & ~n20575 ) | ( n20570 & n21143 ) | ( ~n20575 & n21143 ) ;
  assign n21261 = n20583 &  n21143 ;
  assign n21263 = ( n21143 & ~n21262 ) | ( n21143 & n21261 ) | ( ~n21262 & n21261 ) ;
  assign n21264 = ( n21261 & ~n20570 ) | ( n21261 & n21262 ) | ( ~n20570 & n21262 ) ;
  assign n21265 = ( n20575 & ~n21263 ) | ( n20575 & n21264 ) | ( ~n21263 & n21264 ) ;
  assign n21266 = ( n21260 & ~n14341 ) | ( n21260 & n21265 ) | ( ~n14341 & n21265 ) ;
  assign n21267 = ( n13784 & ~n21266 ) | ( n13784 & 1'b0 ) | ( ~n21266 & 1'b0 ) ;
  assign n21268 = n20603 | n21143 ;
  assign n21269 = ( n20590 & ~n20603 ) | ( n20590 & n20599 ) | ( ~n20603 & n20599 ) ;
  assign n21271 = ( n20603 & n21268 ) | ( n20603 & n21269 ) | ( n21268 & n21269 ) ;
  assign n21270 = ( n20599 & ~n21269 ) | ( n20599 & n21268 ) | ( ~n21269 & n21268 ) ;
  assign n21272 = ( n20590 & ~n21271 ) | ( n20590 & n21270 ) | ( ~n21271 & n21270 ) ;
  assign n21273 = n14341 | n21245 ;
  assign n21274 = ( n21259 & ~n21273 ) | ( n21259 & 1'b0 ) | ( ~n21273 & 1'b0 ) ;
  assign n21275 = n21265 | n21274 ;
  assign n21276 = ( n21253 & ~n21256 ) | ( n21253 & 1'b0 ) | ( ~n21256 & 1'b0 ) ;
  assign n21277 = ( n21250 & ~n14905 ) | ( n21250 & n21276 ) | ( ~n14905 & n21276 ) ;
  assign n21278 = ( n14341 & ~n21277 ) | ( n14341 & 1'b0 ) | ( ~n21277 & 1'b0 ) ;
  assign n21279 = n13784 | n21278 ;
  assign n21280 = ( n21275 & ~n21279 ) | ( n21275 & 1'b0 ) | ( ~n21279 & 1'b0 ) ;
  assign n21281 = n21272 | n21280 ;
  assign n21282 = ~n21267 & n21281 ;
  assign n21283 = n20605 &  n21143 ;
  assign n21284 = ( n20592 & n20597 ) | ( n20592 & n21143 ) | ( n20597 & n21143 ) ;
  assign n21286 = ( n21283 & ~n20592 ) | ( n21283 & n21284 ) | ( ~n20592 & n21284 ) ;
  assign n21285 = ( n21143 & ~n21284 ) | ( n21143 & n21283 ) | ( ~n21284 & n21283 ) ;
  assign n21287 = ( n20597 & ~n21286 ) | ( n20597 & n21285 ) | ( ~n21286 & n21285 ) ;
  assign n21288 = ( n21282 & ~n13242 ) | ( n21282 & n21287 ) | ( ~n13242 & n21287 ) ;
  assign n21289 = ( n12707 & ~n21288 ) | ( n12707 & 1'b0 ) | ( ~n21288 & 1'b0 ) ;
  assign n21290 = n20625 | n21143 ;
  assign n21291 = ( n20612 & ~n20625 ) | ( n20612 & n20621 ) | ( ~n20625 & n20621 ) ;
  assign n21293 = ( n20625 & n21290 ) | ( n20625 & n21291 ) | ( n21290 & n21291 ) ;
  assign n21292 = ( n20621 & ~n21291 ) | ( n20621 & n21290 ) | ( ~n21291 & n21290 ) ;
  assign n21294 = ( n20612 & ~n21293 ) | ( n20612 & n21292 ) | ( ~n21293 & n21292 ) ;
  assign n21295 = n13242 | n21267 ;
  assign n21296 = ( n21281 & ~n21295 ) | ( n21281 & 1'b0 ) | ( ~n21295 & 1'b0 ) ;
  assign n21297 = n21287 | n21296 ;
  assign n21298 = ( n21275 & ~n21278 ) | ( n21275 & 1'b0 ) | ( ~n21278 & 1'b0 ) ;
  assign n21299 = ( n21272 & ~n13784 ) | ( n21272 & n21298 ) | ( ~n13784 & n21298 ) ;
  assign n21300 = ( n13242 & ~n21299 ) | ( n13242 & 1'b0 ) | ( ~n21299 & 1'b0 ) ;
  assign n21301 = n12707 | n21300 ;
  assign n21302 = ( n21297 & ~n21301 ) | ( n21297 & 1'b0 ) | ( ~n21301 & 1'b0 ) ;
  assign n21303 = n21294 | n21302 ;
  assign n21304 = ~n21289 & n21303 ;
  assign n21305 = n20627 &  n21143 ;
  assign n21306 = ( n20614 & n20619 ) | ( n20614 & n21143 ) | ( n20619 & n21143 ) ;
  assign n21308 = ( n21305 & ~n20614 ) | ( n21305 & n21306 ) | ( ~n20614 & n21306 ) ;
  assign n21307 = ( n21143 & ~n21306 ) | ( n21143 & n21305 ) | ( ~n21306 & n21305 ) ;
  assign n21309 = ( n20619 & ~n21308 ) | ( n20619 & n21307 ) | ( ~n21308 & n21307 ) ;
  assign n21310 = ( n21304 & ~n12187 ) | ( n21304 & n21309 ) | ( ~n12187 & n21309 ) ;
  assign n21311 = ( n11674 & ~n21310 ) | ( n11674 & 1'b0 ) | ( ~n21310 & 1'b0 ) ;
  assign n21312 = n20647 | n21143 ;
  assign n21313 = ( n20634 & ~n20647 ) | ( n20634 & n20643 ) | ( ~n20647 & n20643 ) ;
  assign n21315 = ( n20647 & n21312 ) | ( n20647 & n21313 ) | ( n21312 & n21313 ) ;
  assign n21314 = ( n20643 & ~n21313 ) | ( n20643 & n21312 ) | ( ~n21313 & n21312 ) ;
  assign n21316 = ( n20634 & ~n21315 ) | ( n20634 & n21314 ) | ( ~n21315 & n21314 ) ;
  assign n21317 = n12187 | n21289 ;
  assign n21318 = ( n21303 & ~n21317 ) | ( n21303 & 1'b0 ) | ( ~n21317 & 1'b0 ) ;
  assign n21319 = n21309 | n21318 ;
  assign n21320 = ( n21297 & ~n21300 ) | ( n21297 & 1'b0 ) | ( ~n21300 & 1'b0 ) ;
  assign n21321 = ( n21294 & ~n12707 ) | ( n21294 & n21320 ) | ( ~n12707 & n21320 ) ;
  assign n21322 = ( n12187 & ~n21321 ) | ( n12187 & 1'b0 ) | ( ~n21321 & 1'b0 ) ;
  assign n21323 = n11674 | n21322 ;
  assign n21324 = ( n21319 & ~n21323 ) | ( n21319 & 1'b0 ) | ( ~n21323 & 1'b0 ) ;
  assign n21325 = n21316 | n21324 ;
  assign n21326 = ~n21311 & n21325 ;
  assign n21328 = ( n20636 & ~n20641 ) | ( n20636 & n21143 ) | ( ~n20641 & n21143 ) ;
  assign n21327 = n20649 &  n21143 ;
  assign n21329 = ( n21143 & ~n21328 ) | ( n21143 & n21327 ) | ( ~n21328 & n21327 ) ;
  assign n21330 = ( n21327 & ~n20636 ) | ( n21327 & n21328 ) | ( ~n20636 & n21328 ) ;
  assign n21331 = ( n20641 & ~n21329 ) | ( n20641 & n21330 ) | ( ~n21329 & n21330 ) ;
  assign n21332 = ( n21326 & ~n11176 ) | ( n21326 & n21331 ) | ( ~n11176 & n21331 ) ;
  assign n21333 = ( n10685 & ~n21332 ) | ( n10685 & 1'b0 ) | ( ~n21332 & 1'b0 ) ;
  assign n21334 = n20669 | n21143 ;
  assign n21335 = ( n20656 & ~n20669 ) | ( n20656 & n20665 ) | ( ~n20669 & n20665 ) ;
  assign n21337 = ( n20669 & n21334 ) | ( n20669 & n21335 ) | ( n21334 & n21335 ) ;
  assign n21336 = ( n20665 & ~n21335 ) | ( n20665 & n21334 ) | ( ~n21335 & n21334 ) ;
  assign n21338 = ( n20656 & ~n21337 ) | ( n20656 & n21336 ) | ( ~n21337 & n21336 ) ;
  assign n21339 = n11176 | n21311 ;
  assign n21340 = ( n21325 & ~n21339 ) | ( n21325 & 1'b0 ) | ( ~n21339 & 1'b0 ) ;
  assign n21341 = n21331 | n21340 ;
  assign n21342 = ( n21319 & ~n21322 ) | ( n21319 & 1'b0 ) | ( ~n21322 & 1'b0 ) ;
  assign n21343 = ( n21316 & ~n11674 ) | ( n21316 & n21342 ) | ( ~n11674 & n21342 ) ;
  assign n21344 = ( n11176 & ~n21343 ) | ( n11176 & 1'b0 ) | ( ~n21343 & 1'b0 ) ;
  assign n21345 = n10685 | n21344 ;
  assign n21346 = ( n21341 & ~n21345 ) | ( n21341 & 1'b0 ) | ( ~n21345 & 1'b0 ) ;
  assign n21347 = n21338 | n21346 ;
  assign n21348 = ~n21333 & n21347 ;
  assign n21349 = n20671 &  n21143 ;
  assign n21350 = ( n20658 & n20663 ) | ( n20658 & n21143 ) | ( n20663 & n21143 ) ;
  assign n21352 = ( n21349 & ~n20658 ) | ( n21349 & n21350 ) | ( ~n20658 & n21350 ) ;
  assign n21351 = ( n21143 & ~n21350 ) | ( n21143 & n21349 ) | ( ~n21350 & n21349 ) ;
  assign n21353 = ( n20663 & ~n21352 ) | ( n20663 & n21351 ) | ( ~n21352 & n21351 ) ;
  assign n21354 = ( n21348 & ~n10209 ) | ( n21348 & n21353 ) | ( ~n10209 & n21353 ) ;
  assign n21355 = n9740 | n21354 ;
  assign n21356 = n20691 | n21143 ;
  assign n21357 = ( n20678 & ~n20687 ) | ( n20678 & n20691 ) | ( ~n20687 & n20691 ) ;
  assign n21358 = ( n20687 & n21356 ) | ( n20687 & n21357 ) | ( n21356 & n21357 ) ;
  assign n21359 = ( n20691 & ~n21357 ) | ( n20691 & n21356 ) | ( ~n21357 & n21356 ) ;
  assign n21360 = ( n20678 & ~n21358 ) | ( n20678 & n21359 ) | ( ~n21358 & n21359 ) ;
  assign n21361 = n10209 | n21333 ;
  assign n21362 = ( n21347 & ~n21361 ) | ( n21347 & 1'b0 ) | ( ~n21361 & 1'b0 ) ;
  assign n21363 = n21353 | n21362 ;
  assign n21364 = ( n21341 & ~n21344 ) | ( n21341 & 1'b0 ) | ( ~n21344 & 1'b0 ) ;
  assign n21365 = ( n21338 & ~n10685 ) | ( n21338 & n21364 ) | ( ~n10685 & n21364 ) ;
  assign n21366 = ( n10209 & ~n21365 ) | ( n10209 & 1'b0 ) | ( ~n21365 & 1'b0 ) ;
  assign n21367 = ( n9740 & ~n21366 ) | ( n9740 & 1'b0 ) | ( ~n21366 & 1'b0 ) ;
  assign n21368 = n21363 &  n21367 ;
  assign n21369 = n21360 | n21368 ;
  assign n21370 = n21355 &  n21369 ;
  assign n21371 = ( n20680 & ~n21143 ) | ( n20680 & 1'b0 ) | ( ~n21143 & 1'b0 ) ;
  assign n21372 = ( n20680 & n20685 ) | ( n20680 & n20693 ) | ( n20685 & n20693 ) ;
  assign n21373 = ( n21371 & ~n20693 ) | ( n21371 & n21372 ) | ( ~n20693 & n21372 ) ;
  assign n21374 = ( n20680 & ~n21372 ) | ( n20680 & n21371 ) | ( ~n21372 & n21371 ) ;
  assign n21375 = ( n20685 & ~n21373 ) | ( n20685 & n21374 ) | ( ~n21373 & n21374 ) ;
  assign n21376 = ( n21370 & ~n9286 ) | ( n21370 & n21375 ) | ( ~n9286 & n21375 ) ;
  assign n21377 = ( n8839 & ~n21376 ) | ( n8839 & 1'b0 ) | ( ~n21376 & 1'b0 ) ;
  assign n21378 = n20713 | n21143 ;
  assign n21379 = ( n20700 & ~n20709 ) | ( n20700 & n20713 ) | ( ~n20709 & n20713 ) ;
  assign n21380 = ( n20709 & n21378 ) | ( n20709 & n21379 ) | ( n21378 & n21379 ) ;
  assign n21381 = ( n20713 & ~n21379 ) | ( n20713 & n21378 ) | ( ~n21379 & n21378 ) ;
  assign n21382 = ( n20700 & ~n21380 ) | ( n20700 & n21381 ) | ( ~n21380 & n21381 ) ;
  assign n21383 = ~n9286 & n21355 ;
  assign n21384 = n21369 &  n21383 ;
  assign n21385 = n21375 | n21384 ;
  assign n21386 = ( n21363 & ~n21366 ) | ( n21363 & 1'b0 ) | ( ~n21366 & 1'b0 ) ;
  assign n21387 = ( n9740 & n21360 ) | ( n9740 & n21386 ) | ( n21360 & n21386 ) ;
  assign n21388 = ( n9286 & ~n21387 ) | ( n9286 & 1'b0 ) | ( ~n21387 & 1'b0 ) ;
  assign n21389 = n8839 | n21388 ;
  assign n21390 = ( n21385 & ~n21389 ) | ( n21385 & 1'b0 ) | ( ~n21389 & 1'b0 ) ;
  assign n21391 = n21382 | n21390 ;
  assign n21392 = ~n21377 & n21391 ;
  assign n21393 = n20702 | n21143 ;
  assign n21394 = ( n20702 & ~n20715 ) | ( n20702 & n20707 ) | ( ~n20715 & n20707 ) ;
  assign n21395 = ( n20715 & n21393 ) | ( n20715 & n21394 ) | ( n21393 & n21394 ) ;
  assign n21396 = ( n20702 & ~n21394 ) | ( n20702 & n21393 ) | ( ~n21394 & n21393 ) ;
  assign n21397 = ( n20707 & ~n21395 ) | ( n20707 & n21396 ) | ( ~n21395 & n21396 ) ;
  assign n21398 = ( n21392 & ~n8407 ) | ( n21392 & n21397 ) | ( ~n8407 & n21397 ) ;
  assign n21399 = ( n7982 & ~n21398 ) | ( n7982 & 1'b0 ) | ( ~n21398 & 1'b0 ) ;
  assign n21400 = n20735 | n21143 ;
  assign n21401 = ( n20722 & ~n20735 ) | ( n20722 & n20731 ) | ( ~n20735 & n20731 ) ;
  assign n21403 = ( n20735 & n21400 ) | ( n20735 & n21401 ) | ( n21400 & n21401 ) ;
  assign n21402 = ( n20731 & ~n21401 ) | ( n20731 & n21400 ) | ( ~n21401 & n21400 ) ;
  assign n21404 = ( n20722 & ~n21403 ) | ( n20722 & n21402 ) | ( ~n21403 & n21402 ) ;
  assign n21405 = n8407 | n21377 ;
  assign n21406 = ( n21391 & ~n21405 ) | ( n21391 & 1'b0 ) | ( ~n21405 & 1'b0 ) ;
  assign n21407 = n21397 | n21406 ;
  assign n21408 = ( n21385 & ~n21388 ) | ( n21385 & 1'b0 ) | ( ~n21388 & 1'b0 ) ;
  assign n21409 = ( n21382 & ~n8839 ) | ( n21382 & n21408 ) | ( ~n8839 & n21408 ) ;
  assign n21410 = ( n8407 & ~n21409 ) | ( n8407 & 1'b0 ) | ( ~n21409 & 1'b0 ) ;
  assign n21411 = n7982 | n21410 ;
  assign n21412 = ( n21407 & ~n21411 ) | ( n21407 & 1'b0 ) | ( ~n21411 & 1'b0 ) ;
  assign n21413 = n21404 | n21412 ;
  assign n21414 = ~n21399 & n21413 ;
  assign n21415 = n20724 | n21143 ;
  assign n21416 = ( n20729 & ~n20724 ) | ( n20729 & n20737 ) | ( ~n20724 & n20737 ) ;
  assign n21418 = ( n20724 & n21415 ) | ( n20724 & n21416 ) | ( n21415 & n21416 ) ;
  assign n21417 = ( n20737 & ~n21416 ) | ( n20737 & n21415 ) | ( ~n21416 & n21415 ) ;
  assign n21419 = ( n20729 & ~n21418 ) | ( n20729 & n21417 ) | ( ~n21418 & n21417 ) ;
  assign n21420 = ( n7572 & n21414 ) | ( n7572 & n21419 ) | ( n21414 & n21419 ) ;
  assign n21421 = n7169 | n21420 ;
  assign n21423 = ( n20753 & ~n20744 ) | ( n20753 & n20757 ) | ( ~n20744 & n20757 ) ;
  assign n21422 = ( n20757 & ~n21143 ) | ( n20757 & 1'b0 ) | ( ~n21143 & 1'b0 ) ;
  assign n21425 = ( n20757 & ~n21423 ) | ( n20757 & n21422 ) | ( ~n21423 & n21422 ) ;
  assign n21424 = ( n21422 & ~n20753 ) | ( n21422 & n21423 ) | ( ~n20753 & n21423 ) ;
  assign n21426 = ( n20744 & ~n21425 ) | ( n20744 & n21424 ) | ( ~n21425 & n21424 ) ;
  assign n21427 = ( n7572 & ~n21399 ) | ( n7572 & 1'b0 ) | ( ~n21399 & 1'b0 ) ;
  assign n21428 = n21413 &  n21427 ;
  assign n21429 = n21419 | n21428 ;
  assign n21430 = ( n21407 & ~n21410 ) | ( n21407 & 1'b0 ) | ( ~n21410 & 1'b0 ) ;
  assign n21431 = ( n21404 & ~n7982 ) | ( n21404 & n21430 ) | ( ~n7982 & n21430 ) ;
  assign n21432 = n7572 | n21431 ;
  assign n21433 = n7169 &  n21432 ;
  assign n21434 = n21429 &  n21433 ;
  assign n21435 = n21426 | n21434 ;
  assign n21436 = n21421 &  n21435 ;
  assign n21437 = ( n20746 & ~n21143 ) | ( n20746 & 1'b0 ) | ( ~n21143 & 1'b0 ) ;
  assign n21438 = ( n20746 & n20751 ) | ( n20746 & n20759 ) | ( n20751 & n20759 ) ;
  assign n21439 = ( n21437 & ~n20759 ) | ( n21437 & n21438 ) | ( ~n20759 & n21438 ) ;
  assign n21440 = ( n20746 & ~n21438 ) | ( n20746 & n21437 ) | ( ~n21438 & n21437 ) ;
  assign n21441 = ( n20751 & ~n21439 ) | ( n20751 & n21440 ) | ( ~n21439 & n21440 ) ;
  assign n21442 = ( n21436 & ~n6781 ) | ( n21436 & n21441 ) | ( ~n6781 & n21441 ) ;
  assign n21443 = n6399 | n21442 ;
  assign n21444 = n20779 | n21143 ;
  assign n21445 = ( n20766 & ~n20775 ) | ( n20766 & n20779 ) | ( ~n20775 & n20779 ) ;
  assign n21446 = ( n20775 & n21444 ) | ( n20775 & n21445 ) | ( n21444 & n21445 ) ;
  assign n21447 = ( n20779 & ~n21445 ) | ( n20779 & n21444 ) | ( ~n21445 & n21444 ) ;
  assign n21448 = ( n20766 & ~n21446 ) | ( n20766 & n21447 ) | ( ~n21446 & n21447 ) ;
  assign n21449 = ~n6781 & n21421 ;
  assign n21450 = n21435 &  n21449 ;
  assign n21451 = n21441 | n21450 ;
  assign n21452 = n21429 &  n21432 ;
  assign n21453 = ( n7169 & n21426 ) | ( n7169 & n21452 ) | ( n21426 & n21452 ) ;
  assign n21454 = ( n6781 & ~n21453 ) | ( n6781 & 1'b0 ) | ( ~n21453 & 1'b0 ) ;
  assign n21455 = ( n6399 & ~n21454 ) | ( n6399 & 1'b0 ) | ( ~n21454 & 1'b0 ) ;
  assign n21456 = n21451 &  n21455 ;
  assign n21457 = n21448 | n21456 ;
  assign n21458 = n21443 &  n21457 ;
  assign n21459 = ( n20768 & ~n21143 ) | ( n20768 & 1'b0 ) | ( ~n21143 & 1'b0 ) ;
  assign n21460 = ( n20768 & n20773 ) | ( n20768 & n20781 ) | ( n20773 & n20781 ) ;
  assign n21461 = ( n21459 & ~n20781 ) | ( n21459 & n21460 ) | ( ~n20781 & n21460 ) ;
  assign n21462 = ( n20768 & ~n21460 ) | ( n20768 & n21459 ) | ( ~n21460 & n21459 ) ;
  assign n21463 = ( n20773 & ~n21461 ) | ( n20773 & n21462 ) | ( ~n21461 & n21462 ) ;
  assign n21464 = ( n21458 & ~n6032 ) | ( n21458 & n21463 ) | ( ~n6032 & n21463 ) ;
  assign n21465 = n5672 | n21464 ;
  assign n21466 = n20801 | n21143 ;
  assign n21467 = ( n20788 & ~n20797 ) | ( n20788 & n20801 ) | ( ~n20797 & n20801 ) ;
  assign n21468 = ( n20797 & n21466 ) | ( n20797 & n21467 ) | ( n21466 & n21467 ) ;
  assign n21469 = ( n20801 & ~n21467 ) | ( n20801 & n21466 ) | ( ~n21467 & n21466 ) ;
  assign n21470 = ( n20788 & ~n21468 ) | ( n20788 & n21469 ) | ( ~n21468 & n21469 ) ;
  assign n21471 = ~n6032 & n21443 ;
  assign n21472 = n21457 &  n21471 ;
  assign n21473 = n21463 | n21472 ;
  assign n21474 = ( n21451 & ~n21454 ) | ( n21451 & 1'b0 ) | ( ~n21454 & 1'b0 ) ;
  assign n21475 = ( n6399 & n21448 ) | ( n6399 & n21474 ) | ( n21448 & n21474 ) ;
  assign n21476 = ( n6032 & ~n21475 ) | ( n6032 & 1'b0 ) | ( ~n21475 & 1'b0 ) ;
  assign n21477 = ( n5672 & ~n21476 ) | ( n5672 & 1'b0 ) | ( ~n21476 & 1'b0 ) ;
  assign n21478 = n21473 &  n21477 ;
  assign n21479 = n21470 | n21478 ;
  assign n21480 = n21465 &  n21479 ;
  assign n21481 = ( n20790 & ~n21143 ) | ( n20790 & 1'b0 ) | ( ~n21143 & 1'b0 ) ;
  assign n21482 = ( n20790 & n20795 ) | ( n20790 & n20803 ) | ( n20795 & n20803 ) ;
  assign n21483 = ( n21481 & ~n20803 ) | ( n21481 & n21482 ) | ( ~n20803 & n21482 ) ;
  assign n21484 = ( n20790 & ~n21482 ) | ( n20790 & n21481 ) | ( ~n21482 & n21481 ) ;
  assign n21485 = ( n20795 & ~n21483 ) | ( n20795 & n21484 ) | ( ~n21483 & n21484 ) ;
  assign n21486 = ( n21480 & ~n5327 ) | ( n21480 & n21485 ) | ( ~n5327 & n21485 ) ;
  assign n21487 = ( n4990 & ~n21486 ) | ( n4990 & 1'b0 ) | ( ~n21486 & 1'b0 ) ;
  assign n21488 = n20823 | n21143 ;
  assign n21489 = ( n20810 & ~n20819 ) | ( n20810 & n20823 ) | ( ~n20819 & n20823 ) ;
  assign n21490 = ( n20819 & n21488 ) | ( n20819 & n21489 ) | ( n21488 & n21489 ) ;
  assign n21491 = ( n20823 & ~n21489 ) | ( n20823 & n21488 ) | ( ~n21489 & n21488 ) ;
  assign n21492 = ( n20810 & ~n21490 ) | ( n20810 & n21491 ) | ( ~n21490 & n21491 ) ;
  assign n21493 = ~n5327 & n21465 ;
  assign n21494 = n21479 &  n21493 ;
  assign n21495 = n21485 | n21494 ;
  assign n21496 = ( n21473 & ~n21476 ) | ( n21473 & 1'b0 ) | ( ~n21476 & 1'b0 ) ;
  assign n21497 = ( n5672 & n21470 ) | ( n5672 & n21496 ) | ( n21470 & n21496 ) ;
  assign n21498 = ( n5327 & ~n21497 ) | ( n5327 & 1'b0 ) | ( ~n21497 & 1'b0 ) ;
  assign n21499 = n4990 | n21498 ;
  assign n21500 = ( n21495 & ~n21499 ) | ( n21495 & 1'b0 ) | ( ~n21499 & 1'b0 ) ;
  assign n21501 = n21492 | n21500 ;
  assign n21502 = ~n21487 & n21501 ;
  assign n21503 = n20812 | n21143 ;
  assign n21504 = ( n20817 & ~n20812 ) | ( n20817 & n20825 ) | ( ~n20812 & n20825 ) ;
  assign n21506 = ( n20812 & n21503 ) | ( n20812 & n21504 ) | ( n21503 & n21504 ) ;
  assign n21505 = ( n20825 & ~n21504 ) | ( n20825 & n21503 ) | ( ~n21504 & n21503 ) ;
  assign n21507 = ( n20817 & ~n21506 ) | ( n20817 & n21505 ) | ( ~n21506 & n21505 ) ;
  assign n21508 = ( n21502 & ~n4668 ) | ( n21502 & n21507 ) | ( ~n4668 & n21507 ) ;
  assign n21509 = ( n4353 & ~n21508 ) | ( n4353 & 1'b0 ) | ( ~n21508 & 1'b0 ) ;
  assign n21510 = n20845 | n21143 ;
  assign n21511 = ( n20832 & ~n20841 ) | ( n20832 & n20845 ) | ( ~n20841 & n20845 ) ;
  assign n21512 = ( n20841 & n21510 ) | ( n20841 & n21511 ) | ( n21510 & n21511 ) ;
  assign n21513 = ( n20845 & ~n21511 ) | ( n20845 & n21510 ) | ( ~n21511 & n21510 ) ;
  assign n21514 = ( n20832 & ~n21512 ) | ( n20832 & n21513 ) | ( ~n21512 & n21513 ) ;
  assign n21515 = n4668 | n21487 ;
  assign n21516 = ( n21501 & ~n21515 ) | ( n21501 & 1'b0 ) | ( ~n21515 & 1'b0 ) ;
  assign n21517 = n21507 | n21516 ;
  assign n21518 = ( n21495 & ~n21498 ) | ( n21495 & 1'b0 ) | ( ~n21498 & 1'b0 ) ;
  assign n21519 = ( n21492 & ~n4990 ) | ( n21492 & n21518 ) | ( ~n4990 & n21518 ) ;
  assign n21520 = ( n4668 & ~n21519 ) | ( n4668 & 1'b0 ) | ( ~n21519 & 1'b0 ) ;
  assign n21521 = n4353 | n21520 ;
  assign n21522 = ( n21517 & ~n21521 ) | ( n21517 & 1'b0 ) | ( ~n21521 & 1'b0 ) ;
  assign n21523 = n21514 | n21522 ;
  assign n21524 = ~n21509 & n21523 ;
  assign n21525 = n20834 | n21143 ;
  assign n21526 = ( n20839 & ~n20834 ) | ( n20839 & n20847 ) | ( ~n20834 & n20847 ) ;
  assign n21528 = ( n20834 & n21525 ) | ( n20834 & n21526 ) | ( n21525 & n21526 ) ;
  assign n21527 = ( n20847 & ~n21526 ) | ( n20847 & n21525 ) | ( ~n21526 & n21525 ) ;
  assign n21529 = ( n20839 & ~n21528 ) | ( n20839 & n21527 ) | ( ~n21528 & n21527 ) ;
  assign n21530 = ( n21524 & ~n4053 ) | ( n21524 & n21529 ) | ( ~n4053 & n21529 ) ;
  assign n21531 = ( n3760 & ~n21530 ) | ( n3760 & 1'b0 ) | ( ~n21530 & 1'b0 ) ;
  assign n21532 = n20867 | n21143 ;
  assign n21533 = ( n20854 & ~n20863 ) | ( n20854 & n20867 ) | ( ~n20863 & n20867 ) ;
  assign n21534 = ( n20863 & n21532 ) | ( n20863 & n21533 ) | ( n21532 & n21533 ) ;
  assign n21535 = ( n20867 & ~n21533 ) | ( n20867 & n21532 ) | ( ~n21533 & n21532 ) ;
  assign n21536 = ( n20854 & ~n21534 ) | ( n20854 & n21535 ) | ( ~n21534 & n21535 ) ;
  assign n21537 = n4053 | n21509 ;
  assign n21538 = ( n21523 & ~n21537 ) | ( n21523 & 1'b0 ) | ( ~n21537 & 1'b0 ) ;
  assign n21539 = n21529 | n21538 ;
  assign n21540 = ( n21517 & ~n21520 ) | ( n21517 & 1'b0 ) | ( ~n21520 & 1'b0 ) ;
  assign n21541 = ( n21514 & ~n4353 ) | ( n21514 & n21540 ) | ( ~n4353 & n21540 ) ;
  assign n21542 = ( n4053 & ~n21541 ) | ( n4053 & 1'b0 ) | ( ~n21541 & 1'b0 ) ;
  assign n21543 = n3760 | n21542 ;
  assign n21544 = ( n21539 & ~n21543 ) | ( n21539 & 1'b0 ) | ( ~n21543 & 1'b0 ) ;
  assign n21545 = n21536 | n21544 ;
  assign n21546 = ~n21531 & n21545 ;
  assign n21547 = n20856 | n21143 ;
  assign n21548 = ( n20861 & ~n20856 ) | ( n20861 & n20869 ) | ( ~n20856 & n20869 ) ;
  assign n21550 = ( n20856 & n21547 ) | ( n20856 & n21548 ) | ( n21547 & n21548 ) ;
  assign n21549 = ( n20869 & ~n21548 ) | ( n20869 & n21547 ) | ( ~n21548 & n21547 ) ;
  assign n21551 = ( n20861 & ~n21550 ) | ( n20861 & n21549 ) | ( ~n21550 & n21549 ) ;
  assign n21552 = ( n21546 & ~n3482 ) | ( n21546 & n21551 ) | ( ~n3482 & n21551 ) ;
  assign n21553 = ( n3211 & ~n21552 ) | ( n3211 & 1'b0 ) | ( ~n21552 & 1'b0 ) ;
  assign n21554 = n20889 | n21143 ;
  assign n21555 = ( n20876 & ~n20885 ) | ( n20876 & n20889 ) | ( ~n20885 & n20889 ) ;
  assign n21556 = ( n20885 & n21554 ) | ( n20885 & n21555 ) | ( n21554 & n21555 ) ;
  assign n21557 = ( n20889 & ~n21555 ) | ( n20889 & n21554 ) | ( ~n21555 & n21554 ) ;
  assign n21558 = ( n20876 & ~n21556 ) | ( n20876 & n21557 ) | ( ~n21556 & n21557 ) ;
  assign n21559 = n3482 | n21531 ;
  assign n21560 = ( n21545 & ~n21559 ) | ( n21545 & 1'b0 ) | ( ~n21559 & 1'b0 ) ;
  assign n21561 = n21551 | n21560 ;
  assign n21562 = ( n21539 & ~n21542 ) | ( n21539 & 1'b0 ) | ( ~n21542 & 1'b0 ) ;
  assign n21563 = ( n21536 & ~n3760 ) | ( n21536 & n21562 ) | ( ~n3760 & n21562 ) ;
  assign n21564 = ( n3482 & ~n21563 ) | ( n3482 & 1'b0 ) | ( ~n21563 & 1'b0 ) ;
  assign n21565 = n3211 | n21564 ;
  assign n21566 = ( n21561 & ~n21565 ) | ( n21561 & 1'b0 ) | ( ~n21565 & 1'b0 ) ;
  assign n21567 = n21558 | n21566 ;
  assign n21568 = ~n21553 & n21567 ;
  assign n21569 = n20878 | n21143 ;
  assign n21570 = ( n20883 & ~n20878 ) | ( n20883 & n20891 ) | ( ~n20878 & n20891 ) ;
  assign n21572 = ( n20878 & n21569 ) | ( n20878 & n21570 ) | ( n21569 & n21570 ) ;
  assign n21571 = ( n20891 & ~n21570 ) | ( n20891 & n21569 ) | ( ~n21570 & n21569 ) ;
  assign n21573 = ( n20883 & ~n21572 ) | ( n20883 & n21571 ) | ( ~n21572 & n21571 ) ;
  assign n21574 = ( n21568 & ~n2955 ) | ( n21568 & n21573 ) | ( ~n2955 & n21573 ) ;
  assign n21575 = ( n2706 & ~n21574 ) | ( n2706 & 1'b0 ) | ( ~n21574 & 1'b0 ) ;
  assign n21576 = n20911 | n21143 ;
  assign n21577 = ( n20898 & ~n20907 ) | ( n20898 & n20911 ) | ( ~n20907 & n20911 ) ;
  assign n21578 = ( n20907 & n21576 ) | ( n20907 & n21577 ) | ( n21576 & n21577 ) ;
  assign n21579 = ( n20911 & ~n21577 ) | ( n20911 & n21576 ) | ( ~n21577 & n21576 ) ;
  assign n21580 = ( n20898 & ~n21578 ) | ( n20898 & n21579 ) | ( ~n21578 & n21579 ) ;
  assign n21581 = n2955 | n21553 ;
  assign n21582 = ( n21567 & ~n21581 ) | ( n21567 & 1'b0 ) | ( ~n21581 & 1'b0 ) ;
  assign n21583 = n21573 | n21582 ;
  assign n21584 = ( n21561 & ~n21564 ) | ( n21561 & 1'b0 ) | ( ~n21564 & 1'b0 ) ;
  assign n21585 = ( n21558 & ~n3211 ) | ( n21558 & n21584 ) | ( ~n3211 & n21584 ) ;
  assign n21586 = ( n2955 & ~n21585 ) | ( n2955 & 1'b0 ) | ( ~n21585 & 1'b0 ) ;
  assign n21587 = n2706 | n21586 ;
  assign n21588 = ( n21583 & ~n21587 ) | ( n21583 & 1'b0 ) | ( ~n21587 & 1'b0 ) ;
  assign n21589 = n21580 | n21588 ;
  assign n21590 = ~n21575 & n21589 ;
  assign n21591 = n20900 | n21143 ;
  assign n21592 = ( n20900 & ~n20913 ) | ( n20900 & n20905 ) | ( ~n20913 & n20905 ) ;
  assign n21593 = ( n20913 & n21591 ) | ( n20913 & n21592 ) | ( n21591 & n21592 ) ;
  assign n21594 = ( n20900 & ~n21592 ) | ( n20900 & n21591 ) | ( ~n21592 & n21591 ) ;
  assign n21595 = ( n20905 & ~n21593 ) | ( n20905 & n21594 ) | ( ~n21593 & n21594 ) ;
  assign n21596 = ( n2472 & ~n21590 ) | ( n2472 & n21595 ) | ( ~n21590 & n21595 ) ;
  assign n21597 = n2245 &  n21596 ;
  assign n21599 = ( n20929 & ~n20920 ) | ( n20929 & n20933 ) | ( ~n20920 & n20933 ) ;
  assign n21598 = n20933 | n21143 ;
  assign n21601 = ( n20933 & ~n21599 ) | ( n20933 & n21598 ) | ( ~n21599 & n21598 ) ;
  assign n21600 = ( n21598 & ~n20929 ) | ( n21598 & n21599 ) | ( ~n20929 & n21599 ) ;
  assign n21602 = ( n20920 & ~n21601 ) | ( n20920 & n21600 ) | ( ~n21601 & n21600 ) ;
  assign n21603 = n2472 | n21575 ;
  assign n21604 = ( n21589 & ~n21603 ) | ( n21589 & 1'b0 ) | ( ~n21603 & 1'b0 ) ;
  assign n21605 = ( n21595 & ~n21604 ) | ( n21595 & 1'b0 ) | ( ~n21604 & 1'b0 ) ;
  assign n21606 = ( n21583 & ~n21586 ) | ( n21583 & 1'b0 ) | ( ~n21586 & 1'b0 ) ;
  assign n21607 = ( n21580 & ~n2706 ) | ( n21580 & n21606 ) | ( ~n2706 & n21606 ) ;
  assign n21608 = ( n2472 & ~n21607 ) | ( n2472 & 1'b0 ) | ( ~n21607 & 1'b0 ) ;
  assign n21609 = n2245 | n21608 ;
  assign n21610 = n21605 | n21609 ;
  assign n21611 = n21602 &  n21610 ;
  assign n21612 = n21597 | n21611 ;
  assign n21613 = n20922 | n21143 ;
  assign n21614 = ( n20922 & n20927 ) | ( n20922 & n20935 ) | ( n20927 & n20935 ) ;
  assign n21615 = ( n21613 & ~n20935 ) | ( n21613 & n21614 ) | ( ~n20935 & n21614 ) ;
  assign n21616 = ( n20922 & ~n21614 ) | ( n20922 & n21613 ) | ( ~n21614 & n21613 ) ;
  assign n21617 = ( n20927 & ~n21615 ) | ( n20927 & n21616 ) | ( ~n21615 & n21616 ) ;
  assign n21618 = ( n21612 & ~n2033 ) | ( n21612 & n21617 ) | ( ~n2033 & n21617 ) ;
  assign n21619 = n1827 &  n21618 ;
  assign n21620 = n20955 | n21143 ;
  assign n21621 = ( n20942 & ~n20955 ) | ( n20942 & n20951 ) | ( ~n20955 & n20951 ) ;
  assign n21623 = ( n20955 & n21620 ) | ( n20955 & n21621 ) | ( n21620 & n21621 ) ;
  assign n21622 = ( n20951 & ~n21621 ) | ( n20951 & n21620 ) | ( ~n21621 & n21620 ) ;
  assign n21624 = ( n20942 & ~n21623 ) | ( n20942 & n21622 ) | ( ~n21623 & n21622 ) ;
  assign n21625 = ( n2033 & ~n21597 ) | ( n2033 & 1'b0 ) | ( ~n21597 & 1'b0 ) ;
  assign n21626 = ~n21611 & n21625 ;
  assign n21627 = ( n21617 & ~n21626 ) | ( n21617 & 1'b0 ) | ( ~n21626 & 1'b0 ) ;
  assign n21628 = n21605 | n21608 ;
  assign n21629 = ( n2245 & n21602 ) | ( n2245 & n21628 ) | ( n21602 & n21628 ) ;
  assign n21630 = ~n2033 & n21629 ;
  assign n21631 = n1827 | n21630 ;
  assign n21632 = n21627 | n21631 ;
  assign n21633 = n21624 &  n21632 ;
  assign n21634 = n21619 | n21633 ;
  assign n21635 = n20944 | n21143 ;
  assign n21636 = ( n20944 & n20949 ) | ( n20944 & n20957 ) | ( n20949 & n20957 ) ;
  assign n21637 = ( n21635 & ~n20957 ) | ( n21635 & n21636 ) | ( ~n20957 & n21636 ) ;
  assign n21638 = ( n20944 & ~n21636 ) | ( n20944 & n21635 ) | ( ~n21636 & n21635 ) ;
  assign n21639 = ( n20949 & ~n21637 ) | ( n20949 & n21638 ) | ( ~n21637 & n21638 ) ;
  assign n21640 = ( n21634 & ~n1636 ) | ( n21634 & n21639 ) | ( ~n1636 & n21639 ) ;
  assign n21641 = ~n1452 & n21640 ;
  assign n21642 = n20977 | n21143 ;
  assign n21643 = ( n20964 & ~n20973 ) | ( n20964 & n20977 ) | ( ~n20973 & n20977 ) ;
  assign n21644 = ( n20973 & n21642 ) | ( n20973 & n21643 ) | ( n21642 & n21643 ) ;
  assign n21645 = ( n20977 & ~n21643 ) | ( n20977 & n21642 ) | ( ~n21643 & n21642 ) ;
  assign n21646 = ( n20964 & ~n21644 ) | ( n20964 & n21645 ) | ( ~n21644 & n21645 ) ;
  assign n21647 = ( n1636 & ~n21619 ) | ( n1636 & 1'b0 ) | ( ~n21619 & 1'b0 ) ;
  assign n21648 = ~n21633 & n21647 ;
  assign n21649 = ( n21639 & ~n21648 ) | ( n21639 & 1'b0 ) | ( ~n21648 & 1'b0 ) ;
  assign n21650 = n21627 | n21630 ;
  assign n21651 = ( n1827 & n21624 ) | ( n1827 & n21650 ) | ( n21624 & n21650 ) ;
  assign n21652 = ~n1636 & n21651 ;
  assign n21653 = ( n1452 & ~n21652 ) | ( n1452 & 1'b0 ) | ( ~n21652 & 1'b0 ) ;
  assign n21654 = ~n21649 & n21653 ;
  assign n21655 = n21646 | n21654 ;
  assign n21656 = ~n21641 & n21655 ;
  assign n21657 = ( n20966 & ~n21143 ) | ( n20966 & 1'b0 ) | ( ~n21143 & 1'b0 ) ;
  assign n21658 = ( n20966 & n20971 ) | ( n20966 & n20979 ) | ( n20971 & n20979 ) ;
  assign n21659 = ( n21657 & ~n20979 ) | ( n21657 & n21658 ) | ( ~n20979 & n21658 ) ;
  assign n21660 = ( n20966 & ~n21658 ) | ( n20966 & n21657 ) | ( ~n21658 & n21657 ) ;
  assign n21661 = ( n20971 & ~n21659 ) | ( n20971 & n21660 ) | ( ~n21659 & n21660 ) ;
  assign n21662 = ( n21656 & ~n1283 ) | ( n21656 & n21661 ) | ( ~n1283 & n21661 ) ;
  assign n21663 = n1122 | n21662 ;
  assign n21664 = n20999 | n21143 ;
  assign n21665 = ( n20986 & ~n20999 ) | ( n20986 & n20995 ) | ( ~n20999 & n20995 ) ;
  assign n21667 = ( n20999 & n21664 ) | ( n20999 & n21665 ) | ( n21664 & n21665 ) ;
  assign n21666 = ( n20995 & ~n21665 ) | ( n20995 & n21664 ) | ( ~n21665 & n21664 ) ;
  assign n21668 = ( n20986 & ~n21667 ) | ( n20986 & n21666 ) | ( ~n21667 & n21666 ) ;
  assign n21669 = n1283 | n21641 ;
  assign n21670 = ( n21655 & ~n21669 ) | ( n21655 & 1'b0 ) | ( ~n21669 & 1'b0 ) ;
  assign n21671 = n21661 | n21670 ;
  assign n21672 = n21649 | n21652 ;
  assign n21673 = ( n1452 & ~n21672 ) | ( n1452 & n21646 ) | ( ~n21672 & n21646 ) ;
  assign n21674 = ( n1283 & ~n21673 ) | ( n1283 & 1'b0 ) | ( ~n21673 & 1'b0 ) ;
  assign n21675 = ( n1122 & ~n21674 ) | ( n1122 & 1'b0 ) | ( ~n21674 & 1'b0 ) ;
  assign n21676 = n21671 &  n21675 ;
  assign n21677 = ( n21668 & ~n21676 ) | ( n21668 & 1'b0 ) | ( ~n21676 & 1'b0 ) ;
  assign n21678 = ( n21663 & ~n21677 ) | ( n21663 & 1'b0 ) | ( ~n21677 & 1'b0 ) ;
  assign n21679 = n20988 | n21143 ;
  assign n21680 = ( n20993 & ~n20988 ) | ( n20993 & n21001 ) | ( ~n20988 & n21001 ) ;
  assign n21682 = ( n20988 & n21679 ) | ( n20988 & n21680 ) | ( n21679 & n21680 ) ;
  assign n21681 = ( n21001 & ~n21680 ) | ( n21001 & n21679 ) | ( ~n21680 & n21679 ) ;
  assign n21683 = ( n20993 & ~n21682 ) | ( n20993 & n21681 ) | ( ~n21682 & n21681 ) ;
  assign n21684 = ( n976 & n21678 ) | ( n976 & n21683 ) | ( n21678 & n21683 ) ;
  assign n21685 = ( n837 & ~n21684 ) | ( n837 & 1'b0 ) | ( ~n21684 & 1'b0 ) ;
  assign n21686 = ( n21021 & ~n21143 ) | ( n21021 & 1'b0 ) | ( ~n21143 & 1'b0 ) ;
  assign n21687 = ( n21008 & n21017 ) | ( n21008 & n21021 ) | ( n21017 & n21021 ) ;
  assign n21688 = ( n21686 & ~n21017 ) | ( n21686 & n21687 ) | ( ~n21017 & n21687 ) ;
  assign n21689 = ( n21021 & ~n21687 ) | ( n21021 & n21686 ) | ( ~n21687 & n21686 ) ;
  assign n21690 = ( n21008 & ~n21688 ) | ( n21008 & n21689 ) | ( ~n21688 & n21689 ) ;
  assign n21691 = n976 &  n21663 ;
  assign n21692 = ~n21677 & n21691 ;
  assign n21693 = n21683 | n21692 ;
  assign n21694 = ( n21671 & ~n21674 ) | ( n21671 & 1'b0 ) | ( ~n21674 & 1'b0 ) ;
  assign n21695 = ( n1122 & ~n21668 ) | ( n1122 & n21694 ) | ( ~n21668 & n21694 ) ;
  assign n21696 = n976 | n21695 ;
  assign n21697 = ~n837 & n21696 ;
  assign n21698 = n21693 &  n21697 ;
  assign n21699 = ( n21690 & ~n21698 ) | ( n21690 & 1'b0 ) | ( ~n21698 & 1'b0 ) ;
  assign n21700 = n21685 | n21699 ;
  assign n21701 = n21010 | n21143 ;
  assign n21702 = ( n21010 & ~n21023 ) | ( n21010 & n21015 ) | ( ~n21023 & n21015 ) ;
  assign n21703 = ( n21023 & n21701 ) | ( n21023 & n21702 ) | ( n21701 & n21702 ) ;
  assign n21704 = ( n21010 & ~n21702 ) | ( n21010 & n21701 ) | ( ~n21702 & n21701 ) ;
  assign n21705 = ( n21015 & ~n21703 ) | ( n21015 & n21704 ) | ( ~n21703 & n21704 ) ;
  assign n21706 = ( n713 & n21700 ) | ( n713 & n21705 ) | ( n21700 & n21705 ) ;
  assign n21707 = n595 &  n21706 ;
  assign n21708 = n21043 | n21143 ;
  assign n21709 = ( n21030 & n21039 ) | ( n21030 & n21043 ) | ( n21039 & n21043 ) ;
  assign n21710 = ( n21708 & ~n21039 ) | ( n21708 & n21709 ) | ( ~n21039 & n21709 ) ;
  assign n21711 = ( n21043 & ~n21709 ) | ( n21043 & n21708 ) | ( ~n21709 & n21708 ) ;
  assign n21712 = ( n21030 & ~n21710 ) | ( n21030 & n21711 ) | ( ~n21710 & n21711 ) ;
  assign n21713 = n713 | n21685 ;
  assign n21714 = n21699 | n21713 ;
  assign n21715 = n21705 &  n21714 ;
  assign n21716 = n21693 &  n21696 ;
  assign n21717 = ( n837 & ~n21716 ) | ( n837 & n21690 ) | ( ~n21716 & n21690 ) ;
  assign n21718 = n713 &  n21717 ;
  assign n21719 = n595 | n21718 ;
  assign n21720 = n21715 | n21719 ;
  assign n21721 = ~n21712 & n21720 ;
  assign n21722 = n21707 | n21721 ;
  assign n21728 = ( n492 & ~n21727 ) | ( n492 & n21722 ) | ( ~n21727 & n21722 ) ;
  assign n21729 = n396 &  n21728 ;
  assign n21730 = n21065 | n21143 ;
  assign n21731 = ( n21052 & n21061 ) | ( n21052 & n21065 ) | ( n21061 & n21065 ) ;
  assign n21732 = ( n21730 & ~n21061 ) | ( n21730 & n21731 ) | ( ~n21061 & n21731 ) ;
  assign n21733 = ( n21065 & ~n21731 ) | ( n21065 & n21730 ) | ( ~n21731 & n21730 ) ;
  assign n21734 = ( n21052 & ~n21732 ) | ( n21052 & n21733 ) | ( ~n21732 & n21733 ) ;
  assign n21735 = n492 | n21707 ;
  assign n21736 = n21721 | n21735 ;
  assign n21737 = ~n21727 & n21736 ;
  assign n21738 = n21715 | n21718 ;
  assign n21739 = ( n595 & ~n21712 ) | ( n595 & n21738 ) | ( ~n21712 & n21738 ) ;
  assign n21740 = n492 &  n21739 ;
  assign n21741 = n396 | n21740 ;
  assign n21742 = n21737 | n21741 ;
  assign n21743 = ~n21734 & n21742 ;
  assign n21744 = n21729 | n21743 ;
  assign n21750 = ( n315 & ~n21749 ) | ( n315 & n21744 ) | ( ~n21749 & n21744 ) ;
  assign n21751 = n240 &  n21750 ;
  assign n21752 = n21087 | n21143 ;
  assign n21753 = ( n21074 & n21083 ) | ( n21074 & n21087 ) | ( n21083 & n21087 ) ;
  assign n21754 = ( n21752 & ~n21083 ) | ( n21752 & n21753 ) | ( ~n21083 & n21753 ) ;
  assign n21755 = ( n21087 & ~n21753 ) | ( n21087 & n21752 ) | ( ~n21753 & n21752 ) ;
  assign n21756 = ( n21074 & ~n21754 ) | ( n21074 & n21755 ) | ( ~n21754 & n21755 ) ;
  assign n21757 = n315 | n21729 ;
  assign n21758 = n21743 | n21757 ;
  assign n21759 = ~n21749 & n21758 ;
  assign n21760 = n21737 | n21740 ;
  assign n21761 = ( n396 & ~n21734 ) | ( n396 & n21760 ) | ( ~n21734 & n21760 ) ;
  assign n21762 = n315 &  n21761 ;
  assign n21763 = n240 | n21762 ;
  assign n21764 = n21759 | n21763 ;
  assign n21765 = ~n21756 & n21764 ;
  assign n21766 = n21751 | n21765 ;
  assign n21767 = n21076 | n21143 ;
  assign n21768 = ( n21076 & n21081 ) | ( n21076 & n21089 ) | ( n21081 & n21089 ) ;
  assign n21769 = ( n21767 & ~n21089 ) | ( n21767 & n21768 ) | ( ~n21089 & n21768 ) ;
  assign n21770 = ( n21076 & ~n21768 ) | ( n21076 & n21767 ) | ( ~n21768 & n21767 ) ;
  assign n21771 = ( n21081 & ~n21769 ) | ( n21081 & n21770 ) | ( ~n21769 & n21770 ) ;
  assign n21772 = ( n181 & n21766 ) | ( n181 & n21771 ) | ( n21766 & n21771 ) ;
  assign n21773 = ~n145 & n21772 ;
  assign n21779 = n181 | n21751 ;
  assign n21780 = n21765 | n21779 ;
  assign n21781 = n21771 &  n21780 ;
  assign n21782 = n21759 | n21762 ;
  assign n21783 = ( n240 & ~n21756 ) | ( n240 & n21782 ) | ( ~n21756 & n21782 ) ;
  assign n21784 = n181 &  n21783 ;
  assign n21785 = ( n145 & ~n21784 ) | ( n145 & 1'b0 ) | ( ~n21784 & 1'b0 ) ;
  assign n21786 = ~n21781 & n21785 ;
  assign n21787 = n21778 | n21786 ;
  assign n21788 = ~n21773 & n21787 ;
  assign n21789 = ( n21098 & ~n21106 ) | ( n21098 & n21110 ) | ( ~n21106 & n21110 ) ;
  assign n21790 = ( n21106 & n21143 ) | ( n21106 & n21789 ) | ( n21143 & n21789 ) ;
  assign n21791 = ( n21098 & ~n21789 ) | ( n21098 & n21143 ) | ( ~n21789 & n21143 ) ;
  assign n21792 = ( n21110 & ~n21790 ) | ( n21110 & n21791 ) | ( ~n21790 & n21791 ) ;
  assign n21793 = ( n21788 & ~n150 ) | ( n21788 & n21792 ) | ( ~n150 & n21792 ) ;
  assign n21794 = n21134 | n21143 ;
  assign n21795 = ( n21117 & ~n21131 ) | ( n21117 & n21134 ) | ( ~n21131 & n21134 ) ;
  assign n21796 = ( n21131 & n21794 ) | ( n21131 & n21795 ) | ( n21794 & n21795 ) ;
  assign n21797 = ( n21134 & ~n21795 ) | ( n21134 & n21794 ) | ( ~n21795 & n21794 ) ;
  assign n21798 = ( n21117 & ~n21796 ) | ( n21117 & n21797 ) | ( ~n21796 & n21797 ) ;
  assign n21799 = ( n21118 & ~n21123 ) | ( n21118 & 1'b0 ) | ( ~n21123 & 1'b0 ) ;
  assign n21800 = ~n21143 & n21799 ;
  assign n21801 = ( n21137 & ~n21800 ) | ( n21137 & n21799 ) | ( ~n21800 & n21799 ) ;
  assign n21802 = ( n21798 & ~n21801 ) | ( n21798 & 1'b0 ) | ( ~n21801 & 1'b0 ) ;
  assign n21803 = n21793 &  n21802 ;
  assign n21804 = ( n133 & ~n21803 ) | ( n133 & n21802 ) | ( ~n21803 & n21802 ) ;
  assign n21807 = n21781 | n21784 ;
  assign n21808 = ( n145 & ~n21807 ) | ( n145 & n21778 ) | ( ~n21807 & n21778 ) ;
  assign n21809 = ( n150 & ~n21808 ) | ( n150 & 1'b0 ) | ( ~n21808 & 1'b0 ) ;
  assign n21810 = n21798 | n21809 ;
  assign n21805 = n150 | n21773 ;
  assign n21806 = ( n21787 & ~n21805 ) | ( n21787 & 1'b0 ) | ( ~n21805 & 1'b0 ) ;
  assign n21811 = ~n21792 & n21806 ;
  assign n21812 = ( n21792 & ~n21810 ) | ( n21792 & n21811 ) | ( ~n21810 & n21811 ) ;
  assign n21814 = ( n133 & ~n21123 ) | ( n133 & n21118 ) | ( ~n21123 & n21118 ) ;
  assign n21813 = ( n21123 & ~n21118 ) | ( n21123 & n21143 ) | ( ~n21118 & n21143 ) ;
  assign n21815 = ~n21123 & n21813 ;
  assign n21816 = ( n21123 & n21814 ) | ( n21123 & n21815 ) | ( n21814 & n21815 ) ;
  assign n21817 = n21812 | n21816 ;
  assign n21818 = ~n21804 |  n21817 ;
  assign n22483 = ( n21773 & ~n21778 ) | ( n21773 & n21818 ) | ( ~n21778 & n21818 ) ;
  assign n22482 = n21786 &  n21818 ;
  assign n22484 = ( n21818 & ~n22483 ) | ( n21818 & n22482 ) | ( ~n22483 & n22482 ) ;
  assign n22485 = ( n22482 & ~n21773 ) | ( n22482 & n22483 ) | ( ~n21773 & n22483 ) ;
  assign n22486 = ( n21778 & ~n22484 ) | ( n21778 & n22485 ) | ( ~n22484 & n22485 ) ;
  assign n22468 = ( n21780 & ~n21771 ) | ( n21780 & n21784 ) | ( ~n21771 & n21784 ) ;
  assign n22467 = n21784 | n21818 ;
  assign n22470 = ( n21784 & ~n22468 ) | ( n21784 & n22467 ) | ( ~n22468 & n22467 ) ;
  assign n22469 = ( n22467 & ~n21780 ) | ( n22467 & n22468 ) | ( ~n21780 & n22468 ) ;
  assign n22471 = ( n21771 & ~n22470 ) | ( n21771 & n22469 ) | ( ~n22470 & n22469 ) ;
  assign n22461 = ( n21751 & ~n21756 ) | ( n21751 & n21764 ) | ( ~n21756 & n21764 ) ;
  assign n22460 = n21751 | n21818 ;
  assign n22463 = ( n21751 & ~n22461 ) | ( n21751 & n22460 ) | ( ~n22461 & n22460 ) ;
  assign n22462 = ( n22460 & ~n21764 ) | ( n22460 & n22461 ) | ( ~n21764 & n22461 ) ;
  assign n22464 = ( n21756 & ~n22463 ) | ( n21756 & n22462 ) | ( ~n22463 & n22462 ) ;
  assign n22445 = n21762 | n21818 ;
  assign n22446 = ( n21749 & n21758 ) | ( n21749 & n21762 ) | ( n21758 & n21762 ) ;
  assign n22447 = ( n22445 & ~n21758 ) | ( n22445 & n22446 ) | ( ~n21758 & n22446 ) ;
  assign n22448 = ( n21762 & ~n22446 ) | ( n21762 & n22445 ) | ( ~n22446 & n22445 ) ;
  assign n22449 = ( n21749 & ~n22447 ) | ( n21749 & n22448 ) | ( ~n22447 & n22448 ) ;
  assign n22439 = ( n21729 & ~n21734 ) | ( n21729 & n21742 ) | ( ~n21734 & n21742 ) ;
  assign n22438 = n21729 | n21818 ;
  assign n22441 = ( n21729 & ~n22439 ) | ( n21729 & n22438 ) | ( ~n22439 & n22438 ) ;
  assign n22440 = ( n22438 & ~n21742 ) | ( n22438 & n22439 ) | ( ~n21742 & n22439 ) ;
  assign n22442 = ( n21734 & ~n22441 ) | ( n21734 & n22440 ) | ( ~n22441 & n22440 ) ;
  assign n22423 = n21740 | n21818 ;
  assign n22424 = ( n21727 & n21736 ) | ( n21727 & n21740 ) | ( n21736 & n21740 ) ;
  assign n22425 = ( n22423 & ~n21736 ) | ( n22423 & n22424 ) | ( ~n21736 & n22424 ) ;
  assign n22426 = ( n21740 & ~n22424 ) | ( n21740 & n22423 ) | ( ~n22424 & n22423 ) ;
  assign n22427 = ( n21727 & ~n22425 ) | ( n21727 & n22426 ) | ( ~n22425 & n22426 ) ;
  assign n22417 = ( n21707 & ~n21712 ) | ( n21707 & n21720 ) | ( ~n21712 & n21720 ) ;
  assign n22416 = n21707 | n21818 ;
  assign n22419 = ( n21707 & ~n22417 ) | ( n21707 & n22416 ) | ( ~n22417 & n22416 ) ;
  assign n22418 = ( n22416 & ~n21720 ) | ( n22416 & n22417 ) | ( ~n21720 & n22417 ) ;
  assign n22420 = ( n21712 & ~n22419 ) | ( n21712 & n22418 ) | ( ~n22419 & n22418 ) ;
  assign n22402 = ( n21714 & ~n21705 ) | ( n21714 & n21718 ) | ( ~n21705 & n21718 ) ;
  assign n22401 = n21718 | n21818 ;
  assign n22404 = ( n21718 & ~n22402 ) | ( n21718 & n22401 ) | ( ~n22402 & n22401 ) ;
  assign n22403 = ( n22401 & ~n21714 ) | ( n22401 & n22402 ) | ( ~n21714 & n22402 ) ;
  assign n22405 = ( n21705 & ~n22404 ) | ( n21705 & n22403 ) | ( ~n22404 & n22403 ) ;
  assign n22394 = n21685 | n21818 ;
  assign n22395 = ( n21685 & ~n21698 ) | ( n21685 & n21690 ) | ( ~n21698 & n21690 ) ;
  assign n22396 = ( n21698 & n22394 ) | ( n21698 & n22395 ) | ( n22394 & n22395 ) ;
  assign n22397 = ( n21685 & ~n22395 ) | ( n21685 & n22394 ) | ( ~n22395 & n22394 ) ;
  assign n22398 = ( n21690 & ~n22396 ) | ( n21690 & n22397 ) | ( ~n22396 & n22397 ) ;
  assign n22380 = ( n21692 & ~n21683 ) | ( n21692 & n21696 ) | ( ~n21683 & n21696 ) ;
  assign n22379 = ( n21696 & ~n21818 ) | ( n21696 & 1'b0 ) | ( ~n21818 & 1'b0 ) ;
  assign n22382 = ( n21696 & ~n22380 ) | ( n21696 & n22379 ) | ( ~n22380 & n22379 ) ;
  assign n22381 = ( n22379 & ~n21692 ) | ( n22379 & n22380 ) | ( ~n21692 & n22380 ) ;
  assign n22383 = ( n21683 & ~n22382 ) | ( n21683 & n22381 ) | ( ~n22382 & n22381 ) ;
  assign n22373 = ( n21663 & ~n21668 ) | ( n21663 & n21676 ) | ( ~n21668 & n21676 ) ;
  assign n22372 = ( n21663 & ~n21818 ) | ( n21663 & 1'b0 ) | ( ~n21818 & 1'b0 ) ;
  assign n22375 = ( n21663 & ~n22373 ) | ( n21663 & n22372 ) | ( ~n22373 & n22372 ) ;
  assign n22374 = ( n22372 & ~n21676 ) | ( n22372 & n22373 ) | ( ~n21676 & n22373 ) ;
  assign n22376 = ( n21668 & ~n22375 ) | ( n21668 & n22374 ) | ( ~n22375 & n22374 ) ;
  assign n22357 = n21674 | n21818 ;
  assign n22358 = ( n21661 & ~n21670 ) | ( n21661 & n21674 ) | ( ~n21670 & n21674 ) ;
  assign n22359 = ( n21670 & n22357 ) | ( n21670 & n22358 ) | ( n22357 & n22358 ) ;
  assign n22360 = ( n21674 & ~n22358 ) | ( n21674 & n22357 ) | ( ~n22358 & n22357 ) ;
  assign n22361 = ( n21661 & ~n22359 ) | ( n21661 & n22360 ) | ( ~n22359 & n22360 ) ;
  assign n22350 = n21641 | n21818 ;
  assign n22351 = ( n21646 & ~n21641 ) | ( n21646 & n21654 ) | ( ~n21641 & n21654 ) ;
  assign n22353 = ( n21641 & n22350 ) | ( n21641 & n22351 ) | ( n22350 & n22351 ) ;
  assign n22352 = ( n21654 & ~n22351 ) | ( n21654 & n22350 ) | ( ~n22351 & n22350 ) ;
  assign n22354 = ( n21646 & ~n22353 ) | ( n21646 & n22352 ) | ( ~n22353 & n22352 ) ;
  assign n22335 = n21652 | n21818 ;
  assign n22336 = ( n21639 & ~n21652 ) | ( n21639 & n21648 ) | ( ~n21652 & n21648 ) ;
  assign n22338 = ( n21652 & n22335 ) | ( n21652 & n22336 ) | ( n22335 & n22336 ) ;
  assign n22337 = ( n21648 & ~n22336 ) | ( n21648 & n22335 ) | ( ~n22336 & n22335 ) ;
  assign n22339 = ( n21639 & ~n22338 ) | ( n21639 & n22337 ) | ( ~n22338 & n22337 ) ;
  assign n22328 = n21619 | n21818 ;
  assign n22329 = ( n21619 & n21624 ) | ( n21619 & n21632 ) | ( n21624 & n21632 ) ;
  assign n22330 = ( n22328 & ~n21632 ) | ( n22328 & n22329 ) | ( ~n21632 & n22329 ) ;
  assign n22331 = ( n21619 & ~n22329 ) | ( n21619 & n22328 ) | ( ~n22329 & n22328 ) ;
  assign n22332 = ( n21624 & ~n22330 ) | ( n21624 & n22331 ) | ( ~n22330 & n22331 ) ;
  assign n22313 = n21630 | n21818 ;
  assign n22314 = ( n21617 & ~n21630 ) | ( n21617 & n21626 ) | ( ~n21630 & n21626 ) ;
  assign n22316 = ( n21630 & n22313 ) | ( n21630 & n22314 ) | ( n22313 & n22314 ) ;
  assign n22315 = ( n21626 & ~n22314 ) | ( n21626 & n22313 ) | ( ~n22314 & n22313 ) ;
  assign n22317 = ( n21617 & ~n22316 ) | ( n21617 & n22315 ) | ( ~n22316 & n22315 ) ;
  assign n22306 = n21597 | n21818 ;
  assign n22307 = ( n21597 & n21602 ) | ( n21597 & n21610 ) | ( n21602 & n21610 ) ;
  assign n22308 = ( n22306 & ~n21610 ) | ( n22306 & n22307 ) | ( ~n21610 & n22307 ) ;
  assign n22309 = ( n21597 & ~n22307 ) | ( n21597 & n22306 ) | ( ~n22307 & n22306 ) ;
  assign n22310 = ( n21602 & ~n22308 ) | ( n21602 & n22309 ) | ( ~n22308 & n22309 ) ;
  assign n22291 = n21608 | n21818 ;
  assign n22292 = ( n21595 & ~n21608 ) | ( n21595 & n21604 ) | ( ~n21608 & n21604 ) ;
  assign n22294 = ( n21608 & n22291 ) | ( n21608 & n22292 ) | ( n22291 & n22292 ) ;
  assign n22293 = ( n21604 & ~n22292 ) | ( n21604 & n22291 ) | ( ~n22292 & n22291 ) ;
  assign n22295 = ( n21595 & ~n22294 ) | ( n21595 & n22293 ) | ( ~n22294 & n22293 ) ;
  assign n22284 = n21575 | n21818 ;
  assign n22285 = ( n21580 & ~n21575 ) | ( n21580 & n21588 ) | ( ~n21575 & n21588 ) ;
  assign n22287 = ( n21575 & n22284 ) | ( n21575 & n22285 ) | ( n22284 & n22285 ) ;
  assign n22286 = ( n21588 & ~n22285 ) | ( n21588 & n22284 ) | ( ~n22285 & n22284 ) ;
  assign n22288 = ( n21580 & ~n22287 ) | ( n21580 & n22286 ) | ( ~n22287 & n22286 ) ;
  assign n22269 = n21586 | n21818 ;
  assign n22270 = ( n21573 & ~n21582 ) | ( n21573 & n21586 ) | ( ~n21582 & n21586 ) ;
  assign n22271 = ( n21582 & n22269 ) | ( n21582 & n22270 ) | ( n22269 & n22270 ) ;
  assign n22272 = ( n21586 & ~n22270 ) | ( n21586 & n22269 ) | ( ~n22270 & n22269 ) ;
  assign n22273 = ( n21573 & ~n22271 ) | ( n21573 & n22272 ) | ( ~n22271 & n22272 ) ;
  assign n22262 = n21553 | n21818 ;
  assign n22263 = ( n21558 & ~n21553 ) | ( n21558 & n21566 ) | ( ~n21553 & n21566 ) ;
  assign n22265 = ( n21553 & n22262 ) | ( n21553 & n22263 ) | ( n22262 & n22263 ) ;
  assign n22264 = ( n21566 & ~n22263 ) | ( n21566 & n22262 ) | ( ~n22263 & n22262 ) ;
  assign n22266 = ( n21558 & ~n22265 ) | ( n21558 & n22264 ) | ( ~n22265 & n22264 ) ;
  assign n22247 = n21564 | n21818 ;
  assign n22248 = ( n21551 & ~n21560 ) | ( n21551 & n21564 ) | ( ~n21560 & n21564 ) ;
  assign n22249 = ( n21560 & n22247 ) | ( n21560 & n22248 ) | ( n22247 & n22248 ) ;
  assign n22250 = ( n21564 & ~n22248 ) | ( n21564 & n22247 ) | ( ~n22248 & n22247 ) ;
  assign n22251 = ( n21551 & ~n22249 ) | ( n21551 & n22250 ) | ( ~n22249 & n22250 ) ;
  assign n22240 = n21531 | n21818 ;
  assign n22241 = ( n21536 & ~n21531 ) | ( n21536 & n21544 ) | ( ~n21531 & n21544 ) ;
  assign n22243 = ( n21531 & n22240 ) | ( n21531 & n22241 ) | ( n22240 & n22241 ) ;
  assign n22242 = ( n21544 & ~n22241 ) | ( n21544 & n22240 ) | ( ~n22241 & n22240 ) ;
  assign n22244 = ( n21536 & ~n22243 ) | ( n21536 & n22242 ) | ( ~n22243 & n22242 ) ;
  assign n22225 = n21542 | n21818 ;
  assign n22226 = ( n21529 & ~n21538 ) | ( n21529 & n21542 ) | ( ~n21538 & n21542 ) ;
  assign n22227 = ( n21538 & n22225 ) | ( n21538 & n22226 ) | ( n22225 & n22226 ) ;
  assign n22228 = ( n21542 & ~n22226 ) | ( n21542 & n22225 ) | ( ~n22226 & n22225 ) ;
  assign n22229 = ( n21529 & ~n22227 ) | ( n21529 & n22228 ) | ( ~n22227 & n22228 ) ;
  assign n22218 = n21509 | n21818 ;
  assign n22219 = ( n21514 & ~n21509 ) | ( n21514 & n21522 ) | ( ~n21509 & n21522 ) ;
  assign n22221 = ( n21509 & n22218 ) | ( n21509 & n22219 ) | ( n22218 & n22219 ) ;
  assign n22220 = ( n21522 & ~n22219 ) | ( n21522 & n22218 ) | ( ~n22219 & n22218 ) ;
  assign n22222 = ( n21514 & ~n22221 ) | ( n21514 & n22220 ) | ( ~n22221 & n22220 ) ;
  assign n22203 = n21520 | n21818 ;
  assign n22204 = ( n21507 & ~n21516 ) | ( n21507 & n21520 ) | ( ~n21516 & n21520 ) ;
  assign n22205 = ( n21516 & n22203 ) | ( n21516 & n22204 ) | ( n22203 & n22204 ) ;
  assign n22206 = ( n21520 & ~n22204 ) | ( n21520 & n22203 ) | ( ~n22204 & n22203 ) ;
  assign n22207 = ( n21507 & ~n22205 ) | ( n21507 & n22206 ) | ( ~n22205 & n22206 ) ;
  assign n22196 = n21487 | n21818 ;
  assign n22197 = ( n21492 & ~n21487 ) | ( n21492 & n21500 ) | ( ~n21487 & n21500 ) ;
  assign n22199 = ( n21487 & n22196 ) | ( n21487 & n22197 ) | ( n22196 & n22197 ) ;
  assign n22198 = ( n21500 & ~n22197 ) | ( n21500 & n22196 ) | ( ~n22197 & n22196 ) ;
  assign n22200 = ( n21492 & ~n22199 ) | ( n21492 & n22198 ) | ( ~n22199 & n22198 ) ;
  assign n22181 = n21498 | n21818 ;
  assign n22182 = ( n21485 & ~n21494 ) | ( n21485 & n21498 ) | ( ~n21494 & n21498 ) ;
  assign n22183 = ( n21494 & n22181 ) | ( n21494 & n22182 ) | ( n22181 & n22182 ) ;
  assign n22184 = ( n21498 & ~n22182 ) | ( n21498 & n22181 ) | ( ~n22182 & n22181 ) ;
  assign n22185 = ( n21485 & ~n22183 ) | ( n21485 & n22184 ) | ( ~n22183 & n22184 ) ;
  assign n22174 = ( n21465 & ~n21818 ) | ( n21465 & 1'b0 ) | ( ~n21818 & 1'b0 ) ;
  assign n22175 = ( n21465 & n21470 ) | ( n21465 & n21478 ) | ( n21470 & n21478 ) ;
  assign n22176 = ( n22174 & ~n21478 ) | ( n22174 & n22175 ) | ( ~n21478 & n22175 ) ;
  assign n22177 = ( n21465 & ~n22175 ) | ( n21465 & n22174 ) | ( ~n22175 & n22174 ) ;
  assign n22178 = ( n21470 & ~n22176 ) | ( n21470 & n22177 ) | ( ~n22176 & n22177 ) ;
  assign n22159 = n21476 | n21818 ;
  assign n22160 = ( n21463 & ~n21472 ) | ( n21463 & n21476 ) | ( ~n21472 & n21476 ) ;
  assign n22161 = ( n21472 & n22159 ) | ( n21472 & n22160 ) | ( n22159 & n22160 ) ;
  assign n22162 = ( n21476 & ~n22160 ) | ( n21476 & n22159 ) | ( ~n22160 & n22159 ) ;
  assign n22163 = ( n21463 & ~n22161 ) | ( n21463 & n22162 ) | ( ~n22161 & n22162 ) ;
  assign n22152 = ( n21443 & ~n21818 ) | ( n21443 & 1'b0 ) | ( ~n21818 & 1'b0 ) ;
  assign n22153 = ( n21443 & n21448 ) | ( n21443 & n21456 ) | ( n21448 & n21456 ) ;
  assign n22154 = ( n22152 & ~n21456 ) | ( n22152 & n22153 ) | ( ~n21456 & n22153 ) ;
  assign n22155 = ( n21443 & ~n22153 ) | ( n21443 & n22152 ) | ( ~n22153 & n22152 ) ;
  assign n22156 = ( n21448 & ~n22154 ) | ( n21448 & n22155 ) | ( ~n22154 & n22155 ) ;
  assign n22137 = n21454 | n21818 ;
  assign n22138 = ( n21441 & ~n21450 ) | ( n21441 & n21454 ) | ( ~n21450 & n21454 ) ;
  assign n22139 = ( n21450 & n22137 ) | ( n21450 & n22138 ) | ( n22137 & n22138 ) ;
  assign n22140 = ( n21454 & ~n22138 ) | ( n21454 & n22137 ) | ( ~n22138 & n22137 ) ;
  assign n22141 = ( n21441 & ~n22139 ) | ( n21441 & n22140 ) | ( ~n22139 & n22140 ) ;
  assign n22130 = ( n21421 & ~n21818 ) | ( n21421 & 1'b0 ) | ( ~n21818 & 1'b0 ) ;
  assign n22131 = ( n21421 & n21426 ) | ( n21421 & n21434 ) | ( n21426 & n21434 ) ;
  assign n22132 = ( n22130 & ~n21434 ) | ( n22130 & n22131 ) | ( ~n21434 & n22131 ) ;
  assign n22133 = ( n21421 & ~n22131 ) | ( n21421 & n22130 ) | ( ~n22131 & n22130 ) ;
  assign n22134 = ( n21426 & ~n22132 ) | ( n21426 & n22133 ) | ( ~n22132 & n22133 ) ;
  assign n22116 = ( n21428 & ~n21419 ) | ( n21428 & n21432 ) | ( ~n21419 & n21432 ) ;
  assign n22115 = ( n21432 & ~n21818 ) | ( n21432 & 1'b0 ) | ( ~n21818 & 1'b0 ) ;
  assign n22118 = ( n21432 & ~n22116 ) | ( n21432 & n22115 ) | ( ~n22116 & n22115 ) ;
  assign n22117 = ( n22115 & ~n21428 ) | ( n22115 & n22116 ) | ( ~n21428 & n22116 ) ;
  assign n22119 = ( n21419 & ~n22118 ) | ( n21419 & n22117 ) | ( ~n22118 & n22117 ) ;
  assign n22108 = n21399 | n21818 ;
  assign n22109 = ( n21404 & ~n21399 ) | ( n21404 & n21412 ) | ( ~n21399 & n21412 ) ;
  assign n22111 = ( n21399 & n22108 ) | ( n21399 & n22109 ) | ( n22108 & n22109 ) ;
  assign n22110 = ( n21412 & ~n22109 ) | ( n21412 & n22108 ) | ( ~n22109 & n22108 ) ;
  assign n22112 = ( n21404 & ~n22111 ) | ( n21404 & n22110 ) | ( ~n22111 & n22110 ) ;
  assign n22093 = n21410 | n21818 ;
  assign n22094 = ( n21397 & ~n21410 ) | ( n21397 & n21406 ) | ( ~n21410 & n21406 ) ;
  assign n22096 = ( n21410 & n22093 ) | ( n21410 & n22094 ) | ( n22093 & n22094 ) ;
  assign n22095 = ( n21406 & ~n22094 ) | ( n21406 & n22093 ) | ( ~n22094 & n22093 ) ;
  assign n22097 = ( n21397 & ~n22096 ) | ( n21397 & n22095 ) | ( ~n22096 & n22095 ) ;
  assign n22086 = n21390 &  n21818 ;
  assign n22087 = ( n21377 & n21382 ) | ( n21377 & n21818 ) | ( n21382 & n21818 ) ;
  assign n22089 = ( n22086 & ~n21377 ) | ( n22086 & n22087 ) | ( ~n21377 & n22087 ) ;
  assign n22088 = ( n21818 & ~n22087 ) | ( n21818 & n22086 ) | ( ~n22087 & n22086 ) ;
  assign n22090 = ( n21382 & ~n22089 ) | ( n21382 & n22088 ) | ( ~n22089 & n22088 ) ;
  assign n22071 = n21388 | n21818 ;
  assign n22072 = ( n21375 & ~n21384 ) | ( n21375 & n21388 ) | ( ~n21384 & n21388 ) ;
  assign n22073 = ( n21384 & n22071 ) | ( n21384 & n22072 ) | ( n22071 & n22072 ) ;
  assign n22074 = ( n21388 & ~n22072 ) | ( n21388 & n22071 ) | ( ~n22072 & n22071 ) ;
  assign n22075 = ( n21375 & ~n22073 ) | ( n21375 & n22074 ) | ( ~n22073 & n22074 ) ;
  assign n22064 = n21368 &  n21818 ;
  assign n22065 = ( n21360 & ~n21355 ) | ( n21360 & n21818 ) | ( ~n21355 & n21818 ) ;
  assign n22067 = ( n22064 & n21355 ) | ( n22064 & n22065 ) | ( n21355 & n22065 ) ;
  assign n22066 = ( n21818 & ~n22065 ) | ( n21818 & n22064 ) | ( ~n22065 & n22064 ) ;
  assign n22068 = ( n21360 & ~n22067 ) | ( n21360 & n22066 ) | ( ~n22067 & n22066 ) ;
  assign n22049 = n21366 | n21818 ;
  assign n22050 = ( n21353 & ~n21366 ) | ( n21353 & n21362 ) | ( ~n21366 & n21362 ) ;
  assign n22052 = ( n21366 & n22049 ) | ( n21366 & n22050 ) | ( n22049 & n22050 ) ;
  assign n22051 = ( n21362 & ~n22050 ) | ( n21362 & n22049 ) | ( ~n22050 & n22049 ) ;
  assign n22053 = ( n21353 & ~n22052 ) | ( n21353 & n22051 ) | ( ~n22052 & n22051 ) ;
  assign n22043 = ( n21333 & ~n21338 ) | ( n21333 & n21818 ) | ( ~n21338 & n21818 ) ;
  assign n22042 = n21346 &  n21818 ;
  assign n22044 = ( n21818 & ~n22043 ) | ( n21818 & n22042 ) | ( ~n22043 & n22042 ) ;
  assign n22045 = ( n22042 & ~n21333 ) | ( n22042 & n22043 ) | ( ~n21333 & n22043 ) ;
  assign n22046 = ( n21338 & ~n22044 ) | ( n21338 & n22045 ) | ( ~n22044 & n22045 ) ;
  assign n22027 = n21344 | n21818 ;
  assign n22028 = ( n21331 & ~n21344 ) | ( n21331 & n21340 ) | ( ~n21344 & n21340 ) ;
  assign n22030 = ( n21344 & n22027 ) | ( n21344 & n22028 ) | ( n22027 & n22028 ) ;
  assign n22029 = ( n21340 & ~n22028 ) | ( n21340 & n22027 ) | ( ~n22028 & n22027 ) ;
  assign n22031 = ( n21331 & ~n22030 ) | ( n21331 & n22029 ) | ( ~n22030 & n22029 ) ;
  assign n22021 = ( n21311 & ~n21316 ) | ( n21311 & n21818 ) | ( ~n21316 & n21818 ) ;
  assign n22020 = n21324 &  n21818 ;
  assign n22022 = ( n21818 & ~n22021 ) | ( n21818 & n22020 ) | ( ~n22021 & n22020 ) ;
  assign n22023 = ( n22020 & ~n21311 ) | ( n22020 & n22021 ) | ( ~n21311 & n22021 ) ;
  assign n22024 = ( n21316 & ~n22022 ) | ( n21316 & n22023 ) | ( ~n22022 & n22023 ) ;
  assign n22005 = n21322 | n21818 ;
  assign n22006 = ( n21309 & ~n21322 ) | ( n21309 & n21318 ) | ( ~n21322 & n21318 ) ;
  assign n22008 = ( n21322 & n22005 ) | ( n21322 & n22006 ) | ( n22005 & n22006 ) ;
  assign n22007 = ( n21318 & ~n22006 ) | ( n21318 & n22005 ) | ( ~n22006 & n22005 ) ;
  assign n22009 = ( n21309 & ~n22008 ) | ( n21309 & n22007 ) | ( ~n22008 & n22007 ) ;
  assign n21999 = ( n21289 & ~n21294 ) | ( n21289 & n21818 ) | ( ~n21294 & n21818 ) ;
  assign n21998 = n21302 &  n21818 ;
  assign n22000 = ( n21818 & ~n21999 ) | ( n21818 & n21998 ) | ( ~n21999 & n21998 ) ;
  assign n22001 = ( n21998 & ~n21289 ) | ( n21998 & n21999 ) | ( ~n21289 & n21999 ) ;
  assign n22002 = ( n21294 & ~n22000 ) | ( n21294 & n22001 ) | ( ~n22000 & n22001 ) ;
  assign n21983 = n21300 | n21818 ;
  assign n21984 = ( n21287 & ~n21300 ) | ( n21287 & n21296 ) | ( ~n21300 & n21296 ) ;
  assign n21986 = ( n21300 & n21983 ) | ( n21300 & n21984 ) | ( n21983 & n21984 ) ;
  assign n21985 = ( n21296 & ~n21984 ) | ( n21296 & n21983 ) | ( ~n21984 & n21983 ) ;
  assign n21987 = ( n21287 & ~n21986 ) | ( n21287 & n21985 ) | ( ~n21986 & n21985 ) ;
  assign n21977 = ( n21267 & ~n21272 ) | ( n21267 & n21818 ) | ( ~n21272 & n21818 ) ;
  assign n21976 = n21280 &  n21818 ;
  assign n21978 = ( n21818 & ~n21977 ) | ( n21818 & n21976 ) | ( ~n21977 & n21976 ) ;
  assign n21979 = ( n21976 & ~n21267 ) | ( n21976 & n21977 ) | ( ~n21267 & n21977 ) ;
  assign n21980 = ( n21272 & ~n21978 ) | ( n21272 & n21979 ) | ( ~n21978 & n21979 ) ;
  assign n21961 = n21278 | n21818 ;
  assign n21962 = ( n21265 & ~n21278 ) | ( n21265 & n21274 ) | ( ~n21278 & n21274 ) ;
  assign n21964 = ( n21278 & n21961 ) | ( n21278 & n21962 ) | ( n21961 & n21962 ) ;
  assign n21963 = ( n21274 & ~n21962 ) | ( n21274 & n21961 ) | ( ~n21962 & n21961 ) ;
  assign n21965 = ( n21265 & ~n21964 ) | ( n21265 & n21963 ) | ( ~n21964 & n21963 ) ;
  assign n21955 = ( n21245 & ~n21250 ) | ( n21245 & n21818 ) | ( ~n21250 & n21818 ) ;
  assign n21954 = n21258 &  n21818 ;
  assign n21956 = ( n21818 & ~n21955 ) | ( n21818 & n21954 ) | ( ~n21955 & n21954 ) ;
  assign n21957 = ( n21954 & ~n21245 ) | ( n21954 & n21955 ) | ( ~n21245 & n21955 ) ;
  assign n21958 = ( n21250 & ~n21956 ) | ( n21250 & n21957 ) | ( ~n21956 & n21957 ) ;
  assign n21939 = n21256 | n21818 ;
  assign n21940 = ( n21243 & ~n21256 ) | ( n21243 & n21252 ) | ( ~n21256 & n21252 ) ;
  assign n21942 = ( n21256 & n21939 ) | ( n21256 & n21940 ) | ( n21939 & n21940 ) ;
  assign n21941 = ( n21252 & ~n21940 ) | ( n21252 & n21939 ) | ( ~n21940 & n21939 ) ;
  assign n21943 = ( n21243 & ~n21942 ) | ( n21243 & n21941 ) | ( ~n21942 & n21941 ) ;
  assign n21932 = n21236 &  n21818 ;
  assign n21933 = ( n21223 & n21228 ) | ( n21223 & n21818 ) | ( n21228 & n21818 ) ;
  assign n21935 = ( n21932 & ~n21223 ) | ( n21932 & n21933 ) | ( ~n21223 & n21933 ) ;
  assign n21934 = ( n21818 & ~n21933 ) | ( n21818 & n21932 ) | ( ~n21933 & n21932 ) ;
  assign n21936 = ( n21228 & ~n21935 ) | ( n21228 & n21934 ) | ( ~n21935 & n21934 ) ;
  assign n21917 = n21234 | n21818 ;
  assign n21918 = ( n21221 & ~n21234 ) | ( n21221 & n21230 ) | ( ~n21234 & n21230 ) ;
  assign n21920 = ( n21234 & n21917 ) | ( n21234 & n21918 ) | ( n21917 & n21918 ) ;
  assign n21919 = ( n21230 & ~n21918 ) | ( n21230 & n21917 ) | ( ~n21918 & n21917 ) ;
  assign n21921 = ( n21221 & ~n21920 ) | ( n21221 & n21919 ) | ( ~n21920 & n21919 ) ;
  assign n21910 = n21214 &  n21818 ;
  assign n21911 = ( n21201 & n21206 ) | ( n21201 & n21818 ) | ( n21206 & n21818 ) ;
  assign n21913 = ( n21910 & ~n21201 ) | ( n21910 & n21911 ) | ( ~n21201 & n21911 ) ;
  assign n21912 = ( n21818 & ~n21911 ) | ( n21818 & n21910 ) | ( ~n21911 & n21910 ) ;
  assign n21914 = ( n21206 & ~n21913 ) | ( n21206 & n21912 ) | ( ~n21913 & n21912 ) ;
  assign n21895 = n21212 | n21818 ;
  assign n21896 = ( n21199 & ~n21212 ) | ( n21199 & n21208 ) | ( ~n21212 & n21208 ) ;
  assign n21898 = ( n21212 & n21895 ) | ( n21212 & n21896 ) | ( n21895 & n21896 ) ;
  assign n21897 = ( n21208 & ~n21896 ) | ( n21208 & n21895 ) | ( ~n21896 & n21895 ) ;
  assign n21899 = ( n21199 & ~n21898 ) | ( n21199 & n21897 ) | ( ~n21898 & n21897 ) ;
  assign n21889 = ( n21179 & ~n21184 ) | ( n21179 & n21818 ) | ( ~n21184 & n21818 ) ;
  assign n21888 = n21192 &  n21818 ;
  assign n21890 = ( n21818 & ~n21889 ) | ( n21818 & n21888 ) | ( ~n21889 & n21888 ) ;
  assign n21891 = ( n21888 & ~n21179 ) | ( n21888 & n21889 ) | ( ~n21179 & n21889 ) ;
  assign n21892 = ( n21184 & ~n21890 ) | ( n21184 & n21891 ) | ( ~n21890 & n21891 ) ;
  assign n21873 = n21190 | n21818 ;
  assign n21874 = ( n21177 & ~n21190 ) | ( n21177 & n21186 ) | ( ~n21190 & n21186 ) ;
  assign n21876 = ( n21190 & n21873 ) | ( n21190 & n21874 ) | ( n21873 & n21874 ) ;
  assign n21875 = ( n21186 & ~n21874 ) | ( n21186 & n21873 ) | ( ~n21874 & n21873 ) ;
  assign n21877 = ( n21177 & ~n21876 ) | ( n21177 & n21875 ) | ( ~n21876 & n21875 ) ;
  assign n21866 = ( n21154 & ~n21156 ) | ( n21154 & 1'b0 ) | ( ~n21156 & 1'b0 ) ;
  assign n21867 = ( n21156 & ~n21866 ) | ( n21156 & n21165 ) | ( ~n21866 & n21165 ) ;
  assign n21869 = ( n21818 & n21866 ) | ( n21818 & n21867 ) | ( n21866 & n21867 ) ;
  assign n21868 = ( n21156 & ~n21867 ) | ( n21156 & n21818 ) | ( ~n21867 & n21818 ) ;
  assign n21870 = ( n21165 & ~n21869 ) | ( n21165 & n21868 ) | ( ~n21869 & n21868 ) ;
  assign n21850 = ~x6 & n21143 ;
  assign n21851 = ( x7 & ~n21850 ) | ( x7 & 1'b0 ) | ( ~n21850 & 1'b0 ) ;
  assign n21852 = n21157 | n21851 ;
  assign n21847 = ( n21143 & ~x6 ) | ( n21143 & n21149 ) | ( ~x6 & n21149 ) ;
  assign n21848 = x6 &  n21847 ;
  assign n21849 = ( n21145 & ~n21848 ) | ( n21145 & n21149 ) | ( ~n21848 & n21149 ) ;
  assign n21853 = ( n21818 & ~n21852 ) | ( n21818 & n21849 ) | ( ~n21852 & n21849 ) ;
  assign n21855 = ( n21818 & ~n21853 ) | ( n21818 & 1'b0 ) | ( ~n21853 & 1'b0 ) ;
  assign n21854 = ~n21849 & n21853 ;
  assign n21856 = ( n21852 & ~n21855 ) | ( n21852 & n21854 ) | ( ~n21855 & n21854 ) ;
  assign n21837 = ( n21143 & ~n21816 ) | ( n21143 & 1'b0 ) | ( ~n21816 & 1'b0 ) ;
  assign n21838 = ( n21804 & ~n21837 ) | ( n21804 & n21812 ) | ( ~n21837 & n21812 ) ;
  assign n21839 = ( n21804 & ~n21838 ) | ( n21804 & 1'b0 ) | ( ~n21838 & 1'b0 ) ;
  assign n21830 = ~n20476 & n21818 ;
  assign n21840 = ( n21830 & ~n21839 ) | ( n21830 & 1'b0 ) | ( ~n21839 & 1'b0 ) ;
  assign n21841 = ( x6 & n21839 ) | ( x6 & n21840 ) | ( n21839 & n21840 ) ;
  assign n21842 = x6 | n21839 ;
  assign n21843 = n21830 | n21842 ;
  assign n21844 = ~n21841 & n21843 ;
  assign n21832 = ( x4 & ~n21818 ) | ( x4 & x5 ) | ( ~n21818 & x5 ) ;
  assign n21834 = ( x4 & ~x5 ) | ( x4 & 1'b0 ) | ( ~x5 & 1'b0 ) ;
  assign n21820 = x2 | x3 ;
  assign n21821 = ~x4 & n21820 ;
  assign n21822 = ( x4 & ~n21142 ) | ( x4 & n21821 ) | ( ~n21142 & n21821 ) ;
  assign n21823 = n21129 &  n21822 ;
  assign n21833 = ( n21818 & ~x5 ) | ( n21818 & n21823 ) | ( ~x5 & n21823 ) ;
  assign n21835 = ( n21832 & ~n21834 ) | ( n21832 & n21833 ) | ( ~n21834 & n21833 ) ;
  assign n21824 = x4 | n21820 ;
  assign n21819 = x4 &  n21818 ;
  assign n21825 = ( n21143 & ~n21824 ) | ( n21143 & n21819 ) | ( ~n21824 & n21819 ) ;
  assign n21857 = n20475 | n21825 ;
  assign n21858 = ( n21835 & ~n21857 ) | ( n21835 & 1'b0 ) | ( ~n21857 & 1'b0 ) ;
  assign n21859 = n21844 | n21858 ;
  assign n21860 = n21825 &  n21835 ;
  assign n21861 = ( n20475 & ~n21835 ) | ( n20475 & n21860 ) | ( ~n21835 & n21860 ) ;
  assign n21862 = n19819 | n21861 ;
  assign n21863 = ( n21859 & ~n21862 ) | ( n21859 & 1'b0 ) | ( ~n21862 & 1'b0 ) ;
  assign n21864 = n21856 | n21863 ;
  assign n21836 = ~n21825 & n21835 ;
  assign n21845 = ( n21836 & ~n20475 ) | ( n21836 & n21844 ) | ( ~n20475 & n21844 ) ;
  assign n21846 = ( n19819 & ~n21845 ) | ( n19819 & 1'b0 ) | ( ~n21845 & 1'b0 ) ;
  assign n21878 = n19175 | n21846 ;
  assign n21879 = ( n21864 & ~n21878 ) | ( n21864 & 1'b0 ) | ( ~n21878 & 1'b0 ) ;
  assign n21880 = n21870 | n21879 ;
  assign n21881 = ( n21859 & ~n21861 ) | ( n21859 & 1'b0 ) | ( ~n21861 & 1'b0 ) ;
  assign n21882 = ( n21856 & ~n19819 ) | ( n21856 & n21881 ) | ( ~n19819 & n21881 ) ;
  assign n21883 = ( n19175 & ~n21882 ) | ( n19175 & 1'b0 ) | ( ~n21882 & 1'b0 ) ;
  assign n21884 = n18532 | n21883 ;
  assign n21885 = ( n21880 & ~n21884 ) | ( n21880 & 1'b0 ) | ( ~n21884 & 1'b0 ) ;
  assign n21886 = n21877 | n21885 ;
  assign n21865 = ~n21846 & n21864 ;
  assign n21871 = ( n21865 & ~n19175 ) | ( n21865 & n21870 ) | ( ~n19175 & n21870 ) ;
  assign n21872 = ( n18532 & ~n21871 ) | ( n18532 & 1'b0 ) | ( ~n21871 & 1'b0 ) ;
  assign n21900 = n17902 | n21872 ;
  assign n21901 = ( n21886 & ~n21900 ) | ( n21886 & 1'b0 ) | ( ~n21900 & 1'b0 ) ;
  assign n21902 = n21892 | n21901 ;
  assign n21903 = ( n21880 & ~n21883 ) | ( n21880 & 1'b0 ) | ( ~n21883 & 1'b0 ) ;
  assign n21904 = ( n21877 & ~n18532 ) | ( n21877 & n21903 ) | ( ~n18532 & n21903 ) ;
  assign n21905 = ( n17902 & ~n21904 ) | ( n17902 & 1'b0 ) | ( ~n21904 & 1'b0 ) ;
  assign n21906 = n17279 | n21905 ;
  assign n21907 = ( n21902 & ~n21906 ) | ( n21902 & 1'b0 ) | ( ~n21906 & 1'b0 ) ;
  assign n21908 = n21899 | n21907 ;
  assign n21887 = ~n21872 & n21886 ;
  assign n21893 = ( n21887 & ~n17902 ) | ( n21887 & n21892 ) | ( ~n17902 & n21892 ) ;
  assign n21894 = ( n17279 & ~n21893 ) | ( n17279 & 1'b0 ) | ( ~n21893 & 1'b0 ) ;
  assign n21922 = n16671 | n21894 ;
  assign n21923 = ( n21908 & ~n21922 ) | ( n21908 & 1'b0 ) | ( ~n21922 & 1'b0 ) ;
  assign n21924 = n21914 | n21923 ;
  assign n21925 = ( n21902 & ~n21905 ) | ( n21902 & 1'b0 ) | ( ~n21905 & 1'b0 ) ;
  assign n21926 = ( n21899 & ~n17279 ) | ( n21899 & n21925 ) | ( ~n17279 & n21925 ) ;
  assign n21927 = ( n16671 & ~n21926 ) | ( n16671 & 1'b0 ) | ( ~n21926 & 1'b0 ) ;
  assign n21928 = n16070 | n21927 ;
  assign n21929 = ( n21924 & ~n21928 ) | ( n21924 & 1'b0 ) | ( ~n21928 & 1'b0 ) ;
  assign n21930 = n21921 | n21929 ;
  assign n21909 = ~n21894 & n21908 ;
  assign n21915 = ( n21909 & ~n16671 ) | ( n21909 & n21914 ) | ( ~n16671 & n21914 ) ;
  assign n21916 = ( n16070 & ~n21915 ) | ( n16070 & 1'b0 ) | ( ~n21915 & 1'b0 ) ;
  assign n21944 = n15484 | n21916 ;
  assign n21945 = ( n21930 & ~n21944 ) | ( n21930 & 1'b0 ) | ( ~n21944 & 1'b0 ) ;
  assign n21946 = n21936 | n21945 ;
  assign n21947 = ( n21924 & ~n21927 ) | ( n21924 & 1'b0 ) | ( ~n21927 & 1'b0 ) ;
  assign n21948 = ( n21921 & ~n16070 ) | ( n21921 & n21947 ) | ( ~n16070 & n21947 ) ;
  assign n21949 = ( n15484 & ~n21948 ) | ( n15484 & 1'b0 ) | ( ~n21948 & 1'b0 ) ;
  assign n21950 = n14905 | n21949 ;
  assign n21951 = ( n21946 & ~n21950 ) | ( n21946 & 1'b0 ) | ( ~n21950 & 1'b0 ) ;
  assign n21952 = n21943 | n21951 ;
  assign n21931 = ~n21916 & n21930 ;
  assign n21937 = ( n21931 & ~n15484 ) | ( n21931 & n21936 ) | ( ~n15484 & n21936 ) ;
  assign n21938 = ( n14905 & ~n21937 ) | ( n14905 & 1'b0 ) | ( ~n21937 & 1'b0 ) ;
  assign n21966 = n14341 | n21938 ;
  assign n21967 = ( n21952 & ~n21966 ) | ( n21952 & 1'b0 ) | ( ~n21966 & 1'b0 ) ;
  assign n21968 = n21958 | n21967 ;
  assign n21969 = ( n21946 & ~n21949 ) | ( n21946 & 1'b0 ) | ( ~n21949 & 1'b0 ) ;
  assign n21970 = ( n21943 & ~n14905 ) | ( n21943 & n21969 ) | ( ~n14905 & n21969 ) ;
  assign n21971 = ( n14341 & ~n21970 ) | ( n14341 & 1'b0 ) | ( ~n21970 & 1'b0 ) ;
  assign n21972 = n13784 | n21971 ;
  assign n21973 = ( n21968 & ~n21972 ) | ( n21968 & 1'b0 ) | ( ~n21972 & 1'b0 ) ;
  assign n21974 = n21965 | n21973 ;
  assign n21953 = ~n21938 & n21952 ;
  assign n21959 = ( n21953 & ~n14341 ) | ( n21953 & n21958 ) | ( ~n14341 & n21958 ) ;
  assign n21960 = ( n13784 & ~n21959 ) | ( n13784 & 1'b0 ) | ( ~n21959 & 1'b0 ) ;
  assign n21988 = n13242 | n21960 ;
  assign n21989 = ( n21974 & ~n21988 ) | ( n21974 & 1'b0 ) | ( ~n21988 & 1'b0 ) ;
  assign n21990 = n21980 | n21989 ;
  assign n21991 = ( n21968 & ~n21971 ) | ( n21968 & 1'b0 ) | ( ~n21971 & 1'b0 ) ;
  assign n21992 = ( n21965 & ~n13784 ) | ( n21965 & n21991 ) | ( ~n13784 & n21991 ) ;
  assign n21993 = ( n13242 & ~n21992 ) | ( n13242 & 1'b0 ) | ( ~n21992 & 1'b0 ) ;
  assign n21994 = n12707 | n21993 ;
  assign n21995 = ( n21990 & ~n21994 ) | ( n21990 & 1'b0 ) | ( ~n21994 & 1'b0 ) ;
  assign n21996 = n21987 | n21995 ;
  assign n21975 = ~n21960 & n21974 ;
  assign n21981 = ( n21975 & ~n13242 ) | ( n21975 & n21980 ) | ( ~n13242 & n21980 ) ;
  assign n21982 = ( n12707 & ~n21981 ) | ( n12707 & 1'b0 ) | ( ~n21981 & 1'b0 ) ;
  assign n22010 = n12187 | n21982 ;
  assign n22011 = ( n21996 & ~n22010 ) | ( n21996 & 1'b0 ) | ( ~n22010 & 1'b0 ) ;
  assign n22012 = n22002 | n22011 ;
  assign n22013 = ( n21990 & ~n21993 ) | ( n21990 & 1'b0 ) | ( ~n21993 & 1'b0 ) ;
  assign n22014 = ( n21987 & ~n12707 ) | ( n21987 & n22013 ) | ( ~n12707 & n22013 ) ;
  assign n22015 = ( n12187 & ~n22014 ) | ( n12187 & 1'b0 ) | ( ~n22014 & 1'b0 ) ;
  assign n22016 = n11674 | n22015 ;
  assign n22017 = ( n22012 & ~n22016 ) | ( n22012 & 1'b0 ) | ( ~n22016 & 1'b0 ) ;
  assign n22018 = n22009 | n22017 ;
  assign n21997 = ~n21982 & n21996 ;
  assign n22003 = ( n21997 & ~n12187 ) | ( n21997 & n22002 ) | ( ~n12187 & n22002 ) ;
  assign n22004 = ( n11674 & ~n22003 ) | ( n11674 & 1'b0 ) | ( ~n22003 & 1'b0 ) ;
  assign n22032 = n11176 | n22004 ;
  assign n22033 = ( n22018 & ~n22032 ) | ( n22018 & 1'b0 ) | ( ~n22032 & 1'b0 ) ;
  assign n22034 = n22024 | n22033 ;
  assign n22035 = ( n22012 & ~n22015 ) | ( n22012 & 1'b0 ) | ( ~n22015 & 1'b0 ) ;
  assign n22036 = ( n22009 & ~n11674 ) | ( n22009 & n22035 ) | ( ~n11674 & n22035 ) ;
  assign n22037 = ( n11176 & ~n22036 ) | ( n11176 & 1'b0 ) | ( ~n22036 & 1'b0 ) ;
  assign n22038 = n10685 | n22037 ;
  assign n22039 = ( n22034 & ~n22038 ) | ( n22034 & 1'b0 ) | ( ~n22038 & 1'b0 ) ;
  assign n22040 = n22031 | n22039 ;
  assign n22019 = ~n22004 & n22018 ;
  assign n22025 = ( n22019 & ~n11176 ) | ( n22019 & n22024 ) | ( ~n11176 & n22024 ) ;
  assign n22026 = ( n10685 & ~n22025 ) | ( n10685 & 1'b0 ) | ( ~n22025 & 1'b0 ) ;
  assign n22054 = n10209 | n22026 ;
  assign n22055 = ( n22040 & ~n22054 ) | ( n22040 & 1'b0 ) | ( ~n22054 & 1'b0 ) ;
  assign n22056 = n22046 | n22055 ;
  assign n22057 = ( n22034 & ~n22037 ) | ( n22034 & 1'b0 ) | ( ~n22037 & 1'b0 ) ;
  assign n22058 = ( n22031 & ~n10685 ) | ( n22031 & n22057 ) | ( ~n10685 & n22057 ) ;
  assign n22059 = ( n10209 & ~n22058 ) | ( n10209 & 1'b0 ) | ( ~n22058 & 1'b0 ) ;
  assign n22060 = ( n9740 & ~n22059 ) | ( n9740 & 1'b0 ) | ( ~n22059 & 1'b0 ) ;
  assign n22061 = n22056 &  n22060 ;
  assign n22062 = n22053 | n22061 ;
  assign n22041 = ~n22026 & n22040 ;
  assign n22047 = ( n22041 & ~n10209 ) | ( n22041 & n22046 ) | ( ~n10209 & n22046 ) ;
  assign n22048 = n9740 | n22047 ;
  assign n22076 = ~n9286 & n22048 ;
  assign n22077 = n22062 &  n22076 ;
  assign n22078 = n22068 | n22077 ;
  assign n22079 = ( n22056 & ~n22059 ) | ( n22056 & 1'b0 ) | ( ~n22059 & 1'b0 ) ;
  assign n22080 = ( n9740 & n22053 ) | ( n9740 & n22079 ) | ( n22053 & n22079 ) ;
  assign n22081 = ( n9286 & ~n22080 ) | ( n9286 & 1'b0 ) | ( ~n22080 & 1'b0 ) ;
  assign n22082 = n8839 | n22081 ;
  assign n22083 = ( n22078 & ~n22082 ) | ( n22078 & 1'b0 ) | ( ~n22082 & 1'b0 ) ;
  assign n22084 = n22075 | n22083 ;
  assign n22063 = n22048 &  n22062 ;
  assign n22069 = ( n22063 & ~n9286 ) | ( n22063 & n22068 ) | ( ~n9286 & n22068 ) ;
  assign n22070 = ( n8839 & ~n22069 ) | ( n8839 & 1'b0 ) | ( ~n22069 & 1'b0 ) ;
  assign n22098 = n8407 | n22070 ;
  assign n22099 = ( n22084 & ~n22098 ) | ( n22084 & 1'b0 ) | ( ~n22098 & 1'b0 ) ;
  assign n22100 = n22090 | n22099 ;
  assign n22101 = ( n22078 & ~n22081 ) | ( n22078 & 1'b0 ) | ( ~n22081 & 1'b0 ) ;
  assign n22102 = ( n22075 & ~n8839 ) | ( n22075 & n22101 ) | ( ~n8839 & n22101 ) ;
  assign n22103 = ( n8407 & ~n22102 ) | ( n8407 & 1'b0 ) | ( ~n22102 & 1'b0 ) ;
  assign n22104 = n7982 | n22103 ;
  assign n22105 = ( n22100 & ~n22104 ) | ( n22100 & 1'b0 ) | ( ~n22104 & 1'b0 ) ;
  assign n22106 = n22097 | n22105 ;
  assign n22085 = ~n22070 & n22084 ;
  assign n22091 = ( n22085 & ~n8407 ) | ( n22085 & n22090 ) | ( ~n8407 & n22090 ) ;
  assign n22092 = ( n7982 & ~n22091 ) | ( n7982 & 1'b0 ) | ( ~n22091 & 1'b0 ) ;
  assign n22120 = ( n7572 & ~n22092 ) | ( n7572 & 1'b0 ) | ( ~n22092 & 1'b0 ) ;
  assign n22121 = n22106 &  n22120 ;
  assign n22122 = n22112 | n22121 ;
  assign n22123 = ( n22100 & ~n22103 ) | ( n22100 & 1'b0 ) | ( ~n22103 & 1'b0 ) ;
  assign n22124 = ( n22097 & ~n7982 ) | ( n22097 & n22123 ) | ( ~n7982 & n22123 ) ;
  assign n22125 = n7572 | n22124 ;
  assign n22126 = n7169 &  n22125 ;
  assign n22127 = n22122 &  n22126 ;
  assign n22128 = n22119 | n22127 ;
  assign n22107 = ~n22092 & n22106 ;
  assign n22113 = ( n7572 & n22107 ) | ( n7572 & n22112 ) | ( n22107 & n22112 ) ;
  assign n22114 = n7169 | n22113 ;
  assign n22142 = ~n6781 & n22114 ;
  assign n22143 = n22128 &  n22142 ;
  assign n22144 = n22134 | n22143 ;
  assign n22145 = n22122 &  n22125 ;
  assign n22146 = ( n7169 & n22119 ) | ( n7169 & n22145 ) | ( n22119 & n22145 ) ;
  assign n22147 = ( n6781 & ~n22146 ) | ( n6781 & 1'b0 ) | ( ~n22146 & 1'b0 ) ;
  assign n22148 = ( n6399 & ~n22147 ) | ( n6399 & 1'b0 ) | ( ~n22147 & 1'b0 ) ;
  assign n22149 = n22144 &  n22148 ;
  assign n22150 = n22141 | n22149 ;
  assign n22129 = n22114 &  n22128 ;
  assign n22135 = ( n22129 & ~n6781 ) | ( n22129 & n22134 ) | ( ~n6781 & n22134 ) ;
  assign n22136 = n6399 | n22135 ;
  assign n22164 = ~n6032 & n22136 ;
  assign n22165 = n22150 &  n22164 ;
  assign n22166 = n22156 | n22165 ;
  assign n22167 = ( n22144 & ~n22147 ) | ( n22144 & 1'b0 ) | ( ~n22147 & 1'b0 ) ;
  assign n22168 = ( n6399 & n22141 ) | ( n6399 & n22167 ) | ( n22141 & n22167 ) ;
  assign n22169 = ( n6032 & ~n22168 ) | ( n6032 & 1'b0 ) | ( ~n22168 & 1'b0 ) ;
  assign n22170 = ( n5672 & ~n22169 ) | ( n5672 & 1'b0 ) | ( ~n22169 & 1'b0 ) ;
  assign n22171 = n22166 &  n22170 ;
  assign n22172 = n22163 | n22171 ;
  assign n22151 = n22136 &  n22150 ;
  assign n22157 = ( n22151 & ~n6032 ) | ( n22151 & n22156 ) | ( ~n6032 & n22156 ) ;
  assign n22158 = n5672 | n22157 ;
  assign n22186 = ~n5327 & n22158 ;
  assign n22187 = n22172 &  n22186 ;
  assign n22188 = n22178 | n22187 ;
  assign n22189 = ( n22166 & ~n22169 ) | ( n22166 & 1'b0 ) | ( ~n22169 & 1'b0 ) ;
  assign n22190 = ( n5672 & n22163 ) | ( n5672 & n22189 ) | ( n22163 & n22189 ) ;
  assign n22191 = ( n5327 & ~n22190 ) | ( n5327 & 1'b0 ) | ( ~n22190 & 1'b0 ) ;
  assign n22192 = n4990 | n22191 ;
  assign n22193 = ( n22188 & ~n22192 ) | ( n22188 & 1'b0 ) | ( ~n22192 & 1'b0 ) ;
  assign n22194 = n22185 | n22193 ;
  assign n22173 = n22158 &  n22172 ;
  assign n22179 = ( n22173 & ~n5327 ) | ( n22173 & n22178 ) | ( ~n5327 & n22178 ) ;
  assign n22180 = ( n4990 & ~n22179 ) | ( n4990 & 1'b0 ) | ( ~n22179 & 1'b0 ) ;
  assign n22208 = n4668 | n22180 ;
  assign n22209 = ( n22194 & ~n22208 ) | ( n22194 & 1'b0 ) | ( ~n22208 & 1'b0 ) ;
  assign n22210 = n22200 | n22209 ;
  assign n22211 = ( n22188 & ~n22191 ) | ( n22188 & 1'b0 ) | ( ~n22191 & 1'b0 ) ;
  assign n22212 = ( n22185 & ~n4990 ) | ( n22185 & n22211 ) | ( ~n4990 & n22211 ) ;
  assign n22213 = ( n4668 & ~n22212 ) | ( n4668 & 1'b0 ) | ( ~n22212 & 1'b0 ) ;
  assign n22214 = n4353 | n22213 ;
  assign n22215 = ( n22210 & ~n22214 ) | ( n22210 & 1'b0 ) | ( ~n22214 & 1'b0 ) ;
  assign n22216 = n22207 | n22215 ;
  assign n22195 = ~n22180 & n22194 ;
  assign n22201 = ( n22195 & ~n4668 ) | ( n22195 & n22200 ) | ( ~n4668 & n22200 ) ;
  assign n22202 = ( n4353 & ~n22201 ) | ( n4353 & 1'b0 ) | ( ~n22201 & 1'b0 ) ;
  assign n22230 = n4053 | n22202 ;
  assign n22231 = ( n22216 & ~n22230 ) | ( n22216 & 1'b0 ) | ( ~n22230 & 1'b0 ) ;
  assign n22232 = n22222 | n22231 ;
  assign n22233 = ( n22210 & ~n22213 ) | ( n22210 & 1'b0 ) | ( ~n22213 & 1'b0 ) ;
  assign n22234 = ( n22207 & ~n4353 ) | ( n22207 & n22233 ) | ( ~n4353 & n22233 ) ;
  assign n22235 = ( n4053 & ~n22234 ) | ( n4053 & 1'b0 ) | ( ~n22234 & 1'b0 ) ;
  assign n22236 = n3760 | n22235 ;
  assign n22237 = ( n22232 & ~n22236 ) | ( n22232 & 1'b0 ) | ( ~n22236 & 1'b0 ) ;
  assign n22238 = n22229 | n22237 ;
  assign n22217 = ~n22202 & n22216 ;
  assign n22223 = ( n22217 & ~n4053 ) | ( n22217 & n22222 ) | ( ~n4053 & n22222 ) ;
  assign n22224 = ( n3760 & ~n22223 ) | ( n3760 & 1'b0 ) | ( ~n22223 & 1'b0 ) ;
  assign n22252 = n3482 | n22224 ;
  assign n22253 = ( n22238 & ~n22252 ) | ( n22238 & 1'b0 ) | ( ~n22252 & 1'b0 ) ;
  assign n22254 = n22244 | n22253 ;
  assign n22255 = ( n22232 & ~n22235 ) | ( n22232 & 1'b0 ) | ( ~n22235 & 1'b0 ) ;
  assign n22256 = ( n22229 & ~n3760 ) | ( n22229 & n22255 ) | ( ~n3760 & n22255 ) ;
  assign n22257 = ( n3482 & ~n22256 ) | ( n3482 & 1'b0 ) | ( ~n22256 & 1'b0 ) ;
  assign n22258 = n3211 | n22257 ;
  assign n22259 = ( n22254 & ~n22258 ) | ( n22254 & 1'b0 ) | ( ~n22258 & 1'b0 ) ;
  assign n22260 = n22251 | n22259 ;
  assign n22239 = ~n22224 & n22238 ;
  assign n22245 = ( n22239 & ~n3482 ) | ( n22239 & n22244 ) | ( ~n3482 & n22244 ) ;
  assign n22246 = ( n3211 & ~n22245 ) | ( n3211 & 1'b0 ) | ( ~n22245 & 1'b0 ) ;
  assign n22274 = n2955 | n22246 ;
  assign n22275 = ( n22260 & ~n22274 ) | ( n22260 & 1'b0 ) | ( ~n22274 & 1'b0 ) ;
  assign n22276 = n22266 | n22275 ;
  assign n22277 = ( n22254 & ~n22257 ) | ( n22254 & 1'b0 ) | ( ~n22257 & 1'b0 ) ;
  assign n22278 = ( n22251 & ~n3211 ) | ( n22251 & n22277 ) | ( ~n3211 & n22277 ) ;
  assign n22279 = ( n2955 & ~n22278 ) | ( n2955 & 1'b0 ) | ( ~n22278 & 1'b0 ) ;
  assign n22280 = n2706 | n22279 ;
  assign n22281 = ( n22276 & ~n22280 ) | ( n22276 & 1'b0 ) | ( ~n22280 & 1'b0 ) ;
  assign n22282 = n22273 | n22281 ;
  assign n22261 = ~n22246 & n22260 ;
  assign n22267 = ( n22261 & ~n2955 ) | ( n22261 & n22266 ) | ( ~n2955 & n22266 ) ;
  assign n22268 = ( n2706 & ~n22267 ) | ( n2706 & 1'b0 ) | ( ~n22267 & 1'b0 ) ;
  assign n22296 = n2472 | n22268 ;
  assign n22297 = ( n22282 & ~n22296 ) | ( n22282 & 1'b0 ) | ( ~n22296 & 1'b0 ) ;
  assign n22298 = n22288 | n22297 ;
  assign n22299 = ( n22276 & ~n22279 ) | ( n22276 & 1'b0 ) | ( ~n22279 & 1'b0 ) ;
  assign n22300 = ( n22273 & ~n2706 ) | ( n22273 & n22299 ) | ( ~n2706 & n22299 ) ;
  assign n22301 = ( n2472 & ~n22300 ) | ( n2472 & 1'b0 ) | ( ~n22300 & 1'b0 ) ;
  assign n22302 = n2245 | n22301 ;
  assign n22303 = ( n22298 & ~n22302 ) | ( n22298 & 1'b0 ) | ( ~n22302 & 1'b0 ) ;
  assign n22304 = ( n22295 & ~n22303 ) | ( n22295 & 1'b0 ) | ( ~n22303 & 1'b0 ) ;
  assign n22283 = ~n22268 & n22282 ;
  assign n22289 = ( n22283 & ~n2472 ) | ( n22283 & n22288 ) | ( ~n2472 & n22288 ) ;
  assign n22290 = ( n2245 & ~n22289 ) | ( n2245 & 1'b0 ) | ( ~n22289 & 1'b0 ) ;
  assign n22318 = ( n2033 & ~n22290 ) | ( n2033 & 1'b0 ) | ( ~n22290 & 1'b0 ) ;
  assign n22319 = ~n22304 & n22318 ;
  assign n22320 = ( n22310 & ~n22319 ) | ( n22310 & 1'b0 ) | ( ~n22319 & 1'b0 ) ;
  assign n22321 = ( n22298 & ~n22301 ) | ( n22298 & 1'b0 ) | ( ~n22301 & 1'b0 ) ;
  assign n22322 = ( n2245 & ~n22321 ) | ( n2245 & n22295 ) | ( ~n22321 & n22295 ) ;
  assign n22323 = ~n2033 & n22322 ;
  assign n22324 = n1827 | n22323 ;
  assign n22325 = n22320 | n22324 ;
  assign n22326 = n22317 &  n22325 ;
  assign n22305 = n22290 | n22304 ;
  assign n22311 = ( n22305 & ~n2033 ) | ( n22305 & n22310 ) | ( ~n2033 & n22310 ) ;
  assign n22312 = n1827 &  n22311 ;
  assign n22340 = ( n1636 & ~n22312 ) | ( n1636 & 1'b0 ) | ( ~n22312 & 1'b0 ) ;
  assign n22341 = ~n22326 & n22340 ;
  assign n22342 = ( n22332 & ~n22341 ) | ( n22332 & 1'b0 ) | ( ~n22341 & 1'b0 ) ;
  assign n22343 = n22320 | n22323 ;
  assign n22344 = ( n1827 & n22317 ) | ( n1827 & n22343 ) | ( n22317 & n22343 ) ;
  assign n22345 = ~n1636 & n22344 ;
  assign n22346 = ( n1452 & ~n22345 ) | ( n1452 & 1'b0 ) | ( ~n22345 & 1'b0 ) ;
  assign n22347 = ~n22342 & n22346 ;
  assign n22348 = ( n22339 & ~n22347 ) | ( n22339 & 1'b0 ) | ( ~n22347 & 1'b0 ) ;
  assign n22327 = n22312 | n22326 ;
  assign n22333 = ( n22327 & ~n1636 ) | ( n22327 & n22332 ) | ( ~n1636 & n22332 ) ;
  assign n22334 = ~n1452 & n22333 ;
  assign n22362 = n1283 | n22334 ;
  assign n22363 = n22348 | n22362 ;
  assign n22364 = ~n22354 & n22363 ;
  assign n22365 = n22342 | n22345 ;
  assign n22366 = ( n22339 & ~n1452 ) | ( n22339 & n22365 ) | ( ~n1452 & n22365 ) ;
  assign n22367 = n1283 &  n22366 ;
  assign n22368 = ( n1122 & ~n22367 ) | ( n1122 & 1'b0 ) | ( ~n22367 & 1'b0 ) ;
  assign n22369 = ~n22364 & n22368 ;
  assign n22370 = n22361 | n22369 ;
  assign n22349 = n22334 | n22348 ;
  assign n22355 = ( n1283 & ~n22354 ) | ( n1283 & n22349 ) | ( ~n22354 & n22349 ) ;
  assign n22356 = ~n1122 & n22355 ;
  assign n22384 = ( n976 & ~n22356 ) | ( n976 & 1'b0 ) | ( ~n22356 & 1'b0 ) ;
  assign n22385 = n22370 &  n22384 ;
  assign n22386 = ( n22376 & ~n22385 ) | ( n22376 & 1'b0 ) | ( ~n22385 & 1'b0 ) ;
  assign n22387 = n22364 | n22367 ;
  assign n22388 = ( n1122 & ~n22387 ) | ( n1122 & n22361 ) | ( ~n22387 & n22361 ) ;
  assign n22389 = n976 | n22388 ;
  assign n22390 = ~n837 & n22389 ;
  assign n22391 = ~n22386 & n22390 ;
  assign n22392 = n22383 | n22391 ;
  assign n22371 = ~n22356 & n22370 ;
  assign n22377 = ( n976 & ~n22376 ) | ( n976 & n22371 ) | ( ~n22376 & n22371 ) ;
  assign n22378 = ( n837 & ~n22377 ) | ( n837 & 1'b0 ) | ( ~n22377 & 1'b0 ) ;
  assign n22406 = n713 | n22378 ;
  assign n22407 = ( n22392 & ~n22406 ) | ( n22392 & 1'b0 ) | ( ~n22406 & 1'b0 ) ;
  assign n22408 = ( n22398 & ~n22407 ) | ( n22398 & 1'b0 ) | ( ~n22407 & 1'b0 ) ;
  assign n22409 = ~n22386 & n22389 ;
  assign n22410 = ( n22383 & ~n837 ) | ( n22383 & n22409 ) | ( ~n837 & n22409 ) ;
  assign n22411 = ( n713 & ~n22410 ) | ( n713 & 1'b0 ) | ( ~n22410 & 1'b0 ) ;
  assign n22412 = n595 | n22411 ;
  assign n22413 = n22408 | n22412 ;
  assign n22414 = n22405 &  n22413 ;
  assign n22393 = ~n22378 & n22392 ;
  assign n22399 = ( n713 & ~n22393 ) | ( n713 & n22398 ) | ( ~n22393 & n22398 ) ;
  assign n22400 = n595 &  n22399 ;
  assign n22428 = n492 | n22400 ;
  assign n22429 = n22414 | n22428 ;
  assign n22430 = ~n22420 & n22429 ;
  assign n22431 = n22408 | n22411 ;
  assign n22432 = ( n595 & n22405 ) | ( n595 & n22431 ) | ( n22405 & n22431 ) ;
  assign n22433 = n492 &  n22432 ;
  assign n22434 = n396 | n22433 ;
  assign n22435 = n22430 | n22434 ;
  assign n22436 = ~n22427 & n22435 ;
  assign n22415 = n22400 | n22414 ;
  assign n22421 = ( n492 & ~n22420 ) | ( n492 & n22415 ) | ( ~n22420 & n22415 ) ;
  assign n22422 = n396 &  n22421 ;
  assign n22450 = n315 | n22422 ;
  assign n22451 = n22436 | n22450 ;
  assign n22452 = ~n22442 & n22451 ;
  assign n22453 = n22430 | n22433 ;
  assign n22454 = ( n396 & ~n22427 ) | ( n396 & n22453 ) | ( ~n22427 & n22453 ) ;
  assign n22455 = n315 &  n22454 ;
  assign n22456 = n240 | n22455 ;
  assign n22457 = n22452 | n22456 ;
  assign n22458 = ~n22449 & n22457 ;
  assign n22437 = n22422 | n22436 ;
  assign n22443 = ( n315 & ~n22442 ) | ( n315 & n22437 ) | ( ~n22442 & n22437 ) ;
  assign n22444 = n240 &  n22443 ;
  assign n22472 = n181 | n22444 ;
  assign n22473 = n22458 | n22472 ;
  assign n22474 = ~n22464 & n22473 ;
  assign n22475 = n22452 | n22455 ;
  assign n22476 = ( n240 & ~n22449 ) | ( n240 & n22475 ) | ( ~n22449 & n22475 ) ;
  assign n22477 = n181 &  n22476 ;
  assign n22500 = n22474 | n22477 ;
  assign n22501 = ( n22471 & ~n145 ) | ( n22471 & n22500 ) | ( ~n145 & n22500 ) ;
  assign n22502 = n150 &  n22501 ;
  assign n22478 = ( n145 & ~n22477 ) | ( n145 & 1'b0 ) | ( ~n22477 & 1'b0 ) ;
  assign n22479 = ~n22474 & n22478 ;
  assign n22480 = ( n22471 & ~n22479 ) | ( n22471 & 1'b0 ) | ( ~n22479 & 1'b0 ) ;
  assign n22459 = n22444 | n22458 ;
  assign n22465 = ( n181 & ~n22464 ) | ( n181 & n22459 ) | ( ~n22464 & n22459 ) ;
  assign n22466 = ~n145 & n22465 ;
  assign n22498 = n150 | n22466 ;
  assign n22499 = n22480 | n22498 ;
  assign n23183 = ( n22499 & ~n22486 ) | ( n22499 & n22502 ) | ( ~n22486 & n22502 ) ;
  assign n22488 = ( n21792 & ~n21809 ) | ( n21792 & n21806 ) | ( ~n21809 & n21806 ) ;
  assign n22489 = ( n21809 & n21818 ) | ( n21809 & n22488 ) | ( n21818 & n22488 ) ;
  assign n22490 = ( n21806 & ~n22488 ) | ( n21806 & n21818 ) | ( ~n22488 & n21818 ) ;
  assign n22491 = ( n21792 & ~n22489 ) | ( n21792 & n22490 ) | ( ~n22489 & n22490 ) ;
  assign n22492 = ~n21793 & n21798 ;
  assign n22493 = ~n21818 & n22492 ;
  assign n22494 = ( n21812 & ~n22493 ) | ( n21812 & n22492 ) | ( ~n22493 & n22492 ) ;
  assign n22495 = n22491 | n22494 ;
  assign n22481 = n22466 | n22480 ;
  assign n22487 = ( n150 & ~n22486 ) | ( n150 & n22481 ) | ( ~n22486 & n22481 ) ;
  assign n22496 = n22487 | n22495 ;
  assign n22497 = ( n133 & ~n22495 ) | ( n133 & n22496 ) | ( ~n22495 & n22496 ) ;
  assign n22504 = n22486 | n22499 ;
  assign n22503 = ( n22491 & ~n22502 ) | ( n22491 & 1'b0 ) | ( ~n22502 & 1'b0 ) ;
  assign n22505 = ( n22486 & ~n22504 ) | ( n22486 & n22503 ) | ( ~n22504 & n22503 ) ;
  assign n22507 = ( n133 & ~n21793 ) | ( n133 & n21798 ) | ( ~n21793 & n21798 ) ;
  assign n22506 = ( n21793 & ~n21798 ) | ( n21793 & n21818 ) | ( ~n21798 & n21818 ) ;
  assign n22508 = n21798 &  n22506 ;
  assign n22509 = ( n22507 & ~n21798 ) | ( n22507 & n22508 ) | ( ~n21798 & n22508 ) ;
  assign n22510 = n22505 | n22509 ;
  assign n22511 = ~n22497 |  n22510 ;
  assign n23182 = n22502 | n22511 ;
  assign n23185 = ( n22502 & ~n23183 ) | ( n22502 & n23182 ) | ( ~n23183 & n23182 ) ;
  assign n23184 = ( n23182 & ~n22499 ) | ( n23182 & n23183 ) | ( ~n22499 & n23183 ) ;
  assign n23186 = ( n22486 & ~n23185 ) | ( n22486 & n23184 ) | ( ~n23185 & n23184 ) ;
  assign n23145 = ~n22457 & n22511 ;
  assign n23146 = ( n22444 & ~n23145 ) | ( n22444 & n22511 ) | ( ~n23145 & n22511 ) ;
  assign n23147 = ( n22449 & ~n22444 ) | ( n22449 & n23146 ) | ( ~n22444 & n23146 ) ;
  assign n23148 = ( n22444 & ~n23146 ) | ( n22444 & n22449 ) | ( ~n23146 & n22449 ) ;
  assign n23149 = ( n23147 & ~n22449 ) | ( n23147 & n23148 ) | ( ~n22449 & n23148 ) ;
  assign n23136 = n22455 | n22511 ;
  assign n23137 = ( n22442 & n22451 ) | ( n22442 & n22455 ) | ( n22451 & n22455 ) ;
  assign n23138 = ( n23136 & ~n22451 ) | ( n23136 & n23137 ) | ( ~n22451 & n23137 ) ;
  assign n23139 = ( n22455 & ~n23137 ) | ( n22455 & n23136 ) | ( ~n23137 & n23136 ) ;
  assign n23140 = ( n22442 & ~n23138 ) | ( n22442 & n23139 ) | ( ~n23138 & n23139 ) ;
  assign n23122 = ~n22435 & n22511 ;
  assign n23123 = ( n22422 & ~n23122 ) | ( n22422 & n22511 ) | ( ~n23122 & n22511 ) ;
  assign n23124 = ( n22427 & ~n22422 ) | ( n22427 & n23123 ) | ( ~n22422 & n23123 ) ;
  assign n23125 = ( n22422 & ~n23123 ) | ( n22422 & n22427 ) | ( ~n23123 & n22427 ) ;
  assign n23126 = ( n23124 & ~n22427 ) | ( n23124 & n23125 ) | ( ~n22427 & n23125 ) ;
  assign n23113 = n22433 | n22511 ;
  assign n23114 = ( n22420 & n22429 ) | ( n22420 & n22433 ) | ( n22429 & n22433 ) ;
  assign n23115 = ( n23113 & ~n22429 ) | ( n23113 & n23114 ) | ( ~n22429 & n23114 ) ;
  assign n23116 = ( n22433 & ~n23114 ) | ( n22433 & n23113 ) | ( ~n23114 & n23113 ) ;
  assign n23117 = ( n22420 & ~n23115 ) | ( n22420 & n23116 ) | ( ~n23115 & n23116 ) ;
  assign n23099 = ~n22413 & n22511 ;
  assign n23100 = ( n22400 & ~n23099 ) | ( n22400 & n22511 ) | ( ~n23099 & n22511 ) ;
  assign n23101 = ( n22400 & ~n23100 ) | ( n22400 & n22405 ) | ( ~n23100 & n22405 ) ;
  assign n23102 = ( n22405 & ~n22400 ) | ( n22405 & n23100 ) | ( ~n22400 & n23100 ) ;
  assign n23103 = ( n23101 & ~n22405 ) | ( n23101 & n23102 ) | ( ~n22405 & n23102 ) ;
  assign n23090 = n22411 | n22511 ;
  assign n23091 = ( n22398 & ~n22411 ) | ( n22398 & n22407 ) | ( ~n22411 & n22407 ) ;
  assign n23093 = ( n22411 & n23090 ) | ( n22411 & n23091 ) | ( n23090 & n23091 ) ;
  assign n23092 = ( n22407 & ~n23091 ) | ( n22407 & n23090 ) | ( ~n23091 & n23090 ) ;
  assign n23094 = ( n22398 & ~n23093 ) | ( n22398 & n23092 ) | ( ~n23093 & n23092 ) ;
  assign n23076 = n22391 &  n22511 ;
  assign n23077 = ( n22378 & ~n23076 ) | ( n22378 & n22511 ) | ( ~n23076 & n22511 ) ;
  assign n23078 = ( n22383 & ~n22378 ) | ( n22383 & n23077 ) | ( ~n22378 & n23077 ) ;
  assign n23079 = ( n22378 & ~n23077 ) | ( n22378 & n22383 ) | ( ~n23077 & n22383 ) ;
  assign n23080 = ( n23078 & ~n22383 ) | ( n23078 & n23079 ) | ( ~n22383 & n23079 ) ;
  assign n23053 = n22369 &  n22511 ;
  assign n23054 = ( n22356 & ~n23053 ) | ( n22356 & n22511 ) | ( ~n23053 & n22511 ) ;
  assign n23055 = ( n22361 & ~n22356 ) | ( n22361 & n23054 ) | ( ~n22356 & n23054 ) ;
  assign n23056 = ( n22356 & ~n23054 ) | ( n22356 & n22361 ) | ( ~n23054 & n22361 ) ;
  assign n23057 = ( n23055 & ~n22361 ) | ( n23055 & n23056 ) | ( ~n22361 & n23056 ) ;
  assign n23030 = n22347 &  n22511 ;
  assign n23031 = ( n22334 & ~n23030 ) | ( n22334 & n22511 ) | ( ~n23030 & n22511 ) ;
  assign n23032 = ( n22334 & ~n23031 ) | ( n22334 & n22339 ) | ( ~n23031 & n22339 ) ;
  assign n23033 = ( n22339 & ~n22334 ) | ( n22339 & n23031 ) | ( ~n22334 & n23031 ) ;
  assign n23034 = ( n23032 & ~n22339 ) | ( n23032 & n23033 ) | ( ~n22339 & n23033 ) ;
  assign n23021 = n22345 | n22511 ;
  assign n23022 = ( n22332 & ~n22345 ) | ( n22332 & n22341 ) | ( ~n22345 & n22341 ) ;
  assign n23024 = ( n22345 & n23021 ) | ( n22345 & n23022 ) | ( n23021 & n23022 ) ;
  assign n23023 = ( n22341 & ~n23022 ) | ( n22341 & n23021 ) | ( ~n23022 & n23021 ) ;
  assign n23025 = ( n22332 & ~n23024 ) | ( n22332 & n23023 ) | ( ~n23024 & n23023 ) ;
  assign n23007 = ~n22325 & n22511 ;
  assign n23008 = ( n22312 & n22317 ) | ( n22312 & n22511 ) | ( n22317 & n22511 ) ;
  assign n23010 = ( n23007 & ~n22312 ) | ( n23007 & n23008 ) | ( ~n22312 & n23008 ) ;
  assign n23009 = ( n22511 & ~n23008 ) | ( n22511 & n23007 ) | ( ~n23008 & n23007 ) ;
  assign n23011 = ( n22317 & ~n23010 ) | ( n22317 & n23009 ) | ( ~n23010 & n23009 ) ;
  assign n22984 = n22303 &  n22511 ;
  assign n22985 = ( n22290 & ~n22984 ) | ( n22290 & n22511 ) | ( ~n22984 & n22511 ) ;
  assign n22986 = ( n22290 & ~n22985 ) | ( n22290 & n22295 ) | ( ~n22985 & n22295 ) ;
  assign n22987 = ( n22295 & ~n22290 ) | ( n22295 & n22985 ) | ( ~n22290 & n22985 ) ;
  assign n22988 = ( n22986 & ~n22295 ) | ( n22986 & n22987 ) | ( ~n22295 & n22987 ) ;
  assign n22975 = n22301 | n22511 ;
  assign n22976 = ( n22288 & ~n22297 ) | ( n22288 & n22301 ) | ( ~n22297 & n22301 ) ;
  assign n22977 = ( n22297 & n22975 ) | ( n22297 & n22976 ) | ( n22975 & n22976 ) ;
  assign n22978 = ( n22301 & ~n22976 ) | ( n22301 & n22975 ) | ( ~n22976 & n22975 ) ;
  assign n22979 = ( n22288 & ~n22977 ) | ( n22288 & n22978 ) | ( ~n22977 & n22978 ) ;
  assign n22961 = n22281 &  n22511 ;
  assign n22962 = ( n22268 & ~n22961 ) | ( n22268 & n22511 ) | ( ~n22961 & n22511 ) ;
  assign n22963 = ( n22273 & ~n22268 ) | ( n22273 & n22962 ) | ( ~n22268 & n22962 ) ;
  assign n22964 = ( n22268 & ~n22962 ) | ( n22268 & n22273 ) | ( ~n22962 & n22273 ) ;
  assign n22965 = ( n22963 & ~n22273 ) | ( n22963 & n22964 ) | ( ~n22273 & n22964 ) ;
  assign n22952 = n22279 | n22511 ;
  assign n22953 = ( n22266 & ~n22275 ) | ( n22266 & n22279 ) | ( ~n22275 & n22279 ) ;
  assign n22954 = ( n22275 & n22952 ) | ( n22275 & n22953 ) | ( n22952 & n22953 ) ;
  assign n22955 = ( n22279 & ~n22953 ) | ( n22279 & n22952 ) | ( ~n22953 & n22952 ) ;
  assign n22956 = ( n22266 & ~n22954 ) | ( n22266 & n22955 ) | ( ~n22954 & n22955 ) ;
  assign n22938 = n22259 &  n22511 ;
  assign n22939 = ( n22246 & n22251 ) | ( n22246 & n22511 ) | ( n22251 & n22511 ) ;
  assign n22941 = ( n22938 & ~n22246 ) | ( n22938 & n22939 ) | ( ~n22246 & n22939 ) ;
  assign n22940 = ( n22511 & ~n22939 ) | ( n22511 & n22938 ) | ( ~n22939 & n22938 ) ;
  assign n22942 = ( n22251 & ~n22941 ) | ( n22251 & n22940 ) | ( ~n22941 & n22940 ) ;
  assign n22929 = n22257 | n22511 ;
  assign n22930 = ( n22244 & ~n22253 ) | ( n22244 & n22257 ) | ( ~n22253 & n22257 ) ;
  assign n22931 = ( n22253 & n22929 ) | ( n22253 & n22930 ) | ( n22929 & n22930 ) ;
  assign n22932 = ( n22257 & ~n22930 ) | ( n22257 & n22929 ) | ( ~n22930 & n22929 ) ;
  assign n22933 = ( n22244 & ~n22931 ) | ( n22244 & n22932 ) | ( ~n22931 & n22932 ) ;
  assign n22915 = n22237 &  n22511 ;
  assign n22916 = ( n22224 & ~n22915 ) | ( n22224 & n22511 ) | ( ~n22915 & n22511 ) ;
  assign n22917 = ( n22229 & ~n22224 ) | ( n22229 & n22916 ) | ( ~n22224 & n22916 ) ;
  assign n22918 = ( n22224 & ~n22916 ) | ( n22224 & n22229 ) | ( ~n22916 & n22229 ) ;
  assign n22919 = ( n22917 & ~n22229 ) | ( n22917 & n22918 ) | ( ~n22229 & n22918 ) ;
  assign n22906 = n22235 | n22511 ;
  assign n22907 = ( n22222 & ~n22231 ) | ( n22222 & n22235 ) | ( ~n22231 & n22235 ) ;
  assign n22908 = ( n22231 & n22906 ) | ( n22231 & n22907 ) | ( n22906 & n22907 ) ;
  assign n22909 = ( n22235 & ~n22907 ) | ( n22235 & n22906 ) | ( ~n22907 & n22906 ) ;
  assign n22910 = ( n22222 & ~n22908 ) | ( n22222 & n22909 ) | ( ~n22908 & n22909 ) ;
  assign n22892 = n22215 &  n22511 ;
  assign n22893 = ( n22202 & ~n22892 ) | ( n22202 & n22511 ) | ( ~n22892 & n22511 ) ;
  assign n22894 = ( n22207 & ~n22202 ) | ( n22207 & n22893 ) | ( ~n22202 & n22893 ) ;
  assign n22895 = ( n22202 & ~n22893 ) | ( n22202 & n22207 ) | ( ~n22893 & n22207 ) ;
  assign n22896 = ( n22894 & ~n22207 ) | ( n22894 & n22895 ) | ( ~n22207 & n22895 ) ;
  assign n22883 = n22213 | n22511 ;
  assign n22884 = ( n22200 & ~n22209 ) | ( n22200 & n22213 ) | ( ~n22209 & n22213 ) ;
  assign n22885 = ( n22209 & n22883 ) | ( n22209 & n22884 ) | ( n22883 & n22884 ) ;
  assign n22886 = ( n22213 & ~n22884 ) | ( n22213 & n22883 ) | ( ~n22884 & n22883 ) ;
  assign n22887 = ( n22200 & ~n22885 ) | ( n22200 & n22886 ) | ( ~n22885 & n22886 ) ;
  assign n22869 = n22193 &  n22511 ;
  assign n22870 = ( n22180 & ~n22869 ) | ( n22180 & n22511 ) | ( ~n22869 & n22511 ) ;
  assign n22871 = ( n22185 & ~n22180 ) | ( n22185 & n22870 ) | ( ~n22180 & n22870 ) ;
  assign n22872 = ( n22180 & ~n22870 ) | ( n22180 & n22185 ) | ( ~n22870 & n22185 ) ;
  assign n22873 = ( n22871 & ~n22185 ) | ( n22871 & n22872 ) | ( ~n22185 & n22872 ) ;
  assign n22860 = n22191 | n22511 ;
  assign n22861 = ( n22178 & ~n22187 ) | ( n22178 & n22191 ) | ( ~n22187 & n22191 ) ;
  assign n22862 = ( n22187 & n22860 ) | ( n22187 & n22861 ) | ( n22860 & n22861 ) ;
  assign n22863 = ( n22191 & ~n22861 ) | ( n22191 & n22860 ) | ( ~n22861 & n22860 ) ;
  assign n22864 = ( n22178 & ~n22862 ) | ( n22178 & n22863 ) | ( ~n22862 & n22863 ) ;
  assign n22846 = n22171 &  n22511 ;
  assign n22847 = ( n22158 & ~n22511 ) | ( n22158 & n22163 ) | ( ~n22511 & n22163 ) ;
  assign n22848 = ( n22511 & n22846 ) | ( n22511 & n22847 ) | ( n22846 & n22847 ) ;
  assign n22849 = ( n22158 & ~n22847 ) | ( n22158 & n22846 ) | ( ~n22847 & n22846 ) ;
  assign n22850 = ( n22163 & ~n22848 ) | ( n22163 & n22849 ) | ( ~n22848 & n22849 ) ;
  assign n22837 = n22169 | n22511 ;
  assign n22838 = ( n22156 & ~n22165 ) | ( n22156 & n22169 ) | ( ~n22165 & n22169 ) ;
  assign n22839 = ( n22165 & n22837 ) | ( n22165 & n22838 ) | ( n22837 & n22838 ) ;
  assign n22840 = ( n22169 & ~n22838 ) | ( n22169 & n22837 ) | ( ~n22838 & n22837 ) ;
  assign n22841 = ( n22156 & ~n22839 ) | ( n22156 & n22840 ) | ( ~n22839 & n22840 ) ;
  assign n22823 = n22149 &  n22511 ;
  assign n22824 = ( n22136 & ~n22511 ) | ( n22136 & n22823 ) | ( ~n22511 & n22823 ) ;
  assign n22825 = ( n22136 & ~n22824 ) | ( n22136 & n22141 ) | ( ~n22824 & n22141 ) ;
  assign n22826 = ( n22141 & ~n22136 ) | ( n22141 & n22824 ) | ( ~n22136 & n22824 ) ;
  assign n22827 = ( n22825 & ~n22141 ) | ( n22825 & n22826 ) | ( ~n22141 & n22826 ) ;
  assign n22814 = n22147 | n22511 ;
  assign n22815 = ( n22134 & ~n22143 ) | ( n22134 & n22147 ) | ( ~n22143 & n22147 ) ;
  assign n22816 = ( n22143 & n22814 ) | ( n22143 & n22815 ) | ( n22814 & n22815 ) ;
  assign n22817 = ( n22147 & ~n22815 ) | ( n22147 & n22814 ) | ( ~n22815 & n22814 ) ;
  assign n22818 = ( n22134 & ~n22816 ) | ( n22134 & n22817 ) | ( ~n22816 & n22817 ) ;
  assign n22800 = n22127 &  n22511 ;
  assign n22801 = ( n22114 & ~n22511 ) | ( n22114 & n22800 ) | ( ~n22511 & n22800 ) ;
  assign n22802 = ( n22114 & ~n22801 ) | ( n22114 & n22119 ) | ( ~n22801 & n22119 ) ;
  assign n22803 = ( n22119 & ~n22114 ) | ( n22119 & n22801 ) | ( ~n22114 & n22801 ) ;
  assign n22804 = ( n22802 & ~n22119 ) | ( n22802 & n22803 ) | ( ~n22119 & n22803 ) ;
  assign n22792 = ( n22121 & ~n22112 ) | ( n22121 & n22125 ) | ( ~n22112 & n22125 ) ;
  assign n22791 = ( n22125 & ~n22511 ) | ( n22125 & 1'b0 ) | ( ~n22511 & 1'b0 ) ;
  assign n22794 = ( n22125 & ~n22792 ) | ( n22125 & n22791 ) | ( ~n22792 & n22791 ) ;
  assign n22793 = ( n22791 & ~n22121 ) | ( n22791 & n22792 ) | ( ~n22121 & n22792 ) ;
  assign n22795 = ( n22112 & ~n22794 ) | ( n22112 & n22793 ) | ( ~n22794 & n22793 ) ;
  assign n22778 = ( n22092 & ~n22097 ) | ( n22092 & n22511 ) | ( ~n22097 & n22511 ) ;
  assign n22777 = n22105 &  n22511 ;
  assign n22779 = ( n22511 & ~n22778 ) | ( n22511 & n22777 ) | ( ~n22778 & n22777 ) ;
  assign n22780 = ( n22777 & ~n22092 ) | ( n22777 & n22778 ) | ( ~n22092 & n22778 ) ;
  assign n22781 = ( n22097 & ~n22779 ) | ( n22097 & n22780 ) | ( ~n22779 & n22780 ) ;
  assign n22768 = n22103 | n22511 ;
  assign n22769 = ( n22090 & ~n22099 ) | ( n22090 & n22103 ) | ( ~n22099 & n22103 ) ;
  assign n22770 = ( n22099 & n22768 ) | ( n22099 & n22769 ) | ( n22768 & n22769 ) ;
  assign n22771 = ( n22103 & ~n22769 ) | ( n22103 & n22768 ) | ( ~n22769 & n22768 ) ;
  assign n22772 = ( n22090 & ~n22770 ) | ( n22090 & n22771 ) | ( ~n22770 & n22771 ) ;
  assign n22754 = n22083 &  n22511 ;
  assign n22755 = ( n22070 & n22075 ) | ( n22070 & n22511 ) | ( n22075 & n22511 ) ;
  assign n22757 = ( n22754 & ~n22070 ) | ( n22754 & n22755 ) | ( ~n22070 & n22755 ) ;
  assign n22756 = ( n22511 & ~n22755 ) | ( n22511 & n22754 ) | ( ~n22755 & n22754 ) ;
  assign n22758 = ( n22075 & ~n22757 ) | ( n22075 & n22756 ) | ( ~n22757 & n22756 ) ;
  assign n22745 = n22081 | n22511 ;
  assign n22746 = ( n22068 & ~n22081 ) | ( n22068 & n22077 ) | ( ~n22081 & n22077 ) ;
  assign n22748 = ( n22081 & n22745 ) | ( n22081 & n22746 ) | ( n22745 & n22746 ) ;
  assign n22747 = ( n22077 & ~n22746 ) | ( n22077 & n22745 ) | ( ~n22746 & n22745 ) ;
  assign n22749 = ( n22068 & ~n22748 ) | ( n22068 & n22747 ) | ( ~n22748 & n22747 ) ;
  assign n22732 = ( n22048 & ~n22511 ) | ( n22048 & n22053 ) | ( ~n22511 & n22053 ) ;
  assign n22731 = n22061 &  n22511 ;
  assign n22733 = ( n22511 & n22732 ) | ( n22511 & n22731 ) | ( n22732 & n22731 ) ;
  assign n22734 = ( n22731 & ~n22732 ) | ( n22731 & n22048 ) | ( ~n22732 & n22048 ) ;
  assign n22735 = ( n22053 & ~n22733 ) | ( n22053 & n22734 ) | ( ~n22733 & n22734 ) ;
  assign n22722 = n22059 | n22511 ;
  assign n22723 = ( n22046 & ~n22059 ) | ( n22046 & n22055 ) | ( ~n22059 & n22055 ) ;
  assign n22725 = ( n22059 & n22722 ) | ( n22059 & n22723 ) | ( n22722 & n22723 ) ;
  assign n22724 = ( n22055 & ~n22723 ) | ( n22055 & n22722 ) | ( ~n22723 & n22722 ) ;
  assign n22726 = ( n22046 & ~n22725 ) | ( n22046 & n22724 ) | ( ~n22725 & n22724 ) ;
  assign n22709 = ( n22026 & ~n22031 ) | ( n22026 & n22511 ) | ( ~n22031 & n22511 ) ;
  assign n22708 = n22039 &  n22511 ;
  assign n22710 = ( n22511 & ~n22709 ) | ( n22511 & n22708 ) | ( ~n22709 & n22708 ) ;
  assign n22711 = ( n22708 & ~n22026 ) | ( n22708 & n22709 ) | ( ~n22026 & n22709 ) ;
  assign n22712 = ( n22031 & ~n22710 ) | ( n22031 & n22711 ) | ( ~n22710 & n22711 ) ;
  assign n22699 = n22037 | n22511 ;
  assign n22700 = ( n22024 & ~n22037 ) | ( n22024 & n22033 ) | ( ~n22037 & n22033 ) ;
  assign n22702 = ( n22037 & n22699 ) | ( n22037 & n22700 ) | ( n22699 & n22700 ) ;
  assign n22701 = ( n22033 & ~n22700 ) | ( n22033 & n22699 ) | ( ~n22700 & n22699 ) ;
  assign n22703 = ( n22024 & ~n22702 ) | ( n22024 & n22701 ) | ( ~n22702 & n22701 ) ;
  assign n22686 = ( n22004 & ~n22009 ) | ( n22004 & n22511 ) | ( ~n22009 & n22511 ) ;
  assign n22685 = n22017 &  n22511 ;
  assign n22687 = ( n22511 & ~n22686 ) | ( n22511 & n22685 ) | ( ~n22686 & n22685 ) ;
  assign n22688 = ( n22685 & ~n22004 ) | ( n22685 & n22686 ) | ( ~n22004 & n22686 ) ;
  assign n22689 = ( n22009 & ~n22687 ) | ( n22009 & n22688 ) | ( ~n22687 & n22688 ) ;
  assign n22676 = n22015 | n22511 ;
  assign n22677 = ( n22002 & ~n22015 ) | ( n22002 & n22011 ) | ( ~n22015 & n22011 ) ;
  assign n22679 = ( n22015 & n22676 ) | ( n22015 & n22677 ) | ( n22676 & n22677 ) ;
  assign n22678 = ( n22011 & ~n22677 ) | ( n22011 & n22676 ) | ( ~n22677 & n22676 ) ;
  assign n22680 = ( n22002 & ~n22679 ) | ( n22002 & n22678 ) | ( ~n22679 & n22678 ) ;
  assign n22663 = ( n21982 & ~n21987 ) | ( n21982 & n22511 ) | ( ~n21987 & n22511 ) ;
  assign n22662 = n21995 &  n22511 ;
  assign n22664 = ( n22511 & ~n22663 ) | ( n22511 & n22662 ) | ( ~n22663 & n22662 ) ;
  assign n22665 = ( n22662 & ~n21982 ) | ( n22662 & n22663 ) | ( ~n21982 & n22663 ) ;
  assign n22666 = ( n21987 & ~n22664 ) | ( n21987 & n22665 ) | ( ~n22664 & n22665 ) ;
  assign n22653 = n21993 | n22511 ;
  assign n22654 = ( n21980 & ~n21993 ) | ( n21980 & n21989 ) | ( ~n21993 & n21989 ) ;
  assign n22656 = ( n21993 & n22653 ) | ( n21993 & n22654 ) | ( n22653 & n22654 ) ;
  assign n22655 = ( n21989 & ~n22654 ) | ( n21989 & n22653 ) | ( ~n22654 & n22653 ) ;
  assign n22657 = ( n21980 & ~n22656 ) | ( n21980 & n22655 ) | ( ~n22656 & n22655 ) ;
  assign n22639 = n21973 &  n22511 ;
  assign n22640 = ( n21960 & n21965 ) | ( n21960 & n22511 ) | ( n21965 & n22511 ) ;
  assign n22642 = ( n22639 & ~n21960 ) | ( n22639 & n22640 ) | ( ~n21960 & n22640 ) ;
  assign n22641 = ( n22511 & ~n22640 ) | ( n22511 & n22639 ) | ( ~n22640 & n22639 ) ;
  assign n22643 = ( n21965 & ~n22642 ) | ( n21965 & n22641 ) | ( ~n22642 & n22641 ) ;
  assign n22630 = n21971 | n22511 ;
  assign n22631 = ( n21958 & ~n21971 ) | ( n21958 & n21967 ) | ( ~n21971 & n21967 ) ;
  assign n22633 = ( n21971 & n22630 ) | ( n21971 & n22631 ) | ( n22630 & n22631 ) ;
  assign n22632 = ( n21967 & ~n22631 ) | ( n21967 & n22630 ) | ( ~n22631 & n22630 ) ;
  assign n22634 = ( n21958 & ~n22633 ) | ( n21958 & n22632 ) | ( ~n22633 & n22632 ) ;
  assign n22617 = ( n21938 & ~n21943 ) | ( n21938 & n22511 ) | ( ~n21943 & n22511 ) ;
  assign n22616 = n21951 &  n22511 ;
  assign n22618 = ( n22511 & ~n22617 ) | ( n22511 & n22616 ) | ( ~n22617 & n22616 ) ;
  assign n22619 = ( n22616 & ~n21938 ) | ( n22616 & n22617 ) | ( ~n21938 & n22617 ) ;
  assign n22620 = ( n21943 & ~n22618 ) | ( n21943 & n22619 ) | ( ~n22618 & n22619 ) ;
  assign n22607 = n21949 | n22511 ;
  assign n22608 = ( n21936 & ~n21949 ) | ( n21936 & n21945 ) | ( ~n21949 & n21945 ) ;
  assign n22610 = ( n21949 & n22607 ) | ( n21949 & n22608 ) | ( n22607 & n22608 ) ;
  assign n22609 = ( n21945 & ~n22608 ) | ( n21945 & n22607 ) | ( ~n22608 & n22607 ) ;
  assign n22611 = ( n21936 & ~n22610 ) | ( n21936 & n22609 ) | ( ~n22610 & n22609 ) ;
  assign n22594 = ( n21916 & ~n21921 ) | ( n21916 & n22511 ) | ( ~n21921 & n22511 ) ;
  assign n22593 = n21929 &  n22511 ;
  assign n22595 = ( n22511 & ~n22594 ) | ( n22511 & n22593 ) | ( ~n22594 & n22593 ) ;
  assign n22596 = ( n22593 & ~n21916 ) | ( n22593 & n22594 ) | ( ~n21916 & n22594 ) ;
  assign n22597 = ( n21921 & ~n22595 ) | ( n21921 & n22596 ) | ( ~n22595 & n22596 ) ;
  assign n22584 = n21927 | n22511 ;
  assign n22585 = ( n21914 & ~n21927 ) | ( n21914 & n21923 ) | ( ~n21927 & n21923 ) ;
  assign n22587 = ( n21927 & n22584 ) | ( n21927 & n22585 ) | ( n22584 & n22585 ) ;
  assign n22586 = ( n21923 & ~n22585 ) | ( n21923 & n22584 ) | ( ~n22585 & n22584 ) ;
  assign n22588 = ( n21914 & ~n22587 ) | ( n21914 & n22586 ) | ( ~n22587 & n22586 ) ;
  assign n22571 = n21907 &  n22511 ;
  assign n22572 = ( n21894 & n21899 ) | ( n21894 & n22511 ) | ( n21899 & n22511 ) ;
  assign n22574 = ( n22571 & ~n21894 ) | ( n22571 & n22572 ) | ( ~n21894 & n22572 ) ;
  assign n22573 = ( n22511 & ~n22572 ) | ( n22511 & n22571 ) | ( ~n22572 & n22571 ) ;
  assign n22575 = ( n21899 & ~n22574 ) | ( n21899 & n22573 ) | ( ~n22574 & n22573 ) ;
  assign n22562 = n21905 | n22511 ;
  assign n22563 = ( n21892 & ~n21905 ) | ( n21892 & n21901 ) | ( ~n21905 & n21901 ) ;
  assign n22565 = ( n21905 & n22562 ) | ( n21905 & n22563 ) | ( n22562 & n22563 ) ;
  assign n22564 = ( n21901 & ~n22563 ) | ( n21901 & n22562 ) | ( ~n22563 & n22562 ) ;
  assign n22566 = ( n21892 & ~n22565 ) | ( n21892 & n22564 ) | ( ~n22565 & n22564 ) ;
  assign n22555 = ( n21872 & ~n21877 ) | ( n21872 & n22511 ) | ( ~n21877 & n22511 ) ;
  assign n22554 = n21885 &  n22511 ;
  assign n22556 = ( n22511 & ~n22555 ) | ( n22511 & n22554 ) | ( ~n22555 & n22554 ) ;
  assign n22557 = ( n22554 & ~n21872 ) | ( n22554 & n22555 ) | ( ~n21872 & n22555 ) ;
  assign n22558 = ( n21877 & ~n22556 ) | ( n21877 & n22557 ) | ( ~n22556 & n22557 ) ;
  assign n22548 = n21883 | n22511 ;
  assign n22549 = ( n21870 & ~n21883 ) | ( n21870 & n21879 ) | ( ~n21883 & n21879 ) ;
  assign n22551 = ( n21883 & n22548 ) | ( n21883 & n22549 ) | ( n22548 & n22549 ) ;
  assign n22550 = ( n21879 & ~n22549 ) | ( n21879 & n22548 ) | ( ~n22549 & n22548 ) ;
  assign n22552 = ( n21870 & ~n22551 ) | ( n21870 & n22550 ) | ( ~n22551 & n22550 ) ;
  assign n22542 = n21846 | n22511 ;
  assign n22543 = ( n21856 & ~n21846 ) | ( n21856 & n21863 ) | ( ~n21846 & n21863 ) ;
  assign n22545 = ( n21846 & n22542 ) | ( n21846 & n22543 ) | ( n22542 & n22543 ) ;
  assign n22544 = ( n21863 & ~n22543 ) | ( n21863 & n22542 ) | ( ~n22543 & n22542 ) ;
  assign n22546 = ( n21856 & ~n22545 ) | ( n21856 & n22544 ) | ( ~n22545 & n22544 ) ;
  assign n22536 = ~n21858 & n21861 ;
  assign n22537 = ( n21844 & ~n21858 ) | ( n21844 & n22536 ) | ( ~n21858 & n22536 ) ;
  assign n22539 = ( n21858 & n22511 ) | ( n21858 & n22537 ) | ( n22511 & n22537 ) ;
  assign n22538 = ( n22511 & ~n22537 ) | ( n22511 & n22536 ) | ( ~n22537 & n22536 ) ;
  assign n22540 = ( n21844 & ~n22539 ) | ( n21844 & n22538 ) | ( ~n22539 & n22538 ) ;
  assign n21828 = ~x4 & n21818 ;
  assign n21829 = ( x5 & ~n21828 ) | ( x5 & 1'b0 ) | ( ~n21828 & 1'b0 ) ;
  assign n21831 = n21829 | n21830 ;
  assign n21826 = n21819 | n21823 ;
  assign n21827 = ( n21825 & ~n21819 ) | ( n21825 & n21826 ) | ( ~n21819 & n21826 ) ;
  assign n22512 = ( n21827 & ~n21831 ) | ( n21827 & n22511 ) | ( ~n21831 & n22511 ) ;
  assign n22514 = ( n22511 & ~n22512 ) | ( n22511 & 1'b0 ) | ( ~n22512 & 1'b0 ) ;
  assign n22513 = ~n21827 & n22512 ;
  assign n22515 = ( n21831 & ~n22514 ) | ( n21831 & n22513 ) | ( ~n22514 & n22513 ) ;
  assign n22517 = ( n21818 & ~n22509 ) | ( n21818 & 1'b0 ) | ( ~n22509 & 1'b0 ) ;
  assign n22518 = ( n22497 & ~n22517 ) | ( n22497 & n22505 ) | ( ~n22517 & n22505 ) ;
  assign n22519 = ( n22497 & ~n22518 ) | ( n22497 & 1'b0 ) | ( ~n22518 & 1'b0 ) ;
  assign n22516 = ~n21820 & n22511 ;
  assign n22520 = ~n22519 & n22516 ;
  assign n22521 = ( x4 & n22520 ) | ( x4 & n22519 ) | ( n22520 & n22519 ) ;
  assign n22522 = x4 | n22519 ;
  assign n22523 = n22516 | n22522 ;
  assign n22524 = ~n22521 & n22523 ;
  assign n22525 = x0 | x1 ;
  assign n22526 = ~x2 & n22525 ;
  assign n22527 = ( x2 & ~n22509 ) | ( x2 & 1'b0 ) | ( ~n22509 & 1'b0 ) ;
  assign n22528 = ( n22497 & ~n22527 ) | ( n22497 & n22505 ) | ( ~n22527 & n22505 ) ;
  assign n22529 = ( n22497 & ~n22528 ) | ( n22497 & 1'b0 ) | ( ~n22528 & 1'b0 ) ;
  assign n22530 = n22526 | n22529 ;
  assign n22531 = ~x2 & n22511 ;
  assign n22532 = ( x3 & ~n22531 ) | ( x3 & 1'b0 ) | ( ~n22531 & 1'b0 ) ;
  assign n22533 = n22516 | n22532 ;
  assign n22534 = ( n22530 & ~n21818 ) | ( n22530 & n22533 ) | ( ~n21818 & n22533 ) ;
  assign n22535 = ( n22524 & ~n21143 ) | ( n22524 & n22534 ) | ( ~n21143 & n22534 ) ;
  assign n22541 = ( n22515 & ~n20475 ) | ( n22515 & n22535 ) | ( ~n20475 & n22535 ) ;
  assign n22547 = ( n22540 & ~n19819 ) | ( n22540 & n22541 ) | ( ~n19819 & n22541 ) ;
  assign n22553 = ( n22546 & ~n19175 ) | ( n22546 & n22547 ) | ( ~n19175 & n22547 ) ;
  assign n22559 = ( n22552 & ~n18532 ) | ( n22552 & n22553 ) | ( ~n18532 & n22553 ) ;
  assign n22561 = n22558 &  n22559 ;
  assign n22560 = n22558 | n22559 ;
  assign n22580 = ~n17902 & n22560 ;
  assign n22581 = n22561 | n22580 ;
  assign n22582 = ( n22566 & ~n17279 ) | ( n22566 & n22581 ) | ( ~n17279 & n22581 ) ;
  assign n22583 = n22575 &  n22582 ;
  assign n22567 = n22561 | n22566 ;
  assign n22568 = n17902 | n22560 ;
  assign n22569 = ( n22567 & ~n17902 ) | ( n22567 & n22568 ) | ( ~n17902 & n22568 ) ;
  assign n22570 = ~n17279 & n22569 ;
  assign n22576 = ( n22558 & ~n17902 ) | ( n22558 & n22559 ) | ( ~n17902 & n22559 ) ;
  assign n22577 = n22566 &  n22576 ;
  assign n22578 = n22575 | n22577 ;
  assign n22579 = n22570 | n22578 ;
  assign n22603 = ~n16671 & n22579 ;
  assign n22604 = n22583 | n22603 ;
  assign n22605 = ( n22588 & ~n16070 ) | ( n22588 & n22604 ) | ( ~n16070 & n22604 ) ;
  assign n22606 = n22597 &  n22605 ;
  assign n22589 = n22583 | n22588 ;
  assign n22590 = n16671 | n22579 ;
  assign n22591 = ( n22589 & ~n16671 ) | ( n22589 & n22590 ) | ( ~n16671 & n22590 ) ;
  assign n22592 = ~n16070 & n22591 ;
  assign n22598 = n22570 | n22577 ;
  assign n22599 = ( n22575 & ~n16671 ) | ( n22575 & n22598 ) | ( ~n16671 & n22598 ) ;
  assign n22600 = n22588 &  n22599 ;
  assign n22601 = n22597 | n22600 ;
  assign n22602 = n22592 | n22601 ;
  assign n22626 = ~n15484 & n22602 ;
  assign n22627 = n22606 | n22626 ;
  assign n22628 = ( n22611 & ~n14905 ) | ( n22611 & n22627 ) | ( ~n14905 & n22627 ) ;
  assign n22629 = n22620 &  n22628 ;
  assign n22612 = n22606 | n22611 ;
  assign n22613 = n15484 | n22602 ;
  assign n22614 = ( n22612 & ~n15484 ) | ( n22612 & n22613 ) | ( ~n15484 & n22613 ) ;
  assign n22615 = ~n14905 & n22614 ;
  assign n22621 = n22592 | n22600 ;
  assign n22622 = ( n22597 & ~n15484 ) | ( n22597 & n22621 ) | ( ~n15484 & n22621 ) ;
  assign n22623 = n22611 &  n22622 ;
  assign n22624 = n22620 | n22623 ;
  assign n22625 = n22615 | n22624 ;
  assign n22649 = ~n14341 & n22625 ;
  assign n22650 = n22629 | n22649 ;
  assign n22651 = ( n22634 & ~n13784 ) | ( n22634 & n22650 ) | ( ~n13784 & n22650 ) ;
  assign n22652 = n22643 &  n22651 ;
  assign n22635 = n22629 | n22634 ;
  assign n22636 = n14341 | n22625 ;
  assign n22637 = ( n22635 & ~n14341 ) | ( n22635 & n22636 ) | ( ~n14341 & n22636 ) ;
  assign n22638 = ~n13784 & n22637 ;
  assign n22644 = n22615 | n22623 ;
  assign n22645 = ( n22620 & ~n14341 ) | ( n22620 & n22644 ) | ( ~n14341 & n22644 ) ;
  assign n22646 = n22634 &  n22645 ;
  assign n22647 = n22643 | n22646 ;
  assign n22648 = n22638 | n22647 ;
  assign n22672 = ~n13242 & n22648 ;
  assign n22673 = n22652 | n22672 ;
  assign n22674 = ( n22657 & ~n12707 ) | ( n22657 & n22673 ) | ( ~n12707 & n22673 ) ;
  assign n22675 = n22666 &  n22674 ;
  assign n22658 = n22652 | n22657 ;
  assign n22659 = n13242 | n22648 ;
  assign n22660 = ( n22658 & ~n13242 ) | ( n22658 & n22659 ) | ( ~n13242 & n22659 ) ;
  assign n22661 = ~n12707 & n22660 ;
  assign n22667 = n22638 | n22646 ;
  assign n22668 = ( n22643 & ~n13242 ) | ( n22643 & n22667 ) | ( ~n13242 & n22667 ) ;
  assign n22669 = n22657 &  n22668 ;
  assign n22670 = n22666 | n22669 ;
  assign n22671 = n22661 | n22670 ;
  assign n22695 = ~n12187 & n22671 ;
  assign n22696 = n22675 | n22695 ;
  assign n22697 = ( n22680 & ~n11674 ) | ( n22680 & n22696 ) | ( ~n11674 & n22696 ) ;
  assign n22698 = n22689 &  n22697 ;
  assign n22681 = n22675 | n22680 ;
  assign n22682 = n12187 | n22671 ;
  assign n22683 = ( n22681 & ~n12187 ) | ( n22681 & n22682 ) | ( ~n12187 & n22682 ) ;
  assign n22684 = ~n11674 & n22683 ;
  assign n22690 = n22661 | n22669 ;
  assign n22691 = ( n22666 & ~n12187 ) | ( n22666 & n22690 ) | ( ~n12187 & n22690 ) ;
  assign n22692 = n22680 &  n22691 ;
  assign n22693 = n22689 | n22692 ;
  assign n22694 = n22684 | n22693 ;
  assign n22718 = ~n11176 & n22694 ;
  assign n22719 = n22698 | n22718 ;
  assign n22720 = ( n22703 & ~n10685 ) | ( n22703 & n22719 ) | ( ~n10685 & n22719 ) ;
  assign n22721 = n22712 &  n22720 ;
  assign n22704 = n22698 | n22703 ;
  assign n22705 = n11176 | n22694 ;
  assign n22706 = ( n22704 & ~n11176 ) | ( n22704 & n22705 ) | ( ~n11176 & n22705 ) ;
  assign n22707 = ~n10685 & n22706 ;
  assign n22713 = n22684 | n22692 ;
  assign n22714 = ( n22689 & ~n11176 ) | ( n22689 & n22713 ) | ( ~n11176 & n22713 ) ;
  assign n22715 = n22703 &  n22714 ;
  assign n22716 = n22712 | n22715 ;
  assign n22717 = n22707 | n22716 ;
  assign n22741 = ~n10209 & n22717 ;
  assign n22742 = n22721 | n22741 ;
  assign n22743 = ( n9740 & n22726 ) | ( n9740 & n22742 ) | ( n22726 & n22742 ) ;
  assign n22744 = n22735 &  n22743 ;
  assign n22727 = n22721 | n22726 ;
  assign n22728 = n10209 | n22717 ;
  assign n22729 = ( n22727 & ~n10209 ) | ( n22727 & n22728 ) | ( ~n10209 & n22728 ) ;
  assign n22730 = n9740 &  n22729 ;
  assign n22736 = n22707 | n22715 ;
  assign n22737 = ( n22712 & ~n10209 ) | ( n22712 & n22736 ) | ( ~n10209 & n22736 ) ;
  assign n22738 = n22726 &  n22737 ;
  assign n22739 = n22735 | n22738 ;
  assign n22740 = n22730 | n22739 ;
  assign n22764 = ~n9286 & n22740 ;
  assign n22765 = n22744 | n22764 ;
  assign n22766 = ( n22749 & ~n8839 ) | ( n22749 & n22765 ) | ( ~n8839 & n22765 ) ;
  assign n22767 = n22758 &  n22766 ;
  assign n22750 = n22744 | n22749 ;
  assign n22751 = n9286 | n22740 ;
  assign n22752 = ( n22750 & ~n9286 ) | ( n22750 & n22751 ) | ( ~n9286 & n22751 ) ;
  assign n22753 = ~n8839 & n22752 ;
  assign n22759 = n22730 | n22738 ;
  assign n22760 = ( n22735 & ~n9286 ) | ( n22735 & n22759 ) | ( ~n9286 & n22759 ) ;
  assign n22761 = n22749 &  n22760 ;
  assign n22762 = n22758 | n22761 ;
  assign n22763 = n22753 | n22762 ;
  assign n22787 = ~n8407 & n22763 ;
  assign n22788 = n22767 | n22787 ;
  assign n22789 = ( n22772 & ~n7982 ) | ( n22772 & n22788 ) | ( ~n7982 & n22788 ) ;
  assign n22790 = n22781 &  n22789 ;
  assign n22773 = n22767 | n22772 ;
  assign n22774 = n8407 | n22763 ;
  assign n22775 = ( n22773 & ~n8407 ) | ( n22773 & n22774 ) | ( ~n8407 & n22774 ) ;
  assign n22776 = ~n7982 & n22775 ;
  assign n22782 = n22753 | n22761 ;
  assign n22783 = ( n22758 & ~n8407 ) | ( n22758 & n22782 ) | ( ~n8407 & n22782 ) ;
  assign n22784 = n22772 &  n22783 ;
  assign n22785 = n22781 | n22784 ;
  assign n22786 = n22776 | n22785 ;
  assign n22810 = n7572 &  n22786 ;
  assign n22811 = n22790 | n22810 ;
  assign n22812 = ( n7169 & n22795 ) | ( n7169 & n22811 ) | ( n22795 & n22811 ) ;
  assign n22813 = n22804 &  n22812 ;
  assign n22797 = ( n7572 & ~n22786 ) | ( n7572 & 1'b0 ) | ( ~n22786 & 1'b0 ) ;
  assign n22796 = n22790 | n22795 ;
  assign n22798 = ( n7572 & ~n22797 ) | ( n7572 & n22796 ) | ( ~n22797 & n22796 ) ;
  assign n22799 = n7169 &  n22798 ;
  assign n22805 = n22776 | n22784 ;
  assign n22806 = ( n7572 & n22781 ) | ( n7572 & n22805 ) | ( n22781 & n22805 ) ;
  assign n22807 = n22795 &  n22806 ;
  assign n22808 = n22804 | n22807 ;
  assign n22809 = n22799 | n22808 ;
  assign n22833 = ~n6781 & n22809 ;
  assign n22834 = n22813 | n22833 ;
  assign n22835 = ( n6399 & n22818 ) | ( n6399 & n22834 ) | ( n22818 & n22834 ) ;
  assign n22836 = n22827 &  n22835 ;
  assign n22819 = n22813 | n22818 ;
  assign n22820 = n6781 | n22809 ;
  assign n22821 = ( n22819 & ~n6781 ) | ( n22819 & n22820 ) | ( ~n6781 & n22820 ) ;
  assign n22822 = n6399 &  n22821 ;
  assign n22828 = n22799 | n22807 ;
  assign n22829 = ( n22804 & ~n6781 ) | ( n22804 & n22828 ) | ( ~n6781 & n22828 ) ;
  assign n22830 = n22818 &  n22829 ;
  assign n22831 = n22827 | n22830 ;
  assign n22832 = n22822 | n22831 ;
  assign n22856 = ~n6032 & n22832 ;
  assign n22857 = n22836 | n22856 ;
  assign n22858 = ( n5672 & n22841 ) | ( n5672 & n22857 ) | ( n22841 & n22857 ) ;
  assign n22859 = n22850 &  n22858 ;
  assign n22843 = n22832 | n6032 ;
  assign n22842 = n22836 | n22841 ;
  assign n22844 = ( n22843 & ~n6032 ) | ( n22843 & n22842 ) | ( ~n6032 & n22842 ) ;
  assign n22845 = n5672 &  n22844 ;
  assign n22851 = n22822 | n22830 ;
  assign n22852 = ( n22827 & ~n6032 ) | ( n22827 & n22851 ) | ( ~n6032 & n22851 ) ;
  assign n22853 = n22841 &  n22852 ;
  assign n22854 = n22850 | n22853 ;
  assign n22855 = n22845 | n22854 ;
  assign n22879 = ~n5327 & n22855 ;
  assign n22880 = n22859 | n22879 ;
  assign n22881 = ( n22864 & ~n4990 ) | ( n22864 & n22880 ) | ( ~n4990 & n22880 ) ;
  assign n22882 = n22873 &  n22881 ;
  assign n22866 = n22855 | n5327 ;
  assign n22865 = n22859 | n22864 ;
  assign n22867 = ( n22866 & ~n5327 ) | ( n22866 & n22865 ) | ( ~n5327 & n22865 ) ;
  assign n22868 = ~n4990 & n22867 ;
  assign n22874 = n22845 | n22853 ;
  assign n22875 = ( n22850 & ~n5327 ) | ( n22850 & n22874 ) | ( ~n5327 & n22874 ) ;
  assign n22876 = n22864 &  n22875 ;
  assign n22877 = n22873 | n22876 ;
  assign n22878 = n22868 | n22877 ;
  assign n22902 = ~n4668 & n22878 ;
  assign n22903 = n22882 | n22902 ;
  assign n22904 = ( n22887 & ~n4353 ) | ( n22887 & n22903 ) | ( ~n4353 & n22903 ) ;
  assign n22905 = n22896 &  n22904 ;
  assign n22888 = n22882 | n22887 ;
  assign n22889 = n4668 | n22878 ;
  assign n22890 = ( n22888 & ~n4668 ) | ( n22888 & n22889 ) | ( ~n4668 & n22889 ) ;
  assign n22891 = ~n4353 & n22890 ;
  assign n22897 = n22868 | n22876 ;
  assign n22898 = ( n22873 & ~n4668 ) | ( n22873 & n22897 ) | ( ~n4668 & n22897 ) ;
  assign n22899 = n22887 &  n22898 ;
  assign n22900 = n22896 | n22899 ;
  assign n22901 = n22891 | n22900 ;
  assign n22925 = ~n4053 & n22901 ;
  assign n22926 = n22905 | n22925 ;
  assign n22927 = ( n22910 & ~n3760 ) | ( n22910 & n22926 ) | ( ~n3760 & n22926 ) ;
  assign n22928 = n22919 &  n22927 ;
  assign n22911 = n22905 | n22910 ;
  assign n22912 = n4053 | n22901 ;
  assign n22913 = ( n22911 & ~n4053 ) | ( n22911 & n22912 ) | ( ~n4053 & n22912 ) ;
  assign n22914 = ~n3760 & n22913 ;
  assign n22920 = n22891 | n22899 ;
  assign n22921 = ( n22896 & ~n4053 ) | ( n22896 & n22920 ) | ( ~n4053 & n22920 ) ;
  assign n22922 = n22910 &  n22921 ;
  assign n22923 = n22919 | n22922 ;
  assign n22924 = n22914 | n22923 ;
  assign n22948 = ~n3482 & n22924 ;
  assign n22949 = n22928 | n22948 ;
  assign n22950 = ( n22933 & ~n3211 ) | ( n22933 & n22949 ) | ( ~n3211 & n22949 ) ;
  assign n22951 = n22942 &  n22950 ;
  assign n22934 = n22928 | n22933 ;
  assign n22935 = n3482 | n22924 ;
  assign n22936 = ( n22934 & ~n3482 ) | ( n22934 & n22935 ) | ( ~n3482 & n22935 ) ;
  assign n22937 = ~n3211 & n22936 ;
  assign n22943 = n22914 | n22922 ;
  assign n22944 = ( n22919 & ~n3482 ) | ( n22919 & n22943 ) | ( ~n3482 & n22943 ) ;
  assign n22945 = n22933 &  n22944 ;
  assign n22946 = n22942 | n22945 ;
  assign n22947 = n22937 | n22946 ;
  assign n22971 = ~n2955 & n22947 ;
  assign n22972 = n22951 | n22971 ;
  assign n22973 = ( n22956 & ~n2706 ) | ( n22956 & n22972 ) | ( ~n2706 & n22972 ) ;
  assign n22974 = n22965 &  n22973 ;
  assign n22958 = n22947 | n2955 ;
  assign n22957 = n22951 | n22956 ;
  assign n22959 = ( n22958 & ~n2955 ) | ( n22958 & n22957 ) | ( ~n2955 & n22957 ) ;
  assign n22960 = ~n2706 & n22959 ;
  assign n22966 = n22937 | n22945 ;
  assign n22967 = ( n22942 & ~n2955 ) | ( n22942 & n22966 ) | ( ~n2955 & n22966 ) ;
  assign n22968 = n22956 &  n22967 ;
  assign n22969 = n22965 | n22968 ;
  assign n22970 = n22960 | n22969 ;
  assign n22994 = ~n2472 & n22970 ;
  assign n22995 = n22974 | n22994 ;
  assign n22996 = ( n22979 & ~n2245 ) | ( n22979 & n22995 ) | ( ~n2245 & n22995 ) ;
  assign n22997 = ~n22988 & n22996 ;
  assign n22980 = n22974 | n22979 ;
  assign n22981 = n2472 | n22970 ;
  assign n22982 = ( n22980 & ~n2472 ) | ( n22980 & n22981 ) | ( ~n2472 & n22981 ) ;
  assign n22983 = ~n2245 & n22982 ;
  assign n22989 = n22960 | n22968 ;
  assign n22990 = ( n22965 & ~n2472 ) | ( n22965 & n22989 ) | ( ~n2472 & n22989 ) ;
  assign n22991 = n22979 &  n22990 ;
  assign n22992 = ( n22988 & ~n22991 ) | ( n22988 & 1'b0 ) | ( ~n22991 & 1'b0 ) ;
  assign n22993 = ~n22983 & n22992 ;
  assign n23017 = ( n2033 & ~n22993 ) | ( n2033 & 1'b0 ) | ( ~n22993 & 1'b0 ) ;
  assign n23018 = n22997 | n23017 ;
  assign n22998 = n22323 | n22511 ;
  assign n22999 = ( n22310 & ~n22323 ) | ( n22310 & n22319 ) | ( ~n22323 & n22319 ) ;
  assign n23001 = ( n22323 & n22998 ) | ( n22323 & n22999 ) | ( n22998 & n22999 ) ;
  assign n23000 = ( n22319 & ~n22999 ) | ( n22319 & n22998 ) | ( ~n22999 & n22998 ) ;
  assign n23002 = ( n22310 & ~n23001 ) | ( n22310 & n23000 ) | ( ~n23001 & n23000 ) ;
  assign n23019 = ( n1827 & ~n23018 ) | ( n1827 & n23002 ) | ( ~n23018 & n23002 ) ;
  assign n23020 = n23011 | n23019 ;
  assign n23003 = ~n22997 & n23002 ;
  assign n23004 = n2033 &  n22993 ;
  assign n23005 = ( n23003 & ~n2033 ) | ( n23003 & n23004 ) | ( ~n2033 & n23004 ) ;
  assign n23006 = n1827 | n23005 ;
  assign n23012 = n22983 | n22991 ;
  assign n23013 = ( n2033 & ~n22988 ) | ( n2033 & n23012 ) | ( ~n22988 & n23012 ) ;
  assign n23014 = ~n23002 & n23013 ;
  assign n23015 = ( n23011 & ~n23014 ) | ( n23011 & 1'b0 ) | ( ~n23014 & 1'b0 ) ;
  assign n23016 = n23006 &  n23015 ;
  assign n23040 = ( n1636 & ~n23016 ) | ( n1636 & 1'b0 ) | ( ~n23016 & 1'b0 ) ;
  assign n23041 = ( n23020 & ~n23040 ) | ( n23020 & 1'b0 ) | ( ~n23040 & 1'b0 ) ;
  assign n23042 = ( n23025 & ~n1452 ) | ( n23025 & n23041 ) | ( ~n1452 & n23041 ) ;
  assign n23043 = n23034 | n23042 ;
  assign n23027 = n23016 &  n1636 ;
  assign n23026 = n23020 &  n23025 ;
  assign n23028 = ( n23027 & ~n1636 ) | ( n23027 & n23026 ) | ( ~n1636 & n23026 ) ;
  assign n23029 = ( n1452 & ~n23028 ) | ( n1452 & 1'b0 ) | ( ~n23028 & 1'b0 ) ;
  assign n23035 = ( n23006 & ~n23014 ) | ( n23006 & 1'b0 ) | ( ~n23014 & 1'b0 ) ;
  assign n23036 = ( n23011 & ~n1636 ) | ( n23011 & n23035 ) | ( ~n1636 & n23035 ) ;
  assign n23037 = n23025 | n23036 ;
  assign n23038 = n23034 &  n23037 ;
  assign n23039 = ~n23029 & n23038 ;
  assign n23063 = n1283 | n23039 ;
  assign n23064 = n23043 &  n23063 ;
  assign n23044 = n22367 | n22511 ;
  assign n23045 = ( n22354 & n22363 ) | ( n22354 & n22367 ) | ( n22363 & n22367 ) ;
  assign n23046 = ( n23044 & ~n22363 ) | ( n23044 & n23045 ) | ( ~n22363 & n23045 ) ;
  assign n23047 = ( n22367 & ~n23045 ) | ( n22367 & n23044 ) | ( ~n23045 & n23044 ) ;
  assign n23048 = ( n22354 & ~n23046 ) | ( n22354 & n23047 ) | ( ~n23046 & n23047 ) ;
  assign n23065 = ( n1122 & ~n23064 ) | ( n1122 & n23048 ) | ( ~n23064 & n23048 ) ;
  assign n23066 = n23057 &  n23065 ;
  assign n23049 = ( n23043 & ~n23048 ) | ( n23043 & 1'b0 ) | ( ~n23048 & 1'b0 ) ;
  assign n23050 = ~n1283 & n23039 ;
  assign n23051 = ( n1283 & n23049 ) | ( n1283 & n23050 ) | ( n23049 & n23050 ) ;
  assign n23052 = ( n1122 & ~n23051 ) | ( n1122 & 1'b0 ) | ( ~n23051 & 1'b0 ) ;
  assign n23058 = ~n23029 & n23037 ;
  assign n23059 = ( n1283 & n23034 ) | ( n1283 & n23058 ) | ( n23034 & n23058 ) ;
  assign n23060 = ( n23048 & ~n23059 ) | ( n23048 & 1'b0 ) | ( ~n23059 & 1'b0 ) ;
  assign n23061 = n23057 | n23060 ;
  assign n23062 = n23052 | n23061 ;
  assign n23086 = n976 &  n23062 ;
  assign n23087 = n23066 | n23086 ;
  assign n23067 = ( n22389 & ~n22511 ) | ( n22389 & 1'b0 ) | ( ~n22511 & 1'b0 ) ;
  assign n23068 = ( n22376 & n22385 ) | ( n22376 & n22389 ) | ( n22385 & n22389 ) ;
  assign n23069 = ( n23067 & ~n22385 ) | ( n23067 & n23068 ) | ( ~n22385 & n23068 ) ;
  assign n23070 = ( n22389 & ~n23068 ) | ( n22389 & n23067 ) | ( ~n23068 & n23067 ) ;
  assign n23071 = ( n22376 & ~n23069 ) | ( n22376 & n23070 ) | ( ~n23069 & n23070 ) ;
  assign n23088 = ( n837 & ~n23087 ) | ( n837 & n23071 ) | ( ~n23087 & n23071 ) ;
  assign n23089 = ( n23080 & ~n23088 ) | ( n23080 & 1'b0 ) | ( ~n23088 & 1'b0 ) ;
  assign n23073 = ~n23062 & n976 ;
  assign n23072 = ~n23066 & n23071 ;
  assign n23074 = ( n23073 & ~n976 ) | ( n23073 & n23072 ) | ( ~n976 & n23072 ) ;
  assign n23075 = n837 | n23074 ;
  assign n23081 = n23052 | n23060 ;
  assign n23082 = ( n976 & n23057 ) | ( n976 & n23081 ) | ( n23057 & n23081 ) ;
  assign n23083 = ~n23071 & n23082 ;
  assign n23084 = n23080 | n23083 ;
  assign n23085 = ( n23075 & ~n23084 ) | ( n23075 & 1'b0 ) | ( ~n23084 & 1'b0 ) ;
  assign n23109 = n713 | n23085 ;
  assign n23110 = ~n23089 & n23109 ;
  assign n23111 = ( n595 & n23094 ) | ( n595 & n23110 ) | ( n23094 & n23110 ) ;
  assign n23112 = n23103 | n23111 ;
  assign n23095 = ~n23089 & n23094 ;
  assign n23096 = ~n713 & n23085 ;
  assign n23097 = ( n713 & n23095 ) | ( n713 & n23096 ) | ( n23095 & n23096 ) ;
  assign n23098 = n595 | n23097 ;
  assign n23104 = ( n23075 & ~n23083 ) | ( n23075 & 1'b0 ) | ( ~n23083 & 1'b0 ) ;
  assign n23105 = ( n713 & ~n23080 ) | ( n713 & n23104 ) | ( ~n23080 & n23104 ) ;
  assign n23106 = n23094 | n23105 ;
  assign n23107 = n23103 &  n23106 ;
  assign n23108 = n23098 &  n23107 ;
  assign n23132 = n492 | n23108 ;
  assign n23133 = n23112 &  n23132 ;
  assign n23134 = ( n396 & ~n23117 ) | ( n396 & n23133 ) | ( ~n23117 & n23133 ) ;
  assign n23135 = ( n23126 & ~n23134 ) | ( n23126 & 1'b0 ) | ( ~n23134 & 1'b0 ) ;
  assign n23119 = ~n492 & n23108 ;
  assign n23118 = ( n23112 & ~n23117 ) | ( n23112 & 1'b0 ) | ( ~n23117 & 1'b0 ) ;
  assign n23120 = ( n492 & n23119 ) | ( n492 & n23118 ) | ( n23119 & n23118 ) ;
  assign n23121 = n396 | n23120 ;
  assign n23127 = n23098 &  n23106 ;
  assign n23128 = ( n492 & n23103 ) | ( n492 & n23127 ) | ( n23103 & n23127 ) ;
  assign n23129 = ( n23117 & ~n23128 ) | ( n23117 & 1'b0 ) | ( ~n23128 & 1'b0 ) ;
  assign n23130 = n23126 | n23129 ;
  assign n23131 = ( n23121 & ~n23130 ) | ( n23121 & 1'b0 ) | ( ~n23130 & 1'b0 ) ;
  assign n23155 = n315 | n23131 ;
  assign n23156 = ~n23135 & n23155 ;
  assign n23157 = ( n240 & ~n23140 ) | ( n240 & n23156 ) | ( ~n23140 & n23156 ) ;
  assign n23158 = ( n23149 & ~n23157 ) | ( n23149 & 1'b0 ) | ( ~n23157 & 1'b0 ) ;
  assign n23160 = ( n22473 & ~n22464 ) | ( n22473 & n22477 ) | ( ~n22464 & n22477 ) ;
  assign n23159 = n22477 | n22511 ;
  assign n23162 = ( n22477 & ~n23160 ) | ( n22477 & n23159 ) | ( ~n23160 & n23159 ) ;
  assign n23161 = ( n23159 & ~n22473 ) | ( n23159 & n23160 ) | ( ~n22473 & n23160 ) ;
  assign n23163 = ( n22464 & ~n23162 ) | ( n22464 & n23161 ) | ( ~n23162 & n23161 ) ;
  assign n23164 = n23158 | n23163 ;
  assign n23141 = n23135 | n23140 ;
  assign n23142 = ~n315 & n23131 ;
  assign n23143 = ( n315 & ~n23141 ) | ( n315 & n23142 ) | ( ~n23141 & n23142 ) ;
  assign n23144 = n240 | n23143 ;
  assign n23150 = ( n23121 & ~n23129 ) | ( n23121 & 1'b0 ) | ( ~n23129 & 1'b0 ) ;
  assign n23151 = ( n315 & ~n23126 ) | ( n315 & n23150 ) | ( ~n23126 & n23150 ) ;
  assign n23152 = ( n23140 & ~n23151 ) | ( n23140 & 1'b0 ) | ( ~n23151 & 1'b0 ) ;
  assign n23153 = n23149 | n23152 ;
  assign n23154 = ( n23144 & ~n23153 ) | ( n23144 & 1'b0 ) | ( ~n23153 & 1'b0 ) ;
  assign n23165 = ~n181 & n23154 ;
  assign n23166 = ( n181 & ~n23164 ) | ( n181 & n23165 ) | ( ~n23164 & n23165 ) ;
  assign n23167 = ( n145 & ~n23166 ) | ( n145 & 1'b0 ) | ( ~n23166 & 1'b0 ) ;
  assign n23173 = ( n23144 & ~n23152 ) | ( n23144 & 1'b0 ) | ( ~n23152 & 1'b0 ) ;
  assign n23174 = ( n181 & ~n23149 ) | ( n181 & n23173 ) | ( ~n23149 & n23173 ) ;
  assign n23175 = ( n23163 & ~n23174 ) | ( n23163 & 1'b0 ) | ( ~n23174 & 1'b0 ) ;
  assign n23194 = n23167 | n23175 ;
  assign n23168 = n22466 | n22511 ;
  assign n23169 = ( n22466 & ~n22479 ) | ( n22466 & n22471 ) | ( ~n22479 & n22471 ) ;
  assign n23170 = ( n22479 & n23168 ) | ( n22479 & n23169 ) | ( n23168 & n23169 ) ;
  assign n23171 = ( n22466 & ~n23169 ) | ( n22466 & n23168 ) | ( ~n23169 & n23168 ) ;
  assign n23172 = ( n22471 & ~n23170 ) | ( n22471 & n23171 ) | ( ~n23170 & n23171 ) ;
  assign n23195 = ( n150 & ~n23194 ) | ( n150 & n23172 ) | ( ~n23194 & n23172 ) ;
  assign n23196 = ( n23186 & ~n23195 ) | ( n23186 & 1'b0 ) | ( ~n23195 & 1'b0 ) ;
  assign n23198 = ( n133 & ~n22491 ) | ( n133 & n22487 ) | ( ~n22491 & n22487 ) ;
  assign n23197 = ( n22491 & ~n22487 ) | ( n22491 & n22511 ) | ( ~n22487 & n22511 ) ;
  assign n23199 = ~n22491 & n23197 ;
  assign n23200 = ( n22491 & n23198 ) | ( n22491 & n23199 ) | ( n23198 & n23199 ) ;
  assign n23201 = n23196 | n23200 ;
  assign n23178 = n181 | n23154 ;
  assign n23179 = ~n23158 & n23178 ;
  assign n23180 = ( n145 & ~n23179 ) | ( n145 & n23163 ) | ( ~n23179 & n23163 ) ;
  assign n23181 = ~n23172 & n23180 ;
  assign n23187 = ( n22487 & ~n22491 ) | ( n22487 & 1'b0 ) | ( ~n22491 & 1'b0 ) ;
  assign n23188 = ~n22511 & n23187 ;
  assign n23189 = ( n22505 & ~n23188 ) | ( n22505 & n23187 ) | ( ~n23188 & n23187 ) ;
  assign n23190 = n23186 | n23189 ;
  assign n23191 = n23181 | n23190 ;
  assign n23176 = ( n23172 & ~n23175 ) | ( n23172 & 1'b0 ) | ( ~n23175 & 1'b0 ) ;
  assign n23177 = ~n23167 & n23176 ;
  assign n23192 = ~n150 & n23177 ;
  assign n23193 = ( n150 & ~n23191 ) | ( n150 & n23192 ) | ( ~n23191 & n23192 ) ;
  assign n23202 = ~n133 & n23193 ;
  assign n23203 = ( n133 & ~n23201 ) | ( n133 & n23202 ) | ( ~n23201 & n23202 ) ;
  assign y0 = ~n23203 ;
  assign y1 = n22511 ;
  assign y2 = n21818 ;
  assign y3 = n21143 ;
  assign y4 = n20475 ;
  assign y5 = n19819 ;
  assign y6 = n19175 ;
  assign y7 = n18532 ;
  assign y8 = n17902 ;
  assign y9 = n17279 ;
  assign y10 = n16671 ;
  assign y11 = n16070 ;
  assign y12 = n15484 ;
  assign y13 = n14905 ;
  assign y14 = n14341 ;
  assign y15 = n13784 ;
  assign y16 = n13242 ;
  assign y17 = n12707 ;
  assign y18 = n12187 ;
  assign y19 = n11674 ;
  assign y20 = n11176 ;
  assign y21 = n10685 ;
  assign y22 = n10209 ;
  assign y23 = ~n9740 ;
  assign y24 = n9286 ;
  assign y25 = n8839 ;
  assign y26 = n8407 ;
  assign y27 = n7982 ;
  assign y28 = ~n7572 ;
  assign y29 = ~n7169 ;
  assign y30 = n6781 ;
  assign y31 = ~n6399 ;
  assign y32 = n6032 ;
  assign y33 = ~n5672 ;
  assign y34 = n5327 ;
  assign y35 = n4990 ;
  assign y36 = n4668 ;
  assign y37 = n4353 ;
  assign y38 = n4053 ;
  assign y39 = n3760 ;
  assign y40 = n3482 ;
  assign y41 = n3211 ;
  assign y42 = n2955 ;
  assign y43 = n2706 ;
  assign y44 = n2472 ;
  assign y45 = n2245 ;
  assign y46 = ~n2033 ;
  assign y47 = n1827 ;
  assign y48 = ~n1636 ;
  assign y49 = ~n1452 ;
  assign y50 = n1283 ;
  assign y51 = ~n1122 ;
  assign y52 = ~n976 ;
  assign y53 = n837 ;
  assign y54 = n713 ;
  assign y55 = n595 ;
  assign y56 = n492 ;
  assign y57 = n396 ;
  assign y58 = n315 ;
  assign y59 = n240 ;
  assign y60 = n181 ;
  assign y61 = ~n145 ;
  assign y62 = n150 ;
  assign y63 = n133 ;
endmodule
