module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 ;
  assign n136 = ( x26 & ~x128 ) | ( x26 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n137 = x25 &  x128 ;
  assign n138 = ( x129 & n136 ) | ( x129 & n137 ) | ( n136 & n137 ) ;
  assign n139 = x27 &  x128 ;
  assign n140 = ( x28 & ~x128 ) | ( x28 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n141 = ( n139 & ~x129 ) | ( n139 & n140 ) | ( ~x129 & n140 ) ;
  assign n142 = n138 | n141 ;
  assign n143 = x130 &  n142 ;
  assign n144 = ( x30 & ~x128 ) | ( x30 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n145 = x29 &  x128 ;
  assign n146 = ( x129 & n144 ) | ( x129 & n145 ) | ( n144 & n145 ) ;
  assign n147 = x31 &  x128 ;
  assign n148 = ( x32 & ~x128 ) | ( x32 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n149 = ( n147 & ~x129 ) | ( n147 & n148 ) | ( ~x129 & n148 ) ;
  assign n150 = n146 | n149 ;
  assign n151 = ~x130 & n150 ;
  assign n152 = ( n143 & ~x131 ) | ( n143 & n151 ) | ( ~x131 & n151 ) ;
  assign n153 = ( x22 & ~x128 ) | ( x22 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n154 = x21 &  x128 ;
  assign n155 = ( x129 & n153 ) | ( x129 & n154 ) | ( n153 & n154 ) ;
  assign n156 = x23 &  x128 ;
  assign n157 = ( x24 & ~x128 ) | ( x24 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n158 = ( n156 & ~x129 ) | ( n156 & n157 ) | ( ~x129 & n157 ) ;
  assign n159 = n155 | n158 ;
  assign n160 = ~x130 & n159 ;
  assign n161 = ( x18 & ~x128 ) | ( x18 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n162 = x17 &  x128 ;
  assign n163 = ( x129 & n161 ) | ( x129 & n162 ) | ( n161 & n162 ) ;
  assign n164 = x19 &  x128 ;
  assign n165 = ( x20 & ~x128 ) | ( x20 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n166 = ( n164 & ~x129 ) | ( n164 & n165 ) | ( ~x129 & n165 ) ;
  assign n167 = n163 | n166 ;
  assign n168 = x130 &  n167 ;
  assign n169 = ( x131 & n160 ) | ( x131 & n168 ) | ( n160 & n168 ) ;
  assign n170 = n152 | n169 ;
  assign n171 = ~x132 & n170 ;
  assign n172 = ( x10 & ~x128 ) | ( x10 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n173 = x9 &  x128 ;
  assign n174 = ( x129 & n172 ) | ( x129 & n173 ) | ( n172 & n173 ) ;
  assign n175 = x11 &  x128 ;
  assign n176 = ( x12 & ~x128 ) | ( x12 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n177 = ( n175 & ~x129 ) | ( n175 & n176 ) | ( ~x129 & n176 ) ;
  assign n178 = n174 | n177 ;
  assign n179 = x130 &  n178 ;
  assign n180 = ( x14 & ~x128 ) | ( x14 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n181 = x13 &  x128 ;
  assign n182 = ( x129 & n180 ) | ( x129 & n181 ) | ( n180 & n181 ) ;
  assign n183 = x15 &  x128 ;
  assign n184 = ( x16 & ~x128 ) | ( x16 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n185 = ( n183 & ~x129 ) | ( n183 & n184 ) | ( ~x129 & n184 ) ;
  assign n186 = n182 | n185 ;
  assign n187 = ~x130 & n186 ;
  assign n188 = ( n179 & ~x131 ) | ( n179 & n187 ) | ( ~x131 & n187 ) ;
  assign n189 = ( x6 & ~x128 ) | ( x6 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n190 = x5 &  x128 ;
  assign n191 = ( x129 & n189 ) | ( x129 & n190 ) | ( n189 & n190 ) ;
  assign n192 = x7 &  x128 ;
  assign n193 = ( x8 & ~x128 ) | ( x8 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n194 = ( n192 & ~x129 ) | ( n192 & n193 ) | ( ~x129 & n193 ) ;
  assign n195 = n191 | n194 ;
  assign n196 = ~x130 & n195 ;
  assign n197 = ( x2 & ~x128 ) | ( x2 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n198 = x1 &  x128 ;
  assign n199 = ( x129 & n197 ) | ( x129 & n198 ) | ( n197 & n198 ) ;
  assign n200 = x3 &  x128 ;
  assign n201 = ( x4 & ~x128 ) | ( x4 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n202 = ( n200 & ~x129 ) | ( n200 & n201 ) | ( ~x129 & n201 ) ;
  assign n203 = n199 | n202 ;
  assign n204 = x130 &  n203 ;
  assign n205 = ( x131 & n196 ) | ( x131 & n204 ) | ( n196 & n204 ) ;
  assign n206 = n188 | n205 ;
  assign n207 = x132 &  n206 ;
  assign n208 = ( x133 & n171 ) | ( x133 & n207 ) | ( n171 & n207 ) ;
  assign n209 = ( x42 & ~x128 ) | ( x42 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n210 = x41 &  x128 ;
  assign n211 = ( x129 & n209 ) | ( x129 & n210 ) | ( n209 & n210 ) ;
  assign n212 = x43 &  x128 ;
  assign n213 = ( x44 & ~x128 ) | ( x44 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n214 = ( n212 & ~x129 ) | ( n212 & n213 ) | ( ~x129 & n213 ) ;
  assign n215 = n211 | n214 ;
  assign n216 = x130 &  n215 ;
  assign n217 = ( x46 & ~x128 ) | ( x46 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n218 = x45 &  x128 ;
  assign n219 = ( x129 & n217 ) | ( x129 & n218 ) | ( n217 & n218 ) ;
  assign n220 = x47 &  x128 ;
  assign n221 = ( x48 & ~x128 ) | ( x48 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n222 = ( n220 & ~x129 ) | ( n220 & n221 ) | ( ~x129 & n221 ) ;
  assign n223 = n219 | n222 ;
  assign n224 = ~x130 & n223 ;
  assign n225 = ( n216 & ~x131 ) | ( n216 & n224 ) | ( ~x131 & n224 ) ;
  assign n226 = x37 &  x128 ;
  assign n227 = ( x129 & ~n226 ) | ( x129 & 1'b0 ) | ( ~n226 & 1'b0 ) ;
  assign n228 = ( x40 & ~x128 ) | ( x40 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n229 = x129 | n228 ;
  assign n230 = ~n227 & n229 ;
  assign n233 = ( x38 & ~x128 ) | ( x38 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n234 = ( x129 & ~n233 ) | ( x129 & 1'b0 ) | ( ~n233 & 1'b0 ) ;
  assign n231 = x39 &  x128 ;
  assign n232 = x129 | n231 ;
  assign n235 = ( n230 & ~n234 ) | ( n230 & n232 ) | ( ~n234 & n232 ) ;
  assign n236 = ~x130 & n235 ;
  assign n237 = ( x34 & ~x128 ) | ( x34 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n238 = x33 &  x128 ;
  assign n239 = ( x129 & n237 ) | ( x129 & n238 ) | ( n237 & n238 ) ;
  assign n240 = x35 &  x128 ;
  assign n241 = ( x36 & ~x128 ) | ( x36 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n242 = ( n240 & ~x129 ) | ( n240 & n241 ) | ( ~x129 & n241 ) ;
  assign n243 = n239 | n242 ;
  assign n244 = x130 &  n243 ;
  assign n245 = ( x131 & n236 ) | ( x131 & n244 ) | ( n236 & n244 ) ;
  assign n246 = n225 | n245 ;
  assign n247 = x132 &  n246 ;
  assign n248 = ( x58 & ~x128 ) | ( x58 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n249 = x57 &  x128 ;
  assign n250 = ( x129 & n248 ) | ( x129 & n249 ) | ( n248 & n249 ) ;
  assign n251 = x59 &  x128 ;
  assign n252 = ( x60 & ~x128 ) | ( x60 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n253 = ( n251 & ~x129 ) | ( n251 & n252 ) | ( ~x129 & n252 ) ;
  assign n254 = n250 | n253 ;
  assign n255 = x130 &  n254 ;
  assign n256 = ( x62 & ~x128 ) | ( x62 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n257 = x61 &  x128 ;
  assign n258 = ( x129 & n256 ) | ( x129 & n257 ) | ( n256 & n257 ) ;
  assign n259 = x63 &  x128 ;
  assign n260 = ( x64 & ~x128 ) | ( x64 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n261 = ( n259 & ~x129 ) | ( n259 & n260 ) | ( ~x129 & n260 ) ;
  assign n262 = n258 | n261 ;
  assign n263 = ~x130 & n262 ;
  assign n264 = ( n255 & ~x131 ) | ( n255 & n263 ) | ( ~x131 & n263 ) ;
  assign n265 = ( x54 & ~x128 ) | ( x54 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n266 = x53 &  x128 ;
  assign n267 = ( x129 & n265 ) | ( x129 & n266 ) | ( n265 & n266 ) ;
  assign n268 = x55 &  x128 ;
  assign n269 = ( x56 & ~x128 ) | ( x56 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n270 = ( n268 & ~x129 ) | ( n268 & n269 ) | ( ~x129 & n269 ) ;
  assign n271 = n267 | n270 ;
  assign n272 = ~x130 & n271 ;
  assign n273 = ( x50 & ~x128 ) | ( x50 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n274 = x49 &  x128 ;
  assign n275 = ( x129 & n273 ) | ( x129 & n274 ) | ( n273 & n274 ) ;
  assign n276 = x51 &  x128 ;
  assign n277 = ( x52 & ~x128 ) | ( x52 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n278 = ( n276 & ~x129 ) | ( n276 & n277 ) | ( ~x129 & n277 ) ;
  assign n279 = n275 | n278 ;
  assign n280 = x130 &  n279 ;
  assign n281 = ( x131 & n272 ) | ( x131 & n280 ) | ( n272 & n280 ) ;
  assign n282 = n264 | n281 ;
  assign n283 = ~x132 & n282 ;
  assign n284 = ( n247 & ~x133 ) | ( n247 & n283 ) | ( ~x133 & n283 ) ;
  assign n285 = n208 | n284 ;
  assign n286 = x134 &  n285 ;
  assign n287 = ( x90 & ~x128 ) | ( x90 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n288 = x89 &  x128 ;
  assign n289 = ( x129 & n287 ) | ( x129 & n288 ) | ( n287 & n288 ) ;
  assign n290 = x91 &  x128 ;
  assign n291 = ( x92 & ~x128 ) | ( x92 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n292 = ( n290 & ~x129 ) | ( n290 & n291 ) | ( ~x129 & n291 ) ;
  assign n293 = n289 | n292 ;
  assign n294 = x130 &  n293 ;
  assign n295 = ( x94 & ~x128 ) | ( x94 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n296 = x93 &  x128 ;
  assign n297 = ( x129 & n295 ) | ( x129 & n296 ) | ( n295 & n296 ) ;
  assign n298 = x95 &  x128 ;
  assign n299 = ( x96 & ~x128 ) | ( x96 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n300 = ( n298 & ~x129 ) | ( n298 & n299 ) | ( ~x129 & n299 ) ;
  assign n301 = n297 | n300 ;
  assign n302 = ~x130 & n301 ;
  assign n303 = ( n294 & ~x131 ) | ( n294 & n302 ) | ( ~x131 & n302 ) ;
  assign n304 = ( x86 & ~x128 ) | ( x86 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n305 = x85 &  x128 ;
  assign n306 = ( x129 & n304 ) | ( x129 & n305 ) | ( n304 & n305 ) ;
  assign n307 = x87 &  x128 ;
  assign n308 = ( x88 & ~x128 ) | ( x88 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n309 = ( n307 & ~x129 ) | ( n307 & n308 ) | ( ~x129 & n308 ) ;
  assign n310 = n306 | n309 ;
  assign n311 = ~x130 & n310 ;
  assign n312 = ( x82 & ~x128 ) | ( x82 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n313 = x81 &  x128 ;
  assign n314 = ( x129 & n312 ) | ( x129 & n313 ) | ( n312 & n313 ) ;
  assign n315 = x83 &  x128 ;
  assign n316 = ( x84 & ~x128 ) | ( x84 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n317 = ( n315 & ~x129 ) | ( n315 & n316 ) | ( ~x129 & n316 ) ;
  assign n318 = n314 | n317 ;
  assign n319 = x130 &  n318 ;
  assign n320 = ( x131 & n311 ) | ( x131 & n319 ) | ( n311 & n319 ) ;
  assign n321 = n303 | n320 ;
  assign n322 = ~x132 & n321 ;
  assign n323 = ( x74 & ~x128 ) | ( x74 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n324 = x73 &  x128 ;
  assign n325 = ( x129 & n323 ) | ( x129 & n324 ) | ( n323 & n324 ) ;
  assign n326 = x75 &  x128 ;
  assign n327 = ( x76 & ~x128 ) | ( x76 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n328 = ( n326 & ~x129 ) | ( n326 & n327 ) | ( ~x129 & n327 ) ;
  assign n329 = n325 | n328 ;
  assign n330 = x130 &  n329 ;
  assign n331 = ( x78 & ~x128 ) | ( x78 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n332 = x77 &  x128 ;
  assign n333 = ( x129 & n331 ) | ( x129 & n332 ) | ( n331 & n332 ) ;
  assign n334 = x79 &  x128 ;
  assign n335 = ( x80 & ~x128 ) | ( x80 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n336 = ( n334 & ~x129 ) | ( n334 & n335 ) | ( ~x129 & n335 ) ;
  assign n337 = n333 | n336 ;
  assign n338 = ~x130 & n337 ;
  assign n339 = ( n330 & ~x131 ) | ( n330 & n338 ) | ( ~x131 & n338 ) ;
  assign n340 = ( x70 & ~x128 ) | ( x70 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n341 = x69 &  x128 ;
  assign n342 = ( x129 & n340 ) | ( x129 & n341 ) | ( n340 & n341 ) ;
  assign n343 = x71 &  x128 ;
  assign n344 = ( x72 & ~x128 ) | ( x72 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n345 = ( n343 & ~x129 ) | ( n343 & n344 ) | ( ~x129 & n344 ) ;
  assign n346 = n342 | n345 ;
  assign n347 = ~x130 & n346 ;
  assign n348 = ( x66 & ~x128 ) | ( x66 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n349 = x65 &  x128 ;
  assign n350 = ( x129 & n348 ) | ( x129 & n349 ) | ( n348 & n349 ) ;
  assign n351 = x67 &  x128 ;
  assign n352 = ( x68 & ~x128 ) | ( x68 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n353 = ( n351 & ~x129 ) | ( n351 & n352 ) | ( ~x129 & n352 ) ;
  assign n354 = n350 | n353 ;
  assign n355 = x130 &  n354 ;
  assign n356 = ( x131 & n347 ) | ( x131 & n355 ) | ( n347 & n355 ) ;
  assign n357 = n339 | n356 ;
  assign n358 = x132 &  n357 ;
  assign n359 = ( x133 & n322 ) | ( x133 & n358 ) | ( n322 & n358 ) ;
  assign n360 = ( x106 & ~x128 ) | ( x106 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n361 = x105 &  x128 ;
  assign n362 = ( x129 & n360 ) | ( x129 & n361 ) | ( n360 & n361 ) ;
  assign n363 = x107 &  x128 ;
  assign n364 = ( x108 & ~x128 ) | ( x108 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n365 = ( n363 & ~x129 ) | ( n363 & n364 ) | ( ~x129 & n364 ) ;
  assign n366 = n362 | n365 ;
  assign n367 = x130 &  n366 ;
  assign n368 = ( x110 & ~x128 ) | ( x110 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n369 = x109 &  x128 ;
  assign n370 = ( x129 & n368 ) | ( x129 & n369 ) | ( n368 & n369 ) ;
  assign n371 = x111 &  x128 ;
  assign n372 = ( x112 & ~x128 ) | ( x112 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n373 = ( n371 & ~x129 ) | ( n371 & n372 ) | ( ~x129 & n372 ) ;
  assign n374 = n370 | n373 ;
  assign n375 = ~x130 & n374 ;
  assign n376 = ( n367 & ~x131 ) | ( n367 & n375 ) | ( ~x131 & n375 ) ;
  assign n377 = ( x102 & ~x128 ) | ( x102 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n378 = x101 &  x128 ;
  assign n379 = ( x129 & n377 ) | ( x129 & n378 ) | ( n377 & n378 ) ;
  assign n380 = x103 &  x128 ;
  assign n381 = ( x104 & ~x128 ) | ( x104 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n382 = ( n380 & ~x129 ) | ( n380 & n381 ) | ( ~x129 & n381 ) ;
  assign n383 = n379 | n382 ;
  assign n384 = ~x130 & n383 ;
  assign n385 = ( x98 & ~x128 ) | ( x98 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n386 = x97 &  x128 ;
  assign n387 = ( x129 & n385 ) | ( x129 & n386 ) | ( n385 & n386 ) ;
  assign n388 = x99 &  x128 ;
  assign n389 = ( x100 & ~x128 ) | ( x100 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n390 = ( n388 & ~x129 ) | ( n388 & n389 ) | ( ~x129 & n389 ) ;
  assign n391 = n387 | n390 ;
  assign n392 = x130 &  n391 ;
  assign n393 = ( x131 & n384 ) | ( x131 & n392 ) | ( n384 & n392 ) ;
  assign n394 = n376 | n393 ;
  assign n395 = x132 &  n394 ;
  assign n396 = ( x122 & ~x128 ) | ( x122 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n397 = x121 &  x128 ;
  assign n398 = ( x129 & n396 ) | ( x129 & n397 ) | ( n396 & n397 ) ;
  assign n399 = x123 &  x128 ;
  assign n400 = ( x124 & ~x128 ) | ( x124 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n401 = ( n399 & ~x129 ) | ( n399 & n400 ) | ( ~x129 & n400 ) ;
  assign n402 = n398 | n401 ;
  assign n403 = x130 &  n402 ;
  assign n404 = ( x126 & ~x128 ) | ( x126 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n405 = x125 &  x128 ;
  assign n406 = ( x129 & n404 ) | ( x129 & n405 ) | ( n404 & n405 ) ;
  assign n407 = x127 &  x128 ;
  assign n408 = ( x0 & ~x128 ) | ( x0 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n409 = ( n407 & ~x129 ) | ( n407 & n408 ) | ( ~x129 & n408 ) ;
  assign n410 = n406 | n409 ;
  assign n411 = ~x130 & n410 ;
  assign n412 = ( n403 & ~x131 ) | ( n403 & n411 ) | ( ~x131 & n411 ) ;
  assign n413 = ( x118 & ~x128 ) | ( x118 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n414 = x117 &  x128 ;
  assign n415 = ( x129 & n413 ) | ( x129 & n414 ) | ( n413 & n414 ) ;
  assign n416 = x119 &  x128 ;
  assign n417 = ( x120 & ~x128 ) | ( x120 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n418 = ( n416 & ~x129 ) | ( n416 & n417 ) | ( ~x129 & n417 ) ;
  assign n419 = n415 | n418 ;
  assign n420 = ~x130 & n419 ;
  assign n421 = ( x114 & ~x128 ) | ( x114 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n422 = x113 &  x128 ;
  assign n423 = ( x129 & n421 ) | ( x129 & n422 ) | ( n421 & n422 ) ;
  assign n424 = x115 &  x128 ;
  assign n425 = ( x116 & ~x128 ) | ( x116 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n426 = ( n424 & ~x129 ) | ( n424 & n425 ) | ( ~x129 & n425 ) ;
  assign n427 = n423 | n426 ;
  assign n428 = x130 &  n427 ;
  assign n429 = ( x131 & n420 ) | ( x131 & n428 ) | ( n420 & n428 ) ;
  assign n430 = n412 | n429 ;
  assign n431 = ~x132 & n430 ;
  assign n432 = ( n395 & ~x133 ) | ( n395 & n431 ) | ( ~x133 & n431 ) ;
  assign n433 = n359 | n432 ;
  assign n434 = ~x134 & n433 ;
  assign n435 = n286 | n434 ;
  assign n436 = x132 | x133 ;
  assign n437 = x58 &  x128 ;
  assign n438 = ( x129 & ~n437 ) | ( x129 & 1'b0 ) | ( ~n437 & 1'b0 ) ;
  assign n439 = ( x61 & ~x128 ) | ( x61 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n440 = x129 | n439 ;
  assign n441 = ~n438 & n440 ;
  assign n444 = ( x59 & ~x128 ) | ( x59 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n445 = ( x129 & ~n444 ) | ( x129 & 1'b0 ) | ( ~n444 & 1'b0 ) ;
  assign n442 = x60 &  x128 ;
  assign n443 = x129 | n442 ;
  assign n446 = ( n441 & ~n445 ) | ( n441 & n443 ) | ( ~n445 & n443 ) ;
  assign n447 = x130 &  n446 ;
  assign n448 = x62 &  x128 ;
  assign n449 = ( x129 & ~n448 ) | ( x129 & 1'b0 ) | ( ~n448 & 1'b0 ) ;
  assign n450 = ( x65 & ~x128 ) | ( x65 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n451 = x129 | n450 ;
  assign n452 = ~n449 & n451 ;
  assign n455 = ( x63 & ~x128 ) | ( x63 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n456 = ( x129 & ~n455 ) | ( x129 & 1'b0 ) | ( ~n455 & 1'b0 ) ;
  assign n453 = x64 &  x128 ;
  assign n454 = x129 | n453 ;
  assign n457 = ( n452 & ~n456 ) | ( n452 & n454 ) | ( ~n456 & n454 ) ;
  assign n458 = ~x130 & n457 ;
  assign n459 = ( n447 & ~x131 ) | ( n447 & n458 ) | ( ~x131 & n458 ) ;
  assign n460 = x54 &  x128 ;
  assign n461 = ( x129 & ~n460 ) | ( x129 & 1'b0 ) | ( ~n460 & 1'b0 ) ;
  assign n462 = ( x57 & ~x128 ) | ( x57 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n463 = x129 | n462 ;
  assign n464 = ~n461 & n463 ;
  assign n467 = ( x55 & ~x128 ) | ( x55 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n468 = ( x129 & ~n467 ) | ( x129 & 1'b0 ) | ( ~n467 & 1'b0 ) ;
  assign n465 = x56 &  x128 ;
  assign n466 = x129 | n465 ;
  assign n469 = ( n464 & ~n468 ) | ( n464 & n466 ) | ( ~n468 & n466 ) ;
  assign n470 = ~x130 & n469 ;
  assign n471 = x50 &  x128 ;
  assign n472 = ( x129 & ~n471 ) | ( x129 & 1'b0 ) | ( ~n471 & 1'b0 ) ;
  assign n473 = ( x53 & ~x128 ) | ( x53 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n474 = x129 | n473 ;
  assign n475 = ~n472 & n474 ;
  assign n478 = ( x51 & ~x128 ) | ( x51 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n479 = ( x129 & ~n478 ) | ( x129 & 1'b0 ) | ( ~n478 & 1'b0 ) ;
  assign n476 = x52 &  x128 ;
  assign n477 = x129 | n476 ;
  assign n480 = ( n475 & ~n479 ) | ( n475 & n477 ) | ( ~n479 & n477 ) ;
  assign n481 = x130 &  n480 ;
  assign n482 = ( x131 & n470 ) | ( x131 & n481 ) | ( n470 & n481 ) ;
  assign n483 = n459 | n482 ;
  assign n484 = ~n436 & n483 ;
  assign n485 = x132 &  x133 ;
  assign n486 = x10 &  x128 ;
  assign n487 = ( x129 & ~n486 ) | ( x129 & 1'b0 ) | ( ~n486 & 1'b0 ) ;
  assign n488 = ( x13 & ~x128 ) | ( x13 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n489 = x129 | n488 ;
  assign n490 = ~n487 & n489 ;
  assign n493 = ( x11 & ~x128 ) | ( x11 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n494 = ( x129 & ~n493 ) | ( x129 & 1'b0 ) | ( ~n493 & 1'b0 ) ;
  assign n491 = x12 &  x128 ;
  assign n492 = x129 | n491 ;
  assign n495 = ( n490 & ~n494 ) | ( n490 & n492 ) | ( ~n494 & n492 ) ;
  assign n496 = x130 &  n495 ;
  assign n497 = x14 &  x128 ;
  assign n498 = ( x129 & ~n497 ) | ( x129 & 1'b0 ) | ( ~n497 & 1'b0 ) ;
  assign n499 = ( x17 & ~x128 ) | ( x17 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n500 = x129 | n499 ;
  assign n501 = ~n498 & n500 ;
  assign n504 = ( x15 & ~x128 ) | ( x15 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n505 = ( x129 & ~n504 ) | ( x129 & 1'b0 ) | ( ~n504 & 1'b0 ) ;
  assign n502 = x16 &  x128 ;
  assign n503 = x129 | n502 ;
  assign n506 = ( n501 & ~n505 ) | ( n501 & n503 ) | ( ~n505 & n503 ) ;
  assign n507 = ~x130 & n506 ;
  assign n508 = ( n496 & ~x131 ) | ( n496 & n507 ) | ( ~x131 & n507 ) ;
  assign n509 = x6 &  x128 ;
  assign n510 = ( x129 & ~n509 ) | ( x129 & 1'b0 ) | ( ~n509 & 1'b0 ) ;
  assign n511 = ( x9 & ~x128 ) | ( x9 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n512 = x129 | n511 ;
  assign n513 = ~n510 & n512 ;
  assign n516 = ( x7 & ~x128 ) | ( x7 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n517 = ( x129 & ~n516 ) | ( x129 & 1'b0 ) | ( ~n516 & 1'b0 ) ;
  assign n514 = x8 &  x128 ;
  assign n515 = x129 | n514 ;
  assign n518 = ( n513 & ~n517 ) | ( n513 & n515 ) | ( ~n517 & n515 ) ;
  assign n519 = ~x130 & n518 ;
  assign n520 = x2 &  x128 ;
  assign n521 = ( x129 & ~n520 ) | ( x129 & 1'b0 ) | ( ~n520 & 1'b0 ) ;
  assign n522 = ( x5 & ~x128 ) | ( x5 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n523 = x129 | n522 ;
  assign n524 = ~n521 & n523 ;
  assign n527 = ( x3 & ~x128 ) | ( x3 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n528 = ( x129 & ~n527 ) | ( x129 & 1'b0 ) | ( ~n527 & 1'b0 ) ;
  assign n525 = x4 &  x128 ;
  assign n526 = x129 | n525 ;
  assign n529 = ( n524 & ~n528 ) | ( n524 & n526 ) | ( ~n528 & n526 ) ;
  assign n530 = x130 &  n529 ;
  assign n531 = ( x131 & n519 ) | ( x131 & n530 ) | ( n519 & n530 ) ;
  assign n532 = n508 | n531 ;
  assign n533 = n485 &  n532 ;
  assign n534 = n484 | n533 ;
  assign n535 = ~x132 |  x133 ;
  assign n536 = ( x43 & ~x128 ) | ( x43 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n537 = x42 &  x128 ;
  assign n538 = ( x129 & ~n537 ) | ( x129 & n536 ) | ( ~n537 & n536 ) ;
  assign n539 = ~n536 & n538 ;
  assign n540 = x44 &  x128 ;
  assign n541 = ( x45 & ~x128 ) | ( x45 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n542 = ( n540 & ~x129 ) | ( n540 & n541 ) | ( ~x129 & n541 ) ;
  assign n543 = ( x129 & ~n539 ) | ( x129 & n542 ) | ( ~n539 & n542 ) ;
  assign n544 = x130 &  n543 ;
  assign n545 = x46 &  x128 ;
  assign n546 = ( x129 & ~n545 ) | ( x129 & 1'b0 ) | ( ~n545 & 1'b0 ) ;
  assign n547 = ( x49 & ~x128 ) | ( x49 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n548 = x129 | n547 ;
  assign n549 = ~n546 & n548 ;
  assign n552 = ( x47 & ~x128 ) | ( x47 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n553 = ( x129 & ~n552 ) | ( x129 & 1'b0 ) | ( ~n552 & 1'b0 ) ;
  assign n550 = x48 &  x128 ;
  assign n551 = x129 | n550 ;
  assign n554 = ( n549 & ~n553 ) | ( n549 & n551 ) | ( ~n553 & n551 ) ;
  assign n555 = ~x130 & n554 ;
  assign n556 = ( n544 & ~x131 ) | ( n544 & n555 ) | ( ~x131 & n555 ) ;
  assign n557 = ( x39 & ~x128 ) | ( x39 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n558 = x38 &  x128 ;
  assign n559 = ( x129 & ~n558 ) | ( x129 & n557 ) | ( ~n558 & n557 ) ;
  assign n560 = ~n557 & n559 ;
  assign n561 = ( x41 & ~x128 ) | ( x41 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n562 = x40 &  x128 ;
  assign n563 = ( n561 & ~x129 ) | ( n561 & n562 ) | ( ~x129 & n562 ) ;
  assign n564 = ( x129 & ~n560 ) | ( x129 & n563 ) | ( ~n560 & n563 ) ;
  assign n565 = ~x130 & n564 ;
  assign n566 = x34 &  x128 ;
  assign n567 = ( x129 & ~n566 ) | ( x129 & 1'b0 ) | ( ~n566 & 1'b0 ) ;
  assign n568 = ( x37 & ~x128 ) | ( x37 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n569 = x129 | n568 ;
  assign n570 = ~n567 & n569 ;
  assign n573 = ( x35 & ~x128 ) | ( x35 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n574 = ( x129 & ~n573 ) | ( x129 & 1'b0 ) | ( ~n573 & 1'b0 ) ;
  assign n571 = x36 &  x128 ;
  assign n572 = x129 | n571 ;
  assign n575 = ( n570 & ~n574 ) | ( n570 & n572 ) | ( ~n574 & n572 ) ;
  assign n576 = x130 &  n575 ;
  assign n577 = ( x131 & n565 ) | ( x131 & n576 ) | ( n565 & n576 ) ;
  assign n578 = n556 | n577 ;
  assign n579 = ~n535 & n578 ;
  assign n580 = ~x133 |  x132 ;
  assign n581 = x26 &  x128 ;
  assign n582 = ( x129 & ~n581 ) | ( x129 & 1'b0 ) | ( ~n581 & 1'b0 ) ;
  assign n583 = ( x29 & ~x128 ) | ( x29 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n584 = x129 | n583 ;
  assign n585 = ~n582 & n584 ;
  assign n588 = ( x27 & ~x128 ) | ( x27 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n589 = ( x129 & ~n588 ) | ( x129 & 1'b0 ) | ( ~n588 & 1'b0 ) ;
  assign n586 = x28 &  x128 ;
  assign n587 = x129 | n586 ;
  assign n590 = ( n585 & ~n589 ) | ( n585 & n587 ) | ( ~n589 & n587 ) ;
  assign n591 = x130 &  n590 ;
  assign n592 = x30 &  x128 ;
  assign n593 = ( x129 & ~n592 ) | ( x129 & 1'b0 ) | ( ~n592 & 1'b0 ) ;
  assign n594 = ( x33 & ~x128 ) | ( x33 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n595 = x129 | n594 ;
  assign n596 = ~n593 & n595 ;
  assign n599 = ( x31 & ~x128 ) | ( x31 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n600 = ( x129 & ~n599 ) | ( x129 & 1'b0 ) | ( ~n599 & 1'b0 ) ;
  assign n597 = x32 &  x128 ;
  assign n598 = x129 | n597 ;
  assign n601 = ( n596 & ~n600 ) | ( n596 & n598 ) | ( ~n600 & n598 ) ;
  assign n602 = ~x130 & n601 ;
  assign n603 = ( n591 & ~x131 ) | ( n591 & n602 ) | ( ~x131 & n602 ) ;
  assign n604 = x22 &  x128 ;
  assign n605 = ( x129 & ~n604 ) | ( x129 & 1'b0 ) | ( ~n604 & 1'b0 ) ;
  assign n606 = ( x25 & ~x128 ) | ( x25 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n607 = x129 | n606 ;
  assign n608 = ~n605 & n607 ;
  assign n611 = ( x23 & ~x128 ) | ( x23 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n612 = ( x129 & ~n611 ) | ( x129 & 1'b0 ) | ( ~n611 & 1'b0 ) ;
  assign n609 = x24 &  x128 ;
  assign n610 = x129 | n609 ;
  assign n613 = ( n608 & ~n612 ) | ( n608 & n610 ) | ( ~n612 & n610 ) ;
  assign n614 = ~x130 & n613 ;
  assign n615 = x18 &  x128 ;
  assign n616 = ( x129 & ~n615 ) | ( x129 & 1'b0 ) | ( ~n615 & 1'b0 ) ;
  assign n617 = ( x21 & ~x128 ) | ( x21 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n618 = x129 | n617 ;
  assign n619 = ~n616 & n618 ;
  assign n622 = ( x19 & ~x128 ) | ( x19 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n623 = ( x129 & ~n622 ) | ( x129 & 1'b0 ) | ( ~n622 & 1'b0 ) ;
  assign n620 = x20 &  x128 ;
  assign n621 = x129 | n620 ;
  assign n624 = ( n619 & ~n623 ) | ( n619 & n621 ) | ( ~n623 & n621 ) ;
  assign n625 = x130 &  n624 ;
  assign n626 = ( x131 & n614 ) | ( x131 & n625 ) | ( n614 & n625 ) ;
  assign n627 = n603 | n626 ;
  assign n628 = ~n580 & n627 ;
  assign n629 = n579 | n628 ;
  assign n630 = n534 | n629 ;
  assign n631 = x134 &  n630 ;
  assign n632 = x90 &  x128 ;
  assign n633 = ( x129 & ~n632 ) | ( x129 & 1'b0 ) | ( ~n632 & 1'b0 ) ;
  assign n634 = ( x93 & ~x128 ) | ( x93 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n635 = x129 | n634 ;
  assign n636 = ~n633 & n635 ;
  assign n639 = ( x91 & ~x128 ) | ( x91 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n640 = ( x129 & ~n639 ) | ( x129 & 1'b0 ) | ( ~n639 & 1'b0 ) ;
  assign n637 = x92 &  x128 ;
  assign n638 = x129 | n637 ;
  assign n641 = ( n636 & ~n640 ) | ( n636 & n638 ) | ( ~n640 & n638 ) ;
  assign n642 = x130 &  n641 ;
  assign n643 = x94 &  x128 ;
  assign n644 = ( x129 & ~n643 ) | ( x129 & 1'b0 ) | ( ~n643 & 1'b0 ) ;
  assign n645 = ( x97 & ~x128 ) | ( x97 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n646 = x129 | n645 ;
  assign n647 = ~n644 & n646 ;
  assign n650 = ( x95 & ~x128 ) | ( x95 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n651 = ( x129 & ~n650 ) | ( x129 & 1'b0 ) | ( ~n650 & 1'b0 ) ;
  assign n648 = x96 &  x128 ;
  assign n649 = x129 | n648 ;
  assign n652 = ( n647 & ~n651 ) | ( n647 & n649 ) | ( ~n651 & n649 ) ;
  assign n653 = ~x130 & n652 ;
  assign n654 = ( n642 & ~x131 ) | ( n642 & n653 ) | ( ~x131 & n653 ) ;
  assign n655 = x86 &  x128 ;
  assign n656 = ( x129 & ~n655 ) | ( x129 & 1'b0 ) | ( ~n655 & 1'b0 ) ;
  assign n657 = ( x89 & ~x128 ) | ( x89 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n658 = x129 | n657 ;
  assign n659 = ~n656 & n658 ;
  assign n662 = ( x87 & ~x128 ) | ( x87 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n663 = ( x129 & ~n662 ) | ( x129 & 1'b0 ) | ( ~n662 & 1'b0 ) ;
  assign n660 = x88 &  x128 ;
  assign n661 = x129 | n660 ;
  assign n664 = ( n659 & ~n663 ) | ( n659 & n661 ) | ( ~n663 & n661 ) ;
  assign n665 = ~x130 & n664 ;
  assign n666 = x82 &  x128 ;
  assign n667 = ( x129 & ~n666 ) | ( x129 & 1'b0 ) | ( ~n666 & 1'b0 ) ;
  assign n668 = ( x85 & ~x128 ) | ( x85 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n669 = x129 | n668 ;
  assign n670 = ~n667 & n669 ;
  assign n673 = ( x83 & ~x128 ) | ( x83 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n674 = ( x129 & ~n673 ) | ( x129 & 1'b0 ) | ( ~n673 & 1'b0 ) ;
  assign n671 = x84 &  x128 ;
  assign n672 = x129 | n671 ;
  assign n675 = ( n670 & ~n674 ) | ( n670 & n672 ) | ( ~n674 & n672 ) ;
  assign n676 = x130 &  n675 ;
  assign n677 = ( x131 & n665 ) | ( x131 & n676 ) | ( n665 & n676 ) ;
  assign n678 = n654 | n677 ;
  assign n679 = ~x132 & n678 ;
  assign n680 = x74 &  x128 ;
  assign n681 = ( x129 & ~n680 ) | ( x129 & 1'b0 ) | ( ~n680 & 1'b0 ) ;
  assign n682 = ( x77 & ~x128 ) | ( x77 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n683 = x129 | n682 ;
  assign n684 = ~n681 & n683 ;
  assign n687 = ( x75 & ~x128 ) | ( x75 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n688 = ( x129 & ~n687 ) | ( x129 & 1'b0 ) | ( ~n687 & 1'b0 ) ;
  assign n685 = x76 &  x128 ;
  assign n686 = x129 | n685 ;
  assign n689 = ( n684 & ~n688 ) | ( n684 & n686 ) | ( ~n688 & n686 ) ;
  assign n690 = x130 &  n689 ;
  assign n691 = x78 &  x128 ;
  assign n692 = ( x129 & ~n691 ) | ( x129 & 1'b0 ) | ( ~n691 & 1'b0 ) ;
  assign n693 = ( x81 & ~x128 ) | ( x81 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n694 = x129 | n693 ;
  assign n695 = ~n692 & n694 ;
  assign n698 = ( x79 & ~x128 ) | ( x79 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n699 = ( x129 & ~n698 ) | ( x129 & 1'b0 ) | ( ~n698 & 1'b0 ) ;
  assign n696 = x80 &  x128 ;
  assign n697 = x129 | n696 ;
  assign n700 = ( n695 & ~n699 ) | ( n695 & n697 ) | ( ~n699 & n697 ) ;
  assign n701 = ~x130 & n700 ;
  assign n702 = ( n690 & ~x131 ) | ( n690 & n701 ) | ( ~x131 & n701 ) ;
  assign n703 = x70 &  x128 ;
  assign n704 = ( x129 & ~n703 ) | ( x129 & 1'b0 ) | ( ~n703 & 1'b0 ) ;
  assign n705 = ( x73 & ~x128 ) | ( x73 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n706 = x129 | n705 ;
  assign n707 = ~n704 & n706 ;
  assign n710 = ( x71 & ~x128 ) | ( x71 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n711 = ( x129 & ~n710 ) | ( x129 & 1'b0 ) | ( ~n710 & 1'b0 ) ;
  assign n708 = x72 &  x128 ;
  assign n709 = x129 | n708 ;
  assign n712 = ( n707 & ~n711 ) | ( n707 & n709 ) | ( ~n711 & n709 ) ;
  assign n713 = ~x130 & n712 ;
  assign n714 = x66 &  x128 ;
  assign n715 = ( x129 & ~n714 ) | ( x129 & 1'b0 ) | ( ~n714 & 1'b0 ) ;
  assign n716 = ( x69 & ~x128 ) | ( x69 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n717 = x129 | n716 ;
  assign n718 = ~n715 & n717 ;
  assign n721 = ( x67 & ~x128 ) | ( x67 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n722 = ( x129 & ~n721 ) | ( x129 & 1'b0 ) | ( ~n721 & 1'b0 ) ;
  assign n719 = x68 &  x128 ;
  assign n720 = x129 | n719 ;
  assign n723 = ( n718 & ~n722 ) | ( n718 & n720 ) | ( ~n722 & n720 ) ;
  assign n724 = x130 &  n723 ;
  assign n725 = ( x131 & n713 ) | ( x131 & n724 ) | ( n713 & n724 ) ;
  assign n726 = n702 | n725 ;
  assign n727 = x132 &  n726 ;
  assign n728 = ( x133 & n679 ) | ( x133 & n727 ) | ( n679 & n727 ) ;
  assign n729 = x106 &  x128 ;
  assign n730 = ( x129 & ~n729 ) | ( x129 & 1'b0 ) | ( ~n729 & 1'b0 ) ;
  assign n731 = ( x109 & ~x128 ) | ( x109 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n732 = x129 | n731 ;
  assign n733 = ~n730 & n732 ;
  assign n736 = ( x107 & ~x128 ) | ( x107 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n737 = ( x129 & ~n736 ) | ( x129 & 1'b0 ) | ( ~n736 & 1'b0 ) ;
  assign n734 = x108 &  x128 ;
  assign n735 = x129 | n734 ;
  assign n738 = ( n733 & ~n737 ) | ( n733 & n735 ) | ( ~n737 & n735 ) ;
  assign n739 = x130 &  n738 ;
  assign n740 = x110 &  x128 ;
  assign n741 = ( x129 & ~n740 ) | ( x129 & 1'b0 ) | ( ~n740 & 1'b0 ) ;
  assign n742 = ( x113 & ~x128 ) | ( x113 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n743 = x129 | n742 ;
  assign n744 = ~n741 & n743 ;
  assign n747 = ( x111 & ~x128 ) | ( x111 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n748 = ( x129 & ~n747 ) | ( x129 & 1'b0 ) | ( ~n747 & 1'b0 ) ;
  assign n745 = x112 &  x128 ;
  assign n746 = x129 | n745 ;
  assign n749 = ( n744 & ~n748 ) | ( n744 & n746 ) | ( ~n748 & n746 ) ;
  assign n750 = ~x130 & n749 ;
  assign n751 = ( n739 & ~x131 ) | ( n739 & n750 ) | ( ~x131 & n750 ) ;
  assign n752 = x102 &  x128 ;
  assign n753 = ( x129 & ~n752 ) | ( x129 & 1'b0 ) | ( ~n752 & 1'b0 ) ;
  assign n754 = ( x105 & ~x128 ) | ( x105 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n755 = x129 | n754 ;
  assign n756 = ~n753 & n755 ;
  assign n759 = ( x103 & ~x128 ) | ( x103 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n760 = ( x129 & ~n759 ) | ( x129 & 1'b0 ) | ( ~n759 & 1'b0 ) ;
  assign n757 = x104 &  x128 ;
  assign n758 = x129 | n757 ;
  assign n761 = ( n756 & ~n760 ) | ( n756 & n758 ) | ( ~n760 & n758 ) ;
  assign n762 = ~x130 & n761 ;
  assign n763 = x98 &  x128 ;
  assign n764 = ( x129 & ~n763 ) | ( x129 & 1'b0 ) | ( ~n763 & 1'b0 ) ;
  assign n765 = ( x101 & ~x128 ) | ( x101 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n766 = x129 | n765 ;
  assign n767 = ~n764 & n766 ;
  assign n770 = ( x99 & ~x128 ) | ( x99 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n771 = ( x129 & ~n770 ) | ( x129 & 1'b0 ) | ( ~n770 & 1'b0 ) ;
  assign n768 = x100 &  x128 ;
  assign n769 = x129 | n768 ;
  assign n772 = ( n767 & ~n771 ) | ( n767 & n769 ) | ( ~n771 & n769 ) ;
  assign n773 = x130 &  n772 ;
  assign n774 = ( x131 & n762 ) | ( x131 & n773 ) | ( n762 & n773 ) ;
  assign n775 = n751 | n774 ;
  assign n776 = x132 &  n775 ;
  assign n777 = x122 &  x128 ;
  assign n778 = ( x129 & ~n777 ) | ( x129 & 1'b0 ) | ( ~n777 & 1'b0 ) ;
  assign n779 = ( x125 & ~x128 ) | ( x125 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n780 = x129 | n779 ;
  assign n781 = ~n778 & n780 ;
  assign n784 = ( x123 & ~x128 ) | ( x123 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n785 = ( x129 & ~n784 ) | ( x129 & 1'b0 ) | ( ~n784 & 1'b0 ) ;
  assign n782 = x124 &  x128 ;
  assign n783 = x129 | n782 ;
  assign n786 = ( n781 & ~n785 ) | ( n781 & n783 ) | ( ~n785 & n783 ) ;
  assign n787 = x130 &  n786 ;
  assign n788 = x126 &  x128 ;
  assign n789 = ( x129 & ~n788 ) | ( x129 & 1'b0 ) | ( ~n788 & 1'b0 ) ;
  assign n790 = ( x1 & ~x128 ) | ( x1 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n791 = x129 | n790 ;
  assign n792 = ~n789 & n791 ;
  assign n795 = ( x127 & ~x128 ) | ( x127 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n796 = ( x129 & ~n795 ) | ( x129 & 1'b0 ) | ( ~n795 & 1'b0 ) ;
  assign n793 = x0 &  x128 ;
  assign n794 = x129 | n793 ;
  assign n797 = ( n792 & ~n796 ) | ( n792 & n794 ) | ( ~n796 & n794 ) ;
  assign n798 = ~x130 & n797 ;
  assign n799 = ( n787 & ~x131 ) | ( n787 & n798 ) | ( ~x131 & n798 ) ;
  assign n800 = x118 &  x128 ;
  assign n801 = ( x129 & ~n800 ) | ( x129 & 1'b0 ) | ( ~n800 & 1'b0 ) ;
  assign n802 = ( x121 & ~x128 ) | ( x121 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n803 = x129 | n802 ;
  assign n804 = ~n801 & n803 ;
  assign n807 = ( x119 & ~x128 ) | ( x119 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n808 = ( x129 & ~n807 ) | ( x129 & 1'b0 ) | ( ~n807 & 1'b0 ) ;
  assign n805 = x120 &  x128 ;
  assign n806 = x129 | n805 ;
  assign n809 = ( n804 & ~n808 ) | ( n804 & n806 ) | ( ~n808 & n806 ) ;
  assign n810 = ~x130 & n809 ;
  assign n811 = x114 &  x128 ;
  assign n812 = ( x129 & ~n811 ) | ( x129 & 1'b0 ) | ( ~n811 & 1'b0 ) ;
  assign n813 = ( x117 & ~x128 ) | ( x117 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n814 = x129 | n813 ;
  assign n815 = ~n812 & n814 ;
  assign n818 = ( x115 & ~x128 ) | ( x115 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n819 = ( x129 & ~n818 ) | ( x129 & 1'b0 ) | ( ~n818 & 1'b0 ) ;
  assign n816 = x116 &  x128 ;
  assign n817 = x129 | n816 ;
  assign n820 = ( n815 & ~n819 ) | ( n815 & n817 ) | ( ~n819 & n817 ) ;
  assign n821 = x130 &  n820 ;
  assign n822 = ( x131 & n810 ) | ( x131 & n821 ) | ( n810 & n821 ) ;
  assign n823 = n799 | n822 ;
  assign n824 = ~x132 & n823 ;
  assign n825 = ( n776 & ~x133 ) | ( n776 & n824 ) | ( ~x133 & n824 ) ;
  assign n826 = n728 | n825 ;
  assign n827 = ~x134 & n826 ;
  assign n828 = n631 | n827 ;
  assign n829 = ( n256 & ~x129 ) | ( n256 & n257 ) | ( ~x129 & n257 ) ;
  assign n830 = ( x129 & n251 ) | ( x129 & n252 ) | ( n251 & n252 ) ;
  assign n831 = n829 | n830 ;
  assign n832 = x130 &  n831 ;
  assign n833 = ( n348 & ~x129 ) | ( n348 & n349 ) | ( ~x129 & n349 ) ;
  assign n834 = ( x129 & n259 ) | ( x129 & n260 ) | ( n259 & n260 ) ;
  assign n835 = n833 | n834 ;
  assign n836 = ~x130 & n835 ;
  assign n837 = ( n832 & ~x131 ) | ( n832 & n836 ) | ( ~x131 & n836 ) ;
  assign n838 = ( n248 & ~x129 ) | ( n248 & n249 ) | ( ~x129 & n249 ) ;
  assign n839 = ( x129 & n268 ) | ( x129 & n269 ) | ( n268 & n269 ) ;
  assign n840 = n838 | n839 ;
  assign n841 = ~x130 & n840 ;
  assign n842 = ( n265 & ~x129 ) | ( n265 & n266 ) | ( ~x129 & n266 ) ;
  assign n843 = ( x129 & n276 ) | ( x129 & n277 ) | ( n276 & n277 ) ;
  assign n844 = n842 | n843 ;
  assign n845 = x130 &  n844 ;
  assign n846 = ( x131 & n841 ) | ( x131 & n845 ) | ( n841 & n845 ) ;
  assign n847 = n837 | n846 ;
  assign n848 = ~n436 & n847 ;
  assign n849 = ( n180 & ~x129 ) | ( n180 & n181 ) | ( ~x129 & n181 ) ;
  assign n850 = ( x129 & n175 ) | ( x129 & n176 ) | ( n175 & n176 ) ;
  assign n851 = n849 | n850 ;
  assign n852 = x130 &  n851 ;
  assign n853 = ( n161 & ~x129 ) | ( n161 & n162 ) | ( ~x129 & n162 ) ;
  assign n854 = ( x129 & n183 ) | ( x129 & n184 ) | ( n183 & n184 ) ;
  assign n855 = n853 | n854 ;
  assign n856 = ~x130 & n855 ;
  assign n857 = ( n852 & ~x131 ) | ( n852 & n856 ) | ( ~x131 & n856 ) ;
  assign n858 = ( n172 & ~x129 ) | ( n172 & n173 ) | ( ~x129 & n173 ) ;
  assign n859 = ( x129 & n192 ) | ( x129 & n193 ) | ( n192 & n193 ) ;
  assign n860 = n858 | n859 ;
  assign n861 = ~x130 & n860 ;
  assign n862 = ( n189 & ~x129 ) | ( n189 & n190 ) | ( ~x129 & n190 ) ;
  assign n863 = ( x129 & n200 ) | ( x129 & n201 ) | ( n200 & n201 ) ;
  assign n864 = n862 | n863 ;
  assign n865 = x130 &  n864 ;
  assign n866 = ( x131 & n861 ) | ( x131 & n865 ) | ( n861 & n865 ) ;
  assign n867 = n857 | n866 ;
  assign n868 = n485 &  n867 ;
  assign n869 = n848 | n868 ;
  assign n870 = ( x129 & n212 ) | ( x129 & n213 ) | ( n212 & n213 ) ;
  assign n871 = ( n217 & ~x129 ) | ( n217 & n218 ) | ( ~x129 & n218 ) ;
  assign n872 = n870 | n871 ;
  assign n873 = x130 &  n872 ;
  assign n874 = ( n273 & ~x129 ) | ( n273 & n274 ) | ( ~x129 & n274 ) ;
  assign n875 = ( x129 & n220 ) | ( x129 & n221 ) | ( n220 & n221 ) ;
  assign n876 = n874 | n875 ;
  assign n877 = ~x130 & n876 ;
  assign n878 = ( n873 & ~x131 ) | ( n873 & n877 ) | ( ~x131 & n877 ) ;
  assign n879 = ( n209 & ~x129 ) | ( n209 & n210 ) | ( ~x129 & n210 ) ;
  assign n880 = ( x129 & n228 ) | ( x129 & n231 ) | ( n228 & n231 ) ;
  assign n881 = n879 | n880 ;
  assign n882 = ~x130 & n881 ;
  assign n883 = ( n226 & ~x129 ) | ( n226 & n233 ) | ( ~x129 & n233 ) ;
  assign n884 = ( x129 & n240 ) | ( x129 & n241 ) | ( n240 & n241 ) ;
  assign n885 = n883 | n884 ;
  assign n886 = x130 &  n885 ;
  assign n887 = ( x131 & n882 ) | ( x131 & n886 ) | ( n882 & n886 ) ;
  assign n888 = n878 | n887 ;
  assign n889 = ~n535 & n888 ;
  assign n890 = ( n144 & ~x129 ) | ( n144 & n145 ) | ( ~x129 & n145 ) ;
  assign n891 = ( x129 & n139 ) | ( x129 & n140 ) | ( n139 & n140 ) ;
  assign n892 = n890 | n891 ;
  assign n893 = x130 &  n892 ;
  assign n894 = ( n237 & ~x129 ) | ( n237 & n238 ) | ( ~x129 & n238 ) ;
  assign n895 = ( x129 & n147 ) | ( x129 & n148 ) | ( n147 & n148 ) ;
  assign n896 = n894 | n895 ;
  assign n897 = ~x130 & n896 ;
  assign n898 = ( n893 & ~x131 ) | ( n893 & n897 ) | ( ~x131 & n897 ) ;
  assign n899 = ( n136 & ~x129 ) | ( n136 & n137 ) | ( ~x129 & n137 ) ;
  assign n900 = ( x129 & n156 ) | ( x129 & n157 ) | ( n156 & n157 ) ;
  assign n901 = n899 | n900 ;
  assign n902 = ~x130 & n901 ;
  assign n903 = ( n153 & ~x129 ) | ( n153 & n154 ) | ( ~x129 & n154 ) ;
  assign n904 = ( x129 & n164 ) | ( x129 & n165 ) | ( n164 & n165 ) ;
  assign n905 = n903 | n904 ;
  assign n906 = x130 &  n905 ;
  assign n907 = ( x131 & n902 ) | ( x131 & n906 ) | ( n902 & n906 ) ;
  assign n908 = n898 | n907 ;
  assign n909 = ~n580 & n908 ;
  assign n910 = n889 | n909 ;
  assign n911 = n869 | n910 ;
  assign n912 = x134 &  n911 ;
  assign n913 = ( n295 & ~x129 ) | ( n295 & n296 ) | ( ~x129 & n296 ) ;
  assign n914 = ( x129 & n290 ) | ( x129 & n291 ) | ( n290 & n291 ) ;
  assign n915 = n913 | n914 ;
  assign n916 = x130 &  n915 ;
  assign n917 = ( n385 & ~x129 ) | ( n385 & n386 ) | ( ~x129 & n386 ) ;
  assign n918 = ( x129 & n298 ) | ( x129 & n299 ) | ( n298 & n299 ) ;
  assign n919 = n917 | n918 ;
  assign n920 = ~x130 & n919 ;
  assign n921 = ( n916 & ~x131 ) | ( n916 & n920 ) | ( ~x131 & n920 ) ;
  assign n922 = ( n287 & ~x129 ) | ( n287 & n288 ) | ( ~x129 & n288 ) ;
  assign n923 = ( x129 & n307 ) | ( x129 & n308 ) | ( n307 & n308 ) ;
  assign n924 = n922 | n923 ;
  assign n925 = ~x130 & n924 ;
  assign n926 = ( n304 & ~x129 ) | ( n304 & n305 ) | ( ~x129 & n305 ) ;
  assign n927 = ( x129 & n315 ) | ( x129 & n316 ) | ( n315 & n316 ) ;
  assign n928 = n926 | n927 ;
  assign n929 = x130 &  n928 ;
  assign n930 = ( x131 & n925 ) | ( x131 & n929 ) | ( n925 & n929 ) ;
  assign n931 = n921 | n930 ;
  assign n932 = ~x132 & n931 ;
  assign n933 = ( n331 & ~x129 ) | ( n331 & n332 ) | ( ~x129 & n332 ) ;
  assign n934 = ( x129 & n326 ) | ( x129 & n327 ) | ( n326 & n327 ) ;
  assign n935 = n933 | n934 ;
  assign n936 = x130 &  n935 ;
  assign n937 = ( n312 & ~x129 ) | ( n312 & n313 ) | ( ~x129 & n313 ) ;
  assign n938 = ( x129 & n334 ) | ( x129 & n335 ) | ( n334 & n335 ) ;
  assign n939 = n937 | n938 ;
  assign n940 = ~x130 & n939 ;
  assign n941 = ( n936 & ~x131 ) | ( n936 & n940 ) | ( ~x131 & n940 ) ;
  assign n942 = ( n323 & ~x129 ) | ( n323 & n324 ) | ( ~x129 & n324 ) ;
  assign n943 = ( x129 & n343 ) | ( x129 & n344 ) | ( n343 & n344 ) ;
  assign n944 = n942 | n943 ;
  assign n945 = ~x130 & n944 ;
  assign n946 = ( n340 & ~x129 ) | ( n340 & n341 ) | ( ~x129 & n341 ) ;
  assign n947 = ( x129 & n351 ) | ( x129 & n352 ) | ( n351 & n352 ) ;
  assign n948 = n946 | n947 ;
  assign n949 = x130 &  n948 ;
  assign n950 = ( x131 & n945 ) | ( x131 & n949 ) | ( n945 & n949 ) ;
  assign n951 = n941 | n950 ;
  assign n952 = x132 &  n951 ;
  assign n953 = ( x133 & n932 ) | ( x133 & n952 ) | ( n932 & n952 ) ;
  assign n954 = ( n368 & ~x129 ) | ( n368 & n369 ) | ( ~x129 & n369 ) ;
  assign n955 = ( x129 & n363 ) | ( x129 & n364 ) | ( n363 & n364 ) ;
  assign n956 = n954 | n955 ;
  assign n957 = x130 &  n956 ;
  assign n958 = ( n421 & ~x129 ) | ( n421 & n422 ) | ( ~x129 & n422 ) ;
  assign n959 = ( x129 & n371 ) | ( x129 & n372 ) | ( n371 & n372 ) ;
  assign n960 = n958 | n959 ;
  assign n961 = ~x130 & n960 ;
  assign n962 = ( n957 & ~x131 ) | ( n957 & n961 ) | ( ~x131 & n961 ) ;
  assign n963 = ( n360 & ~x129 ) | ( n360 & n361 ) | ( ~x129 & n361 ) ;
  assign n964 = ( x129 & n380 ) | ( x129 & n381 ) | ( n380 & n381 ) ;
  assign n965 = n963 | n964 ;
  assign n966 = ~x130 & n965 ;
  assign n967 = ( n377 & ~x129 ) | ( n377 & n378 ) | ( ~x129 & n378 ) ;
  assign n968 = ( x129 & n388 ) | ( x129 & n389 ) | ( n388 & n389 ) ;
  assign n969 = n967 | n968 ;
  assign n970 = x130 &  n969 ;
  assign n971 = ( x131 & n966 ) | ( x131 & n970 ) | ( n966 & n970 ) ;
  assign n972 = n962 | n971 ;
  assign n973 = x132 &  n972 ;
  assign n974 = ( n404 & ~x129 ) | ( n404 & n405 ) | ( ~x129 & n405 ) ;
  assign n975 = ( x129 & n399 ) | ( x129 & n400 ) | ( n399 & n400 ) ;
  assign n976 = n974 | n975 ;
  assign n977 = x130 &  n976 ;
  assign n978 = ( n197 & ~x129 ) | ( n197 & n198 ) | ( ~x129 & n198 ) ;
  assign n979 = ( x129 & n407 ) | ( x129 & n408 ) | ( n407 & n408 ) ;
  assign n980 = n978 | n979 ;
  assign n981 = ~x130 & n980 ;
  assign n982 = ( n977 & ~x131 ) | ( n977 & n981 ) | ( ~x131 & n981 ) ;
  assign n983 = ( n396 & ~x129 ) | ( n396 & n397 ) | ( ~x129 & n397 ) ;
  assign n984 = ( x129 & n416 ) | ( x129 & n417 ) | ( n416 & n417 ) ;
  assign n985 = n983 | n984 ;
  assign n986 = ~x130 & n985 ;
  assign n987 = ( n413 & ~x129 ) | ( n413 & n414 ) | ( ~x129 & n414 ) ;
  assign n988 = ( x129 & n424 ) | ( x129 & n425 ) | ( n424 & n425 ) ;
  assign n989 = n987 | n988 ;
  assign n990 = x130 &  n989 ;
  assign n991 = ( x131 & n986 ) | ( x131 & n990 ) | ( n986 & n990 ) ;
  assign n992 = n982 | n991 ;
  assign n993 = ~x132 & n992 ;
  assign n994 = ( n973 & ~x133 ) | ( n973 & n993 ) | ( ~x133 & n993 ) ;
  assign n995 = n953 | n994 ;
  assign n996 = ~x134 & n995 ;
  assign n997 = n912 | n996 ;
  assign n998 = ( x129 & n540 ) | ( x129 & n541 ) | ( n540 & n541 ) ;
  assign n999 = ( n545 & ~x129 ) | ( n545 & n552 ) | ( ~x129 & n552 ) ;
  assign n1000 = n998 | n999 ;
  assign n1001 = x130 &  n1000 ;
  assign n1002 = x129 &  n547 ;
  assign n1003 = ~x129 & n471 ;
  assign n1004 = n1002 | n1003 ;
  assign n1006 = ( x129 & ~n550 ) | ( x129 & 1'b0 ) | ( ~n550 & 1'b0 ) ;
  assign n1005 = x129 | n478 ;
  assign n1007 = ( n1004 & ~n1006 ) | ( n1004 & n1005 ) | ( ~n1006 & n1005 ) ;
  assign n1008 = ~x130 & n1007 ;
  assign n1009 = ( n1001 & ~x131 ) | ( n1001 & n1008 ) | ( ~x131 & n1008 ) ;
  assign n1010 = x129 &  n561 ;
  assign n1011 = ~x129 & n537 ;
  assign n1012 = n1010 | n1011 ;
  assign n1014 = ( x129 & ~n562 ) | ( x129 & 1'b0 ) | ( ~n562 & 1'b0 ) ;
  assign n1013 = x129 | n536 ;
  assign n1015 = ( n1012 & ~n1014 ) | ( n1012 & n1013 ) | ( ~n1014 & n1013 ) ;
  assign n1016 = ~x130 & n1015 ;
  assign n1017 = x129 &  n568 ;
  assign n1018 = ~x129 & n558 ;
  assign n1019 = n1017 | n1018 ;
  assign n1021 = ( x129 & ~n571 ) | ( x129 & 1'b0 ) | ( ~n571 & 1'b0 ) ;
  assign n1020 = x129 | n557 ;
  assign n1022 = ( n1019 & ~n1021 ) | ( n1019 & n1020 ) | ( ~n1021 & n1020 ) ;
  assign n1023 = x130 &  n1022 ;
  assign n1024 = ( x131 & n1016 ) | ( x131 & n1023 ) | ( n1016 & n1023 ) ;
  assign n1025 = n1009 | n1024 ;
  assign n1026 = x132 &  n1025 ;
  assign n1027 = x129 &  n439 ;
  assign n1028 = ~x129 & n448 ;
  assign n1029 = n1027 | n1028 ;
  assign n1031 = ( x129 & ~n442 ) | ( x129 & 1'b0 ) | ( ~n442 & 1'b0 ) ;
  assign n1030 = x129 | n455 ;
  assign n1032 = ( n1029 & ~n1031 ) | ( n1029 & n1030 ) | ( ~n1031 & n1030 ) ;
  assign n1033 = x130 &  n1032 ;
  assign n1034 = x129 &  n450 ;
  assign n1035 = ~x129 & n714 ;
  assign n1036 = n1034 | n1035 ;
  assign n1038 = ( x129 & ~n453 ) | ( x129 & 1'b0 ) | ( ~n453 & 1'b0 ) ;
  assign n1037 = x129 | n721 ;
  assign n1039 = ( n1036 & ~n1038 ) | ( n1036 & n1037 ) | ( ~n1038 & n1037 ) ;
  assign n1040 = ~x130 & n1039 ;
  assign n1041 = ( n1033 & ~x131 ) | ( n1033 & n1040 ) | ( ~x131 & n1040 ) ;
  assign n1042 = x129 &  n462 ;
  assign n1043 = ~x129 & n437 ;
  assign n1044 = n1042 | n1043 ;
  assign n1046 = ( x129 & ~n465 ) | ( x129 & 1'b0 ) | ( ~n465 & 1'b0 ) ;
  assign n1045 = x129 | n444 ;
  assign n1047 = ( n1044 & ~n1046 ) | ( n1044 & n1045 ) | ( ~n1046 & n1045 ) ;
  assign n1048 = ~x130 & n1047 ;
  assign n1049 = x129 &  n473 ;
  assign n1050 = ~x129 & n460 ;
  assign n1051 = n1049 | n1050 ;
  assign n1053 = ( x129 & ~n476 ) | ( x129 & 1'b0 ) | ( ~n476 & 1'b0 ) ;
  assign n1052 = x129 | n467 ;
  assign n1054 = ( n1051 & ~n1053 ) | ( n1051 & n1052 ) | ( ~n1053 & n1052 ) ;
  assign n1055 = x130 &  n1054 ;
  assign n1056 = ( x131 & n1048 ) | ( x131 & n1055 ) | ( n1048 & n1055 ) ;
  assign n1057 = n1041 | n1056 ;
  assign n1058 = ~x132 & n1057 ;
  assign n1059 = ( n1026 & ~x133 ) | ( n1026 & n1058 ) | ( ~x133 & n1058 ) ;
  assign n1060 = x129 &  n583 ;
  assign n1061 = ~x129 & n592 ;
  assign n1062 = n1060 | n1061 ;
  assign n1064 = ( x129 & ~n586 ) | ( x129 & 1'b0 ) | ( ~n586 & 1'b0 ) ;
  assign n1063 = x129 | n599 ;
  assign n1065 = ( n1062 & ~n1064 ) | ( n1062 & n1063 ) | ( ~n1064 & n1063 ) ;
  assign n1066 = x130 &  n1065 ;
  assign n1067 = x129 &  n594 ;
  assign n1068 = ~x129 & n566 ;
  assign n1069 = n1067 | n1068 ;
  assign n1071 = ( x129 & ~n597 ) | ( x129 & 1'b0 ) | ( ~n597 & 1'b0 ) ;
  assign n1070 = x129 | n573 ;
  assign n1072 = ( n1069 & ~n1071 ) | ( n1069 & n1070 ) | ( ~n1071 & n1070 ) ;
  assign n1073 = ~x130 & n1072 ;
  assign n1074 = ( n1066 & ~x131 ) | ( n1066 & n1073 ) | ( ~x131 & n1073 ) ;
  assign n1075 = x129 &  n606 ;
  assign n1076 = ~x129 & n581 ;
  assign n1077 = n1075 | n1076 ;
  assign n1079 = ( x129 & ~n609 ) | ( x129 & 1'b0 ) | ( ~n609 & 1'b0 ) ;
  assign n1078 = x129 | n588 ;
  assign n1080 = ( n1077 & ~n1079 ) | ( n1077 & n1078 ) | ( ~n1079 & n1078 ) ;
  assign n1081 = ~x130 & n1080 ;
  assign n1082 = x129 &  n617 ;
  assign n1083 = ~x129 & n604 ;
  assign n1084 = n1082 | n1083 ;
  assign n1086 = ( x129 & ~n620 ) | ( x129 & 1'b0 ) | ( ~n620 & 1'b0 ) ;
  assign n1085 = x129 | n611 ;
  assign n1087 = ( n1084 & ~n1086 ) | ( n1084 & n1085 ) | ( ~n1086 & n1085 ) ;
  assign n1088 = x130 &  n1087 ;
  assign n1089 = ( x131 & n1081 ) | ( x131 & n1088 ) | ( n1081 & n1088 ) ;
  assign n1090 = n1074 | n1089 ;
  assign n1091 = ~x132 & n1090 ;
  assign n1092 = x129 &  n488 ;
  assign n1093 = ~x129 & n497 ;
  assign n1094 = n1092 | n1093 ;
  assign n1096 = ( x129 & ~n491 ) | ( x129 & 1'b0 ) | ( ~n491 & 1'b0 ) ;
  assign n1095 = x129 | n504 ;
  assign n1097 = ( n1094 & ~n1096 ) | ( n1094 & n1095 ) | ( ~n1096 & n1095 ) ;
  assign n1098 = x130 &  n1097 ;
  assign n1099 = x129 &  n499 ;
  assign n1100 = ~x129 & n615 ;
  assign n1101 = n1099 | n1100 ;
  assign n1103 = ( x129 & ~n502 ) | ( x129 & 1'b0 ) | ( ~n502 & 1'b0 ) ;
  assign n1102 = x129 | n622 ;
  assign n1104 = ( n1101 & ~n1103 ) | ( n1101 & n1102 ) | ( ~n1103 & n1102 ) ;
  assign n1105 = ~x130 & n1104 ;
  assign n1106 = ( n1098 & ~x131 ) | ( n1098 & n1105 ) | ( ~x131 & n1105 ) ;
  assign n1107 = x129 &  n511 ;
  assign n1108 = ~x129 & n486 ;
  assign n1109 = n1107 | n1108 ;
  assign n1111 = ( x129 & ~n514 ) | ( x129 & 1'b0 ) | ( ~n514 & 1'b0 ) ;
  assign n1110 = x129 | n493 ;
  assign n1112 = ( n1109 & ~n1111 ) | ( n1109 & n1110 ) | ( ~n1111 & n1110 ) ;
  assign n1113 = ~x130 & n1112 ;
  assign n1114 = x129 &  n522 ;
  assign n1115 = ~x129 & n509 ;
  assign n1116 = n1114 | n1115 ;
  assign n1118 = ( x129 & ~n525 ) | ( x129 & 1'b0 ) | ( ~n525 & 1'b0 ) ;
  assign n1117 = x129 | n516 ;
  assign n1119 = ( n1116 & ~n1118 ) | ( n1116 & n1117 ) | ( ~n1118 & n1117 ) ;
  assign n1120 = x130 &  n1119 ;
  assign n1121 = ( x131 & n1113 ) | ( x131 & n1120 ) | ( n1113 & n1120 ) ;
  assign n1122 = n1106 | n1121 ;
  assign n1123 = x132 &  n1122 ;
  assign n1124 = ( x133 & n1091 ) | ( x133 & n1123 ) | ( n1091 & n1123 ) ;
  assign n1125 = n1059 | n1124 ;
  assign n1126 = x134 &  n1125 ;
  assign n1127 = x129 &  n731 ;
  assign n1128 = ~x129 & n740 ;
  assign n1129 = n1127 | n1128 ;
  assign n1131 = ( x129 & ~n734 ) | ( x129 & 1'b0 ) | ( ~n734 & 1'b0 ) ;
  assign n1130 = x129 | n747 ;
  assign n1132 = ( n1129 & ~n1131 ) | ( n1129 & n1130 ) | ( ~n1131 & n1130 ) ;
  assign n1133 = x130 &  n1132 ;
  assign n1134 = x129 &  n742 ;
  assign n1135 = ~x129 & n811 ;
  assign n1136 = n1134 | n1135 ;
  assign n1138 = ( x129 & ~n745 ) | ( x129 & 1'b0 ) | ( ~n745 & 1'b0 ) ;
  assign n1137 = x129 | n818 ;
  assign n1139 = ( n1136 & ~n1138 ) | ( n1136 & n1137 ) | ( ~n1138 & n1137 ) ;
  assign n1140 = ~x130 & n1139 ;
  assign n1141 = ( n1133 & ~x131 ) | ( n1133 & n1140 ) | ( ~x131 & n1140 ) ;
  assign n1142 = x129 &  n754 ;
  assign n1143 = ~x129 & n729 ;
  assign n1144 = n1142 | n1143 ;
  assign n1146 = ( x129 & ~n757 ) | ( x129 & 1'b0 ) | ( ~n757 & 1'b0 ) ;
  assign n1145 = x129 | n736 ;
  assign n1147 = ( n1144 & ~n1146 ) | ( n1144 & n1145 ) | ( ~n1146 & n1145 ) ;
  assign n1148 = ~x130 & n1147 ;
  assign n1149 = x129 &  n765 ;
  assign n1150 = ~x129 & n752 ;
  assign n1151 = n1149 | n1150 ;
  assign n1153 = ( x129 & ~n768 ) | ( x129 & 1'b0 ) | ( ~n768 & 1'b0 ) ;
  assign n1152 = x129 | n759 ;
  assign n1154 = ( n1151 & ~n1153 ) | ( n1151 & n1152 ) | ( ~n1153 & n1152 ) ;
  assign n1155 = x130 &  n1154 ;
  assign n1156 = ( x131 & n1148 ) | ( x131 & n1155 ) | ( n1148 & n1155 ) ;
  assign n1157 = n1141 | n1156 ;
  assign n1158 = ~n535 & n1157 ;
  assign n1159 = x129 &  n634 ;
  assign n1160 = ~x129 & n643 ;
  assign n1161 = n1159 | n1160 ;
  assign n1163 = ( x129 & ~n637 ) | ( x129 & 1'b0 ) | ( ~n637 & 1'b0 ) ;
  assign n1162 = x129 | n650 ;
  assign n1164 = ( n1161 & ~n1163 ) | ( n1161 & n1162 ) | ( ~n1163 & n1162 ) ;
  assign n1165 = x130 &  n1164 ;
  assign n1166 = x129 &  n645 ;
  assign n1167 = ~x129 & n763 ;
  assign n1168 = n1166 | n1167 ;
  assign n1170 = ( x129 & ~n648 ) | ( x129 & 1'b0 ) | ( ~n648 & 1'b0 ) ;
  assign n1169 = x129 | n770 ;
  assign n1171 = ( n1168 & ~n1170 ) | ( n1168 & n1169 ) | ( ~n1170 & n1169 ) ;
  assign n1172 = ~x130 & n1171 ;
  assign n1173 = ( n1165 & ~x131 ) | ( n1165 & n1172 ) | ( ~x131 & n1172 ) ;
  assign n1174 = x129 &  n657 ;
  assign n1175 = ~x129 & n632 ;
  assign n1176 = n1174 | n1175 ;
  assign n1178 = ( x129 & ~n660 ) | ( x129 & 1'b0 ) | ( ~n660 & 1'b0 ) ;
  assign n1177 = x129 | n639 ;
  assign n1179 = ( n1176 & ~n1178 ) | ( n1176 & n1177 ) | ( ~n1178 & n1177 ) ;
  assign n1180 = ~x130 & n1179 ;
  assign n1181 = x129 &  n668 ;
  assign n1182 = ~x129 & n655 ;
  assign n1183 = n1181 | n1182 ;
  assign n1185 = ( x129 & ~n671 ) | ( x129 & 1'b0 ) | ( ~n671 & 1'b0 ) ;
  assign n1184 = x129 | n662 ;
  assign n1186 = ( n1183 & ~n1185 ) | ( n1183 & n1184 ) | ( ~n1185 & n1184 ) ;
  assign n1187 = x130 &  n1186 ;
  assign n1188 = ( x131 & n1180 ) | ( x131 & n1187 ) | ( n1180 & n1187 ) ;
  assign n1189 = n1173 | n1188 ;
  assign n1190 = ~n580 & n1189 ;
  assign n1191 = n1158 | n1190 ;
  assign n1192 = x129 &  n779 ;
  assign n1193 = ~x129 & n788 ;
  assign n1194 = n1192 | n1193 ;
  assign n1196 = ( x129 & ~n782 ) | ( x129 & 1'b0 ) | ( ~n782 & 1'b0 ) ;
  assign n1195 = x129 | n795 ;
  assign n1197 = ( n1194 & ~n1196 ) | ( n1194 & n1195 ) | ( ~n1196 & n1195 ) ;
  assign n1198 = x130 &  n1197 ;
  assign n1199 = x129 &  n790 ;
  assign n1200 = ~x129 & n520 ;
  assign n1201 = n1199 | n1200 ;
  assign n1203 = ( x129 & ~n793 ) | ( x129 & 1'b0 ) | ( ~n793 & 1'b0 ) ;
  assign n1202 = x129 | n527 ;
  assign n1204 = ( n1201 & ~n1203 ) | ( n1201 & n1202 ) | ( ~n1203 & n1202 ) ;
  assign n1205 = ~x130 & n1204 ;
  assign n1206 = ( n1198 & ~x131 ) | ( n1198 & n1205 ) | ( ~x131 & n1205 ) ;
  assign n1207 = x129 &  n802 ;
  assign n1208 = ~x129 & n777 ;
  assign n1209 = n1207 | n1208 ;
  assign n1211 = ( x129 & ~n805 ) | ( x129 & 1'b0 ) | ( ~n805 & 1'b0 ) ;
  assign n1210 = x129 | n784 ;
  assign n1212 = ( n1209 & ~n1211 ) | ( n1209 & n1210 ) | ( ~n1211 & n1210 ) ;
  assign n1213 = ~x130 & n1212 ;
  assign n1214 = x129 &  n813 ;
  assign n1215 = ~x129 & n800 ;
  assign n1216 = n1214 | n1215 ;
  assign n1218 = ( x129 & ~n816 ) | ( x129 & 1'b0 ) | ( ~n816 & 1'b0 ) ;
  assign n1217 = x129 | n807 ;
  assign n1219 = ( n1216 & ~n1218 ) | ( n1216 & n1217 ) | ( ~n1218 & n1217 ) ;
  assign n1220 = x130 &  n1219 ;
  assign n1221 = ( x131 & n1213 ) | ( x131 & n1220 ) | ( n1213 & n1220 ) ;
  assign n1222 = n1206 | n1221 ;
  assign n1223 = ~n436 & n1222 ;
  assign n1224 = x129 &  n682 ;
  assign n1225 = ~x129 & n691 ;
  assign n1226 = n1224 | n1225 ;
  assign n1228 = ( x129 & ~n685 ) | ( x129 & 1'b0 ) | ( ~n685 & 1'b0 ) ;
  assign n1227 = x129 | n698 ;
  assign n1229 = ( n1226 & ~n1228 ) | ( n1226 & n1227 ) | ( ~n1228 & n1227 ) ;
  assign n1230 = x130 &  n1229 ;
  assign n1231 = x129 &  n693 ;
  assign n1232 = ~x129 & n666 ;
  assign n1233 = n1231 | n1232 ;
  assign n1235 = ( x129 & ~n696 ) | ( x129 & 1'b0 ) | ( ~n696 & 1'b0 ) ;
  assign n1234 = x129 | n673 ;
  assign n1236 = ( n1233 & ~n1235 ) | ( n1233 & n1234 ) | ( ~n1235 & n1234 ) ;
  assign n1237 = ~x130 & n1236 ;
  assign n1238 = ( n1230 & ~x131 ) | ( n1230 & n1237 ) | ( ~x131 & n1237 ) ;
  assign n1239 = x129 &  n705 ;
  assign n1240 = ~x129 & n680 ;
  assign n1241 = n1239 | n1240 ;
  assign n1243 = ( x129 & ~n708 ) | ( x129 & 1'b0 ) | ( ~n708 & 1'b0 ) ;
  assign n1242 = x129 | n687 ;
  assign n1244 = ( n1241 & ~n1243 ) | ( n1241 & n1242 ) | ( ~n1243 & n1242 ) ;
  assign n1245 = ~x130 & n1244 ;
  assign n1246 = x129 &  n716 ;
  assign n1247 = ~x129 & n703 ;
  assign n1248 = n1246 | n1247 ;
  assign n1250 = ( x129 & ~n719 ) | ( x129 & 1'b0 ) | ( ~n719 & 1'b0 ) ;
  assign n1249 = x129 | n710 ;
  assign n1251 = ( n1248 & ~n1250 ) | ( n1248 & n1249 ) | ( ~n1250 & n1249 ) ;
  assign n1252 = x130 &  n1251 ;
  assign n1253 = ( x131 & n1245 ) | ( x131 & n1252 ) | ( n1245 & n1252 ) ;
  assign n1254 = n1238 | n1253 ;
  assign n1255 = n485 &  n1254 ;
  assign n1256 = n1223 | n1255 ;
  assign n1257 = n1191 | n1256 ;
  assign n1258 = ~x134 & n1257 ;
  assign n1259 = n1126 | n1258 ;
  assign n1260 = x130 | x131 ;
  assign n1261 = ( n279 & ~n1260 ) | ( n279 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1262 = ~x130 |  x131 ;
  assign n1263 = ( n223 & ~n1262 ) | ( n223 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1264 = n1261 | n1263 ;
  assign n1265 = x130 &  x131 ;
  assign n1266 = n235 &  n1265 ;
  assign n1267 = ~x131 |  x130 ;
  assign n1268 = ( n215 & ~n1267 ) | ( n215 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1269 = ( n1266 & ~n1264 ) | ( n1266 & n1268 ) | ( ~n1264 & n1268 ) ;
  assign n1270 = n1264 | n1269 ;
  assign n1271 = x132 &  n1270 ;
  assign n1272 = ( n354 & ~n1260 ) | ( n354 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1273 = n271 &  n1265 ;
  assign n1274 = ( n262 & ~n1262 ) | ( n262 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1275 = ( n254 & ~n1267 ) | ( n254 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1276 = ( n1274 & ~n1273 ) | ( n1274 & n1275 ) | ( ~n1273 & n1275 ) ;
  assign n1277 = ( n1273 & ~n1272 ) | ( n1273 & n1276 ) | ( ~n1272 & n1276 ) ;
  assign n1278 = n1272 | n1277 ;
  assign n1279 = ~x132 & n1278 ;
  assign n1280 = ( n1271 & ~x133 ) | ( n1271 & n1279 ) | ( ~x133 & n1279 ) ;
  assign n1281 = ( n243 & ~n1260 ) | ( n243 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1282 = n159 &  n1265 ;
  assign n1283 = ( n150 & ~n1262 ) | ( n150 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1284 = ( n142 & ~n1267 ) | ( n142 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1285 = ( n1283 & ~n1282 ) | ( n1283 & n1284 ) | ( ~n1282 & n1284 ) ;
  assign n1286 = ( n1282 & ~n1281 ) | ( n1282 & n1285 ) | ( ~n1281 & n1285 ) ;
  assign n1287 = n1281 | n1286 ;
  assign n1288 = ~x132 & n1287 ;
  assign n1289 = ( n167 & ~n1260 ) | ( n167 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1290 = n195 &  n1265 ;
  assign n1291 = ( n186 & ~n1262 ) | ( n186 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1292 = ( n178 & ~n1267 ) | ( n178 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1293 = ( n1291 & ~n1290 ) | ( n1291 & n1292 ) | ( ~n1290 & n1292 ) ;
  assign n1294 = ( n1290 & ~n1289 ) | ( n1290 & n1293 ) | ( ~n1289 & n1293 ) ;
  assign n1295 = n1289 | n1294 ;
  assign n1296 = x132 &  n1295 ;
  assign n1297 = ( x133 & n1288 ) | ( x133 & n1296 ) | ( n1288 & n1296 ) ;
  assign n1298 = n1280 | n1297 ;
  assign n1299 = x134 &  n1298 ;
  assign n1300 = ( n391 & ~n1260 ) | ( n391 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1301 = n310 &  n1265 ;
  assign n1302 = ( n301 & ~n1262 ) | ( n301 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1303 = ( n293 & ~n1267 ) | ( n293 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1304 = ( n1302 & ~n1301 ) | ( n1302 & n1303 ) | ( ~n1301 & n1303 ) ;
  assign n1305 = ( n1301 & ~n1300 ) | ( n1301 & n1304 ) | ( ~n1300 & n1304 ) ;
  assign n1306 = n1300 | n1305 ;
  assign n1307 = ~x132 & n1306 ;
  assign n1308 = ( n318 & ~n1260 ) | ( n318 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1309 = n346 &  n1265 ;
  assign n1310 = ( n337 & ~n1262 ) | ( n337 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1311 = ( n329 & ~n1267 ) | ( n329 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1312 = ( n1310 & ~n1309 ) | ( n1310 & n1311 ) | ( ~n1309 & n1311 ) ;
  assign n1313 = ( n1309 & ~n1308 ) | ( n1309 & n1312 ) | ( ~n1308 & n1312 ) ;
  assign n1314 = n1308 | n1313 ;
  assign n1315 = x132 &  n1314 ;
  assign n1316 = ( x133 & n1307 ) | ( x133 & n1315 ) | ( n1307 & n1315 ) ;
  assign n1317 = ( n427 & ~n1260 ) | ( n427 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1318 = n383 &  n1265 ;
  assign n1319 = ( n374 & ~n1262 ) | ( n374 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1320 = ( n366 & ~n1267 ) | ( n366 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1321 = ( n1319 & ~n1318 ) | ( n1319 & n1320 ) | ( ~n1318 & n1320 ) ;
  assign n1322 = ( n1318 & ~n1317 ) | ( n1318 & n1321 ) | ( ~n1317 & n1321 ) ;
  assign n1323 = n1317 | n1322 ;
  assign n1324 = x132 &  n1323 ;
  assign n1325 = ( n203 & ~n1260 ) | ( n203 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1326 = n419 &  n1265 ;
  assign n1327 = ( n410 & ~n1262 ) | ( n410 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1328 = ( n402 & ~n1267 ) | ( n402 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1329 = ( n1327 & ~n1326 ) | ( n1327 & n1328 ) | ( ~n1326 & n1328 ) ;
  assign n1330 = ( n1326 & ~n1325 ) | ( n1326 & n1329 ) | ( ~n1325 & n1329 ) ;
  assign n1331 = n1325 | n1330 ;
  assign n1332 = ~x132 & n1331 ;
  assign n1333 = ( n1324 & ~x133 ) | ( n1324 & n1332 ) | ( ~x133 & n1332 ) ;
  assign n1334 = n1316 | n1333 ;
  assign n1335 = ~x134 & n1334 ;
  assign n1336 = n1299 | n1335 ;
  assign n1337 = ( n480 & ~n1260 ) | ( n480 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1338 = ( n554 & ~n1262 ) | ( n554 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1339 = n1337 | n1338 ;
  assign n1340 = n564 &  n1265 ;
  assign n1341 = ( n543 & ~n1267 ) | ( n543 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1342 = n1340 | n1341 ;
  assign n1343 = n1339 | n1342 ;
  assign n1344 = x132 &  n1343 ;
  assign n1345 = ( n723 & ~n1260 ) | ( n723 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1346 = ( n457 & ~n1262 ) | ( n457 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1347 = n1345 | n1346 ;
  assign n1348 = n469 &  n1265 ;
  assign n1349 = ( n446 & ~n1267 ) | ( n446 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1350 = n1348 | n1349 ;
  assign n1351 = n1347 | n1350 ;
  assign n1352 = ~x132 & n1351 ;
  assign n1353 = ( n1344 & ~x133 ) | ( n1344 & n1352 ) | ( ~x133 & n1352 ) ;
  assign n1354 = ( n575 & ~n1260 ) | ( n575 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1355 = ( n601 & ~n1262 ) | ( n601 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1356 = n1354 | n1355 ;
  assign n1357 = n613 &  n1265 ;
  assign n1358 = ( n590 & ~n1267 ) | ( n590 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1359 = n1357 | n1358 ;
  assign n1360 = n1356 | n1359 ;
  assign n1361 = ~x132 & n1360 ;
  assign n1362 = ( n624 & ~n1260 ) | ( n624 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1363 = ( n506 & ~n1262 ) | ( n506 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1364 = n1362 | n1363 ;
  assign n1365 = n518 &  n1265 ;
  assign n1366 = ( n495 & ~n1267 ) | ( n495 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1367 = n1365 | n1366 ;
  assign n1368 = n1364 | n1367 ;
  assign n1369 = x132 &  n1368 ;
  assign n1370 = ( x133 & n1361 ) | ( x133 & n1369 ) | ( n1361 & n1369 ) ;
  assign n1371 = n1353 | n1370 ;
  assign n1372 = x134 &  n1371 ;
  assign n1373 = ( n772 & ~n1260 ) | ( n772 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1374 = ( n652 & ~n1262 ) | ( n652 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1375 = n1373 | n1374 ;
  assign n1376 = n664 &  n1265 ;
  assign n1377 = ( n641 & ~n1267 ) | ( n641 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1378 = n1376 | n1377 ;
  assign n1379 = n1375 | n1378 ;
  assign n1380 = ~x132 & n1379 ;
  assign n1381 = ( n675 & ~n1260 ) | ( n675 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1382 = ( n700 & ~n1262 ) | ( n700 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1383 = n1381 | n1382 ;
  assign n1384 = n712 &  n1265 ;
  assign n1385 = ( n689 & ~n1267 ) | ( n689 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1386 = n1384 | n1385 ;
  assign n1387 = n1383 | n1386 ;
  assign n1388 = x132 &  n1387 ;
  assign n1389 = ( x133 & n1380 ) | ( x133 & n1388 ) | ( n1380 & n1388 ) ;
  assign n1390 = ( n820 & ~n1260 ) | ( n820 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1391 = ( n749 & ~n1262 ) | ( n749 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1392 = n1390 | n1391 ;
  assign n1393 = n761 &  n1265 ;
  assign n1394 = ( n738 & ~n1267 ) | ( n738 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1395 = n1393 | n1394 ;
  assign n1396 = n1392 | n1395 ;
  assign n1397 = x132 &  n1396 ;
  assign n1398 = ( n529 & ~n1260 ) | ( n529 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1399 = ( n797 & ~n1262 ) | ( n797 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1400 = n1398 | n1399 ;
  assign n1401 = n809 &  n1265 ;
  assign n1402 = ( n786 & ~n1267 ) | ( n786 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1403 = n1401 | n1402 ;
  assign n1404 = n1400 | n1403 ;
  assign n1405 = ~x132 & n1404 ;
  assign n1406 = ( n1397 & ~x133 ) | ( n1397 & n1405 ) | ( ~x133 & n1405 ) ;
  assign n1407 = n1389 | n1406 ;
  assign n1408 = ~x134 & n1407 ;
  assign n1409 = n1372 | n1408 ;
  assign n1410 = ( n844 & ~n1260 ) | ( n844 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1411 = n881 &  n1265 ;
  assign n1412 = ( n876 & ~n1262 ) | ( n876 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1413 = ( n872 & ~n1267 ) | ( n872 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1414 = ( n1412 & ~n1411 ) | ( n1412 & n1413 ) | ( ~n1411 & n1413 ) ;
  assign n1415 = ( n1411 & ~n1410 ) | ( n1411 & n1414 ) | ( ~n1410 & n1414 ) ;
  assign n1416 = n1410 | n1415 ;
  assign n1417 = x132 &  n1416 ;
  assign n1418 = ( n948 & ~n1260 ) | ( n948 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1419 = n840 &  n1265 ;
  assign n1420 = ( n835 & ~n1262 ) | ( n835 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1421 = ( n831 & ~n1267 ) | ( n831 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1422 = ( n1420 & ~n1419 ) | ( n1420 & n1421 ) | ( ~n1419 & n1421 ) ;
  assign n1423 = ( n1419 & ~n1418 ) | ( n1419 & n1422 ) | ( ~n1418 & n1422 ) ;
  assign n1424 = n1418 | n1423 ;
  assign n1425 = ~x132 & n1424 ;
  assign n1426 = ( n1417 & ~x133 ) | ( n1417 & n1425 ) | ( ~x133 & n1425 ) ;
  assign n1427 = ( n885 & ~n1260 ) | ( n885 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1428 = n901 &  n1265 ;
  assign n1429 = ( n896 & ~n1262 ) | ( n896 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1430 = ( n892 & ~n1267 ) | ( n892 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1431 = ( n1429 & ~n1428 ) | ( n1429 & n1430 ) | ( ~n1428 & n1430 ) ;
  assign n1432 = ( n1428 & ~n1427 ) | ( n1428 & n1431 ) | ( ~n1427 & n1431 ) ;
  assign n1433 = n1427 | n1432 ;
  assign n1434 = ~x132 & n1433 ;
  assign n1435 = ( n905 & ~n1260 ) | ( n905 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1436 = n860 &  n1265 ;
  assign n1437 = ( n855 & ~n1262 ) | ( n855 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1438 = ( n851 & ~n1267 ) | ( n851 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1439 = ( n1437 & ~n1436 ) | ( n1437 & n1438 ) | ( ~n1436 & n1438 ) ;
  assign n1440 = ( n1436 & ~n1435 ) | ( n1436 & n1439 ) | ( ~n1435 & n1439 ) ;
  assign n1441 = n1435 | n1440 ;
  assign n1442 = x132 &  n1441 ;
  assign n1443 = ( x133 & n1434 ) | ( x133 & n1442 ) | ( n1434 & n1442 ) ;
  assign n1444 = n1426 | n1443 ;
  assign n1445 = x134 &  n1444 ;
  assign n1446 = ( n969 & ~n1260 ) | ( n969 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1447 = n924 &  n1265 ;
  assign n1448 = ( n919 & ~n1262 ) | ( n919 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1449 = ( n915 & ~n1267 ) | ( n915 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1450 = ( n1448 & ~n1447 ) | ( n1448 & n1449 ) | ( ~n1447 & n1449 ) ;
  assign n1451 = ( n1447 & ~n1446 ) | ( n1447 & n1450 ) | ( ~n1446 & n1450 ) ;
  assign n1452 = n1446 | n1451 ;
  assign n1453 = ~x132 & n1452 ;
  assign n1454 = ( n928 & ~n1260 ) | ( n928 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1455 = n944 &  n1265 ;
  assign n1456 = ( n939 & ~n1262 ) | ( n939 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1457 = ( n935 & ~n1267 ) | ( n935 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1458 = ( n1456 & ~n1455 ) | ( n1456 & n1457 ) | ( ~n1455 & n1457 ) ;
  assign n1459 = ( n1455 & ~n1454 ) | ( n1455 & n1458 ) | ( ~n1454 & n1458 ) ;
  assign n1460 = n1454 | n1459 ;
  assign n1461 = x132 &  n1460 ;
  assign n1462 = ( x133 & n1453 ) | ( x133 & n1461 ) | ( n1453 & n1461 ) ;
  assign n1463 = ( n989 & ~n1260 ) | ( n989 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1464 = n965 &  n1265 ;
  assign n1465 = ( n960 & ~n1262 ) | ( n960 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1466 = ( n956 & ~n1267 ) | ( n956 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1467 = ( n1465 & ~n1464 ) | ( n1465 & n1466 ) | ( ~n1464 & n1466 ) ;
  assign n1468 = ( n1464 & ~n1463 ) | ( n1464 & n1467 ) | ( ~n1463 & n1467 ) ;
  assign n1469 = n1463 | n1468 ;
  assign n1470 = x132 &  n1469 ;
  assign n1471 = ( n864 & ~n1260 ) | ( n864 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1472 = n985 &  n1265 ;
  assign n1473 = ( n980 & ~n1262 ) | ( n980 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1474 = ( n976 & ~n1267 ) | ( n976 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1475 = ( n1473 & ~n1472 ) | ( n1473 & n1474 ) | ( ~n1472 & n1474 ) ;
  assign n1476 = ( n1472 & ~n1471 ) | ( n1472 & n1475 ) | ( ~n1471 & n1475 ) ;
  assign n1477 = n1471 | n1476 ;
  assign n1478 = ~x132 & n1477 ;
  assign n1479 = ( n1470 & ~x133 ) | ( n1470 & n1478 ) | ( ~x133 & n1478 ) ;
  assign n1480 = n1462 | n1479 ;
  assign n1481 = ~x134 & n1480 ;
  assign n1482 = n1445 | n1481 ;
  assign n1483 = ( n1007 & ~n1262 ) | ( n1007 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1484 = ( n1000 & ~n1267 ) | ( n1000 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1485 = n1483 | n1484 ;
  assign n1486 = n1015 &  n1265 ;
  assign n1487 = ( n1054 & ~n1260 ) | ( n1054 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1488 = n1486 | n1487 ;
  assign n1489 = n1485 | n1488 ;
  assign n1490 = x132 &  n1489 ;
  assign n1491 = ( n1251 & ~n1260 ) | ( n1251 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1492 = ( n1039 & ~n1262 ) | ( n1039 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1493 = n1491 | n1492 ;
  assign n1494 = n1047 &  n1265 ;
  assign n1495 = ( n1032 & ~n1267 ) | ( n1032 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1496 = n1494 | n1495 ;
  assign n1497 = n1493 | n1496 ;
  assign n1498 = ~x132 & n1497 ;
  assign n1499 = ( n1490 & ~x133 ) | ( n1490 & n1498 ) | ( ~x133 & n1498 ) ;
  assign n1500 = ( n1022 & ~n1260 ) | ( n1022 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1501 = ( n1072 & ~n1262 ) | ( n1072 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1502 = n1500 | n1501 ;
  assign n1503 = n1080 &  n1265 ;
  assign n1504 = ( n1065 & ~n1267 ) | ( n1065 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1505 = n1503 | n1504 ;
  assign n1506 = n1502 | n1505 ;
  assign n1507 = ~x132 & n1506 ;
  assign n1508 = ( n1087 & ~n1260 ) | ( n1087 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1509 = ( n1104 & ~n1262 ) | ( n1104 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1510 = n1508 | n1509 ;
  assign n1511 = n1112 &  n1265 ;
  assign n1512 = ( n1097 & ~n1267 ) | ( n1097 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1513 = n1511 | n1512 ;
  assign n1514 = n1510 | n1513 ;
  assign n1515 = x132 &  n1514 ;
  assign n1516 = ( x133 & n1507 ) | ( x133 & n1515 ) | ( n1507 & n1515 ) ;
  assign n1517 = n1499 | n1516 ;
  assign n1518 = x134 &  n1517 ;
  assign n1519 = ( n1154 & ~n1260 ) | ( n1154 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1520 = ( n1171 & ~n1262 ) | ( n1171 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1521 = n1519 | n1520 ;
  assign n1522 = n1179 &  n1265 ;
  assign n1523 = ( n1164 & ~n1267 ) | ( n1164 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1524 = n1522 | n1523 ;
  assign n1525 = n1521 | n1524 ;
  assign n1526 = ~x132 & n1525 ;
  assign n1527 = ( n1186 & ~n1260 ) | ( n1186 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1528 = ( n1236 & ~n1262 ) | ( n1236 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1529 = n1527 | n1528 ;
  assign n1530 = n1244 &  n1265 ;
  assign n1531 = ( n1229 & ~n1267 ) | ( n1229 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1532 = n1530 | n1531 ;
  assign n1533 = n1529 | n1532 ;
  assign n1534 = x132 &  n1533 ;
  assign n1535 = ( x133 & n1526 ) | ( x133 & n1534 ) | ( n1526 & n1534 ) ;
  assign n1536 = ( n1219 & ~n1260 ) | ( n1219 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1537 = ( n1139 & ~n1262 ) | ( n1139 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1538 = n1536 | n1537 ;
  assign n1539 = n1147 &  n1265 ;
  assign n1540 = ( n1132 & ~n1267 ) | ( n1132 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1541 = n1539 | n1540 ;
  assign n1542 = n1538 | n1541 ;
  assign n1543 = x132 &  n1542 ;
  assign n1544 = ( n1119 & ~n1260 ) | ( n1119 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1545 = ( n1204 & ~n1262 ) | ( n1204 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1546 = n1544 | n1545 ;
  assign n1547 = n1212 &  n1265 ;
  assign n1548 = ( n1197 & ~n1267 ) | ( n1197 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1549 = n1547 | n1548 ;
  assign n1550 = n1546 | n1549 ;
  assign n1551 = ~x132 & n1550 ;
  assign n1552 = ( n1543 & ~x133 ) | ( n1543 & n1551 ) | ( ~x133 & n1551 ) ;
  assign n1553 = n1535 | n1552 ;
  assign n1554 = ~x134 & n1553 ;
  assign n1555 = n1518 | n1554 ;
  assign n1556 = ( n271 & ~n1260 ) | ( n271 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1557 = n215 &  n1265 ;
  assign n1558 = ( n279 & ~n1262 ) | ( n279 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1559 = ( n223 & ~n1267 ) | ( n223 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1560 = ( n1558 & ~n1557 ) | ( n1558 & n1559 ) | ( ~n1557 & n1559 ) ;
  assign n1561 = ( n1557 & ~n1556 ) | ( n1557 & n1560 ) | ( ~n1556 & n1560 ) ;
  assign n1562 = n1556 | n1561 ;
  assign n1563 = x132 &  n1562 ;
  assign n1564 = ( n346 & ~n1260 ) | ( n346 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1565 = n254 &  n1265 ;
  assign n1566 = ( n354 & ~n1262 ) | ( n354 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1567 = ( n262 & ~n1267 ) | ( n262 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1568 = ( n1566 & ~n1565 ) | ( n1566 & n1567 ) | ( ~n1565 & n1567 ) ;
  assign n1569 = ( n1565 & ~n1564 ) | ( n1565 & n1568 ) | ( ~n1564 & n1568 ) ;
  assign n1570 = n1564 | n1569 ;
  assign n1571 = ~x132 & n1570 ;
  assign n1572 = ( n1563 & ~x133 ) | ( n1563 & n1571 ) | ( ~x133 & n1571 ) ;
  assign n1573 = ( n235 & ~n1260 ) | ( n235 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1574 = n142 &  n1265 ;
  assign n1575 = ( n243 & ~n1262 ) | ( n243 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1576 = ( n150 & ~n1267 ) | ( n150 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1577 = ( n1575 & ~n1574 ) | ( n1575 & n1576 ) | ( ~n1574 & n1576 ) ;
  assign n1578 = ( n1574 & ~n1573 ) | ( n1574 & n1577 ) | ( ~n1573 & n1577 ) ;
  assign n1579 = n1573 | n1578 ;
  assign n1580 = ~x132 & n1579 ;
  assign n1581 = ( n159 & ~n1260 ) | ( n159 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1582 = n178 &  n1265 ;
  assign n1583 = ( n167 & ~n1262 ) | ( n167 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1584 = ( n186 & ~n1267 ) | ( n186 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1585 = ( n1583 & ~n1582 ) | ( n1583 & n1584 ) | ( ~n1582 & n1584 ) ;
  assign n1586 = ( n1582 & ~n1581 ) | ( n1582 & n1585 ) | ( ~n1581 & n1585 ) ;
  assign n1587 = n1581 | n1586 ;
  assign n1588 = x132 &  n1587 ;
  assign n1589 = ( x133 & n1580 ) | ( x133 & n1588 ) | ( n1580 & n1588 ) ;
  assign n1590 = n1572 | n1589 ;
  assign n1591 = x134 &  n1590 ;
  assign n1592 = ( n383 & ~n1260 ) | ( n383 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1593 = n293 &  n1265 ;
  assign n1594 = ( n391 & ~n1262 ) | ( n391 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1595 = ( n301 & ~n1267 ) | ( n301 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1596 = ( n1594 & ~n1593 ) | ( n1594 & n1595 ) | ( ~n1593 & n1595 ) ;
  assign n1597 = ( n1593 & ~n1592 ) | ( n1593 & n1596 ) | ( ~n1592 & n1596 ) ;
  assign n1598 = n1592 | n1597 ;
  assign n1599 = ~x132 & n1598 ;
  assign n1600 = ( n310 & ~n1260 ) | ( n310 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1601 = n329 &  n1265 ;
  assign n1602 = ( n318 & ~n1262 ) | ( n318 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1603 = ( n337 & ~n1267 ) | ( n337 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1604 = ( n1602 & ~n1601 ) | ( n1602 & n1603 ) | ( ~n1601 & n1603 ) ;
  assign n1605 = ( n1601 & ~n1600 ) | ( n1601 & n1604 ) | ( ~n1600 & n1604 ) ;
  assign n1606 = n1600 | n1605 ;
  assign n1607 = x132 &  n1606 ;
  assign n1608 = ( x133 & n1599 ) | ( x133 & n1607 ) | ( n1599 & n1607 ) ;
  assign n1609 = ( n419 & ~n1260 ) | ( n419 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1610 = n366 &  n1265 ;
  assign n1611 = ( n427 & ~n1262 ) | ( n427 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1612 = ( n374 & ~n1267 ) | ( n374 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1613 = ( n1611 & ~n1610 ) | ( n1611 & n1612 ) | ( ~n1610 & n1612 ) ;
  assign n1614 = ( n1610 & ~n1609 ) | ( n1610 & n1613 ) | ( ~n1609 & n1613 ) ;
  assign n1615 = n1609 | n1614 ;
  assign n1616 = x132 &  n1615 ;
  assign n1617 = ( n195 & ~n1260 ) | ( n195 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1618 = n402 &  n1265 ;
  assign n1619 = ( n203 & ~n1262 ) | ( n203 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1620 = ( n410 & ~n1267 ) | ( n410 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1621 = ( n1619 & ~n1618 ) | ( n1619 & n1620 ) | ( ~n1618 & n1620 ) ;
  assign n1622 = ( n1618 & ~n1617 ) | ( n1618 & n1621 ) | ( ~n1617 & n1621 ) ;
  assign n1623 = n1617 | n1622 ;
  assign n1624 = ~x132 & n1623 ;
  assign n1625 = ( n1616 & ~x133 ) | ( n1616 & n1624 ) | ( ~x133 & n1624 ) ;
  assign n1626 = n1608 | n1625 ;
  assign n1627 = ~x134 & n1626 ;
  assign n1628 = n1591 | n1627 ;
  assign n1629 = ( n469 & ~n1260 ) | ( n469 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1630 = ( n480 & ~n1262 ) | ( n480 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1631 = n1629 | n1630 ;
  assign n1632 = n543 &  n1265 ;
  assign n1633 = ( n554 & ~n1267 ) | ( n554 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1634 = n1632 | n1633 ;
  assign n1635 = n1631 | n1634 ;
  assign n1636 = x132 &  n1635 ;
  assign n1637 = ( n712 & ~n1260 ) | ( n712 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1638 = ( n723 & ~n1262 ) | ( n723 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1639 = n1637 | n1638 ;
  assign n1640 = n446 &  n1265 ;
  assign n1641 = ( n457 & ~n1267 ) | ( n457 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1642 = n1640 | n1641 ;
  assign n1643 = n1639 | n1642 ;
  assign n1644 = ~x132 & n1643 ;
  assign n1645 = ( n1636 & ~x133 ) | ( n1636 & n1644 ) | ( ~x133 & n1644 ) ;
  assign n1646 = ( n564 & ~n1260 ) | ( n564 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1647 = ( n575 & ~n1262 ) | ( n575 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1648 = n1646 | n1647 ;
  assign n1649 = n590 &  n1265 ;
  assign n1650 = ( n601 & ~n1267 ) | ( n601 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1651 = n1649 | n1650 ;
  assign n1652 = n1648 | n1651 ;
  assign n1653 = ~x132 & n1652 ;
  assign n1654 = ( n613 & ~n1260 ) | ( n613 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1655 = ( n624 & ~n1262 ) | ( n624 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1656 = n1654 | n1655 ;
  assign n1657 = n495 &  n1265 ;
  assign n1658 = ( n506 & ~n1267 ) | ( n506 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1659 = n1657 | n1658 ;
  assign n1660 = n1656 | n1659 ;
  assign n1661 = x132 &  n1660 ;
  assign n1662 = ( x133 & n1653 ) | ( x133 & n1661 ) | ( n1653 & n1661 ) ;
  assign n1663 = n1645 | n1662 ;
  assign n1664 = x134 &  n1663 ;
  assign n1665 = ( n761 & ~n1260 ) | ( n761 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1666 = ( n772 & ~n1262 ) | ( n772 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1667 = n1665 | n1666 ;
  assign n1668 = n641 &  n1265 ;
  assign n1669 = ( n652 & ~n1267 ) | ( n652 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1670 = n1668 | n1669 ;
  assign n1671 = n1667 | n1670 ;
  assign n1672 = ~x132 & n1671 ;
  assign n1673 = ( n664 & ~n1260 ) | ( n664 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1674 = ( n675 & ~n1262 ) | ( n675 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1675 = n1673 | n1674 ;
  assign n1676 = n689 &  n1265 ;
  assign n1677 = ( n700 & ~n1267 ) | ( n700 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1678 = n1676 | n1677 ;
  assign n1679 = n1675 | n1678 ;
  assign n1680 = x132 &  n1679 ;
  assign n1681 = ( x133 & n1672 ) | ( x133 & n1680 ) | ( n1672 & n1680 ) ;
  assign n1682 = ( n809 & ~n1260 ) | ( n809 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1683 = ( n820 & ~n1262 ) | ( n820 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1684 = n1682 | n1683 ;
  assign n1685 = n738 &  n1265 ;
  assign n1686 = ( n749 & ~n1267 ) | ( n749 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1687 = n1685 | n1686 ;
  assign n1688 = n1684 | n1687 ;
  assign n1689 = x132 &  n1688 ;
  assign n1690 = ( n518 & ~n1260 ) | ( n518 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1691 = ( n529 & ~n1262 ) | ( n529 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1692 = n1690 | n1691 ;
  assign n1693 = n786 &  n1265 ;
  assign n1694 = ( n797 & ~n1267 ) | ( n797 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1695 = n1693 | n1694 ;
  assign n1696 = n1692 | n1695 ;
  assign n1697 = ~x132 & n1696 ;
  assign n1698 = ( n1689 & ~x133 ) | ( n1689 & n1697 ) | ( ~x133 & n1697 ) ;
  assign n1699 = n1681 | n1698 ;
  assign n1700 = ~x134 & n1699 ;
  assign n1701 = n1664 | n1700 ;
  assign n1702 = ( n840 & ~n1260 ) | ( n840 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1703 = n872 &  n1265 ;
  assign n1704 = ( n844 & ~n1262 ) | ( n844 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1705 = ( n876 & ~n1267 ) | ( n876 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1706 = ( n1704 & ~n1703 ) | ( n1704 & n1705 ) | ( ~n1703 & n1705 ) ;
  assign n1707 = ( n1703 & ~n1702 ) | ( n1703 & n1706 ) | ( ~n1702 & n1706 ) ;
  assign n1708 = n1702 | n1707 ;
  assign n1709 = x132 &  n1708 ;
  assign n1710 = ( n944 & ~n1260 ) | ( n944 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1711 = n831 &  n1265 ;
  assign n1712 = ( n948 & ~n1262 ) | ( n948 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1713 = ( n835 & ~n1267 ) | ( n835 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1714 = ( n1712 & ~n1711 ) | ( n1712 & n1713 ) | ( ~n1711 & n1713 ) ;
  assign n1715 = ( n1711 & ~n1710 ) | ( n1711 & n1714 ) | ( ~n1710 & n1714 ) ;
  assign n1716 = n1710 | n1715 ;
  assign n1717 = ~x132 & n1716 ;
  assign n1718 = ( n1709 & ~x133 ) | ( n1709 & n1717 ) | ( ~x133 & n1717 ) ;
  assign n1719 = ( n881 & ~n1260 ) | ( n881 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1720 = n892 &  n1265 ;
  assign n1721 = ( n885 & ~n1262 ) | ( n885 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1722 = ( n896 & ~n1267 ) | ( n896 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1723 = ( n1721 & ~n1720 ) | ( n1721 & n1722 ) | ( ~n1720 & n1722 ) ;
  assign n1724 = ( n1720 & ~n1719 ) | ( n1720 & n1723 ) | ( ~n1719 & n1723 ) ;
  assign n1725 = n1719 | n1724 ;
  assign n1726 = ~x132 & n1725 ;
  assign n1727 = ( n901 & ~n1260 ) | ( n901 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1728 = n851 &  n1265 ;
  assign n1729 = ( n905 & ~n1262 ) | ( n905 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1730 = ( n855 & ~n1267 ) | ( n855 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1731 = ( n1729 & ~n1728 ) | ( n1729 & n1730 ) | ( ~n1728 & n1730 ) ;
  assign n1732 = ( n1728 & ~n1727 ) | ( n1728 & n1731 ) | ( ~n1727 & n1731 ) ;
  assign n1733 = n1727 | n1732 ;
  assign n1734 = x132 &  n1733 ;
  assign n1735 = ( x133 & n1726 ) | ( x133 & n1734 ) | ( n1726 & n1734 ) ;
  assign n1736 = n1718 | n1735 ;
  assign n1737 = x134 &  n1736 ;
  assign n1738 = ( n965 & ~n1260 ) | ( n965 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1739 = n915 &  n1265 ;
  assign n1740 = ( n969 & ~n1262 ) | ( n969 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1741 = ( n919 & ~n1267 ) | ( n919 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1742 = ( n1740 & ~n1739 ) | ( n1740 & n1741 ) | ( ~n1739 & n1741 ) ;
  assign n1743 = ( n1739 & ~n1738 ) | ( n1739 & n1742 ) | ( ~n1738 & n1742 ) ;
  assign n1744 = n1738 | n1743 ;
  assign n1745 = ~x132 & n1744 ;
  assign n1746 = ( n924 & ~n1260 ) | ( n924 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1747 = n935 &  n1265 ;
  assign n1748 = ( n928 & ~n1262 ) | ( n928 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1749 = ( n939 & ~n1267 ) | ( n939 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1750 = ( n1748 & ~n1747 ) | ( n1748 & n1749 ) | ( ~n1747 & n1749 ) ;
  assign n1751 = ( n1747 & ~n1746 ) | ( n1747 & n1750 ) | ( ~n1746 & n1750 ) ;
  assign n1752 = n1746 | n1751 ;
  assign n1753 = x132 &  n1752 ;
  assign n1754 = ( x133 & n1745 ) | ( x133 & n1753 ) | ( n1745 & n1753 ) ;
  assign n1755 = ( n985 & ~n1260 ) | ( n985 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1756 = n956 &  n1265 ;
  assign n1757 = ( n989 & ~n1262 ) | ( n989 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1758 = ( n960 & ~n1267 ) | ( n960 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1759 = ( n1757 & ~n1756 ) | ( n1757 & n1758 ) | ( ~n1756 & n1758 ) ;
  assign n1760 = ( n1756 & ~n1755 ) | ( n1756 & n1759 ) | ( ~n1755 & n1759 ) ;
  assign n1761 = n1755 | n1760 ;
  assign n1762 = x132 &  n1761 ;
  assign n1763 = ( n860 & ~n1260 ) | ( n860 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1764 = n976 &  n1265 ;
  assign n1765 = ( n864 & ~n1262 ) | ( n864 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1766 = ( n980 & ~n1267 ) | ( n980 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1767 = ( n1765 & ~n1764 ) | ( n1765 & n1766 ) | ( ~n1764 & n1766 ) ;
  assign n1768 = ( n1764 & ~n1763 ) | ( n1764 & n1767 ) | ( ~n1763 & n1767 ) ;
  assign n1769 = n1763 | n1768 ;
  assign n1770 = ~x132 & n1769 ;
  assign n1771 = ( n1762 & ~x133 ) | ( n1762 & n1770 ) | ( ~x133 & n1770 ) ;
  assign n1772 = n1754 | n1771 ;
  assign n1773 = ~x134 & n1772 ;
  assign n1774 = n1737 | n1773 ;
  assign n1775 = ( n1047 & ~n1260 ) | ( n1047 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1776 = ( n1007 & ~n1267 ) | ( n1007 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1777 = n1775 | n1776 ;
  assign n1778 = n1000 &  n1265 ;
  assign n1779 = ( n1054 & ~n1262 ) | ( n1054 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1780 = n1778 | n1779 ;
  assign n1781 = n1777 | n1780 ;
  assign n1782 = x132 &  n1781 ;
  assign n1783 = ( n1244 & ~n1260 ) | ( n1244 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1784 = ( n1251 & ~n1262 ) | ( n1251 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1785 = n1783 | n1784 ;
  assign n1786 = n1032 &  n1265 ;
  assign n1787 = ( n1039 & ~n1267 ) | ( n1039 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1788 = n1786 | n1787 ;
  assign n1789 = n1785 | n1788 ;
  assign n1790 = ~x132 & n1789 ;
  assign n1791 = ( n1782 & ~x133 ) | ( n1782 & n1790 ) | ( ~x133 & n1790 ) ;
  assign n1792 = ( n1015 & ~n1260 ) | ( n1015 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1793 = ( n1022 & ~n1262 ) | ( n1022 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1794 = n1792 | n1793 ;
  assign n1795 = n1065 &  n1265 ;
  assign n1796 = ( n1072 & ~n1267 ) | ( n1072 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1797 = n1795 | n1796 ;
  assign n1798 = n1794 | n1797 ;
  assign n1799 = ~x132 & n1798 ;
  assign n1800 = ( n1080 & ~n1260 ) | ( n1080 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1801 = ( n1087 & ~n1262 ) | ( n1087 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1802 = n1800 | n1801 ;
  assign n1803 = n1097 &  n1265 ;
  assign n1804 = ( n1104 & ~n1267 ) | ( n1104 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1805 = n1803 | n1804 ;
  assign n1806 = n1802 | n1805 ;
  assign n1807 = x132 &  n1806 ;
  assign n1808 = ( x133 & n1799 ) | ( x133 & n1807 ) | ( n1799 & n1807 ) ;
  assign n1809 = n1791 | n1808 ;
  assign n1810 = x134 &  n1809 ;
  assign n1811 = ( n1147 & ~n1260 ) | ( n1147 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1812 = ( n1154 & ~n1262 ) | ( n1154 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1813 = n1811 | n1812 ;
  assign n1814 = n1164 &  n1265 ;
  assign n1815 = ( n1171 & ~n1267 ) | ( n1171 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1816 = n1814 | n1815 ;
  assign n1817 = n1813 | n1816 ;
  assign n1818 = ~x132 & n1817 ;
  assign n1819 = ( n1179 & ~n1260 ) | ( n1179 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1820 = ( n1186 & ~n1262 ) | ( n1186 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1821 = n1819 | n1820 ;
  assign n1822 = n1229 &  n1265 ;
  assign n1823 = ( n1236 & ~n1267 ) | ( n1236 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1824 = n1822 | n1823 ;
  assign n1825 = n1821 | n1824 ;
  assign n1826 = x132 &  n1825 ;
  assign n1827 = ( x133 & n1818 ) | ( x133 & n1826 ) | ( n1818 & n1826 ) ;
  assign n1828 = ( n1212 & ~n1260 ) | ( n1212 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1829 = ( n1219 & ~n1262 ) | ( n1219 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1830 = n1828 | n1829 ;
  assign n1831 = n1132 &  n1265 ;
  assign n1832 = ( n1139 & ~n1267 ) | ( n1139 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1833 = n1831 | n1832 ;
  assign n1834 = n1830 | n1833 ;
  assign n1835 = x132 &  n1834 ;
  assign n1836 = ( n1112 & ~n1260 ) | ( n1112 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1837 = ( n1119 & ~n1262 ) | ( n1119 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1838 = n1836 | n1837 ;
  assign n1839 = n1197 &  n1265 ;
  assign n1840 = ( n1204 & ~n1267 ) | ( n1204 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1841 = n1839 | n1840 ;
  assign n1842 = n1838 | n1841 ;
  assign n1843 = ~x132 & n1842 ;
  assign n1844 = ( n1835 & ~x133 ) | ( n1835 & n1843 ) | ( ~x133 & n1843 ) ;
  assign n1845 = n1827 | n1844 ;
  assign n1846 = ~x134 & n1845 ;
  assign n1847 = n1810 | n1846 ;
  assign n1848 = ( n254 & ~n1260 ) | ( n254 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1849 = n223 &  n1265 ;
  assign n1850 = ( n271 & ~n1262 ) | ( n271 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1851 = ( n279 & ~n1267 ) | ( n279 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1852 = ( n1850 & ~n1849 ) | ( n1850 & n1851 ) | ( ~n1849 & n1851 ) ;
  assign n1853 = ( n1849 & ~n1848 ) | ( n1849 & n1852 ) | ( ~n1848 & n1852 ) ;
  assign n1854 = n1848 | n1853 ;
  assign n1855 = x132 &  n1854 ;
  assign n1856 = ( n329 & ~n1260 ) | ( n329 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1857 = n262 &  n1265 ;
  assign n1858 = ( n346 & ~n1262 ) | ( n346 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1859 = ( n354 & ~n1267 ) | ( n354 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1860 = ( n1858 & ~n1857 ) | ( n1858 & n1859 ) | ( ~n1857 & n1859 ) ;
  assign n1861 = ( n1857 & ~n1856 ) | ( n1857 & n1860 ) | ( ~n1856 & n1860 ) ;
  assign n1862 = n1856 | n1861 ;
  assign n1863 = ~x132 & n1862 ;
  assign n1864 = ( n1855 & ~x133 ) | ( n1855 & n1863 ) | ( ~x133 & n1863 ) ;
  assign n1865 = ( n215 & ~n1260 ) | ( n215 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1866 = ( n235 & ~n1262 ) | ( n235 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1867 = n150 &  n1265 ;
  assign n1868 = ( n243 & ~n1267 ) | ( n243 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1869 = n1867 | n1868 ;
  assign n1870 = ( n1866 & ~n1865 ) | ( n1866 & n1869 ) | ( ~n1865 & n1869 ) ;
  assign n1871 = n1865 | n1870 ;
  assign n1872 = ~x132 & n1871 ;
  assign n1873 = ( n142 & ~n1260 ) | ( n142 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1874 = n186 &  n1265 ;
  assign n1875 = ( n159 & ~n1262 ) | ( n159 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1876 = ( n167 & ~n1267 ) | ( n167 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1877 = ( n1875 & ~n1874 ) | ( n1875 & n1876 ) | ( ~n1874 & n1876 ) ;
  assign n1878 = ( n1874 & ~n1873 ) | ( n1874 & n1877 ) | ( ~n1873 & n1877 ) ;
  assign n1879 = n1873 | n1878 ;
  assign n1880 = x132 &  n1879 ;
  assign n1881 = ( x133 & n1872 ) | ( x133 & n1880 ) | ( n1872 & n1880 ) ;
  assign n1882 = n1864 | n1881 ;
  assign n1883 = x134 &  n1882 ;
  assign n1884 = ( n366 & ~n1260 ) | ( n366 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1885 = n301 &  n1265 ;
  assign n1886 = ( n383 & ~n1262 ) | ( n383 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1887 = ( n391 & ~n1267 ) | ( n391 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1888 = ( n1886 & ~n1885 ) | ( n1886 & n1887 ) | ( ~n1885 & n1887 ) ;
  assign n1889 = ( n1885 & ~n1884 ) | ( n1885 & n1888 ) | ( ~n1884 & n1888 ) ;
  assign n1890 = n1884 | n1889 ;
  assign n1891 = ~x132 & n1890 ;
  assign n1892 = ( n293 & ~n1260 ) | ( n293 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1893 = n337 &  n1265 ;
  assign n1894 = ( n310 & ~n1262 ) | ( n310 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1895 = ( n318 & ~n1267 ) | ( n318 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1896 = ( n1894 & ~n1893 ) | ( n1894 & n1895 ) | ( ~n1893 & n1895 ) ;
  assign n1897 = ( n1893 & ~n1892 ) | ( n1893 & n1896 ) | ( ~n1892 & n1896 ) ;
  assign n1898 = n1892 | n1897 ;
  assign n1899 = x132 &  n1898 ;
  assign n1900 = ( x133 & n1891 ) | ( x133 & n1899 ) | ( n1891 & n1899 ) ;
  assign n1901 = ( n402 & ~n1260 ) | ( n402 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1902 = n374 &  n1265 ;
  assign n1903 = ( n419 & ~n1262 ) | ( n419 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1904 = ( n427 & ~n1267 ) | ( n427 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1905 = ( n1903 & ~n1902 ) | ( n1903 & n1904 ) | ( ~n1902 & n1904 ) ;
  assign n1906 = ( n1902 & ~n1901 ) | ( n1902 & n1905 ) | ( ~n1901 & n1905 ) ;
  assign n1907 = n1901 | n1906 ;
  assign n1908 = x132 &  n1907 ;
  assign n1909 = ( n178 & ~n1260 ) | ( n178 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1910 = n410 &  n1265 ;
  assign n1911 = ( n195 & ~n1262 ) | ( n195 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1912 = ( n203 & ~n1267 ) | ( n203 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1913 = ( n1911 & ~n1910 ) | ( n1911 & n1912 ) | ( ~n1910 & n1912 ) ;
  assign n1914 = ( n1910 & ~n1909 ) | ( n1910 & n1913 ) | ( ~n1909 & n1913 ) ;
  assign n1915 = n1909 | n1914 ;
  assign n1916 = ~x132 & n1915 ;
  assign n1917 = ( n1908 & ~x133 ) | ( n1908 & n1916 ) | ( ~x133 & n1916 ) ;
  assign n1918 = n1900 | n1917 ;
  assign n1919 = ~x134 & n1918 ;
  assign n1920 = n1883 | n1919 ;
  assign n1921 = ( n446 & ~n1260 ) | ( n446 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1922 = ( n469 & ~n1262 ) | ( n469 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1923 = n1921 | n1922 ;
  assign n1924 = n554 &  n1265 ;
  assign n1925 = ( n480 & ~n1267 ) | ( n480 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1926 = n1924 | n1925 ;
  assign n1927 = n1923 | n1926 ;
  assign n1928 = x132 &  n1927 ;
  assign n1929 = ( n689 & ~n1260 ) | ( n689 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1930 = ( n712 & ~n1262 ) | ( n712 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1931 = n1929 | n1930 ;
  assign n1932 = n457 &  n1265 ;
  assign n1933 = ( n723 & ~n1267 ) | ( n723 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1934 = n1932 | n1933 ;
  assign n1935 = n1931 | n1934 ;
  assign n1936 = ~x132 & n1935 ;
  assign n1937 = ( n1928 & ~x133 ) | ( n1928 & n1936 ) | ( ~x133 & n1936 ) ;
  assign n1938 = ( n543 & ~n1260 ) | ( n543 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1939 = ( n564 & ~n1262 ) | ( n564 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1940 = n1938 | n1939 ;
  assign n1941 = n601 &  n1265 ;
  assign n1942 = ( n575 & ~n1267 ) | ( n575 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1943 = n1941 | n1942 ;
  assign n1944 = n1940 | n1943 ;
  assign n1945 = ~x132 & n1944 ;
  assign n1946 = ( n590 & ~n1260 ) | ( n590 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1947 = ( n613 & ~n1262 ) | ( n613 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1948 = n1946 | n1947 ;
  assign n1949 = n506 &  n1265 ;
  assign n1950 = ( n624 & ~n1267 ) | ( n624 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1951 = n1949 | n1950 ;
  assign n1952 = n1948 | n1951 ;
  assign n1953 = x132 &  n1952 ;
  assign n1954 = ( x133 & n1945 ) | ( x133 & n1953 ) | ( n1945 & n1953 ) ;
  assign n1955 = n1937 | n1954 ;
  assign n1956 = x134 &  n1955 ;
  assign n1957 = ( n738 & ~n1260 ) | ( n738 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1958 = ( n761 & ~n1262 ) | ( n761 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1959 = n1957 | n1958 ;
  assign n1960 = n652 &  n1265 ;
  assign n1961 = ( n772 & ~n1267 ) | ( n772 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1962 = n1960 | n1961 ;
  assign n1963 = n1959 | n1962 ;
  assign n1964 = ~x132 & n1963 ;
  assign n1965 = ( n641 & ~n1260 ) | ( n641 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1966 = ( n664 & ~n1262 ) | ( n664 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1967 = n1965 | n1966 ;
  assign n1968 = n700 &  n1265 ;
  assign n1969 = ( n675 & ~n1267 ) | ( n675 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1970 = n1968 | n1969 ;
  assign n1971 = n1967 | n1970 ;
  assign n1972 = x132 &  n1971 ;
  assign n1973 = ( x133 & n1964 ) | ( x133 & n1972 ) | ( n1964 & n1972 ) ;
  assign n1974 = ( n786 & ~n1260 ) | ( n786 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1975 = ( n809 & ~n1262 ) | ( n809 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1976 = n1974 | n1975 ;
  assign n1977 = n749 &  n1265 ;
  assign n1978 = ( n820 & ~n1267 ) | ( n820 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1979 = n1977 | n1978 ;
  assign n1980 = n1976 | n1979 ;
  assign n1981 = x132 &  n1980 ;
  assign n1982 = ( n495 & ~n1260 ) | ( n495 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1983 = ( n518 & ~n1262 ) | ( n518 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1984 = n1982 | n1983 ;
  assign n1985 = n797 &  n1265 ;
  assign n1986 = ( n529 & ~n1267 ) | ( n529 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1987 = n1985 | n1986 ;
  assign n1988 = n1984 | n1987 ;
  assign n1989 = ~x132 & n1988 ;
  assign n1990 = ( n1981 & ~x133 ) | ( n1981 & n1989 ) | ( ~x133 & n1989 ) ;
  assign n1991 = n1973 | n1990 ;
  assign n1992 = ~x134 & n1991 ;
  assign n1993 = n1956 | n1992 ;
  assign n1994 = ( n831 & ~n1260 ) | ( n831 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n1995 = n876 &  n1265 ;
  assign n1996 = ( n840 & ~n1262 ) | ( n840 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n1997 = ( n844 & ~n1267 ) | ( n844 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n1998 = ( n1996 & ~n1995 ) | ( n1996 & n1997 ) | ( ~n1995 & n1997 ) ;
  assign n1999 = ( n1995 & ~n1994 ) | ( n1995 & n1998 ) | ( ~n1994 & n1998 ) ;
  assign n2000 = n1994 | n1999 ;
  assign n2001 = x132 &  n2000 ;
  assign n2002 = ( n935 & ~n1260 ) | ( n935 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n2003 = n835 &  n1265 ;
  assign n2004 = ( n944 & ~n1262 ) | ( n944 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n2005 = ( n948 & ~n1267 ) | ( n948 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n2006 = ( n2004 & ~n2003 ) | ( n2004 & n2005 ) | ( ~n2003 & n2005 ) ;
  assign n2007 = ( n2003 & ~n2002 ) | ( n2003 & n2006 ) | ( ~n2002 & n2006 ) ;
  assign n2008 = n2002 | n2007 ;
  assign n2009 = ~x132 & n2008 ;
  assign n2010 = ( n2001 & ~x133 ) | ( n2001 & n2009 ) | ( ~x133 & n2009 ) ;
  assign n2011 = ( n872 & ~n1260 ) | ( n872 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n2012 = n896 &  n1265 ;
  assign n2013 = ( n881 & ~n1262 ) | ( n881 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n2014 = ( n885 & ~n1267 ) | ( n885 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n2015 = ( n2013 & ~n2012 ) | ( n2013 & n2014 ) | ( ~n2012 & n2014 ) ;
  assign n2016 = ( n2012 & ~n2011 ) | ( n2012 & n2015 ) | ( ~n2011 & n2015 ) ;
  assign n2017 = n2011 | n2016 ;
  assign n2018 = ~x132 & n2017 ;
  assign n2019 = ( n892 & ~n1260 ) | ( n892 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n2020 = n855 &  n1265 ;
  assign n2021 = ( n901 & ~n1262 ) | ( n901 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n2022 = ( n905 & ~n1267 ) | ( n905 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n2023 = ( n2021 & ~n2020 ) | ( n2021 & n2022 ) | ( ~n2020 & n2022 ) ;
  assign n2024 = ( n2020 & ~n2019 ) | ( n2020 & n2023 ) | ( ~n2019 & n2023 ) ;
  assign n2025 = n2019 | n2024 ;
  assign n2026 = x132 &  n2025 ;
  assign n2027 = ( x133 & n2018 ) | ( x133 & n2026 ) | ( n2018 & n2026 ) ;
  assign n2028 = n2010 | n2027 ;
  assign n2029 = x134 &  n2028 ;
  assign n2030 = ( n956 & ~n1260 ) | ( n956 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n2031 = n919 &  n1265 ;
  assign n2032 = ( n965 & ~n1262 ) | ( n965 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n2033 = ( n969 & ~n1267 ) | ( n969 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n2034 = ( n2032 & ~n2031 ) | ( n2032 & n2033 ) | ( ~n2031 & n2033 ) ;
  assign n2035 = ( n2031 & ~n2030 ) | ( n2031 & n2034 ) | ( ~n2030 & n2034 ) ;
  assign n2036 = n2030 | n2035 ;
  assign n2037 = ~x132 & n2036 ;
  assign n2038 = ( n915 & ~n1260 ) | ( n915 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n2039 = n939 &  n1265 ;
  assign n2040 = ( n924 & ~n1262 ) | ( n924 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n2041 = ( n928 & ~n1267 ) | ( n928 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n2042 = ( n2040 & ~n2039 ) | ( n2040 & n2041 ) | ( ~n2039 & n2041 ) ;
  assign n2043 = ( n2039 & ~n2038 ) | ( n2039 & n2042 ) | ( ~n2038 & n2042 ) ;
  assign n2044 = n2038 | n2043 ;
  assign n2045 = x132 &  n2044 ;
  assign n2046 = ( x133 & n2037 ) | ( x133 & n2045 ) | ( n2037 & n2045 ) ;
  assign n2047 = ( n976 & ~n1260 ) | ( n976 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n2048 = n960 &  n1265 ;
  assign n2049 = ( n985 & ~n1262 ) | ( n985 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n2050 = ( n989 & ~n1267 ) | ( n989 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n2051 = ( n2049 & ~n2048 ) | ( n2049 & n2050 ) | ( ~n2048 & n2050 ) ;
  assign n2052 = ( n2048 & ~n2047 ) | ( n2048 & n2051 ) | ( ~n2047 & n2051 ) ;
  assign n2053 = n2047 | n2052 ;
  assign n2054 = x132 &  n2053 ;
  assign n2055 = ( n851 & ~n1260 ) | ( n851 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n2056 = n980 &  n1265 ;
  assign n2057 = ( n860 & ~n1262 ) | ( n860 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n2058 = ( n864 & ~n1267 ) | ( n864 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n2059 = ( n2057 & ~n2056 ) | ( n2057 & n2058 ) | ( ~n2056 & n2058 ) ;
  assign n2060 = ( n2056 & ~n2055 ) | ( n2056 & n2059 ) | ( ~n2055 & n2059 ) ;
  assign n2061 = n2055 | n2060 ;
  assign n2062 = ~x132 & n2061 ;
  assign n2063 = ( n2054 & ~x133 ) | ( n2054 & n2062 ) | ( ~x133 & n2062 ) ;
  assign n2064 = n2046 | n2063 ;
  assign n2065 = ~x134 & n2064 ;
  assign n2066 = n2029 | n2065 ;
  assign n2067 = ( n1032 & ~n1260 ) | ( n1032 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n2068 = ( n1047 & ~n1262 ) | ( n1047 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n2069 = n2067 | n2068 ;
  assign n2070 = n1007 &  n1265 ;
  assign n2071 = ( n1054 & ~n1267 ) | ( n1054 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n2072 = n2070 | n2071 ;
  assign n2073 = n2069 | n2072 ;
  assign n2074 = x132 &  n2073 ;
  assign n2075 = ( n1229 & ~n1260 ) | ( n1229 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n2076 = ( n1244 & ~n1262 ) | ( n1244 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n2077 = n2075 | n2076 ;
  assign n2078 = n1039 &  n1265 ;
  assign n2079 = ( n1251 & ~n1267 ) | ( n1251 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n2080 = n2078 | n2079 ;
  assign n2081 = n2077 | n2080 ;
  assign n2082 = ~x132 & n2081 ;
  assign n2083 = ( n2074 & ~x133 ) | ( n2074 & n2082 ) | ( ~x133 & n2082 ) ;
  assign n2084 = ( n1000 & ~n1260 ) | ( n1000 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n2085 = ( n1015 & ~n1262 ) | ( n1015 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n2086 = n2084 | n2085 ;
  assign n2087 = n1072 &  n1265 ;
  assign n2088 = ( n1022 & ~n1267 ) | ( n1022 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n2089 = n2087 | n2088 ;
  assign n2090 = n2086 | n2089 ;
  assign n2091 = ~x132 & n2090 ;
  assign n2092 = ( n1065 & ~n1260 ) | ( n1065 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n2093 = ( n1080 & ~n1262 ) | ( n1080 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n2094 = n2092 | n2093 ;
  assign n2095 = n1104 &  n1265 ;
  assign n2096 = ( n1087 & ~n1267 ) | ( n1087 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n2097 = n2095 | n2096 ;
  assign n2098 = n2094 | n2097 ;
  assign n2099 = x132 &  n2098 ;
  assign n2100 = ( x133 & n2091 ) | ( x133 & n2099 ) | ( n2091 & n2099 ) ;
  assign n2101 = n2083 | n2100 ;
  assign n2102 = x134 &  n2101 ;
  assign n2103 = ( n1132 & ~n1260 ) | ( n1132 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n2104 = ( n1147 & ~n1262 ) | ( n1147 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n2105 = n2103 | n2104 ;
  assign n2106 = n1171 &  n1265 ;
  assign n2107 = ( n1154 & ~n1267 ) | ( n1154 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n2108 = n2106 | n2107 ;
  assign n2109 = n2105 | n2108 ;
  assign n2110 = ~x132 & n2109 ;
  assign n2111 = ( n1164 & ~n1260 ) | ( n1164 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n2112 = ( n1179 & ~n1262 ) | ( n1179 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n2113 = n2111 | n2112 ;
  assign n2114 = n1236 &  n1265 ;
  assign n2115 = ( n1186 & ~n1267 ) | ( n1186 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n2116 = n2114 | n2115 ;
  assign n2117 = n2113 | n2116 ;
  assign n2118 = x132 &  n2117 ;
  assign n2119 = ( x133 & n2110 ) | ( x133 & n2118 ) | ( n2110 & n2118 ) ;
  assign n2120 = ( n1197 & ~n1260 ) | ( n1197 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n2121 = ( n1212 & ~n1262 ) | ( n1212 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n2122 = n2120 | n2121 ;
  assign n2123 = n1139 &  n1265 ;
  assign n2124 = ( n1219 & ~n1267 ) | ( n1219 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n2125 = n2123 | n2124 ;
  assign n2126 = n2122 | n2125 ;
  assign n2127 = x132 &  n2126 ;
  assign n2128 = ( n1097 & ~n1260 ) | ( n1097 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n2129 = ( n1112 & ~n1262 ) | ( n1112 & 1'b0 ) | ( ~n1262 & 1'b0 ) ;
  assign n2130 = n2128 | n2129 ;
  assign n2131 = n1204 &  n1265 ;
  assign n2132 = ( n1119 & ~n1267 ) | ( n1119 & 1'b0 ) | ( ~n1267 & 1'b0 ) ;
  assign n2133 = n2131 | n2132 ;
  assign n2134 = n2130 | n2133 ;
  assign n2135 = ~x132 & n2134 ;
  assign n2136 = ( n2127 & ~x133 ) | ( n2127 & n2135 ) | ( ~x133 & n2135 ) ;
  assign n2137 = n2119 | n2136 ;
  assign n2138 = ~x134 & n2137 ;
  assign n2139 = n2102 | n2138 ;
  assign n2140 = ( n357 & ~n436 ) | ( n357 & 1'b0 ) | ( ~n436 & 1'b0 ) ;
  assign n2141 = n170 &  n485 ;
  assign n2142 = n2140 | n2141 ;
  assign n2143 = ( n282 & ~n535 ) | ( n282 & 1'b0 ) | ( ~n535 & 1'b0 ) ;
  assign n2144 = ( n246 & ~n580 ) | ( n246 & 1'b0 ) | ( ~n580 & 1'b0 ) ;
  assign n2145 = ( n2143 & ~n2142 ) | ( n2143 & n2144 ) | ( ~n2142 & n2144 ) ;
  assign n2146 = n2142 | n2145 ;
  assign n2147 = x134 &  n2146 ;
  assign n2148 = n321 &  n485 ;
  assign n2149 = ( n206 & ~n436 ) | ( n206 & 1'b0 ) | ( ~n436 & 1'b0 ) ;
  assign n2150 = ( n394 & ~n580 ) | ( n394 & 1'b0 ) | ( ~n580 & 1'b0 ) ;
  assign n2151 = ( n430 & ~n535 ) | ( n430 & 1'b0 ) | ( ~n535 & 1'b0 ) ;
  assign n2152 = ( n2150 & ~n2149 ) | ( n2150 & n2151 ) | ( ~n2149 & n2151 ) ;
  assign n2153 = ( n2149 & ~n2148 ) | ( n2149 & n2152 ) | ( ~n2148 & n2152 ) ;
  assign n2154 = n2148 | n2153 ;
  assign n2155 = ~x134 & n2154 ;
  assign n2156 = n2147 | n2155 ;
  assign n2157 = ( n483 & ~n535 ) | ( n483 & 1'b0 ) | ( ~n535 & 1'b0 ) ;
  assign n2158 = ~n436 & n726 ;
  assign n2159 = n2157 | n2158 ;
  assign n2160 = ( n578 & ~n580 ) | ( n578 & 1'b0 ) | ( ~n580 & 1'b0 ) ;
  assign n2161 = n485 &  n627 ;
  assign n2162 = n2160 | n2161 ;
  assign n2163 = n2159 | n2162 ;
  assign n2164 = x134 &  n2163 ;
  assign n2165 = n485 &  n678 ;
  assign n2166 = ~n580 & n775 ;
  assign n2167 = n2165 | n2166 ;
  assign n2168 = ~n436 & n532 ;
  assign n2169 = ~n535 & n823 ;
  assign n2170 = n2168 | n2169 ;
  assign n2171 = n2167 | n2170 ;
  assign n2172 = ~x134 & n2171 ;
  assign n2173 = n2164 | n2172 ;
  assign n2174 = ~n535 & n847 ;
  assign n2175 = ~n580 & n888 ;
  assign n2176 = ~n436 & n951 ;
  assign n2177 = n485 &  n908 ;
  assign n2178 = ( n2176 & ~n2175 ) | ( n2176 & n2177 ) | ( ~n2175 & n2177 ) ;
  assign n2179 = ( n2175 & ~n2174 ) | ( n2175 & n2178 ) | ( ~n2174 & n2178 ) ;
  assign n2180 = n2174 | n2179 ;
  assign n2181 = x134 &  n2180 ;
  assign n2182 = n485 &  n931 ;
  assign n2183 = ~n436 & n867 ;
  assign n2184 = ~n580 & n972 ;
  assign n2185 = ~n535 & n992 ;
  assign n2186 = ( n2184 & ~n2183 ) | ( n2184 & n2185 ) | ( ~n2183 & n2185 ) ;
  assign n2187 = ( n2183 & ~n2182 ) | ( n2183 & n2186 ) | ( ~n2182 & n2186 ) ;
  assign n2188 = n2182 | n2187 ;
  assign n2189 = ~x134 & n2188 ;
  assign n2190 = n2181 | n2189 ;
  assign n2191 = ~n535 & n1057 ;
  assign n2192 = ~n436 & n1254 ;
  assign n2193 = n2191 | n2192 ;
  assign n2194 = n485 &  n1090 ;
  assign n2195 = ~n580 & n1025 ;
  assign n2196 = n2194 | n2195 ;
  assign n2197 = n2193 | n2196 ;
  assign n2198 = x134 &  n2197 ;
  assign n2199 = ~n580 & n1157 ;
  assign n2200 = n485 &  n1189 ;
  assign n2201 = n2199 | n2200 ;
  assign n2202 = ~n535 & n1222 ;
  assign n2203 = ~n436 & n1122 ;
  assign n2204 = n2202 | n2203 ;
  assign n2205 = n2201 | n2204 ;
  assign n2206 = ~x134 & n2205 ;
  assign n2207 = n2198 | n2206 ;
  assign n2208 = ~n436 & n1314 ;
  assign n2209 = ~n580 & n1270 ;
  assign n2210 = n2208 | n2209 ;
  assign n2211 = n485 &  n1287 ;
  assign n2212 = ~n535 & n1278 ;
  assign n2213 = n2211 | n2212 ;
  assign n2214 = n2210 | n2213 ;
  assign n2215 = x134 &  n2214 ;
  assign n2216 = n485 &  n1306 ;
  assign n2217 = ~n580 & n1323 ;
  assign n2218 = n2216 | n2217 ;
  assign n2219 = ~n436 & n1295 ;
  assign n2220 = ~n535 & n1331 ;
  assign n2221 = n2219 | n2220 ;
  assign n2222 = n2218 | n2221 ;
  assign n2223 = ~x134 & n2222 ;
  assign n2224 = n2215 | n2223 ;
  assign n2225 = ~n436 & n1387 ;
  assign n2226 = ~n580 & n1343 ;
  assign n2227 = n2225 | n2226 ;
  assign n2228 = n485 &  n1360 ;
  assign n2229 = ~n535 & n1351 ;
  assign n2230 = n2228 | n2229 ;
  assign n2231 = n2227 | n2230 ;
  assign n2232 = x134 &  n2231 ;
  assign n2233 = n485 &  n1379 ;
  assign n2234 = ~n580 & n1396 ;
  assign n2235 = n2233 | n2234 ;
  assign n2236 = ~n436 & n1368 ;
  assign n2237 = ~n535 & n1404 ;
  assign n2238 = n2236 | n2237 ;
  assign n2239 = n2235 | n2238 ;
  assign n2240 = ~x134 & n2239 ;
  assign n2241 = n2232 | n2240 ;
  assign n2242 = ~n436 & n1460 ;
  assign n2243 = ~n580 & n1416 ;
  assign n2244 = n2242 | n2243 ;
  assign n2245 = n485 &  n1433 ;
  assign n2246 = ~n535 & n1424 ;
  assign n2247 = n2245 | n2246 ;
  assign n2248 = n2244 | n2247 ;
  assign n2249 = x134 &  n2248 ;
  assign n2250 = n485 &  n1452 ;
  assign n2251 = ~n580 & n1469 ;
  assign n2252 = n2250 | n2251 ;
  assign n2253 = ~n436 & n1441 ;
  assign n2254 = ~n535 & n1477 ;
  assign n2255 = n2253 | n2254 ;
  assign n2256 = n2252 | n2255 ;
  assign n2257 = ~x134 & n2256 ;
  assign n2258 = n2249 | n2257 ;
  assign n2259 = ~n580 & n1489 ;
  assign n2260 = ~n535 & n1497 ;
  assign n2261 = n2259 | n2260 ;
  assign n2262 = n485 &  n1506 ;
  assign n2263 = ~n436 & n1533 ;
  assign n2264 = n2262 | n2263 ;
  assign n2265 = n2261 | n2264 ;
  assign n2266 = x134 &  n2265 ;
  assign n2267 = n485 &  n1525 ;
  assign n2268 = ~n436 & n1514 ;
  assign n2269 = n2267 | n2268 ;
  assign n2270 = ~n535 & n1550 ;
  assign n2271 = ~n580 & n1542 ;
  assign n2272 = n2270 | n2271 ;
  assign n2273 = n2269 | n2272 ;
  assign n2274 = ~x134 & n2273 ;
  assign n2275 = n2266 | n2274 ;
  assign n2276 = ~n580 & n1562 ;
  assign n2277 = ~n535 & n1570 ;
  assign n2278 = n2276 | n2277 ;
  assign n2279 = n485 &  n1579 ;
  assign n2280 = ~n436 & n1606 ;
  assign n2281 = n2279 | n2280 ;
  assign n2282 = n2278 | n2281 ;
  assign n2283 = x134 &  n2282 ;
  assign n2284 = n485 &  n1598 ;
  assign n2285 = ~n436 & n1587 ;
  assign n2286 = n2284 | n2285 ;
  assign n2287 = ~n535 & n1623 ;
  assign n2288 = ~n580 & n1615 ;
  assign n2289 = n2287 | n2288 ;
  assign n2290 = n2286 | n2289 ;
  assign n2291 = ~x134 & n2290 ;
  assign n2292 = n2283 | n2291 ;
  assign n2293 = ~n580 & n1635 ;
  assign n2294 = ~n535 & n1643 ;
  assign n2295 = n2293 | n2294 ;
  assign n2296 = n485 &  n1652 ;
  assign n2297 = ~n436 & n1679 ;
  assign n2298 = n2296 | n2297 ;
  assign n2299 = n2295 | n2298 ;
  assign n2300 = x134 &  n2299 ;
  assign n2301 = n485 &  n1671 ;
  assign n2302 = ~n436 & n1660 ;
  assign n2303 = n2301 | n2302 ;
  assign n2304 = ~n535 & n1696 ;
  assign n2305 = ~n580 & n1688 ;
  assign n2306 = n2304 | n2305 ;
  assign n2307 = n2303 | n2306 ;
  assign n2308 = ~x134 & n2307 ;
  assign n2309 = n2300 | n2308 ;
  assign n2310 = ~n580 & n1708 ;
  assign n2311 = ~n535 & n1716 ;
  assign n2312 = n2310 | n2311 ;
  assign n2313 = n485 &  n1725 ;
  assign n2314 = ~n436 & n1752 ;
  assign n2315 = n2313 | n2314 ;
  assign n2316 = n2312 | n2315 ;
  assign n2317 = x134 &  n2316 ;
  assign n2318 = n485 &  n1744 ;
  assign n2319 = ~n580 & n1761 ;
  assign n2320 = n2318 | n2319 ;
  assign n2321 = ~n436 & n1733 ;
  assign n2322 = ~n535 & n1769 ;
  assign n2323 = n2321 | n2322 ;
  assign n2324 = n2320 | n2323 ;
  assign n2325 = ~x134 & n2324 ;
  assign n2326 = n2317 | n2325 ;
  assign n2327 = ~n580 & n1781 ;
  assign n2328 = ~n535 & n1789 ;
  assign n2329 = n2327 | n2328 ;
  assign n2330 = n485 &  n1798 ;
  assign n2331 = ~n436 & n1825 ;
  assign n2332 = n2330 | n2331 ;
  assign n2333 = n2329 | n2332 ;
  assign n2334 = x134 &  n2333 ;
  assign n2335 = n485 &  n1817 ;
  assign n2336 = ~n580 & n1834 ;
  assign n2337 = n2335 | n2336 ;
  assign n2338 = ~n436 & n1806 ;
  assign n2339 = ~n535 & n1842 ;
  assign n2340 = n2338 | n2339 ;
  assign n2341 = n2337 | n2340 ;
  assign n2342 = ~x134 & n2341 ;
  assign n2343 = n2334 | n2342 ;
  assign n2344 = ~n580 & n1854 ;
  assign n2345 = ~n535 & n1862 ;
  assign n2346 = n2344 | n2345 ;
  assign n2347 = n485 &  n1871 ;
  assign n2348 = ~n436 & n1898 ;
  assign n2349 = n2347 | n2348 ;
  assign n2350 = n2346 | n2349 ;
  assign n2351 = x134 &  n2350 ;
  assign n2352 = n485 &  n1890 ;
  assign n2353 = ~n580 & n1907 ;
  assign n2354 = n2352 | n2353 ;
  assign n2355 = ~n436 & n1879 ;
  assign n2356 = ~n535 & n1915 ;
  assign n2357 = n2355 | n2356 ;
  assign n2358 = n2354 | n2357 ;
  assign n2359 = ~x134 & n2358 ;
  assign n2360 = n2351 | n2359 ;
  assign n2361 = ~n580 & n1927 ;
  assign n2362 = ~n535 & n1935 ;
  assign n2363 = n2361 | n2362 ;
  assign n2364 = n485 &  n1944 ;
  assign n2365 = ~n436 & n1971 ;
  assign n2366 = n2364 | n2365 ;
  assign n2367 = n2363 | n2366 ;
  assign n2368 = x134 &  n2367 ;
  assign n2369 = n485 &  n1963 ;
  assign n2370 = ~n580 & n1980 ;
  assign n2371 = n2369 | n2370 ;
  assign n2372 = ~n436 & n1952 ;
  assign n2373 = ~n535 & n1988 ;
  assign n2374 = n2372 | n2373 ;
  assign n2375 = n2371 | n2374 ;
  assign n2376 = ~x134 & n2375 ;
  assign n2377 = n2368 | n2376 ;
  assign n2378 = ~n580 & n2000 ;
  assign n2379 = ~n535 & n2008 ;
  assign n2380 = n2378 | n2379 ;
  assign n2381 = n485 &  n2017 ;
  assign n2382 = ~n436 & n2044 ;
  assign n2383 = n2381 | n2382 ;
  assign n2384 = n2380 | n2383 ;
  assign n2385 = x134 &  n2384 ;
  assign n2386 = n485 &  n2036 ;
  assign n2387 = ~n580 & n2053 ;
  assign n2388 = n2386 | n2387 ;
  assign n2389 = ~n436 & n2025 ;
  assign n2390 = ~n535 & n2061 ;
  assign n2391 = n2389 | n2390 ;
  assign n2392 = n2388 | n2391 ;
  assign n2393 = ~x134 & n2392 ;
  assign n2394 = n2385 | n2393 ;
  assign n2395 = ~n580 & n2073 ;
  assign n2396 = ~n535 & n2081 ;
  assign n2397 = n2395 | n2396 ;
  assign n2398 = n485 &  n2090 ;
  assign n2399 = ~n436 & n2117 ;
  assign n2400 = n2398 | n2399 ;
  assign n2401 = n2397 | n2400 ;
  assign n2402 = x134 &  n2401 ;
  assign n2403 = n485 &  n2109 ;
  assign n2404 = ~n580 & n2126 ;
  assign n2405 = n2403 | n2404 ;
  assign n2406 = ~n436 & n2098 ;
  assign n2407 = ~n535 & n2134 ;
  assign n2408 = n2406 | n2407 ;
  assign n2409 = n2405 | n2408 ;
  assign n2410 = ~x134 & n2409 ;
  assign n2411 = n2402 | n2410 ;
  assign n2412 = ( n357 & ~n535 ) | ( n357 & 1'b0 ) | ( ~n535 & 1'b0 ) ;
  assign n2413 = ( n321 & ~n436 ) | ( n321 & 1'b0 ) | ( ~n436 & 1'b0 ) ;
  assign n2414 = n2412 | n2413 ;
  assign n2415 = ( n282 & ~n580 ) | ( n282 & 1'b0 ) | ( ~n580 & 1'b0 ) ;
  assign n2416 = n246 &  n485 ;
  assign n2417 = ( n2415 & ~n2414 ) | ( n2415 & n2416 ) | ( ~n2414 & n2416 ) ;
  assign n2418 = n2414 | n2417 ;
  assign n2419 = x134 &  n2418 ;
  assign n2420 = n394 &  n485 ;
  assign n2421 = ( n170 & ~n436 ) | ( n170 & 1'b0 ) | ( ~n436 & 1'b0 ) ;
  assign n2422 = ( n430 & ~n580 ) | ( n430 & 1'b0 ) | ( ~n580 & 1'b0 ) ;
  assign n2423 = ( n206 & ~n535 ) | ( n206 & 1'b0 ) | ( ~n535 & 1'b0 ) ;
  assign n2424 = ( n2422 & ~n2421 ) | ( n2422 & n2423 ) | ( ~n2421 & n2423 ) ;
  assign n2425 = ( n2421 & ~n2420 ) | ( n2421 & n2424 ) | ( ~n2420 & n2424 ) ;
  assign n2426 = n2420 | n2425 ;
  assign n2427 = ~x134 & n2426 ;
  assign n2428 = n2419 | n2427 ;
  assign n2429 = ( n483 & ~n580 ) | ( n483 & 1'b0 ) | ( ~n580 & 1'b0 ) ;
  assign n2430 = ~n535 & n726 ;
  assign n2431 = n2429 | n2430 ;
  assign n2432 = n485 &  n578 ;
  assign n2433 = ~n436 & n678 ;
  assign n2434 = n2432 | n2433 ;
  assign n2435 = n2431 | n2434 ;
  assign n2436 = x134 &  n2435 ;
  assign n2437 = n485 &  n775 ;
  assign n2438 = ~n580 & n823 ;
  assign n2439 = n2437 | n2438 ;
  assign n2440 = ~n436 & n627 ;
  assign n2441 = ( n532 & ~n535 ) | ( n532 & 1'b0 ) | ( ~n535 & 1'b0 ) ;
  assign n2442 = n2440 | n2441 ;
  assign n2443 = n2439 | n2442 ;
  assign n2444 = ~x134 & n2443 ;
  assign n2445 = n2436 | n2444 ;
  assign n2446 = ~n580 & n847 ;
  assign n2447 = n485 &  n888 ;
  assign n2448 = ~n535 & n951 ;
  assign n2449 = ~n436 & n931 ;
  assign n2450 = ( n2448 & ~n2447 ) | ( n2448 & n2449 ) | ( ~n2447 & n2449 ) ;
  assign n2451 = ( n2447 & ~n2446 ) | ( n2447 & n2450 ) | ( ~n2446 & n2450 ) ;
  assign n2452 = n2446 | n2451 ;
  assign n2453 = x134 &  n2452 ;
  assign n2454 = n485 &  n972 ;
  assign n2455 = ~n436 & n908 ;
  assign n2456 = ~n580 & n992 ;
  assign n2457 = ~n535 & n867 ;
  assign n2458 = ( n2456 & ~n2455 ) | ( n2456 & n2457 ) | ( ~n2455 & n2457 ) ;
  assign n2459 = ( n2455 & ~n2454 ) | ( n2455 & n2458 ) | ( ~n2454 & n2458 ) ;
  assign n2460 = n2454 | n2459 ;
  assign n2461 = ~x134 & n2460 ;
  assign n2462 = n2453 | n2461 ;
  assign n2463 = ~n580 & n1057 ;
  assign n2464 = ~n436 & n1189 ;
  assign n2465 = n2463 | n2464 ;
  assign n2466 = n485 &  n1025 ;
  assign n2467 = ~n535 & n1254 ;
  assign n2468 = n2466 | n2467 ;
  assign n2469 = n2465 | n2468 ;
  assign n2470 = x134 &  n2469 ;
  assign n2471 = n485 &  n1157 ;
  assign n2472 = ~n436 & n1090 ;
  assign n2473 = n2471 | n2472 ;
  assign n2474 = ~n580 & n1222 ;
  assign n2475 = ~n535 & n1122 ;
  assign n2476 = n2474 | n2475 ;
  assign n2477 = n2473 | n2476 ;
  assign n2478 = ~x134 & n2477 ;
  assign n2479 = n2470 | n2478 ;
  assign n2480 = ~n535 & n1314 ;
  assign n2481 = ~n436 & n1306 ;
  assign n2482 = n2480 | n2481 ;
  assign n2483 = ~n580 & n1278 ;
  assign n2484 = n485 &  n1270 ;
  assign n2485 = n2483 | n2484 ;
  assign n2486 = n2482 | n2485 ;
  assign n2487 = x134 &  n2486 ;
  assign n2488 = n485 &  n1323 ;
  assign n2489 = ~n580 & n1331 ;
  assign n2490 = n2488 | n2489 ;
  assign n2491 = ~n436 & n1287 ;
  assign n2492 = ~n535 & n1295 ;
  assign n2493 = n2491 | n2492 ;
  assign n2494 = n2490 | n2493 ;
  assign n2495 = ~x134 & n2494 ;
  assign n2496 = n2487 | n2495 ;
  assign n2497 = ~n535 & n1387 ;
  assign n2498 = ~n436 & n1379 ;
  assign n2499 = n2497 | n2498 ;
  assign n2500 = ~n580 & n1351 ;
  assign n2501 = n485 &  n1343 ;
  assign n2502 = n2500 | n2501 ;
  assign n2503 = n2499 | n2502 ;
  assign n2504 = x134 &  n2503 ;
  assign n2505 = n485 &  n1396 ;
  assign n2506 = ~n580 & n1404 ;
  assign n2507 = n2505 | n2506 ;
  assign n2508 = ~n436 & n1360 ;
  assign n2509 = ~n535 & n1368 ;
  assign n2510 = n2508 | n2509 ;
  assign n2511 = n2507 | n2510 ;
  assign n2512 = ~x134 & n2511 ;
  assign n2513 = n2504 | n2512 ;
  assign n2514 = ~n535 & n1460 ;
  assign n2515 = ~n436 & n1452 ;
  assign n2516 = n2514 | n2515 ;
  assign n2517 = ~n580 & n1424 ;
  assign n2518 = n485 &  n1416 ;
  assign n2519 = n2517 | n2518 ;
  assign n2520 = n2516 | n2519 ;
  assign n2521 = x134 &  n2520 ;
  assign n2522 = n485 &  n1469 ;
  assign n2523 = ~n580 & n1477 ;
  assign n2524 = n2522 | n2523 ;
  assign n2525 = ~n436 & n1433 ;
  assign n2526 = ~n535 & n1441 ;
  assign n2527 = n2525 | n2526 ;
  assign n2528 = n2524 | n2527 ;
  assign n2529 = ~x134 & n2528 ;
  assign n2530 = n2521 | n2529 ;
  assign n2531 = n485 &  n1489 ;
  assign n2532 = ~n580 & n1497 ;
  assign n2533 = n2531 | n2532 ;
  assign n2534 = ~n436 & n1525 ;
  assign n2535 = ~n535 & n1533 ;
  assign n2536 = n2534 | n2535 ;
  assign n2537 = n2533 | n2536 ;
  assign n2538 = x134 &  n2537 ;
  assign n2539 = ~n535 & n1514 ;
  assign n2540 = ~n436 & n1506 ;
  assign n2541 = n2539 | n2540 ;
  assign n2542 = ~n580 & n1550 ;
  assign n2543 = n485 &  n1542 ;
  assign n2544 = n2542 | n2543 ;
  assign n2545 = n2541 | n2544 ;
  assign n2546 = ~x134 & n2545 ;
  assign n2547 = n2538 | n2546 ;
  assign n2548 = n485 &  n1562 ;
  assign n2549 = ~n580 & n1570 ;
  assign n2550 = n2548 | n2549 ;
  assign n2551 = ~n436 & n1598 ;
  assign n2552 = ~n535 & n1606 ;
  assign n2553 = n2551 | n2552 ;
  assign n2554 = n2550 | n2553 ;
  assign n2555 = x134 &  n2554 ;
  assign n2556 = ~n535 & n1587 ;
  assign n2557 = ~n436 & n1579 ;
  assign n2558 = n2556 | n2557 ;
  assign n2559 = ~n580 & n1623 ;
  assign n2560 = n485 &  n1615 ;
  assign n2561 = n2559 | n2560 ;
  assign n2562 = n2558 | n2561 ;
  assign n2563 = ~x134 & n2562 ;
  assign n2564 = n2555 | n2563 ;
  assign n2565 = n485 &  n1635 ;
  assign n2566 = ~n580 & n1643 ;
  assign n2567 = n2565 | n2566 ;
  assign n2568 = ~n436 & n1671 ;
  assign n2569 = ~n535 & n1679 ;
  assign n2570 = n2568 | n2569 ;
  assign n2571 = n2567 | n2570 ;
  assign n2572 = x134 &  n2571 ;
  assign n2573 = ~n535 & n1660 ;
  assign n2574 = ~n436 & n1652 ;
  assign n2575 = n2573 | n2574 ;
  assign n2576 = ~n580 & n1696 ;
  assign n2577 = n485 &  n1688 ;
  assign n2578 = n2576 | n2577 ;
  assign n2579 = n2575 | n2578 ;
  assign n2580 = ~x134 & n2579 ;
  assign n2581 = n2572 | n2580 ;
  assign n2582 = n485 &  n1708 ;
  assign n2583 = ~n580 & n1716 ;
  assign n2584 = n2582 | n2583 ;
  assign n2585 = ~n436 & n1744 ;
  assign n2586 = ~n535 & n1752 ;
  assign n2587 = n2585 | n2586 ;
  assign n2588 = n2584 | n2587 ;
  assign n2589 = x134 &  n2588 ;
  assign n2590 = n485 &  n1761 ;
  assign n2591 = ~n580 & n1769 ;
  assign n2592 = n2590 | n2591 ;
  assign n2593 = ~n436 & n1725 ;
  assign n2594 = ~n535 & n1733 ;
  assign n2595 = n2593 | n2594 ;
  assign n2596 = n2592 | n2595 ;
  assign n2597 = ~x134 & n2596 ;
  assign n2598 = n2589 | n2597 ;
  assign n2599 = n485 &  n1781 ;
  assign n2600 = ~n580 & n1789 ;
  assign n2601 = n2599 | n2600 ;
  assign n2602 = ~n436 & n1817 ;
  assign n2603 = ~n535 & n1825 ;
  assign n2604 = n2602 | n2603 ;
  assign n2605 = n2601 | n2604 ;
  assign n2606 = x134 &  n2605 ;
  assign n2607 = n485 &  n1834 ;
  assign n2608 = ~n580 & n1842 ;
  assign n2609 = n2607 | n2608 ;
  assign n2610 = ~n436 & n1798 ;
  assign n2611 = ~n535 & n1806 ;
  assign n2612 = n2610 | n2611 ;
  assign n2613 = n2609 | n2612 ;
  assign n2614 = ~x134 & n2613 ;
  assign n2615 = n2606 | n2614 ;
  assign n2616 = n485 &  n1854 ;
  assign n2617 = ~n580 & n1862 ;
  assign n2618 = n2616 | n2617 ;
  assign n2619 = ~n436 & n1890 ;
  assign n2620 = ~n535 & n1898 ;
  assign n2621 = n2619 | n2620 ;
  assign n2622 = n2618 | n2621 ;
  assign n2623 = x134 &  n2622 ;
  assign n2624 = n485 &  n1907 ;
  assign n2625 = ~n580 & n1915 ;
  assign n2626 = n2624 | n2625 ;
  assign n2627 = ~n436 & n1871 ;
  assign n2628 = ~n535 & n1879 ;
  assign n2629 = n2627 | n2628 ;
  assign n2630 = n2626 | n2629 ;
  assign n2631 = ~x134 & n2630 ;
  assign n2632 = n2623 | n2631 ;
  assign n2633 = n485 &  n1927 ;
  assign n2634 = ~n580 & n1935 ;
  assign n2635 = n2633 | n2634 ;
  assign n2636 = ~n436 & n1963 ;
  assign n2637 = ~n535 & n1971 ;
  assign n2638 = n2636 | n2637 ;
  assign n2639 = n2635 | n2638 ;
  assign n2640 = x134 &  n2639 ;
  assign n2641 = n485 &  n1980 ;
  assign n2642 = ~n580 & n1988 ;
  assign n2643 = n2641 | n2642 ;
  assign n2644 = ~n436 & n1944 ;
  assign n2645 = ~n535 & n1952 ;
  assign n2646 = n2644 | n2645 ;
  assign n2647 = n2643 | n2646 ;
  assign n2648 = ~x134 & n2647 ;
  assign n2649 = n2640 | n2648 ;
  assign n2650 = n485 &  n2000 ;
  assign n2651 = ~n580 & n2008 ;
  assign n2652 = n2650 | n2651 ;
  assign n2653 = ~n436 & n2036 ;
  assign n2654 = ~n535 & n2044 ;
  assign n2655 = n2653 | n2654 ;
  assign n2656 = n2652 | n2655 ;
  assign n2657 = x134 &  n2656 ;
  assign n2658 = n485 &  n2053 ;
  assign n2659 = ~n580 & n2061 ;
  assign n2660 = n2658 | n2659 ;
  assign n2661 = ~n436 & n2017 ;
  assign n2662 = ~n535 & n2025 ;
  assign n2663 = n2661 | n2662 ;
  assign n2664 = n2660 | n2663 ;
  assign n2665 = ~x134 & n2664 ;
  assign n2666 = n2657 | n2665 ;
  assign n2667 = n485 &  n2073 ;
  assign n2668 = ~n580 & n2081 ;
  assign n2669 = n2667 | n2668 ;
  assign n2670 = ~n436 & n2109 ;
  assign n2671 = ~n535 & n2117 ;
  assign n2672 = n2670 | n2671 ;
  assign n2673 = n2669 | n2672 ;
  assign n2674 = x134 &  n2673 ;
  assign n2675 = n485 &  n2126 ;
  assign n2676 = ~n580 & n2134 ;
  assign n2677 = n2675 | n2676 ;
  assign n2678 = ~n436 & n2090 ;
  assign n2679 = ~n535 & n2098 ;
  assign n2680 = n2678 | n2679 ;
  assign n2681 = n2677 | n2680 ;
  assign n2682 = ~x134 & n2681 ;
  assign n2683 = n2674 | n2682 ;
  assign n2684 = ( n357 & ~n580 ) | ( n357 & 1'b0 ) | ( ~n580 & 1'b0 ) ;
  assign n2685 = n282 &  n485 ;
  assign n2686 = ( n321 & ~n535 ) | ( n321 & 1'b0 ) | ( ~n535 & 1'b0 ) ;
  assign n2687 = ( n394 & ~n436 ) | ( n394 & 1'b0 ) | ( ~n436 & 1'b0 ) ;
  assign n2688 = ( n2686 & ~n2685 ) | ( n2686 & n2687 ) | ( ~n2685 & n2687 ) ;
  assign n2689 = ( n2685 & ~n2684 ) | ( n2685 & n2688 ) | ( ~n2684 & n2688 ) ;
  assign n2690 = n2684 | n2689 ;
  assign n2691 = x134 &  n2690 ;
  assign n2692 = n430 &  n485 ;
  assign n2693 = ( n206 & ~n580 ) | ( n206 & 1'b0 ) | ( ~n580 & 1'b0 ) ;
  assign n2694 = n2692 | n2693 ;
  assign n2695 = ( n246 & ~n436 ) | ( n246 & 1'b0 ) | ( ~n436 & 1'b0 ) ;
  assign n2696 = ( n170 & ~n535 ) | ( n170 & 1'b0 ) | ( ~n535 & 1'b0 ) ;
  assign n2697 = ( n2695 & ~n2694 ) | ( n2695 & n2696 ) | ( ~n2694 & n2696 ) ;
  assign n2698 = n2694 | n2697 ;
  assign n2699 = ~x134 & n2698 ;
  assign n2700 = n2691 | n2699 ;
  assign n2701 = n483 &  n485 ;
  assign n2702 = ~n580 & n726 ;
  assign n2703 = n2701 | n2702 ;
  assign n2704 = ~n436 & n775 ;
  assign n2705 = ~n535 & n678 ;
  assign n2706 = n2704 | n2705 ;
  assign n2707 = n2703 | n2706 ;
  assign n2708 = x134 &  n2707 ;
  assign n2709 = n485 &  n823 ;
  assign n2710 = ( n532 & ~n580 ) | ( n532 & 1'b0 ) | ( ~n580 & 1'b0 ) ;
  assign n2711 = n2709 | n2710 ;
  assign n2712 = ~n436 & n578 ;
  assign n2713 = ~n535 & n627 ;
  assign n2714 = n2712 | n2713 ;
  assign n2715 = n2711 | n2714 ;
  assign n2716 = ~x134 & n2715 ;
  assign n2717 = n2708 | n2716 ;
  assign n2718 = n485 &  n847 ;
  assign n2719 = ~n436 & n972 ;
  assign n2720 = ~n580 & n951 ;
  assign n2721 = ~n535 & n931 ;
  assign n2722 = ( n2720 & ~n2719 ) | ( n2720 & n2721 ) | ( ~n2719 & n2721 ) ;
  assign n2723 = ( n2719 & ~n2718 ) | ( n2719 & n2722 ) | ( ~n2718 & n2722 ) ;
  assign n2724 = n2718 | n2723 ;
  assign n2725 = x134 &  n2724 ;
  assign n2726 = n485 &  n992 ;
  assign n2727 = ~n436 & n888 ;
  assign n2728 = ~n580 & n867 ;
  assign n2729 = ~n535 & n908 ;
  assign n2730 = ( n2728 & ~n2727 ) | ( n2728 & n2729 ) | ( ~n2727 & n2729 ) ;
  assign n2731 = ( n2727 & ~n2726 ) | ( n2727 & n2730 ) | ( ~n2726 & n2730 ) ;
  assign n2732 = n2726 | n2731 ;
  assign n2733 = ~x134 & n2732 ;
  assign n2734 = n2725 | n2733 ;
  assign n2735 = n485 &  n1057 ;
  assign n2736 = ~n436 & n1157 ;
  assign n2737 = n2735 | n2736 ;
  assign n2738 = ~n580 & n1254 ;
  assign n2739 = ~n535 & n1189 ;
  assign n2740 = n2738 | n2739 ;
  assign n2741 = n2737 | n2740 ;
  assign n2742 = x134 &  n2741 ;
  assign n2743 = ~n436 & n1025 ;
  assign n2744 = ~n535 & n1090 ;
  assign n2745 = n2743 | n2744 ;
  assign n2746 = n485 &  n1222 ;
  assign n2747 = ~n580 & n1122 ;
  assign n2748 = n2746 | n2747 ;
  assign n2749 = n2745 | n2748 ;
  assign n2750 = ~x134 & n2749 ;
  assign n2751 = n2742 | n2750 ;
  assign n2752 = ~n580 & n1314 ;
  assign n2753 = ~n535 & n1306 ;
  assign n2754 = n2752 | n2753 ;
  assign n2755 = ~n436 & n1323 ;
  assign n2756 = n485 &  n1278 ;
  assign n2757 = n2755 | n2756 ;
  assign n2758 = n2754 | n2757 ;
  assign n2759 = x134 &  n2758 ;
  assign n2760 = ~n436 & n1270 ;
  assign n2761 = n485 &  n1331 ;
  assign n2762 = n2760 | n2761 ;
  assign n2763 = ~n535 & n1287 ;
  assign n2764 = ~n580 & n1295 ;
  assign n2765 = n2763 | n2764 ;
  assign n2766 = n2762 | n2765 ;
  assign n2767 = ~x134 & n2766 ;
  assign n2768 = n2759 | n2767 ;
  assign n2769 = ~n580 & n1387 ;
  assign n2770 = ~n535 & n1379 ;
  assign n2771 = n2769 | n2770 ;
  assign n2772 = ~n436 & n1396 ;
  assign n2773 = n485 &  n1351 ;
  assign n2774 = n2772 | n2773 ;
  assign n2775 = n2771 | n2774 ;
  assign n2776 = x134 &  n2775 ;
  assign n2777 = ~n436 & n1343 ;
  assign n2778 = n485 &  n1404 ;
  assign n2779 = n2777 | n2778 ;
  assign n2780 = ~n535 & n1360 ;
  assign n2781 = ~n580 & n1368 ;
  assign n2782 = n2780 | n2781 ;
  assign n2783 = n2779 | n2782 ;
  assign n2784 = ~x134 & n2783 ;
  assign n2785 = n2776 | n2784 ;
  assign n2786 = ~n580 & n1460 ;
  assign n2787 = ~n535 & n1452 ;
  assign n2788 = n2786 | n2787 ;
  assign n2789 = ~n436 & n1469 ;
  assign n2790 = n485 &  n1424 ;
  assign n2791 = n2789 | n2790 ;
  assign n2792 = n2788 | n2791 ;
  assign n2793 = x134 &  n2792 ;
  assign n2794 = ~n436 & n1416 ;
  assign n2795 = n485 &  n1477 ;
  assign n2796 = n2794 | n2795 ;
  assign n2797 = ~n535 & n1433 ;
  assign n2798 = ~n580 & n1441 ;
  assign n2799 = n2797 | n2798 ;
  assign n2800 = n2796 | n2799 ;
  assign n2801 = ~x134 & n2800 ;
  assign n2802 = n2793 | n2801 ;
  assign n2803 = n485 &  n1497 ;
  assign n2804 = ~n580 & n1533 ;
  assign n2805 = n2803 | n2804 ;
  assign n2806 = ~n436 & n1542 ;
  assign n2807 = ~n535 & n1525 ;
  assign n2808 = n2806 | n2807 ;
  assign n2809 = n2805 | n2808 ;
  assign n2810 = x134 &  n2809 ;
  assign n2811 = ~n436 & n1489 ;
  assign n2812 = ~n580 & n1514 ;
  assign n2813 = n2811 | n2812 ;
  assign n2814 = n485 &  n1550 ;
  assign n2815 = ~n535 & n1506 ;
  assign n2816 = n2814 | n2815 ;
  assign n2817 = n2813 | n2816 ;
  assign n2818 = ~x134 & n2817 ;
  assign n2819 = n2810 | n2818 ;
  assign n2820 = n485 &  n1570 ;
  assign n2821 = ~n580 & n1606 ;
  assign n2822 = n2820 | n2821 ;
  assign n2823 = ~n436 & n1615 ;
  assign n2824 = ~n535 & n1598 ;
  assign n2825 = n2823 | n2824 ;
  assign n2826 = n2822 | n2825 ;
  assign n2827 = x134 &  n2826 ;
  assign n2828 = ~n436 & n1562 ;
  assign n2829 = ~n580 & n1587 ;
  assign n2830 = n2828 | n2829 ;
  assign n2831 = n485 &  n1623 ;
  assign n2832 = ~n535 & n1579 ;
  assign n2833 = n2831 | n2832 ;
  assign n2834 = n2830 | n2833 ;
  assign n2835 = ~x134 & n2834 ;
  assign n2836 = n2827 | n2835 ;
  assign n2837 = n485 &  n1643 ;
  assign n2838 = ~n580 & n1679 ;
  assign n2839 = n2837 | n2838 ;
  assign n2840 = ~n436 & n1688 ;
  assign n2841 = ~n535 & n1671 ;
  assign n2842 = n2840 | n2841 ;
  assign n2843 = n2839 | n2842 ;
  assign n2844 = x134 &  n2843 ;
  assign n2845 = ~n436 & n1635 ;
  assign n2846 = ~n580 & n1660 ;
  assign n2847 = n2845 | n2846 ;
  assign n2848 = n485 &  n1696 ;
  assign n2849 = ~n535 & n1652 ;
  assign n2850 = n2848 | n2849 ;
  assign n2851 = n2847 | n2850 ;
  assign n2852 = ~x134 & n2851 ;
  assign n2853 = n2844 | n2852 ;
  assign n2854 = n485 &  n1716 ;
  assign n2855 = ~n580 & n1752 ;
  assign n2856 = n2854 | n2855 ;
  assign n2857 = ~n436 & n1761 ;
  assign n2858 = ~n535 & n1744 ;
  assign n2859 = n2857 | n2858 ;
  assign n2860 = n2856 | n2859 ;
  assign n2861 = x134 &  n2860 ;
  assign n2862 = ~n436 & n1708 ;
  assign n2863 = n485 &  n1769 ;
  assign n2864 = n2862 | n2863 ;
  assign n2865 = ~n535 & n1725 ;
  assign n2866 = ~n580 & n1733 ;
  assign n2867 = n2865 | n2866 ;
  assign n2868 = n2864 | n2867 ;
  assign n2869 = ~x134 & n2868 ;
  assign n2870 = n2861 | n2869 ;
  assign n2871 = n485 &  n1789 ;
  assign n2872 = ~n580 & n1825 ;
  assign n2873 = n2871 | n2872 ;
  assign n2874 = ~n436 & n1834 ;
  assign n2875 = ~n535 & n1817 ;
  assign n2876 = n2874 | n2875 ;
  assign n2877 = n2873 | n2876 ;
  assign n2878 = x134 &  n2877 ;
  assign n2879 = ~n436 & n1781 ;
  assign n2880 = n485 &  n1842 ;
  assign n2881 = n2879 | n2880 ;
  assign n2882 = ~n535 & n1798 ;
  assign n2883 = ~n580 & n1806 ;
  assign n2884 = n2882 | n2883 ;
  assign n2885 = n2881 | n2884 ;
  assign n2886 = ~x134 & n2885 ;
  assign n2887 = n2878 | n2886 ;
  assign n2888 = n485 &  n1862 ;
  assign n2889 = ~n580 & n1898 ;
  assign n2890 = n2888 | n2889 ;
  assign n2891 = ~n436 & n1907 ;
  assign n2892 = ~n535 & n1890 ;
  assign n2893 = n2891 | n2892 ;
  assign n2894 = n2890 | n2893 ;
  assign n2895 = x134 &  n2894 ;
  assign n2896 = ~n436 & n1854 ;
  assign n2897 = n485 &  n1915 ;
  assign n2898 = n2896 | n2897 ;
  assign n2899 = ~n535 & n1871 ;
  assign n2900 = ~n580 & n1879 ;
  assign n2901 = n2899 | n2900 ;
  assign n2902 = n2898 | n2901 ;
  assign n2903 = ~x134 & n2902 ;
  assign n2904 = n2895 | n2903 ;
  assign n2905 = n485 &  n1935 ;
  assign n2906 = ~n580 & n1971 ;
  assign n2907 = n2905 | n2906 ;
  assign n2908 = ~n436 & n1980 ;
  assign n2909 = ~n535 & n1963 ;
  assign n2910 = n2908 | n2909 ;
  assign n2911 = n2907 | n2910 ;
  assign n2912 = x134 &  n2911 ;
  assign n2913 = ~n436 & n1927 ;
  assign n2914 = n485 &  n1988 ;
  assign n2915 = n2913 | n2914 ;
  assign n2916 = ~n535 & n1944 ;
  assign n2917 = ~n580 & n1952 ;
  assign n2918 = n2916 | n2917 ;
  assign n2919 = n2915 | n2918 ;
  assign n2920 = ~x134 & n2919 ;
  assign n2921 = n2912 | n2920 ;
  assign n2922 = n485 &  n2008 ;
  assign n2923 = ~n580 & n2044 ;
  assign n2924 = n2922 | n2923 ;
  assign n2925 = ~n436 & n2053 ;
  assign n2926 = ~n535 & n2036 ;
  assign n2927 = n2925 | n2926 ;
  assign n2928 = n2924 | n2927 ;
  assign n2929 = x134 &  n2928 ;
  assign n2930 = ~n436 & n2000 ;
  assign n2931 = n485 &  n2061 ;
  assign n2932 = n2930 | n2931 ;
  assign n2933 = ~n535 & n2017 ;
  assign n2934 = ~n580 & n2025 ;
  assign n2935 = n2933 | n2934 ;
  assign n2936 = n2932 | n2935 ;
  assign n2937 = ~x134 & n2936 ;
  assign n2938 = n2929 | n2937 ;
  assign n2939 = n485 &  n2081 ;
  assign n2940 = ~n580 & n2117 ;
  assign n2941 = n2939 | n2940 ;
  assign n2942 = ~n436 & n2126 ;
  assign n2943 = ~n535 & n2109 ;
  assign n2944 = n2942 | n2943 ;
  assign n2945 = n2941 | n2944 ;
  assign n2946 = x134 &  n2945 ;
  assign n2947 = ~n436 & n2073 ;
  assign n2948 = n485 &  n2134 ;
  assign n2949 = n2947 | n2948 ;
  assign n2950 = ~n535 & n2090 ;
  assign n2951 = ~n580 & n2098 ;
  assign n2952 = n2950 | n2951 ;
  assign n2953 = n2949 | n2952 ;
  assign n2954 = ~x134 & n2953 ;
  assign n2955 = n2946 | n2954 ;
  assign n2956 = ~x134 & n285 ;
  assign n2957 = x134 &  n433 ;
  assign n2958 = n2956 | n2957 ;
  assign n2959 = ~x134 & n630 ;
  assign n2960 = x134 &  n826 ;
  assign n2961 = n2959 | n2960 ;
  assign n2962 = ~x134 & n911 ;
  assign n2963 = x134 &  n995 ;
  assign n2964 = n2962 | n2963 ;
  assign n2965 = ~x134 & n1125 ;
  assign n2966 = x134 &  n1257 ;
  assign n2967 = n2965 | n2966 ;
  assign n2968 = ~x134 & n1298 ;
  assign n2969 = x134 &  n1334 ;
  assign n2970 = n2968 | n2969 ;
  assign n2971 = ~x134 & n1371 ;
  assign n2972 = x134 &  n1407 ;
  assign n2973 = n2971 | n2972 ;
  assign n2974 = ~x134 & n1444 ;
  assign n2975 = x134 &  n1480 ;
  assign n2976 = n2974 | n2975 ;
  assign n2977 = ~x134 & n1517 ;
  assign n2978 = x134 &  n1553 ;
  assign n2979 = n2977 | n2978 ;
  assign n2980 = ~x134 & n1590 ;
  assign n2981 = x134 &  n1626 ;
  assign n2982 = n2980 | n2981 ;
  assign n2983 = ~x134 & n1663 ;
  assign n2984 = x134 &  n1699 ;
  assign n2985 = n2983 | n2984 ;
  assign n2986 = ~x134 & n1736 ;
  assign n2987 = x134 &  n1772 ;
  assign n2988 = n2986 | n2987 ;
  assign n2989 = ~x134 & n1809 ;
  assign n2990 = x134 &  n1845 ;
  assign n2991 = n2989 | n2990 ;
  assign n2992 = ~x134 & n1882 ;
  assign n2993 = x134 &  n1918 ;
  assign n2994 = n2992 | n2993 ;
  assign n2995 = ~x134 & n1955 ;
  assign n2996 = x134 &  n1991 ;
  assign n2997 = n2995 | n2996 ;
  assign n2998 = ~x134 & n2028 ;
  assign n2999 = x134 &  n2064 ;
  assign n3000 = n2998 | n2999 ;
  assign n3001 = ~x134 & n2101 ;
  assign n3002 = x134 &  n2137 ;
  assign n3003 = n3001 | n3002 ;
  assign n3004 = ~x134 & n2146 ;
  assign n3005 = x134 &  n2154 ;
  assign n3006 = n3004 | n3005 ;
  assign n3007 = ~x134 & n2163 ;
  assign n3008 = x134 &  n2171 ;
  assign n3009 = n3007 | n3008 ;
  assign n3010 = ~x134 & n2180 ;
  assign n3011 = x134 &  n2188 ;
  assign n3012 = n3010 | n3011 ;
  assign n3013 = ~x134 & n2197 ;
  assign n3014 = x134 &  n2205 ;
  assign n3015 = n3013 | n3014 ;
  assign n3016 = ~x134 & n2214 ;
  assign n3017 = x134 &  n2222 ;
  assign n3018 = n3016 | n3017 ;
  assign n3019 = ~x134 & n2231 ;
  assign n3020 = x134 &  n2239 ;
  assign n3021 = n3019 | n3020 ;
  assign n3022 = ~x134 & n2248 ;
  assign n3023 = x134 &  n2256 ;
  assign n3024 = n3022 | n3023 ;
  assign n3025 = ~x134 & n2265 ;
  assign n3026 = x134 &  n2273 ;
  assign n3027 = n3025 | n3026 ;
  assign n3028 = ~x134 & n2282 ;
  assign n3029 = x134 &  n2290 ;
  assign n3030 = n3028 | n3029 ;
  assign n3031 = ~x134 & n2299 ;
  assign n3032 = x134 &  n2307 ;
  assign n3033 = n3031 | n3032 ;
  assign n3034 = ~x134 & n2316 ;
  assign n3035 = x134 &  n2324 ;
  assign n3036 = n3034 | n3035 ;
  assign n3037 = ~x134 & n2333 ;
  assign n3038 = x134 &  n2341 ;
  assign n3039 = n3037 | n3038 ;
  assign n3040 = ~x134 & n2350 ;
  assign n3041 = x134 &  n2358 ;
  assign n3042 = n3040 | n3041 ;
  assign n3043 = ~x134 & n2367 ;
  assign n3044 = x134 &  n2375 ;
  assign n3045 = n3043 | n3044 ;
  assign n3046 = ~x134 & n2384 ;
  assign n3047 = x134 &  n2392 ;
  assign n3048 = n3046 | n3047 ;
  assign n3049 = ~x134 & n2401 ;
  assign n3050 = x134 &  n2409 ;
  assign n3051 = n3049 | n3050 ;
  assign n3052 = ~x134 & n2418 ;
  assign n3053 = x134 &  n2426 ;
  assign n3054 = n3052 | n3053 ;
  assign n3055 = ~x134 & n2435 ;
  assign n3056 = x134 &  n2443 ;
  assign n3057 = n3055 | n3056 ;
  assign n3058 = ~x134 & n2452 ;
  assign n3059 = x134 &  n2460 ;
  assign n3060 = n3058 | n3059 ;
  assign n3061 = ~x134 & n2469 ;
  assign n3062 = x134 &  n2477 ;
  assign n3063 = n3061 | n3062 ;
  assign n3064 = ~x134 & n2486 ;
  assign n3065 = x134 &  n2494 ;
  assign n3066 = n3064 | n3065 ;
  assign n3067 = ~x134 & n2503 ;
  assign n3068 = x134 &  n2511 ;
  assign n3069 = n3067 | n3068 ;
  assign n3070 = ~x134 & n2520 ;
  assign n3071 = x134 &  n2528 ;
  assign n3072 = n3070 | n3071 ;
  assign n3073 = ~x134 & n2537 ;
  assign n3074 = x134 &  n2545 ;
  assign n3075 = n3073 | n3074 ;
  assign n3076 = ~x134 & n2554 ;
  assign n3077 = x134 &  n2562 ;
  assign n3078 = n3076 | n3077 ;
  assign n3079 = ~x134 & n2571 ;
  assign n3080 = x134 &  n2579 ;
  assign n3081 = n3079 | n3080 ;
  assign n3082 = ~x134 & n2588 ;
  assign n3083 = x134 &  n2596 ;
  assign n3084 = n3082 | n3083 ;
  assign n3085 = ~x134 & n2605 ;
  assign n3086 = x134 &  n2613 ;
  assign n3087 = n3085 | n3086 ;
  assign n3088 = ~x134 & n2622 ;
  assign n3089 = x134 &  n2630 ;
  assign n3090 = n3088 | n3089 ;
  assign n3091 = ~x134 & n2639 ;
  assign n3092 = x134 &  n2647 ;
  assign n3093 = n3091 | n3092 ;
  assign n3094 = ~x134 & n2656 ;
  assign n3095 = x134 &  n2664 ;
  assign n3096 = n3094 | n3095 ;
  assign n3097 = ~x134 & n2673 ;
  assign n3098 = x134 &  n2681 ;
  assign n3099 = n3097 | n3098 ;
  assign n3100 = ~x134 & n2690 ;
  assign n3101 = x134 &  n2698 ;
  assign n3102 = n3100 | n3101 ;
  assign n3103 = ~x134 & n2707 ;
  assign n3104 = x134 &  n2715 ;
  assign n3105 = n3103 | n3104 ;
  assign n3106 = ~x134 & n2724 ;
  assign n3107 = x134 &  n2732 ;
  assign n3108 = n3106 | n3107 ;
  assign n3109 = ~x134 & n2741 ;
  assign n3110 = x134 &  n2749 ;
  assign n3111 = n3109 | n3110 ;
  assign n3112 = ~x134 & n2758 ;
  assign n3113 = x134 &  n2766 ;
  assign n3114 = n3112 | n3113 ;
  assign n3115 = ~x134 & n2775 ;
  assign n3116 = x134 &  n2783 ;
  assign n3117 = n3115 | n3116 ;
  assign n3118 = ~x134 & n2792 ;
  assign n3119 = x134 &  n2800 ;
  assign n3120 = n3118 | n3119 ;
  assign n3121 = ~x134 & n2809 ;
  assign n3122 = x134 &  n2817 ;
  assign n3123 = n3121 | n3122 ;
  assign n3124 = ~x134 & n2826 ;
  assign n3125 = x134 &  n2834 ;
  assign n3126 = n3124 | n3125 ;
  assign n3127 = ~x134 & n2843 ;
  assign n3128 = x134 &  n2851 ;
  assign n3129 = n3127 | n3128 ;
  assign n3130 = ~x134 & n2860 ;
  assign n3131 = x134 &  n2868 ;
  assign n3132 = n3130 | n3131 ;
  assign n3133 = ~x134 & n2877 ;
  assign n3134 = x134 &  n2885 ;
  assign n3135 = n3133 | n3134 ;
  assign n3136 = ~x134 & n2894 ;
  assign n3137 = x134 &  n2902 ;
  assign n3138 = n3136 | n3137 ;
  assign n3139 = ~x134 & n2911 ;
  assign n3140 = x134 &  n2919 ;
  assign n3141 = n3139 | n3140 ;
  assign n3142 = ~x134 & n2928 ;
  assign n3143 = x134 &  n2936 ;
  assign n3144 = n3142 | n3143 ;
  assign n3145 = ~x134 & n2945 ;
  assign n3146 = x134 &  n2953 ;
  assign n3147 = n3145 | n3146 ;
  assign y0 = n435 ;
  assign y1 = n828 ;
  assign y2 = n997 ;
  assign y3 = n1259 ;
  assign y4 = n1336 ;
  assign y5 = n1409 ;
  assign y6 = n1482 ;
  assign y7 = n1555 ;
  assign y8 = n1628 ;
  assign y9 = n1701 ;
  assign y10 = n1774 ;
  assign y11 = n1847 ;
  assign y12 = n1920 ;
  assign y13 = n1993 ;
  assign y14 = n2066 ;
  assign y15 = n2139 ;
  assign y16 = n2156 ;
  assign y17 = n2173 ;
  assign y18 = n2190 ;
  assign y19 = n2207 ;
  assign y20 = n2224 ;
  assign y21 = n2241 ;
  assign y22 = n2258 ;
  assign y23 = n2275 ;
  assign y24 = n2292 ;
  assign y25 = n2309 ;
  assign y26 = n2326 ;
  assign y27 = n2343 ;
  assign y28 = n2360 ;
  assign y29 = n2377 ;
  assign y30 = n2394 ;
  assign y31 = n2411 ;
  assign y32 = n2428 ;
  assign y33 = n2445 ;
  assign y34 = n2462 ;
  assign y35 = n2479 ;
  assign y36 = n2496 ;
  assign y37 = n2513 ;
  assign y38 = n2530 ;
  assign y39 = n2547 ;
  assign y40 = n2564 ;
  assign y41 = n2581 ;
  assign y42 = n2598 ;
  assign y43 = n2615 ;
  assign y44 = n2632 ;
  assign y45 = n2649 ;
  assign y46 = n2666 ;
  assign y47 = n2683 ;
  assign y48 = n2700 ;
  assign y49 = n2717 ;
  assign y50 = n2734 ;
  assign y51 = n2751 ;
  assign y52 = n2768 ;
  assign y53 = n2785 ;
  assign y54 = n2802 ;
  assign y55 = n2819 ;
  assign y56 = n2836 ;
  assign y57 = n2853 ;
  assign y58 = n2870 ;
  assign y59 = n2887 ;
  assign y60 = n2904 ;
  assign y61 = n2921 ;
  assign y62 = n2938 ;
  assign y63 = n2955 ;
  assign y64 = n2958 ;
  assign y65 = n2961 ;
  assign y66 = n2964 ;
  assign y67 = n2967 ;
  assign y68 = n2970 ;
  assign y69 = n2973 ;
  assign y70 = n2976 ;
  assign y71 = n2979 ;
  assign y72 = n2982 ;
  assign y73 = n2985 ;
  assign y74 = n2988 ;
  assign y75 = n2991 ;
  assign y76 = n2994 ;
  assign y77 = n2997 ;
  assign y78 = n3000 ;
  assign y79 = n3003 ;
  assign y80 = n3006 ;
  assign y81 = n3009 ;
  assign y82 = n3012 ;
  assign y83 = n3015 ;
  assign y84 = n3018 ;
  assign y85 = n3021 ;
  assign y86 = n3024 ;
  assign y87 = n3027 ;
  assign y88 = n3030 ;
  assign y89 = n3033 ;
  assign y90 = n3036 ;
  assign y91 = n3039 ;
  assign y92 = n3042 ;
  assign y93 = n3045 ;
  assign y94 = n3048 ;
  assign y95 = n3051 ;
  assign y96 = n3054 ;
  assign y97 = n3057 ;
  assign y98 = n3060 ;
  assign y99 = n3063 ;
  assign y100 = n3066 ;
  assign y101 = n3069 ;
  assign y102 = n3072 ;
  assign y103 = n3075 ;
  assign y104 = n3078 ;
  assign y105 = n3081 ;
  assign y106 = n3084 ;
  assign y107 = n3087 ;
  assign y108 = n3090 ;
  assign y109 = n3093 ;
  assign y110 = n3096 ;
  assign y111 = n3099 ;
  assign y112 = n3102 ;
  assign y113 = n3105 ;
  assign y114 = n3108 ;
  assign y115 = n3111 ;
  assign y116 = n3114 ;
  assign y117 = n3117 ;
  assign y118 = n3120 ;
  assign y119 = n3123 ;
  assign y120 = n3126 ;
  assign y121 = n3129 ;
  assign y122 = n3132 ;
  assign y123 = n3135 ;
  assign y124 = n3138 ;
  assign y125 = n3141 ;
  assign y126 = n3144 ;
  assign y127 = n3147 ;
endmodule
