module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 ;
  assign n25 = x1 | x2 ;
  assign n26 = x0 | n25 ;
  assign n27 = x3 | n26 ;
  assign n28 = x4 | n27 ;
  assign n29 = x5 | n28 ;
  assign n30 = x6 | n29 ;
  assign n31 = x7 | n30 ;
  assign n245 = ~x22 & n31 ;
  assign n246 = ~x8 & n245 ;
  assign n247 = ( x8 & ~n245 ) | ( x8 & 1'b0 ) | ( ~n245 & 1'b0 ) ;
  assign n248 = n246 | n247 ;
  assign n32 = x8 | n31 ;
  assign n244 = ~x22 & n32 ;
  assign n250 = ( x9 & n244 ) | ( x9 & n248 ) | ( n244 & n248 ) ;
  assign n249 = ( x9 & ~n248 ) | ( x9 & n244 ) | ( ~n248 & n244 ) ;
  assign n251 = ( n248 & ~n250 ) | ( n248 & n249 ) | ( ~n250 & n249 ) ;
  assign n33 = x9 | n32 ;
  assign n253 = ~x22 & n33 ;
  assign n254 = ~x10 & n253 ;
  assign n255 = ( x10 & ~n253 ) | ( x10 & 1'b0 ) | ( ~n253 & 1'b0 ) ;
  assign n256 = n254 | n255 ;
  assign n34 = x10 | n33 ;
  assign n252 = ~x22 & n34 ;
  assign n258 = ( x11 & n252 ) | ( x11 & n256 ) | ( n252 & n256 ) ;
  assign n257 = ( x11 & ~n256 ) | ( x11 & n252 ) | ( ~n256 & n252 ) ;
  assign n259 = ( n256 & ~n258 ) | ( n256 & n257 ) | ( ~n258 & n257 ) ;
  assign n260 = ~n251 |  n259 ;
  assign n35 = x11 | n34 ;
  assign n36 = x12 | n35 ;
  assign n37 = x13 | n36 ;
  assign n38 = x14 | n37 ;
  assign n49 = ~x22 & n38 ;
  assign n50 = ~x15 & n49 ;
  assign n51 = ( x15 & ~n49 ) | ( x15 & 1'b0 ) | ( ~n49 & 1'b0 ) ;
  assign n52 = n50 | n51 ;
  assign n39 = x15 | n38 ;
  assign n40 = x16 | n39 ;
  assign n41 = x17 | n40 ;
  assign n42 = ( x19 & ~x18 ) | ( x19 & n41 ) | ( ~x18 & n41 ) ;
  assign n43 = x18 | n42 ;
  assign n44 = ~x22 & n43 ;
  assign n45 = x21 | n44 ;
  assign n47 = x20 &  n44 ;
  assign n46 = ( x20 & ~x21 ) | ( x20 & 1'b0 ) | ( ~x21 & 1'b0 ) ;
  assign n48 = ( n45 & ~n47 ) | ( n45 & n46 ) | ( ~n47 & n46 ) ;
  assign n106 = ~n52 |  n48 ;
  assign n80 = ( x18 & ~x19 ) | ( x18 & 1'b0 ) | ( ~x19 & 1'b0 ) ;
  assign n79 = ~x22 & n41 ;
  assign n82 = x18 | n79 ;
  assign n81 = x19 | n79 ;
  assign n83 = ( n80 & ~n82 ) | ( n80 & n81 ) | ( ~n82 & n81 ) ;
  assign n59 = ~x22 & n40 ;
  assign n60 = ~x17 & n59 ;
  assign n61 = ( x17 & ~n59 ) | ( x17 & 1'b0 ) | ( ~n59 & 1'b0 ) ;
  assign n62 = n60 | n61 ;
  assign n63 = ~x22 & n39 ;
  assign n64 = ~x16 & n63 ;
  assign n65 = ( x16 & ~n63 ) | ( x16 & 1'b0 ) | ( ~n63 & 1'b0 ) ;
  assign n66 = n64 | n65 ;
  assign n111 = n62 &  n66 ;
  assign n125 = n83 &  n111 ;
  assign n436 = ~n106 & n125 ;
  assign n54 = x22 | n41 ;
  assign n55 = ( x22 & ~x18 ) | ( x22 & n54 ) | ( ~x18 & n54 ) ;
  assign n56 = x19 | x22 ;
  assign n57 = ( x18 & ~n54 ) | ( x18 & x19 ) | ( ~n54 & x19 ) ;
  assign n58 = ( n55 & ~n56 ) | ( n55 & n57 ) | ( ~n56 & n57 ) ;
  assign n70 = n62 | n66 ;
  assign n71 = ( n58 & ~n70 ) | ( n58 & 1'b0 ) | ( ~n70 & 1'b0 ) ;
  assign n487 = ( n71 & ~n106 ) | ( n71 & 1'b0 ) | ( ~n106 & 1'b0 ) ;
  assign n53 = n48 | n52 ;
  assign n67 = ( n62 & ~n66 ) | ( n62 & 1'b0 ) | ( ~n66 & 1'b0 ) ;
  assign n88 = ( x19 & ~x18 ) | ( x19 & n54 ) | ( ~x18 & n54 ) ;
  assign n87 = ( x19 & ~x22 ) | ( x19 & 1'b0 ) | ( ~x22 & 1'b0 ) ;
  assign n89 = ( n55 & ~n88 ) | ( n55 & n87 ) | ( ~n88 & n87 ) ;
  assign n107 = n67 &  n89 ;
  assign n555 = ~n53 & n107 ;
  assign n72 = x22 | n43 ;
  assign n73 = ( x22 & ~x20 ) | ( x22 & n72 ) | ( ~x20 & n72 ) ;
  assign n75 = ( x21 & ~x20 ) | ( x21 & n72 ) | ( ~x20 & n72 ) ;
  assign n74 = ( x21 & ~x22 ) | ( x21 & 1'b0 ) | ( ~x22 & 1'b0 ) ;
  assign n76 = ( n73 & ~n75 ) | ( n73 & n74 ) | ( ~n75 & n74 ) ;
  assign n86 = n52 &  n76 ;
  assign n144 = x18 &  n79 ;
  assign n145 = ( n80 & ~n144 ) | ( n80 & n81 ) | ( ~n144 & n81 ) ;
  assign n161 = ( n111 & ~n145 ) | ( n111 & 1'b0 ) | ( ~n145 & 1'b0 ) ;
  assign n208 = n86 &  n161 ;
  assign n95 = ~n62 & n66 ;
  assign n166 = ( n95 & ~n145 ) | ( n95 & 1'b0 ) | ( ~n145 & 1'b0 ) ;
  assign n230 = ~n53 & n166 ;
  assign n68 = n58 &  n67 ;
  assign n92 = x20 | n44 ;
  assign n93 = ( n45 & ~n92 ) | ( n45 & n46 ) | ( ~n92 & n46 ) ;
  assign n148 = ~n93 |  n52 ;
  assign n311 = ( n68 & ~n148 ) | ( n68 & 1'b0 ) | ( ~n148 & 1'b0 ) ;
  assign n84 = ~n70 & n83 ;
  assign n94 = n52 &  n93 ;
  assign n827 = n84 &  n94 ;
  assign n98 = x21 | x22 ;
  assign n99 = ( x20 & ~n72 ) | ( x20 & x21 ) | ( ~n72 & x21 ) ;
  assign n100 = ( n73 & ~n98 ) | ( n73 & n99 ) | ( ~n98 & n99 ) ;
  assign n101 = ~n52 | ~n100 ;
  assign n380 = ~n101 & n161 ;
  assign n201 = ( n84 & ~n101 ) | ( n84 & 1'b0 ) | ( ~n101 & 1'b0 ) ;
  assign n120 = n68 &  n86 ;
  assign n77 = ~n52 & n76 ;
  assign n121 = n89 &  n95 ;
  assign n122 = n77 &  n121 ;
  assign n123 = n120 | n122 ;
  assign n117 = n58 &  n95 ;
  assign n330 = n86 &  n117 ;
  assign n104 = ~n52 & n100 ;
  assign n331 = ( n58 & ~n66 ) | ( n58 & 1'b0 ) | ( ~n66 & 1'b0 ) ;
  assign n168 = n58 &  n111 ;
  assign n332 = ~n331 & n168 ;
  assign n333 = ( n104 & n332 ) | ( n104 & n331 ) | ( n332 & n331 ) ;
  assign n334 = n330 | n333 ;
  assign n179 = ( n67 & ~n145 ) | ( n67 & 1'b0 ) | ( ~n145 & 1'b0 ) ;
  assign n212 = ~n106 & n179 ;
  assign n69 = ~n53 & n68 ;
  assign n180 = n86 &  n179 ;
  assign n353 = n71 &  n86 ;
  assign n112 = n89 &  n111 ;
  assign n354 = n86 &  n112 ;
  assign n96 = n83 &  n95 ;
  assign n113 = n96 &  n104 ;
  assign n355 = ~n106 & n166 ;
  assign n102 = n67 &  n83 ;
  assign n190 = n77 &  n102 ;
  assign n97 = n94 &  n96 ;
  assign n141 = n94 &  n125 ;
  assign n356 = n97 | n141 ;
  assign n357 = n190 | n356 ;
  assign n358 = n355 | n357 ;
  assign n146 = n70 | n145 ;
  assign n147 = ( n86 & ~n146 ) | ( n86 & 1'b0 ) | ( ~n146 & 1'b0 ) ;
  assign n90 = ~n70 & n89 ;
  assign n165 = n90 &  n94 ;
  assign n191 = n94 &  n121 ;
  assign n359 = n165 | n191 ;
  assign n360 = n147 | n359 ;
  assign n209 = ( n68 & ~n106 ) | ( n68 & 1'b0 ) | ( ~n106 & 1'b0 ) ;
  assign n361 = ~n53 & n84 ;
  assign n362 = n77 &  n96 ;
  assign n363 = n77 &  n107 ;
  assign n310 = n84 &  n104 ;
  assign n364 = n86 &  n166 ;
  assign n365 = n310 | n364 ;
  assign n366 = ( n363 & ~n362 ) | ( n363 & n365 ) | ( ~n362 & n365 ) ;
  assign n367 = n362 | n366 ;
  assign n368 = ( n361 & ~n209 ) | ( n361 & n367 ) | ( ~n209 & n367 ) ;
  assign n369 = n209 | n368 ;
  assign n370 = ( n360 & ~n358 ) | ( n360 & n369 ) | ( ~n358 & n369 ) ;
  assign n371 = ( n358 & ~n113 ) | ( n358 & n370 ) | ( ~n113 & n370 ) ;
  assign n372 = n113 | n371 ;
  assign n373 = ( n354 & ~n353 ) | ( n354 & n372 ) | ( ~n353 & n372 ) ;
  assign n374 = n353 | n373 ;
  assign n375 = ( n180 & ~n69 ) | ( n180 & n374 ) | ( ~n69 & n374 ) ;
  assign n376 = n69 | n375 ;
  assign n377 = n212 | n376 ;
  assign n197 = ( n96 & ~n106 ) | ( n96 & 1'b0 ) | ( ~n106 & 1'b0 ) ;
  assign n612 = ~n53 & n121 ;
  assign n85 = n77 &  n84 ;
  assign n293 = n94 &  n161 ;
  assign n467 = ( n96 & ~n148 ) | ( n96 & 1'b0 ) | ( ~n148 & 1'b0 ) ;
  assign n392 = n104 &  n112 ;
  assign n352 = n90 &  n104 ;
  assign n503 = ~n101 & n107 ;
  assign n756 = ( n352 & ~n392 ) | ( n352 & n503 ) | ( ~n392 & n503 ) ;
  assign n757 = n392 | n756 ;
  assign n758 = n467 | n757 ;
  assign n140 = n77 &  n117 ;
  assign n277 = ( n94 & ~n146 ) | ( n94 & 1'b0 ) | ( ~n146 & 1'b0 ) ;
  assign n438 = n140 | n277 ;
  assign n103 = ~n101 & n102 ;
  assign n200 = ~n101 & n125 ;
  assign n324 = ~n101 & n168 ;
  assign n562 = n200 | n324 ;
  assign n563 = n103 | n562 ;
  assign n316 = ~n53 & n96 ;
  assign n302 = n86 &  n107 ;
  assign n412 = n94 &  n112 ;
  assign n1761 = n302 | n412 ;
  assign n1762 = n316 | n1761 ;
  assign n1763 = n563 | n1762 ;
  assign n1764 = ( n438 & ~n758 ) | ( n438 & n1763 ) | ( ~n758 & n1763 ) ;
  assign n1765 = n758 | n1764 ;
  assign n1766 = ( n293 & ~n85 ) | ( n293 & n1765 ) | ( ~n85 & n1765 ) ;
  assign n1767 = n85 | n1766 ;
  assign n1768 = ( n612 & ~n197 ) | ( n612 & n1767 ) | ( ~n197 & n1767 ) ;
  assign n1769 = n197 | n1768 ;
  assign n160 = n71 &  n94 ;
  assign n468 = ~n53 & n161 ;
  assign n584 = n160 | n468 ;
  assign n198 = n86 &  n102 ;
  assign n261 = ~n53 & n168 ;
  assign n91 = n86 &  n90 ;
  assign n398 = n84 &  n86 ;
  assign n152 = ( n90 & ~n148 ) | ( n90 & 1'b0 ) | ( ~n148 & 1'b0 ) ;
  assign n690 = ( n121 & ~n148 ) | ( n121 & 1'b0 ) | ( ~n148 & 1'b0 ) ;
  assign n691 = n152 | n690 ;
  assign n227 = n94 &  n168 ;
  assign n381 = ( n104 & ~n146 ) | ( n104 & 1'b0 ) | ( ~n146 & 1'b0 ) ;
  assign n755 = n227 | n381 ;
  assign n1770 = n691 | n755 ;
  assign n1771 = ( n398 & ~n91 ) | ( n398 & n1770 ) | ( ~n91 & n1770 ) ;
  assign n1772 = n91 | n1771 ;
  assign n1773 = ( n261 & ~n198 ) | ( n261 & n1772 ) | ( ~n198 & n1772 ) ;
  assign n1774 = n198 | n1773 ;
  assign n1775 = ( n584 & ~n1769 ) | ( n584 & n1774 ) | ( ~n1769 & n1774 ) ;
  assign n1776 = ( n1769 & ~n377 ) | ( n1769 & n1775 ) | ( ~n377 & n1775 ) ;
  assign n1777 = n377 | n1776 ;
  assign n1778 = ( n334 & ~n123 ) | ( n334 & n1777 ) | ( ~n123 & n1777 ) ;
  assign n1779 = n123 | n1778 ;
  assign n1780 = ( n201 & ~n380 ) | ( n201 & n1779 ) | ( ~n380 & n1779 ) ;
  assign n1781 = n380 | n1780 ;
  assign n1782 = ( n827 & ~n311 ) | ( n827 & n1781 ) | ( ~n311 & n1781 ) ;
  assign n1783 = n311 | n1782 ;
  assign n1784 = ( n230 & ~n208 ) | ( n230 & n1783 ) | ( ~n208 & n1783 ) ;
  assign n1785 = n208 | n1784 ;
  assign n1786 = ( n555 & ~n487 ) | ( n555 & n1785 ) | ( ~n487 & n1785 ) ;
  assign n1787 = n487 | n1786 ;
  assign n1788 = n436 | n1787 ;
  assign n229 = ( n84 & ~n148 ) | ( n84 & 1'b0 ) | ( ~n148 & 1'b0 ) ;
  assign n418 = n101 | n146 ;
  assign n315 = n104 &  n179 ;
  assign n108 = ~n106 & n107 ;
  assign n109 = n68 &  n94 ;
  assign n110 = ( n96 & ~n101 ) | ( n96 & 1'b0 ) | ( ~n101 & 1'b0 ) ;
  assign n135 = ~n112 & n100 ;
  assign n114 = n104 &  n107 ;
  assign n115 = n113 | n114 ;
  assign n116 = n68 &  n77 ;
  assign n118 = n104 &  n117 ;
  assign n119 = n116 | n118 ;
  assign n124 = n102 &  n104 ;
  assign n126 = n104 &  n125 ;
  assign n127 = n124 | n126 ;
  assign n128 = ~n106 & n112 ;
  assign n129 = ( n68 & ~n101 ) | ( n68 & 1'b0 ) | ( ~n101 & 1'b0 ) ;
  assign n130 = n128 | n129 ;
  assign n131 = ( n127 & ~n123 ) | ( n127 & n130 ) | ( ~n123 & n130 ) ;
  assign n132 = n123 | n131 ;
  assign n133 = ( n119 & ~n115 ) | ( n119 & n132 ) | ( ~n115 & n132 ) ;
  assign n134 = n115 | n133 ;
  assign n136 = ( n100 & ~n135 ) | ( n100 & n134 ) | ( ~n135 & n134 ) ;
  assign n137 = ( n110 & ~n109 ) | ( n110 & n136 ) | ( ~n109 & n136 ) ;
  assign n138 = n109 | n137 ;
  assign n139 = n108 | n138 ;
  assign n323 = ( n117 & ~n148 ) | ( n117 & 1'b0 ) | ( ~n148 & 1'b0 ) ;
  assign n325 = ~n90 & n166 ;
  assign n326 = ( n90 & n104 ) | ( n90 & n325 ) | ( n104 & n325 ) ;
  assign n327 = ( n324 & ~n201 ) | ( n324 & n326 ) | ( ~n201 & n326 ) ;
  assign n328 = n201 | n327 ;
  assign n329 = n323 | n328 ;
  assign n186 = n86 &  n168 ;
  assign n443 = ~n148 & n168 ;
  assign n195 = ~n101 & n121 ;
  assign n444 = n195 | n412 ;
  assign n275 = n77 &  n161 ;
  assign n445 = n85 | n275 ;
  assign n181 = n94 &  n107 ;
  assign n105 = n68 &  n104 ;
  assign n446 = ~n101 & n179 ;
  assign n447 = n105 | n446 ;
  assign n448 = n181 | n447 ;
  assign n449 = ( n445 & ~n444 ) | ( n445 & n448 ) | ( ~n444 & n448 ) ;
  assign n450 = n444 | n449 ;
  assign n451 = ( n443 & ~n186 ) | ( n443 & n450 ) | ( ~n186 & n450 ) ;
  assign n452 = n186 | n451 ;
  assign n1815 = n354 | n361 ;
  assign n149 = ( n125 & ~n148 ) | ( n125 & 1'b0 ) | ( ~n148 & 1'b0 ) ;
  assign n746 = n149 | n310 ;
  assign n199 = n94 &  n117 ;
  assign n826 = n199 | n467 ;
  assign n1816 = n746 | n826 ;
  assign n1817 = ( n1815 & ~n1774 ) | ( n1815 & n1816 ) | ( ~n1774 & n1816 ) ;
  assign n1818 = n1774 | n1817 ;
  assign n495 = n53 | n146 ;
  assign n496 = ~n97 & n495 ;
  assign n1819 = ( n452 & ~n1818 ) | ( n452 & n496 ) | ( ~n1818 & n496 ) ;
  assign n1820 = ~n452 & n1819 ;
  assign n723 = n77 &  n179 ;
  assign n402 = ~n53 & n117 ;
  assign n290 = n77 &  n90 ;
  assign n317 = n77 &  n168 ;
  assign n318 = ~n148 & n179 ;
  assign n319 = ( n84 & ~n106 ) | ( n84 & 1'b0 ) | ( ~n106 & 1'b0 ) ;
  assign n320 = n318 | n319 ;
  assign n321 = n317 | n320 ;
  assign n322 = n316 | n321 ;
  assign n189 = ( n90 & ~n106 ) | ( n90 & 1'b0 ) | ( ~n106 & 1'b0 ) ;
  assign n600 = n69 | n189 ;
  assign n281 = ( n102 & ~n106 ) | ( n102 & 1'b0 ) | ( ~n106 & 1'b0 ) ;
  assign n282 = ~n106 & n168 ;
  assign n283 = n281 | n282 ;
  assign n643 = ~n106 & n117 ;
  assign n78 = n71 &  n77 ;
  assign n501 = n77 &  n166 ;
  assign n554 = ~n53 & n179 ;
  assign n597 = ~n53 & n90 ;
  assign n1798 = n554 | n597 ;
  assign n1799 = ( n501 & ~n78 ) | ( n501 & n1798 ) | ( ~n78 & n1798 ) ;
  assign n1800 = n78 | n1799 ;
  assign n1801 = n643 | n1800 ;
  assign n211 = ~n106 & n161 ;
  assign n292 = n86 &  n125 ;
  assign n437 = ~n53 & n112 ;
  assign n1802 = n292 | n437 ;
  assign n1803 = n211 | n1802 ;
  assign n1804 = n330 | n436 ;
  assign n1805 = ( n1803 & ~n1801 ) | ( n1803 & n1804 ) | ( ~n1801 & n1804 ) ;
  assign n1806 = ( n1801 & ~n283 ) | ( n1801 & n1805 ) | ( ~n283 & n1805 ) ;
  assign n1807 = n283 | n1806 ;
  assign n378 = n106 | n146 ;
  assign n645 = n146 | n148 ;
  assign n289 = n77 &  n112 ;
  assign n595 = n86 &  n121 ;
  assign n730 = n289 | n595 ;
  assign n731 = n363 | n730 ;
  assign n1691 = ( n645 & ~n731 ) | ( n645 & 1'b0 ) | ( ~n731 & 1'b0 ) ;
  assign n1692 = ( n355 & ~n1691 ) | ( n355 & n378 ) | ( ~n1691 & n378 ) ;
  assign n1693 = ( n378 & ~n1692 ) | ( n378 & 1'b0 ) | ( ~n1692 & 1'b0 ) ;
  assign n1808 = ( n600 & ~n1807 ) | ( n600 & n1693 ) | ( ~n1807 & n1693 ) ;
  assign n1809 = ~n600 & n1808 ;
  assign n1810 = ( n290 & ~n322 ) | ( n290 & n1809 ) | ( ~n322 & n1809 ) ;
  assign n1811 = ~n290 & n1810 ;
  assign n1812 = ( n723 & ~n402 ) | ( n723 & n1811 ) | ( ~n402 & n1811 ) ;
  assign n1813 = ~n723 & n1812 ;
  assign n1814 = ~n197 & n1813 ;
  assign n1821 = ( n329 & ~n1820 ) | ( n329 & n1814 ) | ( ~n1820 & n1814 ) ;
  assign n1822 = ( n139 & ~n1821 ) | ( n139 & n1814 ) | ( ~n1821 & n1814 ) ;
  assign n1823 = ~n139 & n1822 ;
  assign n1824 = ( n315 & ~n1823 ) | ( n315 & n418 ) | ( ~n1823 & n418 ) ;
  assign n1825 = ( n418 & ~n1824 ) | ( n418 & 1'b0 ) | ( ~n1824 & 1'b0 ) ;
  assign n1826 = ( n229 & ~n293 ) | ( n229 & n1825 ) | ( ~n293 & n1825 ) ;
  assign n1827 = ~n229 & n1826 ;
  assign n1828 = ~n212 & n1827 ;
  assign n162 = n104 &  n161 ;
  assign n276 = ( n112 & ~n148 ) | ( n112 & 1'b0 ) | ( ~n148 & 1'b0 ) ;
  assign n169 = n104 &  n168 ;
  assign n887 = n277 | n311 ;
  assign n888 = n554 | n887 ;
  assign n391 = ( n107 & ~n148 ) | ( n107 & 1'b0 ) | ( ~n148 & 1'b0 ) ;
  assign n889 = n364 | n391 ;
  assign n890 = n501 | n889 ;
  assign n892 = n161 | n148 ;
  assign n309 = ( n71 & ~n101 ) | ( n71 & 1'b0 ) | ( ~n101 & 1'b0 ) ;
  assign n891 = n309 | n362 ;
  assign n893 = ( n892 & ~n148 ) | ( n892 & n891 ) | ( ~n148 & n891 ) ;
  assign n894 = n402 | n893 ;
  assign n895 = ( n890 & ~n888 ) | ( n890 & n894 ) | ( ~n888 & n894 ) ;
  assign n896 = ( n888 & ~n329 ) | ( n888 & n895 ) | ( ~n329 & n895 ) ;
  assign n897 = n329 | n896 ;
  assign n898 = ( n169 & ~n123 ) | ( n169 & n897 ) | ( ~n123 & n897 ) ;
  assign n899 = n123 | n898 ;
  assign n900 = ( n276 & ~n186 ) | ( n276 & n899 ) | ( ~n186 & n899 ) ;
  assign n901 = n186 | n900 ;
  assign n902 = n281 | n901 ;
  assign n903 = ( n71 & ~n84 ) | ( n71 & n86 ) | ( ~n84 & n86 ) ;
  assign n904 = ~n71 & n903 ;
  assign n411 = ~n101 & n112 ;
  assign n185 = ~n106 & n121 ;
  assign n422 = n94 &  n179 ;
  assign n830 = n185 | n422 ;
  assign n153 = n71 &  n104 ;
  assign n154 = n152 | n153 ;
  assign n453 = n78 | n302 ;
  assign n905 = ( n154 & ~n830 ) | ( n154 & n453 ) | ( ~n830 & n453 ) ;
  assign n906 = ( n830 & ~n411 ) | ( n830 & n905 ) | ( ~n411 & n905 ) ;
  assign n907 = n411 | n906 ;
  assign n908 = ( n467 & ~n165 ) | ( n467 & n907 ) | ( ~n165 & n907 ) ;
  assign n909 = n165 | n908 ;
  assign n910 = ( n86 & ~n904 ) | ( n86 & n909 ) | ( ~n904 & n909 ) ;
  assign n911 = n436 | n910 ;
  assign n192 = ( n71 & ~n148 ) | ( n71 & 1'b0 ) | ( ~n148 & 1'b0 ) ;
  assign n478 = ~n101 & n117 ;
  assign n678 = n52 &  n161 ;
  assign n679 = ~n52 & n179 ;
  assign n680 = ( n93 & n678 ) | ( n93 & n679 ) | ( n678 & n679 ) ;
  assign n912 = n319 | n680 ;
  assign n913 = ( n418 & ~n912 ) | ( n418 & n478 ) | ( ~n912 & n478 ) ;
  assign n914 = ~n478 & n913 ;
  assign n915 = ( n192 & ~n354 ) | ( n192 & n914 ) | ( ~n354 & n914 ) ;
  assign n916 = ~n192 & n915 ;
  assign n917 = ( n378 & ~n916 ) | ( n378 & n723 ) | ( ~n916 & n723 ) ;
  assign n918 = ( n378 & ~n917 ) | ( n378 & 1'b0 ) | ( ~n917 & 1'b0 ) ;
  assign n558 = ~n121 & n100 ;
  assign n556 = n212 | n555 ;
  assign n557 = n261 | n556 ;
  assign n559 = ( n100 & ~n558 ) | ( n100 & n557 ) | ( ~n558 & n557 ) ;
  assign n267 = ~n90 & n179 ;
  assign n268 = ( n90 & ~n101 ) | ( n90 & n267 ) | ( ~n101 & n267 ) ;
  assign n923 = n197 | n597 ;
  assign n924 = n114 | n827 ;
  assign n925 = ( n923 & ~n268 ) | ( n923 & n924 ) | ( ~n268 & n924 ) ;
  assign n926 = n268 | n925 ;
  assign n927 = ( n496 & n559 ) | ( n496 & n926 ) | ( n559 & n926 ) ;
  assign n928 = ( n496 & ~n927 ) | ( n496 & 1'b0 ) | ( ~n927 & 1'b0 ) ;
  assign n667 = n76 &  n125 ;
  assign n745 = n93 &  n102 ;
  assign n919 = n91 | n745 ;
  assign n920 = n209 | n919 ;
  assign n921 = ( n667 & ~n198 ) | ( n667 & n920 ) | ( ~n198 & n920 ) ;
  assign n922 = n198 | n921 ;
  assign n929 = ( n918 & ~n928 ) | ( n918 & n922 ) | ( ~n928 & n922 ) ;
  assign n930 = ( n911 & ~n929 ) | ( n911 & n918 ) | ( ~n929 & n918 ) ;
  assign n931 = ~n911 & n930 ;
  assign n932 = ( n162 & ~n902 ) | ( n162 & n931 ) | ( ~n902 & n931 ) ;
  assign n933 = ~n162 & n932 ;
  assign n934 = ( n109 & ~n180 ) | ( n109 & n933 ) | ( ~n180 & n933 ) ;
  assign n935 = ~n109 & n934 ;
  assign n936 = ( n140 & ~n437 ) | ( n140 & n935 ) | ( ~n437 & n935 ) ;
  assign n937 = ~n936 |  n140 ;
  assign n143 = n86 &  n96 ;
  assign n829 = n97 | n309 ;
  assign n647 = n94 &  n166 ;
  assign n673 = n422 | n647 ;
  assign n938 = n673 | n923 ;
  assign n939 = ( n829 & ~n503 ) | ( n829 & n938 ) | ( ~n503 & n938 ) ;
  assign n940 = n503 | n939 ;
  assign n941 = n324 | n940 ;
  assign n419 = ( n90 & ~n101 ) | ( n90 & 1'b0 ) | ( ~n101 & 1'b0 ) ;
  assign n497 = n129 | n419 ;
  assign n498 = n361 | n497 ;
  assign n393 = n201 | n392 ;
  assign n644 = n393 | n643 ;
  assign n942 = n498 | n644 ;
  assign n943 = ( n922 & ~n444 ) | ( n922 & n942 ) | ( ~n444 & n942 ) ;
  assign n944 = n444 | n943 ;
  assign n945 = ( n941 & ~n105 ) | ( n941 & n944 ) | ( ~n105 & n944 ) ;
  assign n946 = n105 | n945 ;
  assign n947 = ( n169 & ~n124 ) | ( n169 & n946 ) | ( ~n124 & n946 ) ;
  assign n948 = n124 | n947 ;
  assign n949 = ( n143 & ~n948 ) | ( n143 & n645 ) | ( ~n948 & n645 ) ;
  assign n950 = ~n143 & n949 ;
  assign n951 = ( n275 & ~n612 ) | ( n275 & n950 ) | ( ~n612 & n950 ) ;
  assign n952 = ~n275 & n951 ;
  assign n953 = ( n106 & n112 ) | ( n106 & n146 ) | ( n112 & n146 ) ;
  assign n954 = ( n146 & ~n953 ) | ( n146 & 1'b0 ) | ( ~n953 & 1'b0 ) ;
  assign n955 = ( n84 & ~n125 ) | ( n84 & n94 ) | ( ~n125 & n94 ) ;
  assign n956 = ~n84 & n955 ;
  assign n957 = ( n107 & ~n96 ) | ( n107 & n148 ) | ( ~n96 & n148 ) ;
  assign n958 = n96 | n957 ;
  assign n379 = ~n53 & n71 ;
  assign n454 = n149 | n379 ;
  assign n637 = n381 | n443 ;
  assign n961 = n454 | n637 ;
  assign n959 = ~n62 & n145 ;
  assign n960 = ( n62 & ~n101 ) | ( n62 & n959 ) | ( ~n101 & n959 ) ;
  assign n962 = ( n101 & ~n961 ) | ( n101 & n960 ) | ( ~n961 & n960 ) ;
  assign n963 = ( n148 & ~n958 ) | ( n148 & n962 ) | ( ~n958 & n962 ) ;
  assign n964 = ( n437 & ~n355 ) | ( n437 & n963 ) | ( ~n355 & n963 ) ;
  assign n965 = ~n437 & n964 ;
  assign n278 = ~n53 & n102 ;
  assign n279 = n109 | n229 ;
  assign n280 = n278 | n279 ;
  assign n560 = n93 &  n117 ;
  assign n561 = n436 | n560 ;
  assign n966 = n280 | n561 ;
  assign n967 = ( n495 & ~n966 ) | ( n495 & 1'b0 ) | ( ~n966 & 1'b0 ) ;
  assign n968 = ( n359 & n965 ) | ( n359 & n967 ) | ( n965 & n967 ) ;
  assign n969 = ~n359 & n968 ;
  assign n970 = ( n956 & ~n94 ) | ( n956 & n969 ) | ( ~n94 & n969 ) ;
  assign n971 = ~n230 & n970 ;
  assign n972 = ( n106 & n954 ) | ( n106 & n971 ) | ( n954 & n971 ) ;
  assign n973 = ~n189 & n972 ;
  assign n974 = ( n112 & ~n77 ) | ( n112 & n146 ) | ( ~n77 & n146 ) ;
  assign n975 = ( n146 & ~n974 ) | ( n146 & 1'b0 ) | ( ~n974 & 1'b0 ) ;
  assign n976 = ( n77 & ~n90 ) | ( n77 & n179 ) | ( ~n90 & n179 ) ;
  assign n977 = ~n179 & n976 ;
  assign n596 = n293 | n595 ;
  assign n978 = ( n77 & ~n977 ) | ( n77 & n596 ) | ( ~n977 & n596 ) ;
  assign n979 = ( n77 & ~n975 ) | ( n77 & n978 ) | ( ~n975 & n978 ) ;
  assign n615 = n190 | n354 ;
  assign n668 = n330 | n353 ;
  assign n669 = n140 | n668 ;
  assign n403 = n186 | n402 ;
  assign n182 = n104 &  n121 ;
  assign n980 = n182 | n352 ;
  assign n981 = ( n116 & ~n78 ) | ( n116 & n980 ) | ( ~n78 & n980 ) ;
  assign n982 = n78 | n981 ;
  assign n983 = ( n403 & ~n669 ) | ( n403 & n982 ) | ( ~n669 & n982 ) ;
  assign n984 = n669 | n983 ;
  assign n985 = ( n615 & ~n979 ) | ( n615 & n984 ) | ( ~n979 & n984 ) ;
  assign n986 = n979 | n985 ;
  assign n987 = n115 | n986 ;
  assign n988 = ( n973 & ~n987 ) | ( n973 & 1'b0 ) | ( ~n987 & 1'b0 ) ;
  assign n989 = ( n126 & n952 ) | ( n126 & n988 ) | ( n952 & n988 ) ;
  assign n990 = ~n126 & n989 ;
  assign n991 = ( n380 & ~n501 ) | ( n380 & n990 ) | ( ~n501 & n990 ) ;
  assign n992 = ~n380 & n991 ;
  assign n993 = n937 | n992 ;
  assign n1079 = n937 &  n992 ;
  assign n1080 = ( n993 & ~n1079 ) | ( n993 & 1'b0 ) | ( ~n1079 & 1'b0 ) ;
  assign n521 = ~x22 & n36 ;
  assign n522 = x13 | n521 ;
  assign n523 = ( x13 & ~n521 ) | ( x13 & 1'b0 ) | ( ~n521 & 1'b0 ) ;
  assign n524 = ( x13 & ~n522 ) | ( x13 & ~n523 ) | ( ~n522 & ~n523 ) ;
  assign n434 = ( n53 & ~n179 ) | ( n53 & n166 ) | ( ~n179 & n166 ) ;
  assign n435 = n179 | n434 ;
  assign n439 = ( n437 & ~n119 ) | ( n437 & n438 ) | ( ~n119 & n438 ) ;
  assign n440 = n119 | n439 ;
  assign n441 = ( n436 & ~n212 ) | ( n436 & n440 ) | ( ~n212 & n440 ) ;
  assign n442 = n212 | n441 ;
  assign n196 = n104 &  n166 ;
  assign n291 = ( n102 & ~n148 ) | ( n102 & 1'b0 ) | ( ~n148 & 1'b0 ) ;
  assign n455 = ( n291 & ~n196 ) | ( n291 & n454 ) | ( ~n196 & n454 ) ;
  assign n456 = n196 | n455 ;
  assign n457 = ( n378 & ~n456 ) | ( n378 & 1'b0 ) | ( ~n456 & 1'b0 ) ;
  assign n458 = ~n453 & n457 ;
  assign n459 = ( n442 & ~n452 ) | ( n442 & n458 ) | ( ~n452 & n458 ) ;
  assign n460 = ( n126 & ~n442 ) | ( n126 & n459 ) | ( ~n442 & n459 ) ;
  assign n461 = ~n126 & n460 ;
  assign n462 = ( n160 & ~n169 ) | ( n160 & n461 ) | ( ~n169 & n461 ) ;
  assign n463 = ~n160 & n462 ;
  assign n464 = ( n364 & ~n354 ) | ( n364 & n463 ) | ( ~n354 & n463 ) ;
  assign n465 = ~n364 & n464 ;
  assign n466 = ~n128 & n465 ;
  assign n469 = ~n93 & n84 ;
  assign n470 = ( n84 & ~n469 ) | ( n84 & n411 ) | ( ~n469 & n411 ) ;
  assign n471 = n103 | n470 ;
  assign n472 = ( n468 & ~n190 ) | ( n468 & n471 ) | ( ~n190 & n471 ) ;
  assign n473 = n190 | n472 ;
  assign n474 = n261 | n473 ;
  assign n475 = n113 | n276 ;
  assign n476 = n208 | n282 ;
  assign n477 = n211 | n476 ;
  assign n479 = n362 | n478 ;
  assign n480 = n477 | n479 ;
  assign n481 = ( n475 & ~n474 ) | ( n475 & n480 ) | ( ~n474 & n480 ) ;
  assign n482 = n474 | n481 ;
  assign n483 = ( n322 & ~n380 ) | ( n322 & n482 ) | ( ~n380 & n482 ) ;
  assign n484 = n380 | n483 ;
  assign n485 = ( n467 & ~n122 ) | ( n467 & n484 ) | ( ~n122 & n484 ) ;
  assign n486 = n122 | n485 ;
  assign n488 = n94 &  n102 ;
  assign n489 = ~n152 & n418 ;
  assign n490 = ( n488 & ~n192 ) | ( n488 & n489 ) | ( ~n192 & n489 ) ;
  assign n491 = ~n488 & n490 ;
  assign n492 = ( n109 & ~n355 ) | ( n109 & n491 ) | ( ~n355 & n491 ) ;
  assign n493 = ~n109 & n492 ;
  assign n494 = ~n487 & n493 ;
  assign n164 = n77 &  n125 ;
  assign n499 = n164 | n324 ;
  assign n500 = n209 | n499 ;
  assign n502 = n91 | n501 ;
  assign n504 = n141 | n503 ;
  assign n505 = n165 | n504 ;
  assign n506 = n502 | n505 ;
  assign n507 = ( n500 & ~n498 ) | ( n500 & n506 ) | ( ~n498 & n506 ) ;
  assign n508 = ( n496 & n498 ) | ( n496 & n507 ) | ( n498 & n507 ) ;
  assign n509 = ( n496 & ~n508 ) | ( n496 & 1'b0 ) | ( ~n508 & 1'b0 ) ;
  assign n510 = ( n486 & n494 ) | ( n486 & n509 ) | ( n494 & n509 ) ;
  assign n511 = ~n486 & n510 ;
  assign n512 = ( n422 & n466 ) | ( n422 & n511 ) | ( n466 & n511 ) ;
  assign n513 = ~n422 & n512 ;
  assign n514 = ~n227 & n513 ;
  assign n515 = ( n53 & ~n435 ) | ( n53 & n514 ) | ( ~n435 & n514 ) ;
  assign n1082 = ~n937 & n992 ;
  assign n1083 = ( n515 & ~n1082 ) | ( n515 & 1'b0 ) | ( ~n1082 & 1'b0 ) ;
  assign n1123 = n524 | n1083 ;
  assign n994 = ( n515 & ~n992 ) | ( n515 & n993 ) | ( ~n992 & n993 ) ;
  assign n1124 = n524 &  n994 ;
  assign n1125 = ( n1080 & ~n1123 ) | ( n1080 & n1124 ) | ( ~n1123 & n1124 ) ;
  assign n537 = ~x22 & n37 ;
  assign n538 = ~x14 & n537 ;
  assign n539 = ( x14 & ~n537 ) | ( x14 & 1'b0 ) | ( ~n537 & 1'b0 ) ;
  assign n540 = n538 | n539 ;
  assign n1126 = n1080 | n1083 ;
  assign n1127 = n540 &  n1126 ;
  assign n1081 = ( n994 & ~n1080 ) | ( n994 & 1'b0 ) | ( ~n1080 & 1'b0 ) ;
  assign n1128 = n540 | n1081 ;
  assign n1129 = ( n1125 & ~n1127 ) | ( n1125 & n1128 ) | ( ~n1127 & n1128 ) ;
  assign n787 = ~n168 & n100 ;
  assign n747 = n181 | n276 ;
  assign n748 = ( n746 & ~n444 ) | ( n746 & n747 ) | ( ~n444 & n747 ) ;
  assign n749 = n444 | n748 ;
  assign n750 = ( n182 & ~n115 ) | ( n182 & n749 ) | ( ~n115 & n749 ) ;
  assign n751 = n115 | n750 ;
  assign n752 = ( n201 & ~n745 ) | ( n201 & n751 ) | ( ~n745 & n751 ) ;
  assign n753 = ( n745 & ~n141 ) | ( n745 & n752 ) | ( ~n141 & n752 ) ;
  assign n754 = n141 | n753 ;
  assign n759 = ( n419 & ~n470 ) | ( n419 & n758 ) | ( ~n470 & n758 ) ;
  assign n760 = ( n470 & ~n97 ) | ( n470 & n759 ) | ( ~n97 & n759 ) ;
  assign n761 = n97 | n760 ;
  assign n762 = ( n101 & ~n161 ) | ( n101 & n102 ) | ( ~n161 & n102 ) ;
  assign n763 = n161 | n762 ;
  assign n163 = n160 | n162 ;
  assign n764 = n127 | n163 ;
  assign n765 = ( n763 & ~n101 ) | ( n763 & n764 ) | ( ~n101 & n764 ) ;
  assign n766 = n199 | n765 ;
  assign n767 = ( n323 & ~n192 ) | ( n323 & n766 ) | ( ~n192 & n766 ) ;
  assign n768 = n192 | n767 ;
  assign n769 = ( n761 & ~n755 ) | ( n761 & n768 ) | ( ~n755 & n768 ) ;
  assign n770 = ( n755 & ~n196 ) | ( n755 & n769 ) | ( ~n196 & n769 ) ;
  assign n771 = n196 | n770 ;
  assign n772 = ( n118 & ~n105 ) | ( n118 & n771 ) | ( ~n105 & n771 ) ;
  assign n773 = n105 | n772 ;
  assign n774 = ( n418 & ~n773 ) | ( n418 & n478 ) | ( ~n773 & n478 ) ;
  assign n775 = ~n478 & n774 ;
  assign n776 = ~n110 & n775 ;
  assign n167 = ~n101 & n166 ;
  assign n616 = n129 | n167 ;
  assign n777 = ~n100 & n71 ;
  assign n778 = ( n71 & ~n777 ) | ( n71 & n200 ) | ( ~n777 & n200 ) ;
  assign n779 = ( n311 & ~n443 ) | ( n311 & n778 ) | ( ~n443 & n778 ) ;
  assign n780 = ( n443 & ~n109 ) | ( n443 & n779 ) | ( ~n109 & n779 ) ;
  assign n781 = n109 | n780 ;
  assign n782 = ( n616 & n776 ) | ( n616 & n781 ) | ( n776 & n781 ) ;
  assign n783 = ( n776 & ~n782 ) | ( n776 & 1'b0 ) | ( ~n782 & 1'b0 ) ;
  assign n784 = ( n315 & ~n754 ) | ( n315 & n783 ) | ( ~n754 & n783 ) ;
  assign n785 = ~n315 & n784 ;
  assign n786 = ( n169 & ~n446 ) | ( n169 & n785 ) | ( ~n446 & n785 ) ;
  assign n788 = ( n787 & ~n100 ) | ( n787 & n786 ) | ( ~n100 & n786 ) ;
  assign n1118 = ~x22 & n27 ;
  assign n1119 = ~x4 & n1118 ;
  assign n1120 = ( x4 & ~n1118 ) | ( x4 & 1'b0 ) | ( ~n1118 & 1'b0 ) ;
  assign n1121 = n1119 | n1120 ;
  assign n1122 = ~n788 & n1121 ;
  assign n1130 = ( n937 & ~n1129 ) | ( n937 & n1122 ) | ( ~n1129 & n1122 ) ;
  assign n1288 = ( n937 & ~n1122 ) | ( n937 & n1129 ) | ( ~n1122 & n1129 ) ;
  assign n1289 = ( n1130 & ~n937 ) | ( n1130 & n1288 ) | ( ~n937 & n1288 ) ;
  assign n1177 = ( n53 & ~n166 ) | ( n53 & n90 ) | ( ~n166 & n90 ) ;
  assign n1178 = n166 | n1177 ;
  assign n1179 = n89 | n62 ;
  assign n1180 = ( n62 & ~n1179 ) | ( n62 & n86 ) | ( ~n1179 & n86 ) ;
  assign n1181 = ( n71 & ~n121 ) | ( n71 & n104 ) | ( ~n121 & n104 ) ;
  assign n1182 = ~n71 & n1181 ;
  assign n831 = n468 | n647 ;
  assign n1183 = n195 | n831 ;
  assign n1184 = ( n422 & ~n149 ) | ( n422 & n1183 ) | ( ~n149 & n1183 ) ;
  assign n1185 = n149 | n1184 ;
  assign n1186 = ( n186 & ~n317 ) | ( n186 & n1185 ) | ( ~n317 & n1185 ) ;
  assign n1187 = ( n317 & ~n97 ) | ( n317 & n1186 ) | ( ~n97 & n1186 ) ;
  assign n1188 = n97 | n1187 ;
  assign n1189 = ( n554 & ~n437 ) | ( n554 & n1188 ) | ( ~n437 & n1188 ) ;
  assign n1190 = n437 | n1189 ;
  assign n1191 = n291 | n503 ;
  assign n1192 = n275 | n1191 ;
  assign n576 = ( n71 & ~n161 ) | ( n71 & n121 ) | ( ~n161 & n121 ) ;
  assign n577 = ~n576 & n161 ;
  assign n578 = ( n577 & ~n148 ) | ( n577 & n576 ) | ( ~n148 & n576 ) ;
  assign n579 = n330 | n578 ;
  assign n1193 = n579 | n616 ;
  assign n1194 = ( n1192 & ~n279 ) | ( n1192 & n1193 ) | ( ~n279 & n1193 ) ;
  assign n1195 = n279 | n1194 ;
  assign n646 = ~n402 & n645 ;
  assign n1196 = ( n310 & ~n1195 ) | ( n310 & n646 ) | ( ~n1195 & n646 ) ;
  assign n1197 = ~n310 & n1196 ;
  assign n1198 = ( n323 & ~n1197 ) | ( n323 & n418 ) | ( ~n1197 & n418 ) ;
  assign n1199 = ( n418 & ~n1198 ) | ( n418 & 1'b0 ) | ( ~n1198 & 1'b0 ) ;
  assign n1200 = ( n208 & ~n261 ) | ( n208 & n1199 ) | ( ~n261 & n1199 ) ;
  assign n1201 = ~n208 & n1200 ;
  assign n266 = ( n77 & ~n146 ) | ( n77 & 1'b0 ) | ( ~n146 & 1'b0 ) ;
  assign n1202 = ~n293 & n495 ;
  assign n1203 = ( n147 & ~n277 ) | ( n147 & n1202 ) | ( ~n277 & n1202 ) ;
  assign n1204 = ~n147 & n1203 ;
  assign n1205 = ( n266 & ~n362 ) | ( n266 & n1204 ) | ( ~n362 & n1204 ) ;
  assign n1206 = ~n266 & n1205 ;
  assign n1207 = ( n190 & ~n487 ) | ( n190 & n1206 ) | ( ~n487 & n1206 ) ;
  assign n1208 = ~n190 & n1207 ;
  assign n1209 = ~n128 & n1208 ;
  assign n1210 = ~n600 & n1209 ;
  assign n1211 = ( n766 & n1201 ) | ( n766 & n1210 ) | ( n1201 & n1210 ) ;
  assign n1212 = ~n766 & n1211 ;
  assign n1213 = ~n1190 & n1212 ;
  assign n1214 = ( n1182 & ~n104 ) | ( n1182 & n1213 ) | ( ~n104 & n1213 ) ;
  assign n1215 = ( n1180 & ~n86 ) | ( n1180 & n1214 ) | ( ~n86 & n1214 ) ;
  assign n1216 = ( n53 & ~n1178 ) | ( n53 & n1215 ) | ( ~n1178 & n1215 ) ;
  assign n1217 = ~n185 & n1216 ;
  assign n1255 = n524 &  n937 ;
  assign n1256 = n1217 &  n1255 ;
  assign n1254 = ( n540 & n937 ) | ( n540 & n1217 ) | ( n937 & n1217 ) ;
  assign n1257 = n540 | n937 ;
  assign n1258 = ( n1256 & ~n1254 ) | ( n1256 & n1257 ) | ( ~n1254 & n1257 ) ;
  assign n707 = n96 | n48 ;
  assign n686 = n93 &  n146 ;
  assign n670 = ( n667 & ~n120 ) | ( n667 & n669 ) | ( ~n120 & n669 ) ;
  assign n671 = n120 | n670 ;
  assign n672 = n317 | n391 ;
  assign n226 = ~n148 & n166 ;
  assign n610 = ~n148 & n161 ;
  assign n674 = n226 | n610 ;
  assign n675 = ( n198 & ~n186 ) | ( n198 & n674 ) | ( ~n186 & n674 ) ;
  assign n676 = n186 | n675 ;
  assign n677 = n116 | n676 ;
  assign n681 = ( n677 & ~n673 ) | ( n677 & n680 ) | ( ~n673 & n680 ) ;
  assign n682 = ( n673 & ~n672 ) | ( n673 & n681 ) | ( ~n672 & n681 ) ;
  assign n683 = n672 | n682 ;
  assign n684 = n671 | n683 ;
  assign n685 = n78 | n684 ;
  assign n687 = ( n93 & ~n686 ) | ( n93 & n685 ) | ( ~n686 & n685 ) ;
  assign n142 = ~n53 & n125 ;
  assign n688 = ~n58 & n66 ;
  assign n689 = ( n53 & ~n688 ) | ( n53 & n66 ) | ( ~n688 & n66 ) ;
  assign n692 = n209 | n266 ;
  assign n693 = n487 | n643 ;
  assign n694 = ( n360 & ~n692 ) | ( n360 & n693 ) | ( ~n692 & n693 ) ;
  assign n695 = n692 | n694 ;
  assign n696 = ( n691 & ~n69 ) | ( n691 & n695 ) | ( ~n69 & n695 ) ;
  assign n697 = n69 | n696 ;
  assign n698 = ( n689 & ~n53 ) | ( n689 & n697 ) | ( ~n53 & n697 ) ;
  assign n699 = n282 | n698 ;
  assign n700 = ( n436 & ~n379 ) | ( n436 & n699 ) | ( ~n379 & n699 ) ;
  assign n701 = ( n379 & ~n142 ) | ( n379 & n700 ) | ( ~n142 & n700 ) ;
  assign n702 = n142 | n701 ;
  assign n703 = n281 | n702 ;
  assign n704 = ( n687 & ~n319 ) | ( n687 & n703 ) | ( ~n319 & n703 ) ;
  assign n705 = ( n319 & ~n278 ) | ( n319 & n704 ) | ( ~n278 & n704 ) ;
  assign n706 = n278 | n705 ;
  assign n708 = ( n707 & ~n48 ) | ( n707 & n706 ) | ( ~n48 & n706 ) ;
  assign n724 = ( n502 & ~n364 ) | ( n502 & n723 ) | ( ~n364 & n723 ) ;
  assign n725 = ( n364 & ~n275 ) | ( n364 & n724 ) | ( ~n275 & n724 ) ;
  assign n726 = n275 | n725 ;
  assign n727 = ( n208 & ~n180 ) | ( n208 & n726 ) | ( ~n180 & n726 ) ;
  assign n728 = n180 | n727 ;
  assign n729 = n290 | n728 ;
  assign n571 = n83 | n62 ;
  assign n572 = ( n62 & ~n571 ) | ( n62 & n77 ) | ( ~n571 & n77 ) ;
  assign n732 = ( n615 & ~n302 ) | ( n615 & n731 ) | ( ~n302 & n731 ) ;
  assign n733 = n302 | n732 ;
  assign n734 = ( n398 & ~n143 ) | ( n398 & n733 ) | ( ~n143 & n733 ) ;
  assign n735 = n143 | n734 ;
  assign n736 = ( n77 & ~n572 ) | ( n77 & n735 ) | ( ~n572 & n735 ) ;
  assign n737 = ( n691 & ~n359 ) | ( n691 & n736 ) | ( ~n359 & n736 ) ;
  assign n738 = ( n359 & ~n687 ) | ( n359 & n737 ) | ( ~n687 & n737 ) ;
  assign n739 = n687 | n738 ;
  assign n740 = ( n729 & ~n122 ) | ( n729 & n739 ) | ( ~n122 & n739 ) ;
  assign n741 = n122 | n740 ;
  assign n1172 = ~x22 & n26 ;
  assign n1173 = x3 | n1172 ;
  assign n1174 = ( x3 & ~n1172 ) | ( x3 & 1'b0 ) | ( ~n1172 & 1'b0 ) ;
  assign n1175 = ( n1173 & ~x3 ) | ( n1173 & n1174 ) | ( ~x3 & n1174 ) ;
  assign n1259 = ( n708 & n741 ) | ( n708 & n1175 ) | ( n741 & n1175 ) ;
  assign n1260 = n788 | n1259 ;
  assign n1261 = ( n1258 & ~n1260 ) | ( n1258 & 1'b0 ) | ( ~n1260 & 1'b0 ) ;
  assign n795 = n708 | n741 ;
  assign n796 = n788 &  n795 ;
  assign n1262 = ~n796 & n1121 ;
  assign n742 = n708 &  n741 ;
  assign n743 = ~n708 & n741 ;
  assign n744 = ( n708 & ~n742 ) | ( n708 & n743 ) | ( ~n742 & n743 ) ;
  assign n789 = n742 | n788 ;
  assign n1263 = ( n789 & ~n1121 ) | ( n789 & 1'b0 ) | ( ~n1121 & 1'b0 ) ;
  assign n1264 = ( n1262 & ~n744 ) | ( n1262 & n1263 ) | ( ~n744 & n1263 ) ;
  assign n801 = n744 &  n789 ;
  assign n1074 = ~x22 & n28 ;
  assign n1075 = x5 | n1074 ;
  assign n1076 = ( x5 & ~n1074 ) | ( x5 & 1'b0 ) | ( ~n1074 & 1'b0 ) ;
  assign n1077 = ( x5 & ~n1075 ) | ( x5 & ~n1076 ) | ( ~n1075 & ~n1076 ) ;
  assign n1266 = ~n801 & n1077 ;
  assign n799 = ( n744 & ~n796 ) | ( n744 & 1'b0 ) | ( ~n796 & 1'b0 ) ;
  assign n1265 = n799 | n1077 ;
  assign n1267 = ( n1264 & ~n1266 ) | ( n1264 & n1265 ) | ( ~n1266 & n1265 ) ;
  assign n382 = n196 | n381 ;
  assign n383 = ( n290 & ~n380 ) | ( n290 & n382 ) | ( ~n380 & n382 ) ;
  assign n384 = n380 | n383 ;
  assign n385 = ( n379 & ~n140 ) | ( n379 & n384 ) | ( ~n140 & n384 ) ;
  assign n386 = n140 | n385 ;
  assign n387 = ( n278 & n378 ) | ( n278 & n386 ) | ( n378 & n386 ) ;
  assign n388 = ( n378 & ~n387 ) | ( n378 & 1'b0 ) | ( ~n387 & 1'b0 ) ;
  assign n389 = ( n53 & ~n112 ) | ( n53 & n96 ) | ( ~n112 & n96 ) ;
  assign n390 = n112 | n389 ;
  assign n394 = n391 | n393 ;
  assign n395 = ( n291 & ~n192 ) | ( n291 & n394 ) | ( ~n192 & n394 ) ;
  assign n396 = n192 | n395 ;
  assign n397 = n122 | n396 ;
  assign n399 = n108 | n398 ;
  assign n400 = n152 | n185 ;
  assign n401 = n189 | n400 ;
  assign n404 = n401 | n403 ;
  assign n405 = ( n399 & ~n397 ) | ( n399 & n404 ) | ( ~n397 & n404 ) ;
  assign n406 = ( n397 & ~n162 ) | ( n397 & n405 ) | ( ~n162 & n405 ) ;
  assign n407 = n162 | n406 ;
  assign n408 = ( n229 & ~n116 ) | ( n229 & n407 ) | ( ~n116 & n407 ) ;
  assign n409 = n116 | n408 ;
  assign n410 = ( n390 & ~n53 ) | ( n390 & n409 ) | ( ~n53 & n409 ) ;
  assign n413 = n411 | n412 ;
  assign n414 = ( n292 & ~n275 ) | ( n292 & n413 ) | ( ~n275 & n413 ) ;
  assign n415 = n275 | n414 ;
  assign n416 = ( n282 & ~n142 ) | ( n282 & n415 ) | ( ~n142 & n415 ) ;
  assign n417 = n142 | n416 ;
  assign n423 = n226 | n422 ;
  assign n424 = n199 | n423 ;
  assign n420 = ( n418 & ~n419 ) | ( n418 & 1'b0 ) | ( ~n419 & 1'b0 ) ;
  assign n421 = ~n302 & n420 ;
  assign n425 = ( n417 & ~n424 ) | ( n417 & n421 ) | ( ~n424 & n421 ) ;
  assign n426 = ~n417 & n425 ;
  assign n427 = ~n410 & n426 ;
  assign n428 = ( n377 & n388 ) | ( n377 & n427 ) | ( n388 & n427 ) ;
  assign n429 = ( n352 & ~n377 ) | ( n352 & n428 ) | ( ~n377 & n428 ) ;
  assign n430 = ~n352 & n429 ;
  assign n431 = ~n211 & n430 ;
  assign n432 = ( n68 & ~n93 ) | ( n68 & 1'b0 ) | ( ~n93 & 1'b0 ) ;
  assign n433 = ( n431 & ~n68 ) | ( n431 & n432 ) | ( ~n68 & n432 ) ;
  assign n806 = ( n106 & ~n166 ) | ( n106 & n125 ) | ( ~n166 & n125 ) ;
  assign n807 = n166 | n806 ;
  assign n573 = n91 | n169 ;
  assign n312 = n140 | n311 ;
  assign n808 = ( n312 & ~n211 ) | ( n312 & n643 ) | ( ~n211 & n643 ) ;
  assign n809 = n211 | n808 ;
  assign n810 = n143 | n160 ;
  assign n811 = ( n317 & ~n197 ) | ( n317 & n810 ) | ( ~n197 & n810 ) ;
  assign n812 = n197 | n811 ;
  assign n648 = n103 | n315 ;
  assign n649 = n318 | n648 ;
  assign n813 = n78 | n478 ;
  assign n814 = n379 | n813 ;
  assign n815 = n110 | n153 ;
  assign n816 = n186 | n815 ;
  assign n817 = ( n814 & ~n649 ) | ( n814 & n816 ) | ( ~n649 & n816 ) ;
  assign n818 = n649 | n817 ;
  assign n819 = ( n812 & ~n380 ) | ( n812 & n818 ) | ( ~n380 & n818 ) ;
  assign n820 = n380 | n819 ;
  assign n821 = ( n323 & ~n291 ) | ( n323 & n820 ) | ( ~n291 & n820 ) ;
  assign n822 = n291 | n821 ;
  assign n823 = ( n275 & ~n109 ) | ( n275 & n822 ) | ( ~n109 & n822 ) ;
  assign n824 = n109 | n823 ;
  assign n825 = n69 | n824 ;
  assign n613 = ( n90 & ~n161 ) | ( n90 & n104 ) | ( ~n161 & n104 ) ;
  assign n614 = ~n90 & n613 ;
  assign n264 = ( n121 & ~n107 ) | ( n121 & n148 ) | ( ~n107 & n148 ) ;
  assign n265 = n107 | n264 ;
  assign n270 = n106 &  n68 ;
  assign n269 = n266 | n268 ;
  assign n271 = ( n68 & ~n270 ) | ( n68 & n269 ) | ( ~n270 & n269 ) ;
  assign n272 = n200 | n271 ;
  assign n273 = ( n265 & ~n148 ) | ( n265 & n272 ) | ( ~n148 & n272 ) ;
  assign n274 = n128 | n273 ;
  assign n617 = n127 | n616 ;
  assign n618 = n615 | n617 ;
  assign n619 = n274 | n618 ;
  assign n620 = ( n104 & ~n614 ) | ( n104 & n619 ) | ( ~n614 & n619 ) ;
  assign n621 = ( n191 & ~n105 ) | ( n191 & n620 ) | ( ~n105 & n620 ) ;
  assign n622 = n105 | n621 ;
  assign n623 = ( n289 & ~n612 ) | ( n289 & n622 ) | ( ~n612 & n622 ) ;
  assign n624 = n612 | n623 ;
  assign n625 = ( n324 & ~n361 ) | ( n324 & n624 ) | ( ~n361 & n624 ) ;
  assign n626 = n361 | n625 ;
  assign n828 = n118 | n827 ;
  assign n832 = ( n830 & ~n123 ) | ( n830 & n831 ) | ( ~n123 & n831 ) ;
  assign n833 = n123 | n832 ;
  assign n834 = ( n278 & ~n230 ) | ( n278 & n833 ) | ( ~n230 & n833 ) ;
  assign n835 = n230 | n834 ;
  assign n836 = ( n353 & ~n180 ) | ( n353 & n835 ) | ( ~n180 & n835 ) ;
  assign n837 = n180 | n836 ;
  assign n838 = ( n829 & ~n828 ) | ( n829 & n837 ) | ( ~n828 & n837 ) ;
  assign n839 = ( n828 & ~n626 ) | ( n828 & n838 ) | ( ~n626 & n838 ) ;
  assign n840 = n626 | n839 ;
  assign n841 = ( n826 & ~n825 ) | ( n826 & n840 ) | ( ~n825 & n840 ) ;
  assign n842 = n825 | n841 ;
  assign n843 = ( n809 & ~n147 ) | ( n809 & n842 ) | ( ~n147 & n842 ) ;
  assign n844 = n147 | n843 ;
  assign n845 = ( n573 & ~n723 ) | ( n573 & n844 ) | ( ~n723 & n844 ) ;
  assign n846 = n723 | n845 ;
  assign n847 = ( n807 & ~n106 ) | ( n807 & n846 ) | ( ~n106 & n846 ) ;
  assign n848 = n433 &  n847 ;
  assign n849 = n433 | n847 ;
  assign n850 = ~n848 & n849 ;
  assign n546 = ( n311 & ~n488 ) | ( n311 & n361 ) | ( ~n488 & n361 ) ;
  assign n547 = n488 | n546 ;
  assign n548 = ( n191 & ~n190 ) | ( n191 & n547 ) | ( ~n190 & n547 ) ;
  assign n549 = n190 | n548 ;
  assign n550 = ( n293 & ~n310 ) | ( n293 & n505 ) | ( ~n310 & n505 ) ;
  assign n551 = n310 | n550 ;
  assign n552 = ( n379 & ~n186 ) | ( n379 & n551 ) | ( ~n186 & n551 ) ;
  assign n553 = n186 | n552 ;
  assign n150 = n62 &  n58 ;
  assign n151 = ( n58 & ~n150 ) | ( n58 & n101 ) | ( ~n150 & n101 ) ;
  assign n155 = ( n151 & ~n101 ) | ( n151 & n154 ) | ( ~n101 & n154 ) ;
  assign n156 = ( n149 & ~n147 ) | ( n149 & n155 ) | ( ~n147 & n155 ) ;
  assign n157 = n147 | n156 ;
  assign n158 = ( n143 & ~n142 ) | ( n143 & n157 ) | ( ~n142 & n157 ) ;
  assign n159 = n142 | n158 ;
  assign n564 = ( n477 & ~n561 ) | ( n477 & n563 ) | ( ~n561 & n563 ) ;
  assign n565 = n561 | n564 ;
  assign n566 = ( n559 & ~n159 ) | ( n559 & n565 ) | ( ~n159 & n565 ) ;
  assign n567 = n159 | n566 ;
  assign n568 = ( n391 & ~n105 ) | ( n391 & n567 ) | ( ~n105 & n567 ) ;
  assign n569 = n105 | n568 ;
  assign n570 = n554 | n569 ;
  assign n574 = ( n77 & ~n572 ) | ( n77 & n573 ) | ( ~n572 & n573 ) ;
  assign n575 = n281 | n574 ;
  assign n580 = n317 | n398 ;
  assign n581 = n266 | n580 ;
  assign n582 = n139 | n201 ;
  assign n583 = n290 | n582 ;
  assign n585 = ( n583 & ~n581 ) | ( n583 & n584 ) | ( ~n581 & n584 ) ;
  assign n586 = n581 | n585 ;
  assign n587 = ( n579 & ~n575 ) | ( n579 & n586 ) | ( ~n575 & n586 ) ;
  assign n588 = n575 | n587 ;
  assign n589 = ( n570 & ~n553 ) | ( n570 & n588 ) | ( ~n553 & n588 ) ;
  assign n590 = ( n553 & ~n549 ) | ( n553 & n589 ) | ( ~n549 & n589 ) ;
  assign n591 = n549 | n590 ;
  assign n592 = n437 | n591 ;
  assign n858 = ( n433 & ~n849 ) | ( n433 & n592 ) | ( ~n849 & n592 ) ;
  assign n863 = n850 | n858 ;
  assign n1277 = ~n248 & n863 ;
  assign n790 = ~x22 & n30 ;
  assign n791 = x7 | n790 ;
  assign n792 = ( x7 & ~n790 ) | ( x7 & 1'b0 ) | ( ~n790 & 1'b0 ) ;
  assign n793 = ( x7 & ~n791 ) | ( x7 & ~n792 ) | ( ~n791 & ~n792 ) ;
  assign n1274 = ( n793 & ~n858 ) | ( n793 & 1'b0 ) | ( ~n858 & 1'b0 ) ;
  assign n851 = ( n433 & ~n847 ) | ( n433 & 1'b0 ) | ( ~n847 & 1'b0 ) ;
  assign n852 = n592 | n851 ;
  assign n1275 = ~n793 & n852 ;
  assign n1276 = ( n850 & n1274 ) | ( n850 & n1275 ) | ( n1274 & n1275 ) ;
  assign n861 = ~n850 & n852 ;
  assign n1278 = ( n248 & ~n861 ) | ( n248 & 1'b0 ) | ( ~n861 & 1'b0 ) ;
  assign n1279 = ( n1277 & ~n1276 ) | ( n1277 & n1278 ) | ( ~n1276 & n1278 ) ;
  assign n262 = ( n77 & n96 ) | ( n77 & n148 ) | ( n96 & n148 ) ;
  assign n263 = ~n77 & n262 ;
  assign n284 = ( n280 & ~n118 ) | ( n280 & n283 ) | ( ~n118 & n283 ) ;
  assign n285 = n118 | n284 ;
  assign n286 = ( n277 & ~n276 ) | ( n277 & n285 ) | ( ~n276 & n285 ) ;
  assign n287 = n276 | n286 ;
  assign n288 = n275 | n287 ;
  assign n294 = n143 | n293 ;
  assign n295 = n292 | n294 ;
  assign n296 = ( n291 & ~n129 ) | ( n291 & n295 ) | ( ~n129 & n295 ) ;
  assign n297 = n129 | n296 ;
  assign n298 = ( n208 & ~n192 ) | ( n208 & n297 ) | ( ~n192 & n297 ) ;
  assign n299 = n192 | n298 ;
  assign n300 = ( n290 & ~n289 ) | ( n290 & n299 ) | ( ~n289 & n299 ) ;
  assign n301 = n289 | n300 ;
  assign n303 = n164 | n302 ;
  assign n304 = n149 | n303 ;
  assign n305 = ( n165 & ~n142 ) | ( n165 & n304 ) | ( ~n142 & n304 ) ;
  assign n306 = n142 | n305 ;
  assign n307 = ( n53 & ~n112 ) | ( n53 & n84 ) | ( ~n112 & n84 ) ;
  assign n308 = n112 | n307 ;
  assign n313 = ( n101 & ~n117 ) | ( n101 & n107 ) | ( ~n117 & n107 ) ;
  assign n314 = n117 | n313 ;
  assign n228 = n226 | n227 ;
  assign n335 = n228 | n334 ;
  assign n336 = n329 | n335 ;
  assign n337 = ( n322 & ~n315 ) | ( n322 & n336 ) | ( ~n315 & n336 ) ;
  assign n338 = n315 | n337 ;
  assign n339 = ( n314 & ~n101 ) | ( n314 & n338 ) | ( ~n101 & n338 ) ;
  assign n340 = ( n312 & ~n147 ) | ( n312 & n339 ) | ( ~n147 & n339 ) ;
  assign n341 = n147 | n340 ;
  assign n342 = n197 | n341 ;
  assign n343 = ( n310 & ~n309 ) | ( n310 & n342 ) | ( ~n309 & n342 ) ;
  assign n344 = n309 | n343 ;
  assign n345 = ( n308 & ~n53 ) | ( n308 & n344 ) | ( ~n53 & n344 ) ;
  assign n346 = ( n306 & ~n115 ) | ( n306 & n345 ) | ( ~n115 & n345 ) ;
  assign n347 = n115 | n346 ;
  assign n348 = ( n301 & ~n288 ) | ( n301 & n347 ) | ( ~n288 & n347 ) ;
  assign n349 = ( n288 & ~n274 ) | ( n288 & n348 ) | ( ~n274 & n348 ) ;
  assign n350 = n274 | n349 ;
  assign n351 = ( n96 & ~n263 ) | ( n96 & n350 ) | ( ~n263 & n350 ) ;
  assign n516 = n433 &  n515 ;
  assign n517 = ( n261 & ~n351 ) | ( n261 & n516 ) | ( ~n351 & n516 ) ;
  assign n518 = ~n261 & n517 ;
  assign n519 = n351 | n517 ;
  assign n520 = ( n518 & ~n515 ) | ( n518 & n519 ) | ( ~n515 & n519 ) ;
  assign n710 = x9 | n244 ;
  assign n711 = ( x9 & ~n244 ) | ( x9 & 1'b0 ) | ( ~n244 & 1'b0 ) ;
  assign n712 = ( n710 & ~x9 ) | ( n710 & n711 ) | ( ~x9 & n711 ) ;
  assign n1268 = ( n520 & ~n712 ) | ( n520 & 1'b0 ) | ( ~n712 & 1'b0 ) ;
  assign n526 = n261 | n351 ;
  assign n528 = ~n433 & n526 ;
  assign n527 = n515 &  n526 ;
  assign n529 = ( n515 & ~n526 ) | ( n515 & 1'b0 ) | ( ~n526 & 1'b0 ) ;
  assign n530 = ( n528 & ~n527 ) | ( n528 & n529 ) | ( ~n527 & n529 ) ;
  assign n1269 = n530 &  n712 ;
  assign n1270 = n1268 | n1269 ;
  assign n535 = n529 &  n433 ;
  assign n533 = n515 | n526 ;
  assign n534 = ~n527 & n533 ;
  assign n536 = ( n433 & ~n535 ) | ( n433 & n534 ) | ( ~n535 & n534 ) ;
  assign n1271 = n256 &  n536 ;
  assign n542 = ( n433 & ~n527 ) | ( n433 & n526 ) | ( ~n527 & n526 ) ;
  assign n543 = ~n534 & n542 ;
  assign n1272 = n256 | n543 ;
  assign n1273 = ( n1270 & ~n1271 ) | ( n1270 & n1272 ) | ( ~n1271 & n1272 ) ;
  assign n593 = ( n53 & ~n168 ) | ( n53 & n112 ) | ( ~n168 & n112 ) ;
  assign n594 = n168 | n593 ;
  assign n598 = ( n90 & n94 ) | ( n90 & n146 ) | ( n94 & n146 ) ;
  assign n599 = ~n90 & n598 ;
  assign n601 = n115 | n600 ;
  assign n602 = ( n503 & ~n110 ) | ( n503 & n601 ) | ( ~n110 & n601 ) ;
  assign n603 = n110 | n602 ;
  assign n604 = ( n398 & ~n147 ) | ( n398 & n603 ) | ( ~n147 & n603 ) ;
  assign n605 = n147 | n604 ;
  assign n606 = ( n555 & ~n363 ) | ( n555 & n605 ) | ( ~n363 & n605 ) ;
  assign n607 = n363 | n606 ;
  assign n608 = n196 | n310 ;
  assign n609 = n85 | n608 ;
  assign n611 = n487 | n610 ;
  assign n627 = ~n182 & n418 ;
  assign n628 = ( n411 & ~n143 ) | ( n411 & n627 ) | ( ~n143 & n627 ) ;
  assign n629 = ~n411 & n628 ;
  assign n630 = ( n611 & ~n626 ) | ( n611 & n629 ) | ( ~n626 & n629 ) ;
  assign n631 = ~n611 & n630 ;
  assign n632 = ( n607 & ~n609 ) | ( n607 & n631 ) | ( ~n609 & n631 ) ;
  assign n633 = ~n607 & n632 ;
  assign n634 = ( n599 & ~n94 ) | ( n599 & n633 ) | ( ~n94 & n633 ) ;
  assign n635 = ( n185 & ~n597 ) | ( n185 & n634 ) | ( ~n597 & n634 ) ;
  assign n636 = ~n185 & n635 ;
  assign n638 = ( n479 & ~n169 ) | ( n479 & n637 ) | ( ~n169 & n637 ) ;
  assign n639 = n169 | n638 ;
  assign n640 = ( n422 & ~n309 ) | ( n422 & n639 ) | ( ~n309 & n639 ) ;
  assign n641 = n309 | n640 ;
  assign n642 = n302 | n641 ;
  assign n650 = ( n228 & ~n118 ) | ( n228 & n649 ) | ( ~n118 & n649 ) ;
  assign n651 = n118 | n650 ;
  assign n652 = ( n282 & ~n195 ) | ( n282 & n651 ) | ( ~n195 & n651 ) ;
  assign n653 = n195 | n652 ;
  assign n654 = n108 | n653 ;
  assign n655 = ( n647 & ~n380 ) | ( n647 & n654 ) | ( ~n380 & n654 ) ;
  assign n656 = n380 | n655 ;
  assign n657 = ( n644 & ~n656 ) | ( n644 & n646 ) | ( ~n656 & n646 ) ;
  assign n658 = ( n154 & ~n644 ) | ( n154 & n657 ) | ( ~n644 & n657 ) ;
  assign n659 = ~n154 & n658 ;
  assign n660 = ~n642 & n659 ;
  assign n661 = ( n596 & n636 ) | ( n596 & n660 ) | ( n636 & n660 ) ;
  assign n662 = ~n596 & n661 ;
  assign n663 = ( n53 & ~n594 ) | ( n53 & n662 ) | ( ~n594 & n662 ) ;
  assign n664 = n592 | n663 ;
  assign n665 = n592 &  n663 ;
  assign n666 = ( n664 & ~n665 ) | ( n664 & 1'b0 ) | ( ~n665 & 1'b0 ) ;
  assign n714 = ~n592 & n663 ;
  assign n715 = n708 | n714 ;
  assign n718 = ~n666 & n715 ;
  assign n995 = ~x22 & n29 ;
  assign n996 = ~x6 & n995 ;
  assign n997 = ( x6 & ~n995 ) | ( x6 & 1'b0 ) | ( ~n995 & 1'b0 ) ;
  assign n998 = n996 | n997 ;
  assign n1283 = ~n718 & n998 ;
  assign n1280 = ( n715 & ~n1077 ) | ( n715 & 1'b0 ) | ( ~n1077 & 1'b0 ) ;
  assign n709 = ( n665 & ~n592 ) | ( n665 & n708 ) | ( ~n592 & n708 ) ;
  assign n1281 = ~n709 & n1077 ;
  assign n1282 = ( n666 & n1280 ) | ( n666 & n1281 ) | ( n1280 & n1281 ) ;
  assign n720 = n666 | n709 ;
  assign n1284 = ( n720 & ~n998 ) | ( n720 & 1'b0 ) | ( ~n998 & 1'b0 ) ;
  assign n1285 = ( n1283 & ~n1282 ) | ( n1283 & n1284 ) | ( ~n1282 & n1284 ) ;
  assign n1286 = ( n1279 & ~n1273 ) | ( n1279 & n1285 ) | ( ~n1273 & n1285 ) ;
  assign n1287 = ( n1261 & ~n1267 ) | ( n1261 & n1286 ) | ( ~n1267 & n1286 ) ;
  assign n1134 = ( n256 & ~n861 ) | ( n256 & 1'b0 ) | ( ~n861 & 1'b0 ) ;
  assign n1132 = n712 | n858 ;
  assign n1131 = n712 &  n852 ;
  assign n1133 = ( n850 & ~n1132 ) | ( n850 & n1131 ) | ( ~n1132 & n1131 ) ;
  assign n1135 = ~n256 & n863 ;
  assign n1136 = ( n1134 & ~n1133 ) | ( n1134 & n1135 ) | ( ~n1133 & n1135 ) ;
  assign n1146 = ( n248 & ~n718 ) | ( n248 & 1'b0 ) | ( ~n718 & 1'b0 ) ;
  assign n1143 = ~n709 & n793 ;
  assign n1144 = ( n715 & ~n793 ) | ( n715 & 1'b0 ) | ( ~n793 & 1'b0 ) ;
  assign n1145 = ( n666 & n1143 ) | ( n666 & n1144 ) | ( n1143 & n1144 ) ;
  assign n1147 = ~n248 & n720 ;
  assign n1148 = ( n1146 & ~n1145 ) | ( n1146 & n1147 ) | ( ~n1145 & n1147 ) ;
  assign n881 = x11 | n252 ;
  assign n882 = ( x11 & ~n252 ) | ( x11 & 1'b0 ) | ( ~n252 & 1'b0 ) ;
  assign n883 = ( x11 & ~n881 ) | ( x11 & ~n882 ) | ( ~n881 & ~n882 ) ;
  assign n1137 = n520 &  n883 ;
  assign n1138 = ( n530 & ~n883 ) | ( n530 & 1'b0 ) | ( ~n883 & 1'b0 ) ;
  assign n1139 = n1137 | n1138 ;
  assign n853 = ~x22 & n35 ;
  assign n854 = ~x12 & n853 ;
  assign n855 = ( x12 & ~n853 ) | ( x12 & 1'b0 ) | ( ~n853 & 1'b0 ) ;
  assign n856 = n854 | n855 ;
  assign n1140 = n536 &  n856 ;
  assign n1141 = n543 | n856 ;
  assign n1142 = ( n1139 & ~n1140 ) | ( n1139 & n1141 ) | ( ~n1140 & n1141 ) ;
  assign n1290 = ( n1136 & ~n1148 ) | ( n1136 & n1142 ) | ( ~n1148 & n1142 ) ;
  assign n1291 = ( n1142 & ~n1136 ) | ( n1142 & n1148 ) | ( ~n1136 & n1148 ) ;
  assign n1292 = ( n1290 & ~n1142 ) | ( n1290 & n1291 ) | ( ~n1142 & n1291 ) ;
  assign n1293 = ( n1289 & ~n1287 ) | ( n1289 & n1292 ) | ( ~n1287 & n1292 ) ;
  assign n1078 = n788 | n1077 ;
  assign n1084 = ( n1080 & ~n1083 ) | ( n1080 & 1'b0 ) | ( ~n1083 & 1'b0 ) ;
  assign n1085 = ( n540 & ~n1084 ) | ( n540 & 1'b0 ) | ( ~n1084 & 1'b0 ) ;
  assign n1086 = n540 | n994 ;
  assign n1087 = ( n1081 & ~n1085 ) | ( n1081 & n1086 ) | ( ~n1085 & n1086 ) ;
  assign n1161 = ( n937 & n1078 ) | ( n937 & n1087 ) | ( n1078 & n1087 ) ;
  assign n1088 = ( n1078 & ~n937 ) | ( n1078 & n1087 ) | ( ~n937 & n1087 ) ;
  assign n1162 = ( n937 & ~n1161 ) | ( n937 & n1088 ) | ( ~n1161 & n1088 ) ;
  assign n1167 = n789 &  n1077 ;
  assign n1166 = n796 | n1077 ;
  assign n1168 = ( n744 & ~n1167 ) | ( n744 & n1166 ) | ( ~n1167 & n1166 ) ;
  assign n1170 = n801 | n998 ;
  assign n1169 = ~n799 & n998 ;
  assign n1171 = ( n1168 & ~n1170 ) | ( n1168 & n1169 ) | ( ~n1170 & n1169 ) ;
  assign n1176 = ~n788 & n1175 ;
  assign n1218 = ( n540 & ~n1217 ) | ( n540 & 1'b0 ) | ( ~n1217 & 1'b0 ) ;
  assign n1219 = ( n937 & ~n540 ) | ( n937 & n1218 ) | ( ~n540 & n1218 ) ;
  assign n1223 = ~n524 & n1126 ;
  assign n1220 = ( n856 & ~n1083 ) | ( n856 & 1'b0 ) | ( ~n1083 & 1'b0 ) ;
  assign n1221 = ~n856 & n994 ;
  assign n1222 = ( n1080 & n1220 ) | ( n1080 & n1221 ) | ( n1220 & n1221 ) ;
  assign n1224 = ( n524 & ~n1081 ) | ( n524 & 1'b0 ) | ( ~n1081 & 1'b0 ) ;
  assign n1225 = ( n1223 & ~n1222 ) | ( n1223 & n1224 ) | ( ~n1222 & n1224 ) ;
  assign n1226 = ( n1176 & n1219 ) | ( n1176 & n1225 ) | ( n1219 & n1225 ) ;
  assign n1230 = ( n712 & ~n861 ) | ( n712 & 1'b0 ) | ( ~n861 & 1'b0 ) ;
  assign n1227 = n248 | n858 ;
  assign n1228 = n248 &  n852 ;
  assign n1229 = ( n850 & ~n1227 ) | ( n850 & n1228 ) | ( ~n1227 & n1228 ) ;
  assign n1231 = ~n712 & n863 ;
  assign n1232 = ( n1230 & ~n1229 ) | ( n1230 & n1231 ) | ( ~n1229 & n1231 ) ;
  assign n1239 = n709 | n998 ;
  assign n1240 = n715 &  n998 ;
  assign n1241 = ( n666 & ~n1239 ) | ( n666 & n1240 ) | ( ~n1239 & n1240 ) ;
  assign n1243 = n720 &  n793 ;
  assign n1242 = n718 | n793 ;
  assign n1244 = ( n1241 & ~n1243 ) | ( n1241 & n1242 ) | ( ~n1243 & n1242 ) ;
  assign n1236 = ( n536 & ~n883 ) | ( n536 & 1'b0 ) | ( ~n883 & 1'b0 ) ;
  assign n1233 = ~n256 & n520 ;
  assign n1234 = n256 &  n530 ;
  assign n1235 = n1233 | n1234 ;
  assign n1237 = ~n543 & n883 ;
  assign n1238 = ( n1236 & ~n1235 ) | ( n1236 & n1237 ) | ( ~n1235 & n1237 ) ;
  assign n1245 = ( n1232 & ~n1244 ) | ( n1232 & n1238 ) | ( ~n1244 & n1238 ) ;
  assign n1246 = ( n1171 & n1226 ) | ( n1171 & n1245 ) | ( n1226 & n1245 ) ;
  assign n1093 = ~n524 & n536 ;
  assign n1090 = ( n520 & ~n856 ) | ( n520 & 1'b0 ) | ( ~n856 & 1'b0 ) ;
  assign n1091 = n530 &  n856 ;
  assign n1092 = n1090 | n1091 ;
  assign n1094 = ( n524 & ~n543 ) | ( n524 & 1'b0 ) | ( ~n543 & 1'b0 ) ;
  assign n1095 = ( n1093 & ~n1092 ) | ( n1093 & n1094 ) | ( ~n1092 & n1094 ) ;
  assign n1105 = ( n712 & ~n718 ) | ( n712 & 1'b0 ) | ( ~n718 & 1'b0 ) ;
  assign n1102 = n248 | n709 ;
  assign n1103 = n248 &  n715 ;
  assign n1104 = ( n666 & ~n1102 ) | ( n666 & n1103 ) | ( ~n1102 & n1103 ) ;
  assign n1106 = ~n712 & n720 ;
  assign n1107 = ( n1105 & ~n1104 ) | ( n1105 & n1106 ) | ( ~n1104 & n1106 ) ;
  assign n1097 = n256 | n858 ;
  assign n1096 = n256 &  n852 ;
  assign n1098 = ( n850 & ~n1097 ) | ( n850 & n1096 ) | ( ~n1097 & n1096 ) ;
  assign n1100 = n863 &  n883 ;
  assign n1099 = n861 | n883 ;
  assign n1101 = ( n1098 & ~n1100 ) | ( n1098 & n1099 ) | ( ~n1100 & n1099 ) ;
  assign n1163 = ( n1095 & ~n1107 ) | ( n1095 & n1101 ) | ( ~n1107 & n1101 ) ;
  assign n1164 = ( n1101 & ~n1095 ) | ( n1101 & n1107 ) | ( ~n1095 & n1107 ) ;
  assign n1165 = ( n1163 & ~n1101 ) | ( n1163 & n1164 ) | ( ~n1101 & n1164 ) ;
  assign n1296 = ( n1162 & ~n1246 ) | ( n1162 & n1165 ) | ( ~n1246 & n1165 ) ;
  assign n1297 = ( n1165 & ~n1162 ) | ( n1165 & n1246 ) | ( ~n1162 & n1246 ) ;
  assign n1298 = ( n1296 & ~n1165 ) | ( n1296 & n1297 ) | ( ~n1165 & n1297 ) ;
  assign n1112 = ( n789 & ~n998 ) | ( n789 & 1'b0 ) | ( ~n998 & 1'b0 ) ;
  assign n1113 = ~n796 & n998 ;
  assign n1114 = ( n1112 & ~n744 ) | ( n1112 & n1113 ) | ( ~n744 & n1113 ) ;
  assign n1116 = ( n793 & ~n801 ) | ( n793 & 1'b0 ) | ( ~n801 & 1'b0 ) ;
  assign n1115 = n793 | n799 ;
  assign n1117 = ( n1114 & ~n1116 ) | ( n1114 & n1115 ) | ( ~n1116 & n1115 ) ;
  assign n1149 = ( n1136 & ~n1142 ) | ( n1136 & n1148 ) | ( ~n1142 & n1148 ) ;
  assign n1150 = ( n1130 & ~n1117 ) | ( n1130 & n1149 ) | ( ~n1117 & n1149 ) ;
  assign n1294 = ( n1117 & ~n1149 ) | ( n1117 & n1130 ) | ( ~n1149 & n1130 ) ;
  assign n1295 = ( n1150 & ~n1130 ) | ( n1150 & n1294 ) | ( ~n1130 & n1294 ) ;
  assign n1329 = ( n1293 & ~n1298 ) | ( n1293 & n1295 ) | ( ~n1298 & n1295 ) ;
  assign n1330 = ( n1295 & ~n1293 ) | ( n1295 & n1298 ) | ( ~n1293 & n1298 ) ;
  assign n1331 = ( n1329 & ~n1295 ) | ( n1329 & n1330 ) | ( ~n1295 & n1330 ) ;
  assign n1323 = ( n1171 & ~n1226 ) | ( n1171 & n1245 ) | ( ~n1226 & n1245 ) ;
  assign n1324 = ( n1226 & ~n1246 ) | ( n1226 & n1323 ) | ( ~n1246 & n1323 ) ;
  assign n1302 = n883 | n1083 ;
  assign n1303 = n883 &  n994 ;
  assign n1304 = ( n1080 & ~n1302 ) | ( n1080 & n1303 ) | ( ~n1302 & n1303 ) ;
  assign n1305 = n856 &  n1126 ;
  assign n1306 = n856 | n1081 ;
  assign n1307 = ( n1304 & ~n1305 ) | ( n1304 & n1306 ) | ( ~n1305 & n1306 ) ;
  assign n1308 = ~n796 & n1175 ;
  assign n1309 = ( n789 & ~n1175 ) | ( n789 & 1'b0 ) | ( ~n1175 & 1'b0 ) ;
  assign n1310 = ( n1308 & ~n744 ) | ( n1308 & n1309 ) | ( ~n744 & n1309 ) ;
  assign n1311 = ~n799 & n1121 ;
  assign n1312 = n801 | n1121 ;
  assign n1313 = ( n1310 & ~n1311 ) | ( n1310 & n1312 ) | ( ~n1311 & n1312 ) ;
  assign n1314 = ~n1258 & n1260 ;
  assign n1315 = n1261 | n1314 ;
  assign n1316 = ( n1307 & n1313 ) | ( n1307 & n1315 ) | ( n1313 & n1315 ) ;
  assign n1317 = ( n1176 & ~n1219 ) | ( n1176 & n1225 ) | ( ~n1219 & n1225 ) ;
  assign n1318 = ( n1219 & ~n1226 ) | ( n1219 & n1317 ) | ( ~n1226 & n1317 ) ;
  assign n1320 = ( n1232 & n1238 ) | ( n1232 & n1244 ) | ( n1238 & n1244 ) ;
  assign n1319 = ( n1232 & ~n1238 ) | ( n1232 & n1244 ) | ( ~n1238 & n1244 ) ;
  assign n1321 = ( n1238 & ~n1320 ) | ( n1238 & n1319 ) | ( ~n1320 & n1319 ) ;
  assign n1322 = ( n1316 & ~n1318 ) | ( n1316 & n1321 ) | ( ~n1318 & n1321 ) ;
  assign n1325 = ( n1287 & n1289 ) | ( n1287 & n1292 ) | ( n1289 & n1292 ) ;
  assign n1326 = ( n1287 & ~n1289 ) | ( n1287 & n1292 ) | ( ~n1289 & n1292 ) ;
  assign n1327 = ( n1289 & ~n1325 ) | ( n1289 & n1326 ) | ( ~n1325 & n1326 ) ;
  assign n1328 = ( n1324 & ~n1322 ) | ( n1324 & n1327 ) | ( ~n1322 & n1327 ) ;
  assign n1340 = ~n248 & n520 ;
  assign n1341 = n248 &  n530 ;
  assign n1342 = n1340 | n1341 ;
  assign n1343 = n536 &  n712 ;
  assign n1344 = n543 | n712 ;
  assign n1345 = ( n1342 & ~n1343 ) | ( n1342 & n1344 ) | ( ~n1343 & n1344 ) ;
  assign n1333 = n883 &  n937 ;
  assign n1334 = n1217 &  n1333 ;
  assign n1332 = ( n856 & n937 ) | ( n856 & n1217 ) | ( n937 & n1217 ) ;
  assign n1335 = n856 | n937 ;
  assign n1336 = ( n1334 & ~n1332 ) | ( n1334 & n1335 ) | ( ~n1332 & n1335 ) ;
  assign n1337 = ( n592 & ~n663 ) | ( n592 & n1175 ) | ( ~n663 & n1175 ) ;
  assign n1338 = ( n708 & ~n1337 ) | ( n708 & 1'b0 ) | ( ~n1337 & 1'b0 ) ;
  assign n1339 = n1336 &  n1338 ;
  assign n1346 = n858 | n998 ;
  assign n1347 = n852 &  n998 ;
  assign n1348 = ( n850 & ~n1346 ) | ( n850 & n1347 ) | ( ~n1346 & n1347 ) ;
  assign n1350 = n793 &  n863 ;
  assign n1349 = n793 | n861 ;
  assign n1351 = ( n1348 & ~n1350 ) | ( n1348 & n1349 ) | ( ~n1350 & n1349 ) ;
  assign n1352 = ( n1345 & ~n1339 ) | ( n1345 & n1351 ) | ( ~n1339 & n1351 ) ;
  assign n1354 = n709 | n1121 ;
  assign n1353 = n715 &  n1121 ;
  assign n1355 = ( n666 & ~n1354 ) | ( n666 & n1353 ) | ( ~n1354 & n1353 ) ;
  assign n1357 = n720 &  n1077 ;
  assign n1356 = n718 | n1077 ;
  assign n1358 = ( n1355 & ~n1357 ) | ( n1355 & n1356 ) | ( ~n1357 & n1356 ) ;
  assign n1367 = ~n883 & n1126 ;
  assign n1364 = ( n256 & ~n1083 ) | ( n256 & 1'b0 ) | ( ~n1083 & 1'b0 ) ;
  assign n1365 = ~n256 & n994 ;
  assign n1366 = ( n1080 & n1364 ) | ( n1080 & n1365 ) | ( n1364 & n1365 ) ;
  assign n1368 = ( n883 & ~n1081 ) | ( n883 & 1'b0 ) | ( ~n1081 & 1'b0 ) ;
  assign n1369 = ( n1367 & ~n1366 ) | ( n1367 & n1368 ) | ( ~n1366 & n1368 ) ;
  assign n1359 = ( n937 & ~n524 ) | ( n937 & n1217 ) | ( ~n524 & n1217 ) ;
  assign n1360 = ~n856 & n937 ;
  assign n1361 = n1217 &  n1360 ;
  assign n1362 = ( n524 & ~n937 ) | ( n524 & 1'b0 ) | ( ~n937 & 1'b0 ) ;
  assign n1363 = ( n1359 & ~n1361 ) | ( n1359 & n1362 ) | ( ~n1361 & n1362 ) ;
  assign n1370 = ( n1358 & ~n1369 ) | ( n1358 & n1363 ) | ( ~n1369 & n1363 ) ;
  assign n1372 = ( n1273 & n1279 ) | ( n1273 & n1285 ) | ( n1279 & n1285 ) ;
  assign n1371 = ( n1273 & ~n1285 ) | ( n1273 & n1279 ) | ( ~n1285 & n1279 ) ;
  assign n1373 = ( n1285 & ~n1372 ) | ( n1285 & n1371 ) | ( ~n1372 & n1371 ) ;
  assign n1374 = ( n1352 & n1370 ) | ( n1352 & n1373 ) | ( n1370 & n1373 ) ;
  assign n1378 = ( n1316 & n1318 ) | ( n1316 & n1321 ) | ( n1318 & n1321 ) ;
  assign n1379 = ( n1318 & ~n1378 ) | ( n1318 & n1322 ) | ( ~n1378 & n1322 ) ;
  assign n1375 = ( n1261 & ~n1286 ) | ( n1261 & n1267 ) | ( ~n1286 & n1267 ) ;
  assign n1376 = ( n1267 & ~n1261 ) | ( n1267 & n1286 ) | ( ~n1261 & n1286 ) ;
  assign n1377 = ( n1375 & ~n1267 ) | ( n1375 & n1376 ) | ( ~n1267 & n1376 ) ;
  assign n1380 = ( n1374 & ~n1379 ) | ( n1374 & n1377 ) | ( ~n1379 & n1377 ) ;
  assign n1384 = n1374 | n1377 ;
  assign n1385 = n1374 &  n1377 ;
  assign n1386 = ( n1384 & ~n1385 ) | ( n1384 & 1'b0 ) | ( ~n1385 & 1'b0 ) ;
  assign n1387 = n1379 &  n1386 ;
  assign n1388 = n1379 | n1386 ;
  assign n1389 = ~n1387 & n1388 ;
  assign n1414 = ( n1313 & ~n1307 ) | ( n1313 & n1315 ) | ( ~n1307 & n1315 ) ;
  assign n1415 = ( n1307 & ~n1316 ) | ( n1307 & n1414 ) | ( ~n1316 & n1414 ) ;
  assign n1409 = ( n1339 & ~n1351 ) | ( n1339 & n1345 ) | ( ~n1351 & n1345 ) ;
  assign n1410 = ( n1352 & ~n1345 ) | ( n1352 & n1409 ) | ( ~n1345 & n1409 ) ;
  assign n1390 = n520 &  n793 ;
  assign n1391 = ( n530 & ~n793 ) | ( n530 & 1'b0 ) | ( ~n793 & 1'b0 ) ;
  assign n1392 = n1390 | n1391 ;
  assign n1393 = n248 &  n536 ;
  assign n1394 = n248 | n543 ;
  assign n1395 = ( n1392 & ~n1393 ) | ( n1392 & n1394 ) | ( ~n1393 & n1394 ) ;
  assign n1405 = ~n861 & n998 ;
  assign n1402 = ( n852 & ~n1077 ) | ( n852 & 1'b0 ) | ( ~n1077 & 1'b0 ) ;
  assign n1403 = ~n858 & n1077 ;
  assign n1404 = ( n850 & n1402 ) | ( n850 & n1403 ) | ( n1402 & n1403 ) ;
  assign n1406 = ( n863 & ~n998 ) | ( n863 & 1'b0 ) | ( ~n998 & 1'b0 ) ;
  assign n1407 = ( n1405 & ~n1404 ) | ( n1405 & n1406 ) | ( ~n1404 & n1406 ) ;
  assign n1396 = ( n712 & ~n1083 ) | ( n712 & 1'b0 ) | ( ~n1083 & 1'b0 ) ;
  assign n1397 = ~n712 & n994 ;
  assign n1398 = ( n1080 & n1396 ) | ( n1080 & n1397 ) | ( n1396 & n1397 ) ;
  assign n1399 = n256 &  n1126 ;
  assign n1400 = n256 | n1081 ;
  assign n1401 = ( n1398 & ~n1399 ) | ( n1398 & n1400 ) | ( ~n1399 & n1400 ) ;
  assign n1408 = ( n1395 & ~n1407 ) | ( n1395 & n1401 ) | ( ~n1407 & n1401 ) ;
  assign n1411 = ( n708 & ~n741 ) | ( n708 & 1'b0 ) | ( ~n741 & 1'b0 ) ;
  assign n1412 = ( n1259 & ~n708 ) | ( n1259 & n1411 ) | ( ~n708 & n1411 ) ;
  assign n1413 = ( n1410 & ~n1408 ) | ( n1410 & n1412 ) | ( ~n1408 & n1412 ) ;
  assign n1419 = ( n1352 & ~n1373 ) | ( n1352 & n1370 ) | ( ~n1373 & n1370 ) ;
  assign n1420 = ( n1373 & ~n1374 ) | ( n1373 & n1419 ) | ( ~n1374 & n1419 ) ;
  assign n1421 = ( n1415 & ~n1413 ) | ( n1415 & n1420 ) | ( ~n1413 & n1420 ) ;
  assign n1443 = ~n718 & n1121 ;
  assign n1441 = n709 | n1175 ;
  assign n1440 = n715 &  n1175 ;
  assign n1442 = ( n666 & ~n1441 ) | ( n666 & n1440 ) | ( ~n1441 & n1440 ) ;
  assign n1444 = ( n720 & ~n1121 ) | ( n720 & 1'b0 ) | ( ~n1121 & 1'b0 ) ;
  assign n1445 = ( n1443 & ~n1442 ) | ( n1443 & n1444 ) | ( ~n1442 & n1444 ) ;
  assign n1422 = ( n937 & ~n883 ) | ( n937 & n1217 ) | ( ~n883 & n1217 ) ;
  assign n1423 = ~n256 & n937 ;
  assign n1424 = n1217 &  n1423 ;
  assign n1425 = ( n883 & ~n937 ) | ( n883 & 1'b0 ) | ( ~n937 & 1'b0 ) ;
  assign n1426 = ( n1422 & ~n1424 ) | ( n1422 & n1425 ) | ( ~n1424 & n1425 ) ;
  assign n1436 = ( n536 & ~n793 ) | ( n536 & 1'b0 ) | ( ~n793 & 1'b0 ) ;
  assign n1433 = ( n520 & ~n998 ) | ( n520 & 1'b0 ) | ( ~n998 & 1'b0 ) ;
  assign n1434 = n530 &  n998 ;
  assign n1435 = n1433 | n1434 ;
  assign n1437 = ~n543 & n793 ;
  assign n1438 = ( n1436 & ~n1435 ) | ( n1436 & n1437 ) | ( ~n1435 & n1437 ) ;
  assign n1427 = ( n248 & ~n1083 ) | ( n248 & 1'b0 ) | ( ~n1083 & 1'b0 ) ;
  assign n1428 = ~n248 & n994 ;
  assign n1429 = ( n1080 & n1427 ) | ( n1080 & n1428 ) | ( n1427 & n1428 ) ;
  assign n1430 = n712 &  n1126 ;
  assign n1431 = n712 | n1081 ;
  assign n1432 = ( n1429 & ~n1430 ) | ( n1429 & n1431 ) | ( ~n1430 & n1431 ) ;
  assign n1439 = ( n1426 & ~n1438 ) | ( n1426 & n1432 ) | ( ~n1438 & n1432 ) ;
  assign n1446 = n1336 | n1338 ;
  assign n1447 = ~n1339 & n1446 ;
  assign n1448 = ( n1445 & ~n1439 ) | ( n1445 & n1447 ) | ( ~n1439 & n1447 ) ;
  assign n1452 = ( n1408 & n1410 ) | ( n1408 & n1412 ) | ( n1410 & n1412 ) ;
  assign n1453 = ( n1408 & ~n1452 ) | ( n1408 & n1413 ) | ( ~n1452 & n1413 ) ;
  assign n1416 = n1363 | n1369 ;
  assign n1417 = n1363 &  n1369 ;
  assign n1418 = ( n1416 & ~n1417 ) | ( n1416 & 1'b0 ) | ( ~n1417 & 1'b0 ) ;
  assign n1449 = ( n1358 & ~n1418 ) | ( n1358 & 1'b0 ) | ( ~n1418 & 1'b0 ) ;
  assign n1450 = ~n1358 & n1418 ;
  assign n1451 = n1449 | n1450 ;
  assign n1454 = ( n1448 & ~n1453 ) | ( n1448 & n1451 ) | ( ~n1453 & n1451 ) ;
  assign n1467 = n793 | n1083 ;
  assign n1468 = n793 &  n994 ;
  assign n1469 = ( n1080 & ~n1467 ) | ( n1080 & n1468 ) | ( ~n1467 & n1468 ) ;
  assign n1470 = n248 &  n1126 ;
  assign n1471 = n248 | n1081 ;
  assign n1472 = ( n1469 & ~n1470 ) | ( n1469 & n1471 ) | ( ~n1470 & n1471 ) ;
  assign n1464 = ~n861 & n1121 ;
  assign n1462 = n858 | n1175 ;
  assign n1461 = n852 &  n1175 ;
  assign n1463 = ( n850 & ~n1462 ) | ( n850 & n1461 ) | ( ~n1462 & n1461 ) ;
  assign n1465 = ( n863 & ~n1121 ) | ( n863 & 1'b0 ) | ( ~n1121 & 1'b0 ) ;
  assign n1466 = ( n1464 & ~n1463 ) | ( n1464 & n1465 ) | ( ~n1463 & n1465 ) ;
  assign n1473 = n520 &  n1077 ;
  assign n1474 = ( n530 & ~n1077 ) | ( n530 & 1'b0 ) | ( ~n1077 & 1'b0 ) ;
  assign n1475 = n1473 | n1474 ;
  assign n1476 = n536 &  n998 ;
  assign n1477 = n543 | n998 ;
  assign n1478 = ( n1475 & ~n1476 ) | ( n1475 & n1477 ) | ( ~n1476 & n1477 ) ;
  assign n1479 = ( n1472 & ~n1466 ) | ( n1472 & n1478 ) | ( ~n1466 & n1478 ) ;
  assign n1481 = ( n1426 & n1432 ) | ( n1426 & n1438 ) | ( n1432 & n1438 ) ;
  assign n1480 = ( n1426 & ~n1432 ) | ( n1426 & n1438 ) | ( ~n1432 & n1438 ) ;
  assign n1482 = ( n1432 & ~n1481 ) | ( n1432 & n1480 ) | ( ~n1481 & n1480 ) ;
  assign n1483 = ~n666 & n1175 ;
  assign n1493 = n858 | n1121 ;
  assign n1492 = n852 &  n1121 ;
  assign n1494 = ( n850 & ~n1493 ) | ( n850 & n1492 ) | ( ~n1493 & n1492 ) ;
  assign n1496 = n863 &  n1077 ;
  assign n1495 = n861 | n1077 ;
  assign n1497 = ( n1494 & ~n1496 ) | ( n1494 & n1495 ) | ( ~n1496 & n1495 ) ;
  assign n1485 = ~n712 & n937 ;
  assign n1486 = n1217 &  n1485 ;
  assign n1484 = ( n256 & n937 ) | ( n256 & n1217 ) | ( n937 & n1217 ) ;
  assign n1487 = n256 | n937 ;
  assign n1488 = ( n1486 & ~n1484 ) | ( n1486 & n1487 ) | ( ~n1484 & n1487 ) ;
  assign n1489 = ( n847 & ~n433 ) | ( n847 & n1175 ) | ( ~n433 & n1175 ) ;
  assign n1490 = ( n592 & ~n1489 ) | ( n592 & 1'b0 ) | ( ~n1489 & 1'b0 ) ;
  assign n1491 = n1488 &  n1490 ;
  assign n1498 = ( n1483 & ~n1497 ) | ( n1483 & n1491 ) | ( ~n1497 & n1491 ) ;
  assign n1499 = ( n1483 & ~n1491 ) | ( n1483 & n1497 ) | ( ~n1491 & n1497 ) ;
  assign n1500 = ( n1498 & ~n1483 ) | ( n1498 & n1499 ) | ( ~n1483 & n1499 ) ;
  assign n1501 = ( n1479 & ~n1482 ) | ( n1479 & n1500 ) | ( ~n1482 & n1500 ) ;
  assign n1514 = n793 &  n937 ;
  assign n1515 = n1217 &  n1514 ;
  assign n1513 = ( n248 & n937 ) | ( n248 & n1217 ) | ( n937 & n1217 ) ;
  assign n1516 = n248 | n937 ;
  assign n1517 = ( n1515 & ~n1513 ) | ( n1515 & n1516 ) | ( ~n1513 & n1516 ) ;
  assign n1518 = ( n526 & ~n515 ) | ( n526 & n1175 ) | ( ~n515 & n1175 ) ;
  assign n1519 = n433 | n1518 ;
  assign n1520 = ( n1517 & ~n1519 ) | ( n1517 & 1'b0 ) | ( ~n1519 & 1'b0 ) ;
  assign n1521 = n1077 | n1083 ;
  assign n1522 = n994 &  n1077 ;
  assign n1523 = ( n1080 & ~n1521 ) | ( n1080 & n1522 ) | ( ~n1521 & n1522 ) ;
  assign n1524 = n998 &  n1126 ;
  assign n1525 = n998 | n1081 ;
  assign n1526 = ( n1523 & ~n1524 ) | ( n1523 & n1525 ) | ( ~n1524 & n1525 ) ;
  assign n1527 = ( n520 & ~n1175 ) | ( n520 & 1'b0 ) | ( ~n1175 & 1'b0 ) ;
  assign n1528 = n530 &  n1175 ;
  assign n1529 = n1527 | n1528 ;
  assign n1530 = n536 &  n1121 ;
  assign n1531 = n543 | n1121 ;
  assign n1532 = ( n1529 & ~n1530 ) | ( n1529 & n1531 ) | ( ~n1530 & n1531 ) ;
  assign n1533 = ~n1517 & n1519 ;
  assign n1534 = n1520 | n1533 ;
  assign n1535 = ( n1526 & n1532 ) | ( n1526 & n1534 ) | ( n1532 & n1534 ) ;
  assign n1536 = ( n433 & ~n849 ) | ( n433 & n1489 ) | ( ~n849 & n1489 ) ;
  assign n1537 = ( n1520 & ~n1535 ) | ( n1520 & n1536 ) | ( ~n1535 & n1536 ) ;
  assign n1539 = n937 | n998 ;
  assign n1542 = ( n937 & n998 ) | ( n937 & n1217 ) | ( n998 & n1217 ) ;
  assign n1540 = n937 &  n1077 ;
  assign n1541 = n1217 &  n1540 ;
  assign n1543 = ( n1539 & ~n1542 ) | ( n1539 & n1541 ) | ( ~n1542 & n1541 ) ;
  assign n1544 = ( n937 & ~n992 ) | ( n937 & n1175 ) | ( ~n992 & n1175 ) ;
  assign n1545 = n515 | n1544 ;
  assign n1546 = ( n1543 & ~n1545 ) | ( n1543 & 1'b0 ) | ( ~n1545 & 1'b0 ) ;
  assign n1555 = ~n1077 & n1126 ;
  assign n1552 = ~n1083 & n1121 ;
  assign n1553 = ( n994 & ~n1121 ) | ( n994 & 1'b0 ) | ( ~n1121 & 1'b0 ) ;
  assign n1554 = ( n1080 & n1552 ) | ( n1080 & n1553 ) | ( n1552 & n1553 ) ;
  assign n1556 = ( n1077 & ~n1081 ) | ( n1077 & 1'b0 ) | ( ~n1081 & 1'b0 ) ;
  assign n1557 = ( n1555 & ~n1554 ) | ( n1555 & n1556 ) | ( ~n1554 & n1556 ) ;
  assign n1547 = ( n937 & ~n793 ) | ( n937 & n1217 ) | ( ~n793 & n1217 ) ;
  assign n1548 = n793 | n1547 ;
  assign n1549 = n998 | n1217 ;
  assign n1550 = ( n998 & ~n1549 ) | ( n998 & n1547 ) | ( ~n1549 & n1547 ) ;
  assign n1551 = ( n1548 & ~n937 ) | ( n1548 & n1550 ) | ( ~n937 & n1550 ) ;
  assign n1558 = ( n1546 & ~n1557 ) | ( n1546 & n1551 ) | ( ~n1557 & n1551 ) ;
  assign n1559 = ( n1551 & ~n1546 ) | ( n1551 & n1557 ) | ( ~n1546 & n1557 ) ;
  assign n1560 = ( n1558 & ~n1551 ) | ( n1558 & n1559 ) | ( ~n1551 & n1559 ) ;
  assign n1538 = ~n534 & n1175 ;
  assign n1570 = ( n515 & ~n1544 ) | ( n515 & 1'b0 ) | ( ~n1544 & 1'b0 ) ;
  assign n1571 = ( n937 & ~n1079 ) | ( n937 & n1570 ) | ( ~n1079 & n1570 ) ;
  assign n1561 = ( n937 & ~n1217 ) | ( n937 & n1077 ) | ( ~n1217 & n1077 ) ;
  assign n1562 = n937 &  n1121 ;
  assign n1563 = ( n1217 & ~n937 ) | ( n1217 & n1562 ) | ( ~n937 & n1562 ) ;
  assign n1564 = ( n1561 & ~n1540 ) | ( n1561 & n1563 ) | ( ~n1540 & n1563 ) ;
  assign n1565 = ( n1121 & ~n1217 ) | ( n1121 & 1'b0 ) | ( ~n1217 & 1'b0 ) ;
  assign n1566 = ( n937 & ~n1175 ) | ( n937 & 1'b0 ) | ( ~n1175 & 1'b0 ) ;
  assign n1567 = ~n1565 & n1566 ;
  assign n1568 = n1564 | n1567 ;
  assign n1569 = ( n1545 & ~n1568 ) | ( n1545 & n1567 ) | ( ~n1568 & n1567 ) ;
  assign n1576 = n1571 &  n1569 ;
  assign n1572 = ~n1564 & n1567 ;
  assign n1573 = ~n1543 & n1545 ;
  assign n1574 = n1546 | n1573 ;
  assign n1575 = ~n1572 & n1574 ;
  assign n1577 = ( n1576 & ~n1569 ) | ( n1576 & n1575 ) | ( ~n1569 & n1575 ) ;
  assign n1580 = ~n1084 & n1175 ;
  assign n1578 = n994 &  n1080 ;
  assign n1579 = n1175 | n1578 ;
  assign n1581 = ( n1577 & ~n1580 ) | ( n1577 & n1579 ) | ( ~n1580 & n1579 ) ;
  assign n1582 = n1121 &  n1126 ;
  assign n1583 = n1081 | n1121 ;
  assign n1584 = ( n1581 & ~n1582 ) | ( n1581 & n1583 ) | ( ~n1582 & n1583 ) ;
  assign n1585 = ( n1545 & ~n1571 ) | ( n1545 & 1'b0 ) | ( ~n1571 & 1'b0 ) ;
  assign n1586 = ( n1567 & ~n1564 ) | ( n1567 & n1585 ) | ( ~n1564 & n1585 ) ;
  assign n1587 = ~n1574 & n1586 ;
  assign n1588 = ( n1584 & ~n1587 ) | ( n1584 & 1'b0 ) | ( ~n1587 & 1'b0 ) ;
  assign n1589 = ( n1560 & ~n1538 ) | ( n1560 & n1588 ) | ( ~n1538 & n1588 ) ;
  assign n1592 = ( n1546 & ~n1551 ) | ( n1546 & n1557 ) | ( ~n1551 & n1557 ) ;
  assign n1590 = ( n1532 & ~n1526 ) | ( n1532 & n1534 ) | ( ~n1526 & n1534 ) ;
  assign n1591 = ( n1526 & ~n1535 ) | ( n1526 & n1590 ) | ( ~n1535 & n1590 ) ;
  assign n1593 = ( n1589 & ~n1592 ) | ( n1589 & n1591 ) | ( ~n1592 & n1591 ) ;
  assign n1601 = ~n248 & n937 ;
  assign n1602 = n1217 &  n1601 ;
  assign n1600 = ( n712 & n937 ) | ( n712 & n1217 ) | ( n937 & n1217 ) ;
  assign n1603 = n712 | n937 ;
  assign n1604 = ( n1602 & ~n1600 ) | ( n1602 & n1603 ) | ( ~n1600 & n1603 ) ;
  assign n1597 = ~n793 & n1126 ;
  assign n1594 = ( n998 & ~n1083 ) | ( n998 & 1'b0 ) | ( ~n1083 & 1'b0 ) ;
  assign n1595 = ( n994 & ~n998 ) | ( n994 & 1'b0 ) | ( ~n998 & 1'b0 ) ;
  assign n1596 = ( n1080 & n1594 ) | ( n1080 & n1595 ) | ( n1594 & n1595 ) ;
  assign n1598 = ( n793 & ~n1081 ) | ( n793 & 1'b0 ) | ( ~n1081 & 1'b0 ) ;
  assign n1599 = ( n1597 & ~n1596 ) | ( n1597 & n1598 ) | ( ~n1596 & n1598 ) ;
  assign n1608 = ( n536 & ~n1077 ) | ( n536 & 1'b0 ) | ( ~n1077 & 1'b0 ) ;
  assign n1605 = ( n520 & ~n1121 ) | ( n520 & 1'b0 ) | ( ~n1121 & 1'b0 ) ;
  assign n1606 = n530 &  n1121 ;
  assign n1607 = n1605 | n1606 ;
  assign n1609 = ~n543 & n1077 ;
  assign n1610 = ( n1608 & ~n1607 ) | ( n1608 & n1609 ) | ( ~n1607 & n1609 ) ;
  assign n1611 = ( n1604 & ~n1599 ) | ( n1604 & n1610 ) | ( ~n1599 & n1610 ) ;
  assign n1612 = ( n1599 & ~n1610 ) | ( n1599 & n1604 ) | ( ~n1610 & n1604 ) ;
  assign n1613 = ( n1611 & ~n1604 ) | ( n1611 & n1612 ) | ( ~n1604 & n1612 ) ;
  assign n1614 = ( n1520 & n1535 ) | ( n1520 & n1536 ) | ( n1535 & n1536 ) ;
  assign n1615 = ( n1535 & ~n1520 ) | ( n1535 & n1536 ) | ( ~n1520 & n1536 ) ;
  assign n1616 = ( n1520 & ~n1614 ) | ( n1520 & n1615 ) | ( ~n1614 & n1615 ) ;
  assign n1617 = ( n1593 & ~n1613 ) | ( n1593 & n1616 ) | ( ~n1613 & n1616 ) ;
  assign n1624 = n1472 &  n1478 ;
  assign n1625 = ~n1472 & n1478 ;
  assign n1626 = ( n1472 & ~n1624 ) | ( n1472 & n1625 ) | ( ~n1624 & n1625 ) ;
  assign n1618 = n1488 | n1490 ;
  assign n1619 = ~n1491 & n1618 ;
  assign n1620 = ( n1599 & n1604 ) | ( n1599 & n1610 ) | ( n1604 & n1610 ) ;
  assign n1621 = n1619 &  n1620 ;
  assign n1622 = n1619 | n1620 ;
  assign n1623 = ~n1621 & n1622 ;
  assign n1627 = ( n1466 & ~n1626 ) | ( n1466 & n1623 ) | ( ~n1626 & n1623 ) ;
  assign n1628 = ( n1466 & ~n1623 ) | ( n1466 & n1626 ) | ( ~n1623 & n1626 ) ;
  assign n1629 = ( n1627 & ~n1466 ) | ( n1627 & n1628 ) | ( ~n1466 & n1628 ) ;
  assign n1630 = ( n1537 & ~n1617 ) | ( n1537 & n1629 ) | ( ~n1617 & n1629 ) ;
  assign n1631 = n1466 &  n1626 ;
  assign n1632 = ( n1466 & n1622 ) | ( n1466 & n1626 ) | ( n1622 & n1626 ) ;
  assign n1633 = ( n1621 & ~n1631 ) | ( n1621 & n1632 ) | ( ~n1631 & n1632 ) ;
  assign n1635 = ( n1479 & n1482 ) | ( n1479 & n1500 ) | ( n1482 & n1500 ) ;
  assign n1634 = ( n1479 & ~n1500 ) | ( n1479 & n1482 ) | ( ~n1500 & n1482 ) ;
  assign n1636 = ( n1500 & ~n1635 ) | ( n1500 & n1634 ) | ( ~n1635 & n1634 ) ;
  assign n1637 = ( n1630 & n1633 ) | ( n1630 & n1636 ) | ( n1633 & n1636 ) ;
  assign n1502 = ( n1439 & n1445 ) | ( n1439 & n1447 ) | ( n1445 & n1447 ) ;
  assign n1503 = ( n1439 & ~n1502 ) | ( n1439 & n1448 ) | ( ~n1502 & n1448 ) ;
  assign n1504 = n1395 &  n1401 ;
  assign n1505 = ( n1395 & ~n1401 ) | ( n1395 & 1'b0 ) | ( ~n1401 & 1'b0 ) ;
  assign n1506 = ( n1401 & ~n1504 ) | ( n1401 & n1505 ) | ( ~n1504 & n1505 ) ;
  assign n1507 = ( n1407 & n1498 ) | ( n1407 & n1506 ) | ( n1498 & n1506 ) ;
  assign n1508 = ( n1407 & ~n1506 ) | ( n1407 & n1498 ) | ( ~n1506 & n1498 ) ;
  assign n1509 = ( n1506 & ~n1507 ) | ( n1506 & n1508 ) | ( ~n1507 & n1508 ) ;
  assign n1510 = n1503 &  n1509 ;
  assign n1511 = n1503 | n1509 ;
  assign n1512 = ~n1510 & n1511 ;
  assign n1638 = ( n1501 & ~n1637 ) | ( n1501 & n1512 ) | ( ~n1637 & n1512 ) ;
  assign n1640 = ( n1395 & n1401 ) | ( n1395 & n1407 ) | ( n1401 & n1407 ) ;
  assign n1639 = ( n1395 & ~n1401 ) | ( n1395 & n1407 ) | ( ~n1401 & n1407 ) ;
  assign n1641 = ( n1401 & ~n1640 ) | ( n1401 & n1639 ) | ( ~n1640 & n1639 ) ;
  assign n1642 = ( n1498 & ~n1503 ) | ( n1498 & n1641 ) | ( ~n1503 & n1641 ) ;
  assign n1643 = n1358 &  n1418 ;
  assign n1644 = ( n1418 & ~n1643 ) | ( n1418 & n1449 ) | ( ~n1643 & n1449 ) ;
  assign n1645 = ( n1448 & n1453 ) | ( n1448 & n1644 ) | ( n1453 & n1644 ) ;
  assign n1646 = ( n1448 & ~n1644 ) | ( n1448 & n1453 ) | ( ~n1644 & n1453 ) ;
  assign n1647 = ( n1644 & ~n1645 ) | ( n1644 & n1646 ) | ( ~n1645 & n1646 ) ;
  assign n1648 = ( n1638 & ~n1642 ) | ( n1638 & n1647 ) | ( ~n1642 & n1647 ) ;
  assign n1455 = n1413 &  n1415 ;
  assign n1456 = n1413 | n1415 ;
  assign n1457 = ~n1455 & n1456 ;
  assign n1458 = ~n1420 & n1457 ;
  assign n1459 = ( n1420 & ~n1457 ) | ( n1420 & 1'b0 ) | ( ~n1457 & 1'b0 ) ;
  assign n1460 = n1458 | n1459 ;
  assign n1649 = ( n1454 & ~n1648 ) | ( n1454 & n1460 ) | ( ~n1648 & n1460 ) ;
  assign n1650 = ( n1389 & ~n1421 ) | ( n1389 & n1649 ) | ( ~n1421 & n1649 ) ;
  assign n1381 = ( n1322 & n1324 ) | ( n1322 & n1327 ) | ( n1324 & n1327 ) ;
  assign n1382 = ( n1322 & ~n1324 ) | ( n1322 & n1327 ) | ( ~n1324 & n1327 ) ;
  assign n1383 = ( n1324 & ~n1381 ) | ( n1324 & n1382 ) | ( ~n1381 & n1382 ) ;
  assign n1651 = ( n1380 & ~n1650 ) | ( n1380 & n1383 ) | ( ~n1650 & n1383 ) ;
  assign n1652 = ( n1331 & ~n1328 ) | ( n1331 & n1651 ) | ( ~n1328 & n1651 ) ;
  assign n1829 = ( n1328 & ~n1651 ) | ( n1328 & n1331 ) | ( ~n1651 & n1331 ) ;
  assign n1830 = ( n1652 & ~n1331 ) | ( n1652 & n1829 ) | ( ~n1331 & n1829 ) ;
  assign n1858 = ( n1383 & ~n1380 ) | ( n1383 & n1650 ) | ( ~n1380 & n1650 ) ;
  assign n1859 = ( n1380 & ~n1383 ) | ( n1380 & n1650 ) | ( ~n1383 & n1650 ) ;
  assign n1860 = ( n1858 & ~n1650 ) | ( n1858 & n1859 ) | ( ~n1650 & n1859 ) ;
  assign n1831 = ~n125 & n100 ;
  assign n1832 = ( n100 & ~n1831 ) | ( n100 & n924 ) | ( ~n1831 & n924 ) ;
  assign n1833 = ( n555 & ~n317 ) | ( n555 & n1832 ) | ( ~n317 & n1832 ) ;
  assign n1834 = n317 | n1833 ;
  assign n1835 = n443 | n478 ;
  assign n1836 = ( n318 & ~n595 ) | ( n318 & n1835 ) | ( ~n595 & n1835 ) ;
  assign n1837 = n595 | n1836 ;
  assign n1838 = n108 | n1837 ;
  assign n1839 = ( n1834 & ~n610 ) | ( n1834 & n1838 ) | ( ~n610 & n1838 ) ;
  assign n1840 = n610 | n1839 ;
  assign n1841 = ( n647 & ~n290 ) | ( n647 & n1840 ) | ( ~n290 & n1840 ) ;
  assign n1842 = n290 | n1841 ;
  assign n1843 = n48 | n112 ;
  assign n1844 = ( n1842 & ~n48 ) | ( n1842 & n1843 ) | ( ~n48 & n1843 ) ;
  assign n1694 = n401 | n453 ;
  assign n1695 = ( n475 & ~n143 ) | ( n475 & n1694 ) | ( ~n143 & n1694 ) ;
  assign n1696 = n143 | n1695 ;
  assign n1697 = ( n612 & ~n85 ) | ( n612 & n1696 ) | ( ~n85 & n1696 ) ;
  assign n1698 = n85 | n1697 ;
  assign n1699 = n281 | n1698 ;
  assign n1845 = n228 | n1804 ;
  assign n1846 = ( n1699 & ~n692 ) | ( n1699 & n1845 ) | ( ~n692 & n1845 ) ;
  assign n1847 = n692 | n1846 ;
  assign n1848 = ( n1844 & ~n809 ) | ( n1844 & n1847 ) | ( ~n809 & n1847 ) ;
  assign n1849 = n809 | n1848 ;
  assign n1850 = ( n310 & ~n182 ) | ( n310 & n1849 ) | ( ~n182 & n1849 ) ;
  assign n1851 = n182 | n1850 ;
  assign n1852 = ( n488 & ~n110 ) | ( n488 & n1851 ) | ( ~n110 & n1851 ) ;
  assign n1853 = n110 | n1852 ;
  assign n1854 = ( n198 & ~n97 ) | ( n198 & n1853 ) | ( ~n97 & n1853 ) ;
  assign n1855 = n97 | n1854 ;
  assign n1856 = n289 | n1855 ;
  assign n1857 = n316 | n1856 ;
  assign n1861 = ( n1379 & n1386 ) | ( n1379 & n1421 ) | ( n1386 & n1421 ) ;
  assign n1862 = ( n1379 & ~n1386 ) | ( n1379 & n1421 ) | ( ~n1386 & n1421 ) ;
  assign n1863 = ( n1386 & ~n1861 ) | ( n1386 & n1862 ) | ( ~n1861 & n1862 ) ;
  assign n1864 = ~n381 & n627 ;
  assign n1865 = ( n353 & ~n266 ) | ( n353 & n1864 ) | ( ~n266 & n1864 ) ;
  assign n1866 = ~n353 & n1865 ;
  assign n1867 = n279 | n595 ;
  assign n1868 = n116 | n1867 ;
  assign n1869 = ( n556 & ~n360 ) | ( n556 & n1868 ) | ( ~n360 & n1868 ) ;
  assign n1870 = n360 | n1869 ;
  assign n1871 = ( n890 & n1866 ) | ( n890 & n1870 ) | ( n1866 & n1870 ) ;
  assign n1872 = ( n334 & ~n1871 ) | ( n334 & n1866 ) | ( ~n1871 & n1866 ) ;
  assign n1873 = ~n334 & n1872 ;
  assign n1874 = ( n128 & ~n399 ) | ( n128 & n1873 ) | ( ~n399 & n1873 ) ;
  assign n1875 = ~n128 & n1874 ;
  assign n1876 = n424 | n894 ;
  assign n1877 = ( n457 & ~n1876 ) | ( n457 & n600 ) | ( ~n1876 & n600 ) ;
  assign n1878 = ~n600 & n1877 ;
  assign n1879 = ( n358 & ~n1769 ) | ( n358 & n1878 ) | ( ~n1769 & n1878 ) ;
  assign n1880 = ~n358 & n1879 ;
  assign n1881 = ( n323 & n1875 ) | ( n323 & n1880 ) | ( n1875 & n1880 ) ;
  assign n1882 = ~n323 & n1881 ;
  assign n1883 = ( n488 & ~n723 ) | ( n488 & n1882 ) | ( ~n723 & n1882 ) ;
  assign n1884 = ~n488 & n1883 ;
  assign n1885 = ~n164 & n1884 ;
  assign n1886 = ( n1649 & ~n1863 ) | ( n1649 & n1885 ) | ( ~n1863 & n1885 ) ;
  assign n1887 = ( n597 & ~n1863 ) | ( n597 & n1649 ) | ( ~n1863 & n1649 ) ;
  assign n1888 = ( n1886 & ~n1887 ) | ( n1886 & 1'b0 ) | ( ~n1887 & 1'b0 ) ;
  assign n1889 = ( n1860 & ~n1857 ) | ( n1860 & n1888 ) | ( ~n1857 & n1888 ) ;
  assign n1890 = ( n1828 & n1830 ) | ( n1828 & n1889 ) | ( n1830 & n1889 ) ;
  assign n999 = ~n788 & n998 ;
  assign n1071 = ( n937 & ~n999 ) | ( n937 & n994 ) | ( ~n999 & n994 ) ;
  assign n1072 = ( n937 & ~n994 ) | ( n937 & n999 ) | ( ~n994 & n999 ) ;
  assign n1073 = ( n1071 & ~n937 ) | ( n1071 & n1072 ) | ( ~n937 & n1072 ) ;
  assign n1068 = ( n856 & ~n861 ) | ( n856 & 1'b0 ) | ( ~n861 & 1'b0 ) ;
  assign n1065 = ( n852 & ~n883 ) | ( n852 & 1'b0 ) | ( ~n883 & 1'b0 ) ;
  assign n1066 = ~n858 & n883 ;
  assign n1067 = ( n850 & n1065 ) | ( n850 & n1066 ) | ( n1065 & n1066 ) ;
  assign n1069 = ~n856 & n863 ;
  assign n1070 = ( n1068 & ~n1067 ) | ( n1068 & n1069 ) | ( ~n1067 & n1069 ) ;
  assign n1089 = ( n1073 & ~n1070 ) | ( n1073 & n1088 ) | ( ~n1070 & n1088 ) ;
  assign n1248 = ( n1070 & ~n1088 ) | ( n1070 & n1073 ) | ( ~n1088 & n1073 ) ;
  assign n1249 = ( n1089 & ~n1073 ) | ( n1089 & n1248 ) | ( ~n1073 & n1248 ) ;
  assign n1247 = ( n1162 & ~n1165 ) | ( n1162 & n1246 ) | ( ~n1165 & n1246 ) ;
  assign n1790 = n1247 &  n1249 ;
  assign n1789 = ( n1247 & ~n1249 ) | ( n1247 & 1'b0 ) | ( ~n1249 & 1'b0 ) ;
  assign n1791 = ( n1249 & ~n1790 ) | ( n1249 & n1789 ) | ( ~n1790 & n1789 ) ;
  assign n719 = ( n256 & ~n718 ) | ( n256 & 1'b0 ) | ( ~n718 & 1'b0 ) ;
  assign n713 = n709 | n712 ;
  assign n716 = n712 &  n715 ;
  assign n717 = ( n666 & ~n713 ) | ( n666 & n716 ) | ( ~n713 & n716 ) ;
  assign n721 = ~n256 & n720 ;
  assign n722 = ( n719 & ~n717 ) | ( n719 & n721 ) | ( ~n717 & n721 ) ;
  assign n525 = ~n520 & n524 ;
  assign n531 = n524 | n530 ;
  assign n532 = ~n525 & n531 ;
  assign n541 = n536 &  n540 ;
  assign n544 = n540 | n543 ;
  assign n545 = ( n532 & ~n541 ) | ( n532 & n544 ) | ( ~n541 & n544 ) ;
  assign n794 = n789 &  n793 ;
  assign n797 = n793 | n796 ;
  assign n798 = ( n744 & ~n794 ) | ( n744 & n797 ) | ( ~n794 & n797 ) ;
  assign n802 = n248 | n801 ;
  assign n800 = ( n248 & ~n799 ) | ( n248 & 1'b0 ) | ( ~n799 & 1'b0 ) ;
  assign n803 = ( n798 & ~n802 ) | ( n798 & n800 ) | ( ~n802 & n800 ) ;
  assign n1109 = ( n545 & n722 ) | ( n545 & n803 ) | ( n722 & n803 ) ;
  assign n1110 = ( n545 & ~n722 ) | ( n545 & n803 ) | ( ~n722 & n803 ) ;
  assign n1111 = ( n722 & ~n1109 ) | ( n722 & n1110 ) | ( ~n1109 & n1110 ) ;
  assign n1108 = ( n1095 & ~n1101 ) | ( n1095 & n1107 ) | ( ~n1101 & n1107 ) ;
  assign n1250 = ( n1111 & ~n1108 ) | ( n1111 & n1150 ) | ( ~n1108 & n1150 ) ;
  assign n1251 = ( n1108 & ~n1150 ) | ( n1108 & n1111 ) | ( ~n1150 & n1111 ) ;
  assign n1252 = ( n1250 & ~n1111 ) | ( n1250 & n1251 ) | ( ~n1111 & n1251 ) ;
  assign n1299 = ( n1293 & n1295 ) | ( n1293 & n1298 ) | ( n1295 & n1298 ) ;
  assign n1792 = ( n1252 & n1299 ) | ( n1252 & n1791 ) | ( n1299 & n1791 ) ;
  assign n1793 = ( n1252 & ~n1791 ) | ( n1252 & n1299 ) | ( ~n1791 & n1299 ) ;
  assign n1794 = ( n1791 & ~n1792 ) | ( n1791 & n1793 ) | ( ~n1792 & n1793 ) ;
  assign n1795 = ~n1652 & n1794 ;
  assign n1796 = ( n1652 & ~n1794 ) | ( n1652 & 1'b0 ) | ( ~n1794 & 1'b0 ) ;
  assign n1797 = n1795 | n1796 ;
  assign n1891 = ( n1788 & ~n1890 ) | ( n1788 & n1797 ) | ( ~n1890 & n1797 ) ;
  assign n1718 = ( n323 & ~n412 ) | ( n323 & n443 ) | ( ~n412 & n443 ) ;
  assign n1719 = ( n412 & ~n115 ) | ( n412 & n1718 ) | ( ~n115 & n1718 ) ;
  assign n1720 = n115 | n1719 ;
  assign n1721 = ( n554 & ~n198 ) | ( n554 & n1720 ) | ( ~n198 & n1720 ) ;
  assign n1722 = n198 | n1721 ;
  assign n1723 = n209 | n1722 ;
  assign n1666 = n103 | n278 ;
  assign n1724 = ( n318 & ~n261 ) | ( n318 & n1666 ) | ( ~n261 & n1666 ) ;
  assign n1725 = n261 | n1724 ;
  assign n1726 = ( n600 & ~n979 ) | ( n600 & n1725 ) | ( ~n979 & n1725 ) ;
  assign n1727 = n979 | n1726 ;
  assign n1728 = ( n549 & ~n149 ) | ( n549 & n1727 ) | ( ~n149 & n1727 ) ;
  assign n1729 = n149 | n1728 ;
  assign n1730 = ( n120 & ~n109 ) | ( n120 & n1729 ) | ( ~n109 & n1729 ) ;
  assign n1731 = n109 | n1730 ;
  assign n1732 = n197 | n1731 ;
  assign n1733 = n130 | n1732 ;
  assign n1734 = n291 | n1733 ;
  assign n1735 = n227 | n330 ;
  assign n1736 = n555 | n1735 ;
  assign n1737 = n167 | n211 ;
  assign n1738 = ( n1736 & ~n442 ) | ( n1736 & n1737 ) | ( ~n442 & n1737 ) ;
  assign n1739 = n442 | n1738 ;
  assign n1740 = ( n276 & ~n162 ) | ( n276 & n1739 ) | ( ~n162 & n1739 ) ;
  assign n1741 = n162 | n1740 ;
  assign n1742 = ( n265 & ~n148 ) | ( n265 & n1741 ) | ( ~n148 & n1741 ) ;
  assign n1743 = ( n362 & ~n165 ) | ( n362 & n1742 ) | ( ~n165 & n1742 ) ;
  assign n1744 = n165 | n1743 ;
  assign n1745 = ( n667 & ~n399 ) | ( n667 & n1744 ) | ( ~n399 & n1744 ) ;
  assign n1746 = ( n399 & ~n1734 ) | ( n399 & n1745 ) | ( ~n1734 & n1745 ) ;
  assign n1747 = n1734 | n1746 ;
  assign n1748 = ( n1723 & ~n169 ) | ( n1723 & n1747 ) | ( ~n169 & n1747 ) ;
  assign n1749 = n169 | n1748 ;
  assign n1750 = ( n324 & ~n195 ) | ( n324 & n1749 ) | ( ~n195 & n1749 ) ;
  assign n1751 = n195 | n1750 ;
  assign n1752 = ( n317 & ~n141 ) | ( n317 & n1751 ) | ( ~n141 & n1751 ) ;
  assign n1753 = n141 | n1752 ;
  assign n1754 = n402 | n1753 ;
  assign n1253 = ( n1247 & ~n1252 ) | ( n1247 & n1249 ) | ( ~n1252 & n1249 ) ;
  assign n1300 = ( n1249 & ~n1247 ) | ( n1249 & n1252 ) | ( ~n1247 & n1252 ) ;
  assign n1301 = ( n1253 & ~n1249 ) | ( n1253 & n1300 ) | ( ~n1249 & n1300 ) ;
  assign n1653 = ( n1299 & n1301 ) | ( n1299 & n1652 ) | ( n1301 & n1652 ) ;
  assign n1151 = ( n1108 & ~n1111 ) | ( n1108 & n1150 ) | ( ~n1111 & n1150 ) ;
  assign n866 = ~n530 & n540 ;
  assign n867 = n540 | n542 ;
  assign n868 = ( n543 & ~n866 ) | ( n543 & n867 ) | ( ~n866 & n867 ) ;
  assign n805 = n788 | n793 ;
  assign n859 = n856 | n858 ;
  assign n857 = n852 &  n856 ;
  assign n860 = ( n850 & ~n859 ) | ( n850 & n857 ) | ( ~n859 & n857 ) ;
  assign n864 = n524 &  n863 ;
  assign n862 = n524 | n861 ;
  assign n865 = ( n860 & ~n864 ) | ( n860 & n862 ) | ( ~n864 & n862 ) ;
  assign n870 = ( n805 & n865 ) | ( n805 & n868 ) | ( n865 & n868 ) ;
  assign n869 = ( n805 & ~n868 ) | ( n805 & n865 ) | ( ~n868 & n865 ) ;
  assign n871 = ( n868 & ~n870 ) | ( n868 & n869 ) | ( ~n870 & n869 ) ;
  assign n804 = ( n722 & ~n545 ) | ( n722 & n803 ) | ( ~n545 & n803 ) ;
  assign n872 = ~n248 & n789 ;
  assign n873 = ( n248 & ~n796 ) | ( n248 & 1'b0 ) | ( ~n796 & 1'b0 ) ;
  assign n874 = ( n872 & ~n744 ) | ( n872 & n873 ) | ( ~n744 & n873 ) ;
  assign n875 = ( n712 & ~n799 ) | ( n712 & 1'b0 ) | ( ~n799 & 1'b0 ) ;
  assign n876 = n712 | n801 ;
  assign n877 = ( n874 & ~n875 ) | ( n874 & n876 ) | ( ~n875 & n876 ) ;
  assign n878 = n256 | n709 ;
  assign n879 = n256 &  n715 ;
  assign n880 = ( n666 & ~n878 ) | ( n666 & n879 ) | ( ~n878 & n879 ) ;
  assign n885 = n720 &  n883 ;
  assign n884 = n718 | n883 ;
  assign n886 = ( n880 & ~n885 ) | ( n880 & n884 ) | ( ~n885 & n884 ) ;
  assign n1000 = ( n994 & ~n937 ) | ( n994 & n999 ) | ( ~n937 & n999 ) ;
  assign n1001 = ( n877 & ~n886 ) | ( n877 & n1000 ) | ( ~n886 & n1000 ) ;
  assign n1002 = ( n877 & ~n1000 ) | ( n877 & n886 ) | ( ~n1000 & n886 ) ;
  assign n1003 = ( n1001 & ~n877 ) | ( n1001 & n1002 ) | ( ~n877 & n1002 ) ;
  assign n1004 = ( n804 & n871 ) | ( n804 & n1003 ) | ( n871 & n1003 ) ;
  assign n1152 = ( n804 & ~n871 ) | ( n804 & n1003 ) | ( ~n871 & n1003 ) ;
  assign n1153 = ( n871 & ~n1004 ) | ( n871 & n1152 ) | ( ~n1004 & n1152 ) ;
  assign n1158 = ( n1089 & n1151 ) | ( n1089 & n1153 ) | ( n1151 & n1153 ) ;
  assign n1159 = ( n1089 & ~n1151 ) | ( n1089 & n1153 ) | ( ~n1151 & n1153 ) ;
  assign n1160 = ( n1151 & ~n1158 ) | ( n1151 & n1159 ) | ( ~n1158 & n1159 ) ;
  assign n1755 = n1160 | n1253 ;
  assign n1756 = n1160 &  n1253 ;
  assign n1757 = ( n1755 & ~n1756 ) | ( n1755 & 1'b0 ) | ( ~n1756 & 1'b0 ) ;
  assign n1758 = n1653 | n1757 ;
  assign n1897 = ( n1653 & ~n1757 ) | ( n1653 & 1'b0 ) | ( ~n1757 & 1'b0 ) ;
  assign n1898 = ( n1758 & ~n1653 ) | ( n1758 & n1897 ) | ( ~n1653 & n1897 ) ;
  assign n1899 = ( n1891 & ~n1754 ) | ( n1891 & n1898 ) | ( ~n1754 & n1898 ) ;
  assign n1900 = ( n1754 & ~n1891 ) | ( n1754 & n1898 ) | ( ~n1891 & n1898 ) ;
  assign n1901 = ( n1899 & ~n1898 ) | ( n1899 & n1900 ) | ( ~n1898 & n1900 ) ;
  assign n1903 = ( x10 & n253 ) | ( x10 & n712 ) | ( n253 & n712 ) ;
  assign n1902 = ( x10 & ~n712 ) | ( x10 & n253 ) | ( ~n712 & n253 ) ;
  assign n1904 = ( n712 & ~n1903 ) | ( n712 & n1902 ) | ( ~n1903 & n1902 ) ;
  assign n1905 = ~n251 & n259 ;
  assign n1906 = ~n1904 & n1905 ;
  assign n1907 = ~n1901 & n1906 ;
  assign n1008 = ( n540 & ~n861 ) | ( n540 & 1'b0 ) | ( ~n861 & 1'b0 ) ;
  assign n1005 = ~n524 & n852 ;
  assign n1006 = ( n524 & ~n858 ) | ( n524 & 1'b0 ) | ( ~n858 & 1'b0 ) ;
  assign n1007 = ( n850 & n1005 ) | ( n850 & n1006 ) | ( n1005 & n1006 ) ;
  assign n1009 = ~n540 & n863 ;
  assign n1010 = ( n1008 & ~n1007 ) | ( n1008 & n1009 ) | ( ~n1007 & n1009 ) ;
  assign n1011 = ~n712 & n789 ;
  assign n1012 = ( n712 & ~n796 ) | ( n712 & 1'b0 ) | ( ~n796 & 1'b0 ) ;
  assign n1013 = ( n1011 & ~n744 ) | ( n1011 & n1012 ) | ( ~n744 & n1012 ) ;
  assign n1014 = ( n256 & ~n799 ) | ( n256 & 1'b0 ) | ( ~n799 & 1'b0 ) ;
  assign n1015 = n256 | n801 ;
  assign n1016 = ( n1013 & ~n1014 ) | ( n1013 & n1015 ) | ( ~n1014 & n1015 ) ;
  assign n1020 = ~n718 & n856 ;
  assign n1017 = ( n715 & ~n883 ) | ( n715 & 1'b0 ) | ( ~n883 & 1'b0 ) ;
  assign n1018 = ~n709 & n883 ;
  assign n1019 = ( n666 & n1017 ) | ( n666 & n1018 ) | ( n1017 & n1018 ) ;
  assign n1021 = ( n720 & ~n856 ) | ( n720 & 1'b0 ) | ( ~n856 & 1'b0 ) ;
  assign n1022 = ( n1020 & ~n1019 ) | ( n1020 & n1021 ) | ( ~n1019 & n1021 ) ;
  assign n1023 = ( n1010 & n1016 ) | ( n1010 & n1022 ) | ( n1016 & n1022 ) ;
  assign n1024 = ( n1016 & ~n1010 ) | ( n1016 & n1022 ) | ( ~n1010 & n1022 ) ;
  assign n1025 = ( n1010 & ~n1023 ) | ( n1010 & n1024 ) | ( ~n1023 & n1024 ) ;
  assign n1026 = ( n865 & ~n805 ) | ( n865 & n868 ) | ( ~n805 & n868 ) ;
  assign n1027 = ( n248 & ~n788 ) | ( n248 & 1'b0 ) | ( ~n788 & 1'b0 ) ;
  assign n1028 = ( n542 & ~n805 ) | ( n542 & n1027 ) | ( ~n805 & n1027 ) ;
  assign n1029 = ( n542 & ~n1027 ) | ( n542 & n805 ) | ( ~n1027 & n805 ) ;
  assign n1030 = ( n1028 & ~n542 ) | ( n1028 & n1029 ) | ( ~n542 & n1029 ) ;
  assign n1031 = ( n1026 & ~n1002 ) | ( n1026 & n1030 ) | ( ~n1002 & n1030 ) ;
  assign n1032 = ( n1002 & ~n1030 ) | ( n1002 & n1026 ) | ( ~n1030 & n1026 ) ;
  assign n1033 = ( n1031 & ~n1026 ) | ( n1031 & n1032 ) | ( ~n1026 & n1032 ) ;
  assign n1155 = ( n1004 & n1025 ) | ( n1004 & n1033 ) | ( n1025 & n1033 ) ;
  assign n1156 = ( n1004 & ~n1025 ) | ( n1004 & n1033 ) | ( ~n1025 & n1033 ) ;
  assign n1157 = ( n1025 & ~n1155 ) | ( n1025 & n1156 ) | ( ~n1155 & n1156 ) ;
  assign n1154 = ( n1151 & ~n1089 ) | ( n1151 & n1153 ) | ( ~n1089 & n1153 ) ;
  assign n1654 = ( n1160 & ~n1253 ) | ( n1160 & n1653 ) | ( ~n1253 & n1653 ) ;
  assign n1716 = ( n1154 & n1157 ) | ( n1154 & n1654 ) | ( n1157 & n1654 ) ;
  assign n1715 = ( n1154 & ~n1157 ) | ( n1154 & n1654 ) | ( ~n1157 & n1654 ) ;
  assign n1717 = ( n1157 & ~n1716 ) | ( n1157 & n1715 ) | ( ~n1716 & n1715 ) ;
  assign n1700 = n120 | n392 ;
  assign n1701 = n69 | n391 ;
  assign n1702 = n212 | n1701 ;
  assign n1703 = ( n920 & ~n1700 ) | ( n920 & n1702 ) | ( ~n1700 & n1702 ) ;
  assign n1704 = ( n1700 & ~n616 ) | ( n1700 & n1703 ) | ( ~n616 & n1703 ) ;
  assign n1705 = n616 | n1704 ;
  assign n1706 = ( n611 & ~n444 ) | ( n611 & n1705 ) | ( ~n444 & n1705 ) ;
  assign n1707 = n444 | n1706 ;
  assign n1708 = ( n1699 & ~n342 ) | ( n1699 & n1707 ) | ( ~n342 & n1707 ) ;
  assign n1709 = n342 | n1708 ;
  assign n1710 = ( n474 & n1693 ) | ( n474 & n1709 ) | ( n1693 & n1709 ) ;
  assign n1711 = ( n126 & ~n1710 ) | ( n126 & n1693 ) | ( ~n1710 & n1693 ) ;
  assign n1712 = ~n126 & n1711 ;
  assign n1713 = ( n191 & ~n364 ) | ( n191 & n1712 ) | ( ~n364 & n1712 ) ;
  assign n1714 = ~n191 & n1713 ;
  assign n1759 = n1653 &  n1757 ;
  assign n1760 = ( n1758 & ~n1759 ) | ( n1758 & 1'b0 ) | ( ~n1759 & 1'b0 ) ;
  assign n1892 = ( n1754 & ~n1760 ) | ( n1754 & n1891 ) | ( ~n1760 & n1891 ) ;
  assign n1908 = ( n1714 & n1717 ) | ( n1714 & n1892 ) | ( n1717 & n1892 ) ;
  assign n1909 = ( n1714 & ~n1717 ) | ( n1714 & n1892 ) | ( ~n1717 & n1892 ) ;
  assign n1910 = ( n1717 & ~n1908 ) | ( n1717 & n1909 ) | ( ~n1908 & n1909 ) ;
  assign n1911 = ~n251 & n1904 ;
  assign n1912 = ~n1910 & n1911 ;
  assign n1913 = n1907 | n1912 ;
  assign n1034 = ( n1025 & ~n1004 ) | ( n1025 & n1033 ) | ( ~n1004 & n1033 ) ;
  assign n1655 = ( n1154 & ~n1654 ) | ( n1154 & n1157 ) | ( ~n1654 & n1157 ) ;
  assign n1037 = n709 | n856 ;
  assign n1036 = n715 &  n856 ;
  assign n1038 = ( n666 & ~n1037 ) | ( n666 & n1036 ) | ( ~n1037 & n1036 ) ;
  assign n1040 = n524 &  n720 ;
  assign n1039 = n524 | n718 ;
  assign n1041 = ( n1038 & ~n1040 ) | ( n1038 & n1039 ) | ( ~n1040 & n1039 ) ;
  assign n1035 = ( n712 & ~n788 ) | ( n712 & 1'b0 ) | ( ~n788 & 1'b0 ) ;
  assign n1042 = ~n540 & n850 ;
  assign n1044 = ( n850 & n852 ) | ( n850 & n1042 ) | ( n852 & n1042 ) ;
  assign n1043 = ( n850 & ~n1042 ) | ( n850 & n858 ) | ( ~n1042 & n858 ) ;
  assign n1045 = ( n1042 & ~n1044 ) | ( n1042 & n1043 ) | ( ~n1044 & n1043 ) ;
  assign n1046 = ( n1041 & ~n1035 ) | ( n1041 & n1045 ) | ( ~n1035 & n1045 ) ;
  assign n1047 = ( n1035 & ~n1041 ) | ( n1035 & n1045 ) | ( ~n1041 & n1045 ) ;
  assign n1048 = ( n1046 & ~n1045 ) | ( n1046 & n1047 ) | ( ~n1045 & n1047 ) ;
  assign n1049 = ( n1002 & n1026 ) | ( n1002 & n1030 ) | ( n1026 & n1030 ) ;
  assign n1050 = ( n248 & ~n793 ) | ( n248 & n542 ) | ( ~n793 & n542 ) ;
  assign n1051 = ~n788 & n1050 ;
  assign n1052 = ~n256 & n789 ;
  assign n1053 = ( n256 & ~n796 ) | ( n256 & 1'b0 ) | ( ~n796 & 1'b0 ) ;
  assign n1054 = ( n1052 & ~n744 ) | ( n1052 & n1053 ) | ( ~n744 & n1053 ) ;
  assign n1056 = ~n801 & n883 ;
  assign n1055 = n799 | n883 ;
  assign n1057 = ( n1054 & ~n1056 ) | ( n1054 & n1055 ) | ( ~n1056 & n1055 ) ;
  assign n1058 = ( n1010 & ~n1016 ) | ( n1010 & n1022 ) | ( ~n1016 & n1022 ) ;
  assign n1059 = ( n1051 & ~n1057 ) | ( n1051 & n1058 ) | ( ~n1057 & n1058 ) ;
  assign n1060 = ( n1051 & ~n1058 ) | ( n1051 & n1057 ) | ( ~n1058 & n1057 ) ;
  assign n1061 = ( n1059 & ~n1051 ) | ( n1059 & n1060 ) | ( ~n1051 & n1060 ) ;
  assign n1062 = ( n1048 & ~n1049 ) | ( n1048 & n1061 ) | ( ~n1049 & n1061 ) ;
  assign n1063 = ( n1048 & ~n1061 ) | ( n1048 & n1049 ) | ( ~n1061 & n1049 ) ;
  assign n1064 = ( n1062 & ~n1048 ) | ( n1062 & n1063 ) | ( ~n1048 & n1063 ) ;
  assign n1656 = ( n1034 & ~n1655 ) | ( n1034 & n1064 ) | ( ~n1655 & n1064 ) ;
  assign n1657 = ( n1034 & ~n1064 ) | ( n1034 & n1655 ) | ( ~n1064 & n1655 ) ;
  assign n1658 = ( n1656 & ~n1034 ) | ( n1656 & n1657 ) | ( ~n1034 & n1657 ) ;
  assign n1659 = n200 | n392 ;
  assign n1660 = ( n147 & ~n97 ) | ( n147 & n1659 ) | ( ~n97 & n1659 ) ;
  assign n1661 = n97 | n1660 ;
  assign n1662 = ( n289 & ~n208 ) | ( n289 & n1661 ) | ( ~n208 & n1661 ) ;
  assign n1663 = n208 | n1662 ;
  assign n1664 = ( n190 & ~n142 ) | ( n190 & n1663 ) | ( ~n142 & n1663 ) ;
  assign n1665 = n142 | n1664 ;
  assign n1667 = n115 | n923 ;
  assign n1668 = ( n646 & ~n494 ) | ( n646 & n1667 ) | ( ~n494 & n1667 ) ;
  assign n1669 = ( n646 & ~n1668 ) | ( n646 & 1'b0 ) | ( ~n1668 & 1'b0 ) ;
  assign n1670 = ( n310 & ~n1666 ) | ( n310 & n1669 ) | ( ~n1666 & n1669 ) ;
  assign n1671 = ~n310 & n1670 ;
  assign n1672 = ( n292 & ~n647 ) | ( n292 & n1671 ) | ( ~n647 & n1671 ) ;
  assign n1673 = ~n292 & n1672 ;
  assign n1674 = ~n317 & n1673 ;
  assign n1675 = ~n69 & n466 ;
  assign n1676 = ~n612 & n1675 ;
  assign n1677 = n191 | n201 ;
  assign n1678 = ( n185 & ~n120 ) | ( n185 & n1677 ) | ( ~n120 & n1677 ) ;
  assign n1679 = n120 | n1678 ;
  assign n1680 = n281 | n1679 ;
  assign n1681 = ( n1674 & ~n1676 ) | ( n1674 & n1680 ) | ( ~n1676 & n1680 ) ;
  assign n1682 = ( n1674 & ~n1681 ) | ( n1674 & 1'b0 ) | ( ~n1681 & 1'b0 ) ;
  assign n1683 = ( n315 & ~n1665 ) | ( n315 & n1682 ) | ( ~n1665 & n1682 ) ;
  assign n1684 = ~n315 & n1683 ;
  assign n1685 = ( n167 & ~n352 ) | ( n167 & n1684 ) | ( ~n352 & n1684 ) ;
  assign n1686 = ~n167 & n1685 ;
  assign n1687 = ( n380 & ~n398 ) | ( n380 & n1686 ) | ( ~n398 & n1686 ) ;
  assign n1688 = ~n380 & n1687 ;
  assign n1689 = ( n316 & ~n668 ) | ( n316 & n1688 ) | ( ~n668 & n1688 ) ;
  assign n1690 = ~n316 & n1689 ;
  assign n1893 = ( n1717 & ~n1714 ) | ( n1717 & n1892 ) | ( ~n1714 & n1892 ) ;
  assign n1894 = ( n1658 & n1690 ) | ( n1658 & n1893 ) | ( n1690 & n1893 ) ;
  assign n1895 = ( n1690 & ~n1658 ) | ( n1690 & n1893 ) | ( ~n1658 & n1893 ) ;
  assign n1896 = ( n1658 & ~n1894 ) | ( n1658 & n1895 ) | ( ~n1894 & n1895 ) ;
  assign n1914 = ~n260 & n1896 ;
  assign n1915 = ( n260 & ~n1913 ) | ( n260 & n1914 ) | ( ~n1913 & n1914 ) ;
  assign n1916 = ~n251 | ~n259 ;
  assign n1918 = ( n1652 & n1788 ) | ( n1652 & n1794 ) | ( n1788 & n1794 ) ;
  assign n1917 = ( n1652 & ~n1794 ) | ( n1652 & n1788 ) | ( ~n1794 & n1788 ) ;
  assign n1919 = ( n1794 & ~n1918 ) | ( n1794 & n1917 ) | ( ~n1918 & n1917 ) ;
  assign n1920 = ~n1890 & n1919 ;
  assign n1921 = ( n1890 & ~n1919 ) | ( n1890 & 1'b0 ) | ( ~n1919 & 1'b0 ) ;
  assign n1922 = n1920 | n1921 ;
  assign n1925 = ~n597 & n1885 ;
  assign n1926 = ( n1863 & ~n1649 ) | ( n1863 & n1925 ) | ( ~n1649 & n1925 ) ;
  assign n1927 = ( n1649 & n1863 ) | ( n1649 & n1925 ) | ( n1863 & n1925 ) ;
  assign n1928 = ( ~n1649 & ~n1926 ) | ( ~n1649 & n1927 ) | ( ~n1926 & n1927 ) ;
  assign n1923 = ( n1828 & ~n1830 ) | ( n1828 & n1889 ) | ( ~n1830 & n1889 ) ;
  assign n1924 = ( n1830 & ~n1890 ) | ( n1830 & n1923 ) | ( ~n1890 & n1923 ) ;
  assign n1931 = ~n1928 & n1924 ;
  assign n1929 = ( n1857 & ~n1888 ) | ( n1857 & n1860 ) | ( ~n1888 & n1860 ) ;
  assign n1930 = ( n1889 & ~n1860 ) | ( n1889 & n1929 ) | ( ~n1860 & n1929 ) ;
  assign n1932 = ( n1931 & ~n1924 ) | ( n1931 & n1930 ) | ( ~n1924 & n1930 ) ;
  assign n1933 = ( n1922 & ~n1932 ) | ( n1922 & n1924 ) | ( ~n1932 & n1924 ) ;
  assign n1934 = ( n1901 & n1922 ) | ( n1901 & n1933 ) | ( n1922 & n1933 ) ;
  assign n1935 = ( n1901 & n1910 ) | ( n1901 & n1934 ) | ( n1910 & n1934 ) ;
  assign n1936 = ( n1910 & ~n1896 ) | ( n1910 & n1935 ) | ( ~n1896 & n1935 ) ;
  assign n1937 = ( n1896 & ~n1935 ) | ( n1896 & n1910 ) | ( ~n1935 & n1910 ) ;
  assign n1938 = ( n1936 & ~n1910 ) | ( n1936 & n1937 ) | ( ~n1910 & n1937 ) ;
  assign n1939 = n1916 | n1938 ;
  assign n1940 = n1915 &  n1939 ;
  assign n2061 = n883 &  n1940 ;
  assign n2060 = ( n883 & ~n1940 ) | ( n883 & 1'b0 ) | ( ~n1940 & 1'b0 ) ;
  assign n2062 = ( n1940 & ~n2061 ) | ( n1940 & n2060 ) | ( ~n2061 & n2060 ) ;
  assign n1941 = ( x12 & n853 ) | ( x12 & n883 ) | ( n853 & n883 ) ;
  assign n1942 = ( x12 & ~n883 ) | ( x12 & n853 ) | ( ~n883 & n853 ) ;
  assign n1943 = ( n883 & ~n1941 ) | ( n883 & n1942 ) | ( ~n1941 & n1942 ) ;
  assign n1949 = ( x14 & n524 ) | ( x14 & n537 ) | ( n524 & n537 ) ;
  assign n1950 = ( x14 & ~n524 ) | ( x14 & n537 ) | ( ~n524 & n537 ) ;
  assign n1951 = ( n524 & ~n1949 ) | ( n524 & n1950 ) | ( ~n1949 & n1950 ) ;
  assign n1958 = n1943 | n1951 ;
  assign n1955 = n1928 | n1930 ;
  assign n1956 = n1928 &  n1930 ;
  assign n1957 = ( n1955 & ~n1956 ) | ( n1955 & 1'b0 ) | ( ~n1956 & 1'b0 ) ;
  assign n1959 = ~n1958 & n1957 ;
  assign n1945 = ( x13 & n521 ) | ( x13 & n856 ) | ( n521 & n856 ) ;
  assign n1944 = ( x13 & ~n856 ) | ( x13 & n521 ) | ( ~n856 & n521 ) ;
  assign n1946 = ( n856 & ~n1945 ) | ( n856 & n1944 ) | ( ~n1945 & n1944 ) ;
  assign n1947 = n1943 &  n1946 ;
  assign n1948 = ~n1928 & n1947 ;
  assign n1952 = ~n1943 & n1951 ;
  assign n1953 = n1930 &  n1952 ;
  assign n1954 = n1948 | n1953 ;
  assign n1960 = ( n1959 & ~n1954 ) | ( n1959 & n1958 ) | ( ~n1954 & n1958 ) ;
  assign n1961 = n1928 | n1943 ;
  assign n1965 = ~n1924 & n1952 ;
  assign n1966 = ( n1943 & ~n1951 ) | ( n1943 & 1'b0 ) | ( ~n1951 & 1'b0 ) ;
  assign n1967 = ~n1946 & n1966 ;
  assign n1968 = ~n1928 & n1967 ;
  assign n1969 = n1930 &  n1947 ;
  assign n1970 = n1968 | n1969 ;
  assign n1971 = n1965 | n1970 ;
  assign n1962 = ( n1924 & ~n1956 ) | ( n1924 & 1'b0 ) | ( ~n1956 & 1'b0 ) ;
  assign n1963 = ~n1924 & n1956 ;
  assign n1964 = n1962 | n1963 ;
  assign n1972 = ~n1958 & n1964 ;
  assign n1973 = ( n1958 & ~n1971 ) | ( n1958 & n1972 ) | ( ~n1971 & n1972 ) ;
  assign n1974 = ( n1961 & ~n1960 ) | ( n1961 & n1973 ) | ( ~n1960 & n1973 ) ;
  assign n1975 = ( n1960 & ~n540 ) | ( n1960 & n1974 ) | ( ~n540 & n1974 ) ;
  assign n1976 = n540 &  n1975 ;
  assign n1978 = ~n1924 & n1947 ;
  assign n1979 = n1930 &  n1967 ;
  assign n1980 = n1978 | n1979 ;
  assign n1981 = n1922 | n1952 ;
  assign n1982 = ( n1980 & ~n1922 ) | ( n1980 & n1981 ) | ( ~n1922 & n1981 ) ;
  assign n1983 = ( n1922 & n1924 ) | ( n1922 & n1932 ) | ( n1924 & n1932 ) ;
  assign n1984 = ( n1922 & ~n1924 ) | ( n1922 & n1932 ) | ( ~n1924 & n1932 ) ;
  assign n1985 = ( n1924 & ~n1983 ) | ( n1924 & n1984 ) | ( ~n1983 & n1984 ) ;
  assign n1986 = ~n1958 & n1985 ;
  assign n1987 = n1982 | n1986 ;
  assign n1988 = n540 | n1987 ;
  assign n1989 = n540 &  n1987 ;
  assign n1990 = ( n1988 & ~n1989 ) | ( n1988 & 1'b0 ) | ( ~n1989 & 1'b0 ) ;
  assign n1977 = ( n540 & ~n1928 ) | ( n540 & 1'b0 ) | ( ~n1928 & 1'b0 ) ;
  assign n1991 = ( n1976 & ~n1990 ) | ( n1976 & n1977 ) | ( ~n1990 & n1977 ) ;
  assign n1992 = ( n1976 & ~n1977 ) | ( n1976 & n1990 ) | ( ~n1977 & n1990 ) ;
  assign n1993 = ( n1991 & ~n1976 ) | ( n1991 & n1992 ) | ( ~n1976 & n1992 ) ;
  assign n2041 = ( n1906 & ~n1922 ) | ( n1906 & 1'b0 ) | ( ~n1922 & 1'b0 ) ;
  assign n2042 = ~n1901 & n1911 ;
  assign n2043 = n2041 | n2042 ;
  assign n2044 = ~n260 & n1910 ;
  assign n2045 = ( n260 & ~n2043 ) | ( n260 & n2044 ) | ( ~n2043 & n2044 ) ;
  assign n2046 = ( n1901 & ~n1934 ) | ( n1901 & n1910 ) | ( ~n1934 & n1910 ) ;
  assign n2047 = ( n1901 & ~n1910 ) | ( n1901 & n1934 ) | ( ~n1910 & n1934 ) ;
  assign n2048 = ( n2046 & ~n1901 ) | ( n2046 & n2047 ) | ( ~n1901 & n2047 ) ;
  assign n2049 = n1916 | n2048 ;
  assign n2050 = n2045 &  n2049 ;
  assign n2051 = ( x11 & ~n252 ) | ( x11 & n2050 ) | ( ~n252 & n2050 ) ;
  assign n2052 = ( x11 & ~n2050 ) | ( x11 & n252 ) | ( ~n2050 & n252 ) ;
  assign n2053 = ( n2051 & ~x11 ) | ( n2051 & n2052 ) | ( ~x11 & n2052 ) ;
  assign n2003 = ( n1901 & ~n1922 ) | ( n1901 & n1933 ) | ( ~n1922 & n1933 ) ;
  assign n2004 = ( n1922 & ~n1934 ) | ( n1922 & n2003 ) | ( ~n1934 & n2003 ) ;
  assign n1998 = ( n1906 & ~n1924 ) | ( n1906 & 1'b0 ) | ( ~n1924 & 1'b0 ) ;
  assign n1999 = ( n1911 & ~n1922 ) | ( n1911 & 1'b0 ) | ( ~n1922 & 1'b0 ) ;
  assign n2000 = n1998 | n1999 ;
  assign n2001 = ~n260 & n1901 ;
  assign n2002 = ( n260 & ~n2000 ) | ( n260 & n2001 ) | ( ~n2000 & n2001 ) ;
  assign n2005 = ( n1916 & ~n2004 ) | ( n1916 & n2002 ) | ( ~n2004 & n2002 ) ;
  assign n2006 = ~n1916 & n2005 ;
  assign n2008 = ( n883 & n2002 ) | ( n883 & n2006 ) | ( n2002 & n2006 ) ;
  assign n2007 = ( n883 & ~n2006 ) | ( n883 & n2002 ) | ( ~n2006 & n2002 ) ;
  assign n2009 = ( n2006 & ~n2008 ) | ( n2006 & n2007 ) | ( ~n2008 & n2007 ) ;
  assign n1994 = n540 &  n1961 ;
  assign n1995 = ( n540 & n1960 ) | ( n540 & n1994 ) | ( n1960 & n1994 ) ;
  assign n1996 = ( n540 & ~n1994 ) | ( n540 & n1960 ) | ( ~n1994 & n1960 ) ;
  assign n1997 = ( n1994 & ~n1995 ) | ( n1994 & n1996 ) | ( ~n1995 & n1996 ) ;
  assign n2010 = ( n251 & ~n1928 ) | ( n251 & 1'b0 ) | ( ~n1928 & 1'b0 ) ;
  assign n2011 = ( n1911 & ~n1928 ) | ( n1911 & 1'b0 ) | ( ~n1928 & 1'b0 ) ;
  assign n2012 = ~n260 & n1930 ;
  assign n2013 = n2011 | n2012 ;
  assign n2014 = ~n1916 & n1957 ;
  assign n2015 = ( n1916 & ~n2013 ) | ( n1916 & n2014 ) | ( ~n2013 & n2014 ) ;
  assign n2016 = ( n883 & ~n2010 ) | ( n883 & n2015 ) | ( ~n2010 & n2015 ) ;
  assign n2017 = ~n883 & n2016 ;
  assign n2018 = ( n1906 & ~n1928 ) | ( n1906 & 1'b0 ) | ( ~n1928 & 1'b0 ) ;
  assign n2019 = n1911 &  n1930 ;
  assign n2020 = n2018 | n2019 ;
  assign n2021 = ~n260 & n1924 ;
  assign n2022 = ( n260 & ~n2020 ) | ( n260 & n2021 ) | ( ~n2020 & n2021 ) ;
  assign n2023 = ( n1916 & ~n1964 ) | ( n1916 & n2022 ) | ( ~n1964 & n2022 ) ;
  assign n2024 = ~n1916 & n2023 ;
  assign n2025 = ( n883 & ~n2022 ) | ( n883 & n2024 ) | ( ~n2022 & n2024 ) ;
  assign n2026 = ( n2022 & ~n883 ) | ( n2022 & n2024 ) | ( ~n883 & n2024 ) ;
  assign n2027 = ( n2025 & ~n2024 ) | ( n2025 & n2026 ) | ( ~n2024 & n2026 ) ;
  assign n2028 = n2017 &  n2027 ;
  assign n2029 = ( n1911 & ~n1924 ) | ( n1911 & 1'b0 ) | ( ~n1924 & 1'b0 ) ;
  assign n2030 = n1906 &  n1930 ;
  assign n2031 = n2029 | n2030 ;
  assign n2032 = ~n260 & n1922 ;
  assign n2033 = ( n260 & ~n2031 ) | ( n260 & n2032 ) | ( ~n2031 & n2032 ) ;
  assign n2034 = ( n1916 & n1985 ) | ( n1916 & n2033 ) | ( n1985 & n2033 ) ;
  assign n2035 = ~n1916 & n2034 ;
  assign n2037 = ( n883 & n2033 ) | ( n883 & n2035 ) | ( n2033 & n2035 ) ;
  assign n2036 = ( n883 & ~n2035 ) | ( n883 & n2033 ) | ( ~n2035 & n2033 ) ;
  assign n2038 = ( n2035 & ~n2037 ) | ( n2035 & n2036 ) | ( ~n2037 & n2036 ) ;
  assign n2039 = ( n2028 & ~n1961 ) | ( n2028 & n2038 ) | ( ~n1961 & n2038 ) ;
  assign n2040 = ( n2009 & ~n1997 ) | ( n2009 & n2039 ) | ( ~n1997 & n2039 ) ;
  assign n2054 = ( n540 & ~n1960 ) | ( n540 & n1961 ) | ( ~n1960 & n1961 ) ;
  assign n2055 = n1960 &  n2054 ;
  assign n2056 = ( n1973 & ~n540 ) | ( n1973 & n2055 ) | ( ~n540 & n2055 ) ;
  assign n2057 = ( n540 & ~n1973 ) | ( n540 & n2055 ) | ( ~n1973 & n2055 ) ;
  assign n2058 = ( n2056 & ~n2055 ) | ( n2056 & n2057 ) | ( ~n2055 & n2057 ) ;
  assign n2059 = ( n2053 & ~n2040 ) | ( n2053 & n2058 ) | ( ~n2040 & n2058 ) ;
  assign n2063 = ( n1993 & n2059 ) | ( n1993 & n2062 ) | ( n2059 & n2062 ) ;
  assign n2064 = ( n1993 & ~n2062 ) | ( n1993 & n2059 ) | ( ~n2062 & n2059 ) ;
  assign n2065 = ( n2062 & ~n2063 ) | ( n2062 & n2064 ) | ( ~n2063 & n2064 ) ;
  assign n2066 = ( n2040 & ~n2058 ) | ( n2040 & n2053 ) | ( ~n2058 & n2053 ) ;
  assign n2067 = ( n2059 & ~n2053 ) | ( n2059 & n2066 ) | ( ~n2053 & n2066 ) ;
  assign n2188 = ( x8 & n245 ) | ( x8 & n793 ) | ( n245 & n793 ) ;
  assign n2189 = ( x8 & ~n793 ) | ( x8 & n245 ) | ( ~n793 & n245 ) ;
  assign n2190 = ( n793 & ~n2188 ) | ( n793 & n2189 ) | ( ~n2188 & n2189 ) ;
  assign n2191 = ( x6 & n995 ) | ( x6 & n1077 ) | ( n995 & n1077 ) ;
  assign n2192 = ( x6 & ~n1077 ) | ( x6 & n995 ) | ( ~n1077 & n995 ) ;
  assign n2193 = ( n1077 & ~n2191 ) | ( n1077 & n2192 ) | ( ~n2191 & n2192 ) ;
  assign n2213 = n2190 | n2193 ;
  assign n2082 = ( n256 & ~n788 ) | ( n256 & 1'b0 ) | ( ~n788 & 1'b0 ) ;
  assign n2101 = ( n858 & n1035 ) | ( n858 & n2082 ) | ( n1035 & n2082 ) ;
  assign n2083 = ( n1035 & ~n858 ) | ( n1035 & n2082 ) | ( ~n858 & n2082 ) ;
  assign n2102 = ( n858 & ~n2101 ) | ( n858 & n2083 ) | ( ~n2101 & n2083 ) ;
  assign n2071 = ( n540 & ~n718 ) | ( n540 & 1'b0 ) | ( ~n718 & 1'b0 ) ;
  assign n2068 = ~n524 & n715 ;
  assign n2069 = ( n524 & ~n709 ) | ( n524 & 1'b0 ) | ( ~n709 & 1'b0 ) ;
  assign n2070 = ( n666 & n2068 ) | ( n666 & n2069 ) | ( n2068 & n2069 ) ;
  assign n2072 = ~n540 & n720 ;
  assign n2073 = ( n2071 & ~n2070 ) | ( n2071 & n2072 ) | ( ~n2070 & n2072 ) ;
  assign n2080 = ( n1035 & ~n1045 ) | ( n1035 & n1041 ) | ( ~n1045 & n1041 ) ;
  assign n2074 = n789 &  n883 ;
  assign n2075 = n796 | n883 ;
  assign n2076 = ( n744 & ~n2074 ) | ( n744 & n2075 ) | ( ~n2074 & n2075 ) ;
  assign n2078 = n801 | n856 ;
  assign n2077 = ~n799 & n856 ;
  assign n2079 = ( n2076 & ~n2078 ) | ( n2076 & n2077 ) | ( ~n2078 & n2077 ) ;
  assign n2081 = ( n2073 & ~n2080 ) | ( n2073 & n2079 ) | ( ~n2080 & n2079 ) ;
  assign n2103 = ( n2079 & ~n2073 ) | ( n2079 & n2080 ) | ( ~n2073 & n2080 ) ;
  assign n2104 = ( n2081 & ~n2079 ) | ( n2081 & n2103 ) | ( ~n2079 & n2103 ) ;
  assign n2105 = ( n2102 & ~n1059 ) | ( n2102 & n2104 ) | ( ~n1059 & n2104 ) ;
  assign n2107 = ( n1059 & ~n2104 ) | ( n1059 & n2102 ) | ( ~n2104 & n2102 ) ;
  assign n2108 = ( n2105 & ~n2102 ) | ( n2105 & n2107 ) | ( ~n2102 & n2107 ) ;
  assign n2106 = ( n1049 & ~n1048 ) | ( n1049 & n1061 ) | ( ~n1048 & n1061 ) ;
  assign n2109 = ( n1064 & ~n1034 ) | ( n1064 & n1655 ) | ( ~n1034 & n1655 ) ;
  assign n2181 = ( n2106 & n2108 ) | ( n2106 & n2109 ) | ( n2108 & n2109 ) ;
  assign n2180 = ( n2106 & ~n2108 ) | ( n2106 & n2109 ) | ( ~n2108 & n2109 ) ;
  assign n2182 = ( n2108 & ~n2181 ) | ( n2108 & n2180 ) | ( ~n2181 & n2180 ) ;
  assign n2139 = n153 | n363 ;
  assign n2140 = n282 | n2139 ;
  assign n2151 = n746 | n2140 ;
  assign n2152 = ( n669 & ~n113 ) | ( n669 & n2151 ) | ( ~n113 & n2151 ) ;
  assign n2153 = n113 | n2152 ;
  assign n2154 = ( n162 & ~n105 ) | ( n162 & n2153 ) | ( ~n105 & n2153 ) ;
  assign n2155 = n105 | n2154 ;
  assign n2156 = ( n290 & ~n501 ) | ( n290 & n2155 ) | ( ~n501 & n2155 ) ;
  assign n2157 = n501 | n2156 ;
  assign n2158 = ( n597 & ~n261 ) | ( n597 & n2157 ) | ( ~n261 & n2157 ) ;
  assign n2159 = n261 | n2158 ;
  assign n2160 = n114 | n812 ;
  assign n2161 = ( n647 & ~n467 ) | ( n647 & n2160 ) | ( ~n467 & n2160 ) ;
  assign n2162 = n467 | n2161 ;
  assign n2163 = ( n289 & ~n122 ) | ( n289 & n2162 ) | ( ~n122 & n2162 ) ;
  assign n2164 = n122 | n2163 ;
  assign n2165 = n554 | n2164 ;
  assign n2125 = n110 | n319 ;
  assign n2126 = n380 | n2125 ;
  assign n210 = n208 | n209 ;
  assign n2127 = ( n315 & ~n227 ) | ( n315 & n690 ) | ( ~n227 & n690 ) ;
  assign n2128 = n227 | n2127 ;
  assign n2129 = n1868 | n2128 ;
  assign n2130 = ( n830 & ~n210 ) | ( n830 & n2129 ) | ( ~n210 & n2129 ) ;
  assign n2131 = n210 | n2130 ;
  assign n2132 = ( n2126 & ~n637 ) | ( n2126 & n2131 ) | ( ~n637 & n2131 ) ;
  assign n2133 = n637 | n2132 ;
  assign n2134 = ( n549 & ~n195 ) | ( n549 & n2133 ) | ( ~n195 & n2133 ) ;
  assign n2135 = n195 | n2134 ;
  assign n2136 = ( n324 & ~n199 ) | ( n324 & n2135 ) | ( ~n199 & n2135 ) ;
  assign n2137 = n199 | n2136 ;
  assign n2138 = n180 | n2137 ;
  assign n2166 = n126 | n2138 ;
  assign n2167 = ( n436 & ~n189 ) | ( n436 & n2166 ) | ( ~n189 & n2166 ) ;
  assign n2168 = n189 | n2167 ;
  assign n2169 = ( n1192 & ~n1803 ) | ( n1192 & n2168 ) | ( ~n1803 & n2168 ) ;
  assign n2170 = ( n496 & n1803 ) | ( n496 & n2169 ) | ( n1803 & n2169 ) ;
  assign n2171 = ( n496 & ~n2170 ) | ( n496 & 1'b0 ) | ( ~n2170 & 1'b0 ) ;
  assign n2172 = ( n2159 & ~n2165 ) | ( n2159 & n2171 ) | ( ~n2165 & n2171 ) ;
  assign n2173 = ( n326 & ~n2159 ) | ( n326 & n2172 ) | ( ~n2159 & n2172 ) ;
  assign n2174 = ~n326 & n2173 ;
  assign n2175 = ( n478 & ~n610 ) | ( n478 & n2174 ) | ( ~n610 & n2174 ) ;
  assign n2176 = ~n478 & n2175 ;
  assign n2177 = ( n141 & ~n293 ) | ( n141 & n2176 ) | ( ~n293 & n2176 ) ;
  assign n2178 = ~n141 & n2177 ;
  assign n2179 = ~n412 & n2178 ;
  assign n2183 = ( n1658 & ~n1690 ) | ( n1658 & n1893 ) | ( ~n1690 & n1893 ) ;
  assign n2184 = ( n2182 & ~n2179 ) | ( n2182 & n2183 ) | ( ~n2179 & n2183 ) ;
  assign n2202 = ( n2179 & ~n2183 ) | ( n2179 & n2182 ) | ( ~n2183 & n2182 ) ;
  assign n2203 = ( n2184 & ~n2182 ) | ( n2184 & n2202 ) | ( ~n2182 & n2202 ) ;
  assign n2208 = ( n1896 & n1910 ) | ( n1896 & n1935 ) | ( n1910 & n1935 ) ;
  assign n2224 = ( n1896 & ~n2203 ) | ( n1896 & n2208 ) | ( ~n2203 & n2208 ) ;
  assign n2225 = ( n1896 & ~n2208 ) | ( n1896 & n2203 ) | ( ~n2208 & n2203 ) ;
  assign n2226 = ( n2224 & ~n1896 ) | ( n2224 & n2225 ) | ( ~n1896 & n2225 ) ;
  assign n2194 = ~n2190 |  n2193 ;
  assign n2197 = ( x7 & n790 ) | ( x7 & n998 ) | ( n790 & n998 ) ;
  assign n2196 = ( x7 & ~n998 ) | ( x7 & n790 ) | ( ~n998 & n790 ) ;
  assign n2198 = ( n998 & ~n2197 ) | ( n998 & n2196 ) | ( ~n2197 & n2196 ) ;
  assign n2199 = ~n2190 & n2193 ;
  assign n2200 = ~n2198 & n2199 ;
  assign n2219 = ~n1910 & n2200 ;
  assign n2204 = n2193 &  n2198 ;
  assign n2220 = ~n1896 & n2204 ;
  assign n2221 = n2219 | n2220 ;
  assign n2222 = ~n2194 & n2203 ;
  assign n2223 = ( n2194 & ~n2221 ) | ( n2194 & n2222 ) | ( ~n2221 & n2222 ) ;
  assign n2227 = ( n2213 & ~n2226 ) | ( n2213 & n2223 ) | ( ~n2226 & n2223 ) ;
  assign n2228 = ~n2213 & n2227 ;
  assign n2230 = ( n248 & n2223 ) | ( n248 & n2228 ) | ( n2223 & n2228 ) ;
  assign n2229 = ( n248 & ~n2228 ) | ( n248 & n2223 ) | ( ~n2228 & n2223 ) ;
  assign n2231 = ( n2228 & ~n2230 ) | ( n2228 & n2229 ) | ( ~n2230 & n2229 ) ;
  assign n2232 = ( n1997 & ~n2039 ) | ( n1997 & n2009 ) | ( ~n2039 & n2009 ) ;
  assign n2233 = ( n2040 & ~n2009 ) | ( n2040 & n2232 ) | ( ~n2009 & n2232 ) ;
  assign n2234 = ( n1961 & ~n2028 ) | ( n1961 & n2038 ) | ( ~n2028 & n2038 ) ;
  assign n2235 = ( n2039 & ~n2038 ) | ( n2039 & n2234 ) | ( ~n2038 & n2234 ) ;
  assign n2236 = ~n1901 & n2200 ;
  assign n2237 = ~n1910 & n2204 ;
  assign n2238 = n2236 | n2237 ;
  assign n2239 = ~n1896 & n2194 ;
  assign n2240 = ( n1896 & ~n2238 ) | ( n1896 & n2239 ) | ( ~n2238 & n2239 ) ;
  assign n2241 = ( n2213 & ~n1938 ) | ( n2213 & n2240 ) | ( ~n1938 & n2240 ) ;
  assign n2242 = ~n2213 & n2241 ;
  assign n2244 = ( n248 & n2240 ) | ( n248 & n2242 ) | ( n2240 & n2242 ) ;
  assign n2243 = ( n248 & ~n2242 ) | ( n248 & n2240 ) | ( ~n2242 & n2240 ) ;
  assign n2245 = ( n2242 & ~n2244 ) | ( n2242 & n2243 ) | ( ~n2244 & n2243 ) ;
  assign n2246 = ~n1922 & n2200 ;
  assign n2247 = ~n1901 & n2204 ;
  assign n2248 = n2246 | n2247 ;
  assign n2249 = ~n1910 & n2194 ;
  assign n2250 = ( n1910 & ~n2248 ) | ( n1910 & n2249 ) | ( ~n2248 & n2249 ) ;
  assign n2251 = n2048 | n2213 ;
  assign n2252 = n2250 &  n2251 ;
  assign n2253 = ~n248 & n2252 ;
  assign n2254 = ( n248 & ~n2252 ) | ( n248 & 1'b0 ) | ( ~n2252 & 1'b0 ) ;
  assign n2255 = n2253 | n2254 ;
  assign n2256 = n2017 | n2027 ;
  assign n2257 = ~n2028 & n2256 ;
  assign n2258 = ~n883 & n2010 ;
  assign n2259 = ~n2015 & n2258 ;
  assign n2260 = ( n2015 & ~n2258 ) | ( n2015 & 1'b0 ) | ( ~n2258 & 1'b0 ) ;
  assign n2261 = n2259 | n2260 ;
  assign n2291 = ~n1924 & n2204 ;
  assign n2292 = n1930 &  n2200 ;
  assign n2293 = n2291 | n2292 ;
  assign n2294 = ~n1922 & n2194 ;
  assign n2295 = ( n1922 & ~n2293 ) | ( n1922 & n2294 ) | ( ~n2293 & n2294 ) ;
  assign n2296 = ( n1985 & ~n2213 ) | ( n1985 & 1'b0 ) | ( ~n2213 & 1'b0 ) ;
  assign n2297 = ( n2295 & ~n2296 ) | ( n2295 & 1'b0 ) | ( ~n2296 & 1'b0 ) ;
  assign n2298 = ~n248 & n2297 ;
  assign n2299 = ( n248 & ~n2297 ) | ( n248 & 1'b0 ) | ( ~n2297 & 1'b0 ) ;
  assign n2300 = n2298 | n2299 ;
  assign n2272 = ~n1928 & n2204 ;
  assign n2273 = ( n1930 & ~n2194 ) | ( n1930 & 1'b0 ) | ( ~n2194 & 1'b0 ) ;
  assign n2274 = n2272 | n2273 ;
  assign n2275 = ~n1957 & n2213 ;
  assign n2276 = ( n1957 & ~n2274 ) | ( n1957 & n2275 ) | ( ~n2274 & n2275 ) ;
  assign n2277 = n1928 | n2193 ;
  assign n2278 = ( n2276 & ~n248 ) | ( n2276 & n2277 ) | ( ~n248 & n2277 ) ;
  assign n2279 = n248 &  n2278 ;
  assign n2280 = ~n1928 & n2200 ;
  assign n2281 = n1930 &  n2204 ;
  assign n2282 = n2280 | n2281 ;
  assign n2283 = ~n1924 & n2194 ;
  assign n2284 = ( n1924 & ~n2282 ) | ( n1924 & n2283 ) | ( ~n2282 & n2283 ) ;
  assign n2285 = ( n2213 & ~n1964 ) | ( n2213 & n2284 ) | ( ~n1964 & n2284 ) ;
  assign n2286 = ~n2213 & n2285 ;
  assign n2288 = ( n248 & n2284 ) | ( n248 & n2286 ) | ( n2284 & n2286 ) ;
  assign n2287 = ( n248 & ~n2286 ) | ( n248 & n2284 ) | ( ~n2286 & n2284 ) ;
  assign n2289 = ( n2286 & ~n2288 ) | ( n2286 & n2287 ) | ( ~n2288 & n2287 ) ;
  assign n2290 = ( n2279 & ~n2289 ) | ( n2279 & 1'b0 ) | ( ~n2289 & 1'b0 ) ;
  assign n2301 = ( n2010 & ~n2300 ) | ( n2010 & n2290 ) | ( ~n2300 & n2290 ) ;
  assign n2262 = ~n1924 & n2200 ;
  assign n2263 = ~n1922 & n2204 ;
  assign n2264 = n2262 | n2263 ;
  assign n2265 = ~n1901 & n2194 ;
  assign n2266 = ( n1901 & ~n2264 ) | ( n1901 & n2265 ) | ( ~n2264 & n2265 ) ;
  assign n2267 = ( n2213 & ~n2004 ) | ( n2213 & n2266 ) | ( ~n2004 & n2266 ) ;
  assign n2268 = ~n2213 & n2267 ;
  assign n2269 = ( n248 & ~n2266 ) | ( n248 & n2268 ) | ( ~n2266 & n2268 ) ;
  assign n2270 = ( n2266 & ~n248 ) | ( n2266 & n2268 ) | ( ~n248 & n2268 ) ;
  assign n2271 = ( n2269 & ~n2268 ) | ( n2269 & n2270 ) | ( ~n2268 & n2270 ) ;
  assign n2302 = ( n2261 & ~n2301 ) | ( n2261 & n2271 ) | ( ~n2301 & n2271 ) ;
  assign n2303 = ( n2255 & ~n2257 ) | ( n2255 & n2302 ) | ( ~n2257 & n2302 ) ;
  assign n2304 = ( n2235 & n2245 ) | ( n2235 & n2303 ) | ( n2245 & n2303 ) ;
  assign n2305 = ( n2231 & n2233 ) | ( n2231 & n2304 ) | ( n2233 & n2304 ) ;
  assign n2091 = ~n540 & n666 ;
  assign n2092 = ( n666 & ~n2091 ) | ( n666 & n715 ) | ( ~n2091 & n715 ) ;
  assign n2093 = ( n709 & ~n666 ) | ( n709 & n2091 ) | ( ~n666 & n2091 ) ;
  assign n2094 = ( n2092 & ~n715 ) | ( n2092 & n2093 ) | ( ~n715 & n2093 ) ;
  assign n2084 = n788 | n883 ;
  assign n2085 = ( n789 & ~n856 ) | ( n789 & 1'b0 ) | ( ~n856 & 1'b0 ) ;
  assign n2086 = ~n796 & n856 ;
  assign n2087 = ( n2085 & ~n744 ) | ( n2085 & n2086 ) | ( ~n744 & n2086 ) ;
  assign n2089 = ( n524 & ~n801 ) | ( n524 & 1'b0 ) | ( ~n801 & 1'b0 ) ;
  assign n2088 = n524 | n799 ;
  assign n2090 = ( n2087 & ~n2089 ) | ( n2087 & n2088 ) | ( ~n2089 & n2088 ) ;
  assign n2095 = ( n2084 & n2090 ) | ( n2084 & n2094 ) | ( n2090 & n2094 ) ;
  assign n2096 = ( n2084 & ~n2094 ) | ( n2084 & n2090 ) | ( ~n2094 & n2090 ) ;
  assign n2097 = ( n2094 & ~n2095 ) | ( n2094 & n2096 ) | ( ~n2095 & n2096 ) ;
  assign n2098 = ( n2081 & ~n2083 ) | ( n2081 & n2097 ) | ( ~n2083 & n2097 ) ;
  assign n2099 = ( n2081 & ~n2097 ) | ( n2081 & n2083 ) | ( ~n2097 & n2083 ) ;
  assign n2100 = ( n2098 & ~n2081 ) | ( n2098 & n2099 ) | ( ~n2081 & n2099 ) ;
  assign n2110 = ( n2108 & ~n2106 ) | ( n2108 & n2109 ) | ( ~n2106 & n2109 ) ;
  assign n2112 = ( n2100 & n2105 ) | ( n2100 & n2110 ) | ( n2105 & n2110 ) ;
  assign n2111 = ( n2105 & ~n2100 ) | ( n2105 & n2110 ) | ( ~n2100 & n2110 ) ;
  assign n2113 = ( n2100 & ~n2112 ) | ( n2100 & n2111 ) | ( ~n2112 & n2111 ) ;
  assign n2114 = n226 | n438 ;
  assign n2115 = ( n292 & ~n122 ) | ( n292 & n2114 ) | ( ~n122 & n2114 ) ;
  assign n2116 = n122 | n2115 ;
  assign n2117 = ( n212 & ~n78 ) | ( n212 & n2116 ) | ( ~n78 & n2116 ) ;
  assign n2118 = n78 | n2117 ;
  assign n2119 = ~n575 & n629 ;
  assign n2120 = ( n200 & ~n2118 ) | ( n200 & n2119 ) | ( ~n2118 & n2119 ) ;
  assign n2121 = ~n200 & n2120 ;
  assign n2122 = ( n97 & ~n323 ) | ( n97 & n2121 ) | ( ~n323 & n2121 ) ;
  assign n2123 = ~n97 & n2122 ;
  assign n2124 = ~n355 & n2123 ;
  assign n2141 = ( n693 & ~n2140 ) | ( n693 & n1762 ) | ( ~n2140 & n1762 ) ;
  assign n2142 = ( n2140 & ~n130 ) | ( n2140 & n2141 ) | ( ~n130 & n2141 ) ;
  assign n2143 = n130 | n2142 ;
  assign n2144 = ( n553 & ~n2143 ) | ( n553 & n646 ) | ( ~n2143 & n646 ) ;
  assign n2145 = ~n553 & n2144 ;
  assign n2146 = ( n2124 & ~n2145 ) | ( n2124 & n2138 ) | ( ~n2145 & n2138 ) ;
  assign n2147 = ( n446 & ~n2146 ) | ( n446 & n2124 ) | ( ~n2146 & n2124 ) ;
  assign n2148 = ~n446 & n2147 ;
  assign n2149 = ( n827 & ~n555 ) | ( n827 & n2148 ) | ( ~n555 & n2148 ) ;
  assign n2150 = ~n827 & n2149 ;
  assign n2186 = ( n2113 & n2150 ) | ( n2113 & n2184 ) | ( n2150 & n2184 ) ;
  assign n2185 = ( n2150 & ~n2113 ) | ( n2150 & n2184 ) | ( ~n2113 & n2184 ) ;
  assign n2187 = ( n2113 & ~n2186 ) | ( n2113 & n2185 ) | ( ~n2186 & n2185 ) ;
  assign n2195 = ( n2187 & ~n2194 ) | ( n2187 & 1'b0 ) | ( ~n2194 & 1'b0 ) ;
  assign n2201 = ~n1896 & n2200 ;
  assign n2205 = ~n2203 & n2204 ;
  assign n2206 = n2201 | n2205 ;
  assign n2207 = n2195 | n2206 ;
  assign n2209 = ( n1896 & n2203 ) | ( n1896 & n2208 ) | ( n2203 & n2208 ) ;
  assign n2210 = ( n2203 & ~n2187 ) | ( n2203 & n2209 ) | ( ~n2187 & n2209 ) ;
  assign n2211 = ( n2187 & ~n2209 ) | ( n2187 & n2203 ) | ( ~n2209 & n2203 ) ;
  assign n2212 = ( n2210 & ~n2203 ) | ( n2210 & n2211 ) | ( ~n2203 & n2211 ) ;
  assign n2214 = ( n2212 & ~n2207 ) | ( n2212 & n2213 ) | ( ~n2207 & n2213 ) ;
  assign n2215 = ~n2213 & n2214 ;
  assign n2216 = ( n2207 & ~n248 ) | ( n2207 & n2215 ) | ( ~n248 & n2215 ) ;
  assign n2217 = ( n248 & ~n2207 ) | ( n248 & n2215 ) | ( ~n2207 & n2215 ) ;
  assign n2218 = ( n2216 & ~n2215 ) | ( n2216 & n2217 ) | ( ~n2215 & n2217 ) ;
  assign n2306 = ( n2067 & ~n2305 ) | ( n2067 & n2218 ) | ( ~n2305 & n2218 ) ;
  assign n2307 = ( n2084 & ~n2090 ) | ( n2084 & n2094 ) | ( ~n2090 & n2094 ) ;
  assign n2314 = ~n788 & n856 ;
  assign n2315 = ( n709 & ~n2314 ) | ( n709 & n2084 ) | ( ~n2314 & n2084 ) ;
  assign n2316 = ( n709 & ~n2084 ) | ( n709 & n2314 ) | ( ~n2084 & n2314 ) ;
  assign n2317 = ( n2315 & ~n709 ) | ( n2315 & n2316 ) | ( ~n709 & n2316 ) ;
  assign n2309 = n524 &  n789 ;
  assign n2308 = n524 | n796 ;
  assign n2310 = ( n744 & ~n2309 ) | ( n744 & n2308 ) | ( ~n2309 & n2308 ) ;
  assign n2312 = n540 | n801 ;
  assign n2311 = ( n540 & ~n799 ) | ( n540 & 1'b0 ) | ( ~n799 & 1'b0 ) ;
  assign n2313 = ( n2310 & ~n2312 ) | ( n2310 & n2311 ) | ( ~n2312 & n2311 ) ;
  assign n2318 = ( n2307 & ~n2317 ) | ( n2307 & n2313 ) | ( ~n2317 & n2313 ) ;
  assign n2319 = ( n2307 & ~n2313 ) | ( n2307 & n2317 ) | ( ~n2313 & n2317 ) ;
  assign n2320 = ( n2318 & ~n2307 ) | ( n2318 & n2319 ) | ( ~n2307 & n2319 ) ;
  assign n2321 = ( n2100 & ~n2110 ) | ( n2100 & n2105 ) | ( ~n2110 & n2105 ) ;
  assign n2322 = ( n2099 & n2320 ) | ( n2099 & n2321 ) | ( n2320 & n2321 ) ;
  assign n2323 = ( n2099 & ~n2320 ) | ( n2099 & n2321 ) | ( ~n2320 & n2321 ) ;
  assign n2324 = ( n2320 & ~n2322 ) | ( n2320 & n2323 ) | ( ~n2322 & n2323 ) ;
  assign n2325 = n119 | n814 ;
  assign n2326 = ( n692 & ~n448 ) | ( n692 & n2325 ) | ( ~n448 & n2325 ) ;
  assign n2327 = n448 | n2326 ;
  assign n2328 = ( n358 & ~n637 ) | ( n358 & n2327 ) | ( ~n637 & n2327 ) ;
  assign n2329 = n637 | n2328 ;
  assign n2330 = ( n301 & ~n607 ) | ( n301 & n2329 ) | ( ~n607 & n2329 ) ;
  assign n2331 = n607 | n2330 ;
  assign n2332 = ( n902 & ~n647 ) | ( n902 & n2331 ) | ( ~n647 & n2331 ) ;
  assign n2333 = n647 | n2332 ;
  assign n2334 = ( n723 & ~n353 ) | ( n723 & n2333 ) | ( ~n353 & n2333 ) ;
  assign n2335 = n353 | n2334 ;
  assign n2336 = ( n211 & ~n142 ) | ( n211 & n2335 ) | ( ~n142 & n2335 ) ;
  assign n2337 = n142 | n2336 ;
  assign n2338 = ( n2113 & ~n2184 ) | ( n2113 & n2150 ) | ( ~n2184 & n2150 ) ;
  assign n2340 = ( n2324 & n2337 ) | ( n2324 & n2338 ) | ( n2337 & n2338 ) ;
  assign n2339 = ( n2337 & ~n2324 ) | ( n2337 & n2338 ) | ( ~n2324 & n2338 ) ;
  assign n2341 = ( n2324 & ~n2340 ) | ( n2324 & n2339 ) | ( ~n2340 & n2339 ) ;
  assign n2342 = ( n2187 & ~n2341 ) | ( n2187 & n2210 ) | ( ~n2341 & n2210 ) ;
  assign n2343 = ( n2187 & ~n2210 ) | ( n2187 & n2341 ) | ( ~n2210 & n2341 ) ;
  assign n2344 = ( n2342 & ~n2187 ) | ( n2342 & n2343 ) | ( ~n2187 & n2343 ) ;
  assign n2350 = n2344 | n2213 ;
  assign n2345 = ( n2200 & ~n2203 ) | ( n2200 & 1'b0 ) | ( ~n2203 & 1'b0 ) ;
  assign n2346 = n2187 &  n2204 ;
  assign n2347 = n2345 | n2346 ;
  assign n2348 = ~n2194 & n2341 ;
  assign n2349 = ( n2194 & ~n2347 ) | ( n2194 & n2348 ) | ( ~n2347 & n2348 ) ;
  assign n2351 = ( n2213 & ~n2350 ) | ( n2213 & n2349 ) | ( ~n2350 & n2349 ) ;
  assign n2353 = ( x8 & n245 ) | ( x8 & n2351 ) | ( n245 & n2351 ) ;
  assign n2352 = ( x8 & ~n2351 ) | ( x8 & n245 ) | ( ~n2351 & n245 ) ;
  assign n2354 = ( n2351 & ~n2353 ) | ( n2351 & n2352 ) | ( ~n2353 & n2352 ) ;
  assign n2355 = ( n2065 & ~n2306 ) | ( n2065 & n2354 ) | ( ~n2306 & n2354 ) ;
  assign n2356 = ( n2065 & ~n2354 ) | ( n2065 & n2306 ) | ( ~n2354 & n2306 ) ;
  assign n2357 = ( n2355 & ~n2065 ) | ( n2355 & n2356 ) | ( ~n2065 & n2356 ) ;
  assign n2482 = ( n2218 & ~n2067 ) | ( n2218 & n2305 ) | ( ~n2067 & n2305 ) ;
  assign n2483 = ( n2306 & ~n2218 ) | ( n2306 & n2482 ) | ( ~n2218 & n2482 ) ;
  assign n2359 = ( x5 & n1074 ) | ( x5 & n1121 ) | ( n1074 & n1121 ) ;
  assign n2358 = ( x5 & ~n1121 ) | ( x5 & n1074 ) | ( ~n1121 & n1074 ) ;
  assign n2360 = ( n1121 & ~n2359 ) | ( n1121 & n2358 ) | ( ~n2359 & n2358 ) ;
  assign n2361 = ( x1 & ~x0 ) | ( x1 & x22 ) | ( ~x0 & x22 ) ;
  assign n2362 = x0 | n2361 ;
  assign n2363 = ( x2 & ~x22 ) | ( x2 & n2362 ) | ( ~x22 & n2362 ) ;
  assign n2364 = ( x22 & ~x2 ) | ( x22 & n2362 ) | ( ~x2 & n2362 ) ;
  assign n2365 = ( n2362 & ~n2363 ) | ( n2362 & ~n2364 ) | ( ~n2363 & ~n2364 ) ;
  assign n2366 = ( x3 & n1172 ) | ( x3 & n2365 ) | ( n1172 & n2365 ) ;
  assign n2367 = ( x3 & ~n2365 ) | ( x3 & n1172 ) | ( ~n2365 & n1172 ) ;
  assign n2368 = ( n2365 & ~n2366 ) | ( n2365 & n2367 ) | ( ~n2366 & n2367 ) ;
  assign n2369 = n2360 | n2368 ;
  assign n2456 = ( x4 & n1118 ) | ( x4 & n1175 ) | ( n1118 & n1175 ) ;
  assign n2455 = ( x4 & ~n1175 ) | ( x4 & n1118 ) | ( ~n1175 & n1118 ) ;
  assign n2457 = ( n1175 & ~n2456 ) | ( n1175 & n2455 ) | ( ~n2456 & n2455 ) ;
  assign n2458 = n2360 &  n2368 ;
  assign n2459 = ~n2457 & n2458 ;
  assign n2484 = ~n2341 & n2459 ;
  assign n2406 = n226 | n690 ;
  assign n2407 = ( n723 & ~n612 ) | ( n723 & n2406 ) | ( ~n612 & n2406 ) ;
  assign n2408 = n612 | n2407 ;
  assign n2409 = n487 | n2408 ;
  assign n2410 = ( n403 & ~n311 ) | ( n403 & n2409 ) | ( ~n311 & n2409 ) ;
  assign n2411 = n311 | n2410 ;
  assign n2412 = ( n192 & ~n141 ) | ( n192 & n2411 ) | ( ~n141 & n2411 ) ;
  assign n2413 = n141 | n2412 ;
  assign n2414 = ( n180 & ~n164 ) | ( n180 & n2413 ) | ( ~n164 & n2413 ) ;
  assign n2415 = n164 | n2414 ;
  assign n2416 = ( n355 & ~n468 ) | ( n355 & n2415 ) | ( ~n468 & n2415 ) ;
  assign n2417 = n468 | n2416 ;
  assign n2418 = n127 | n828 ;
  assign n2419 = ( n417 & ~n747 ) | ( n417 & n2418 ) | ( ~n747 & n2418 ) ;
  assign n2420 = n747 | n2419 ;
  assign n2421 = ( n1875 & n2165 ) | ( n1875 & n2420 ) | ( n2165 & n2420 ) ;
  assign n2422 = ( n1875 & ~n2421 ) | ( n1875 & 1'b0 ) | ( ~n2421 & 1'b0 ) ;
  assign n2423 = ( n2417 & ~n2126 ) | ( n2417 & n2422 ) | ( ~n2126 & n2422 ) ;
  assign n2424 = ( n315 & ~n2417 ) | ( n315 & n2423 ) | ( ~n2417 & n2423 ) ;
  assign n2425 = ~n315 & n2424 ;
  assign n2426 = ( n152 & ~n201 ) | ( n152 & n2425 ) | ( ~n201 & n2425 ) ;
  assign n2427 = ~n152 & n2426 ;
  assign n2428 = ( n261 & ~n354 ) | ( n261 & n2427 ) | ( ~n354 & n2427 ) ;
  assign n2429 = ~n261 & n2428 ;
  assign n2430 = ~n189 & n2429 ;
  assign n2434 = ( n2324 & ~n2338 ) | ( n2324 & n2337 ) | ( ~n2338 & n2337 ) ;
  assign n2393 = n524 | n788 ;
  assign n2389 = n540 | n744 ;
  assign n2390 = ( n744 & n789 ) | ( n744 & n2389 ) | ( n789 & n2389 ) ;
  assign n2391 = ( n744 & ~n796 ) | ( n744 & n2389 ) | ( ~n796 & n2389 ) ;
  assign n2392 = ( n789 & ~n2390 ) | ( n789 & n2391 ) | ( ~n2390 & n2391 ) ;
  assign n2394 = ( n2315 & ~n2393 ) | ( n2315 & n2392 ) | ( ~n2393 & n2392 ) ;
  assign n2399 = ( n2392 & ~n2315 ) | ( n2392 & n2393 ) | ( ~n2315 & n2393 ) ;
  assign n2400 = ( n2394 & ~n2392 ) | ( n2394 & n2399 ) | ( ~n2392 & n2399 ) ;
  assign n2398 = ( n2307 & n2313 ) | ( n2307 & n2317 ) | ( n2313 & n2317 ) ;
  assign n2401 = ( n2099 & ~n2321 ) | ( n2099 & n2320 ) | ( ~n2321 & n2320 ) ;
  assign n2431 = ( n2400 & ~n2398 ) | ( n2400 & n2401 ) | ( ~n2398 & n2401 ) ;
  assign n2432 = ( n2398 & ~n2401 ) | ( n2398 & n2400 ) | ( ~n2401 & n2400 ) ;
  assign n2433 = ( n2431 & ~n2400 ) | ( n2431 & n2432 ) | ( ~n2400 & n2432 ) ;
  assign n2435 = ( n2430 & ~n2434 ) | ( n2430 & n2433 ) | ( ~n2434 & n2433 ) ;
  assign n2460 = ( n2433 & ~n2430 ) | ( n2433 & n2434 ) | ( ~n2430 & n2434 ) ;
  assign n2461 = ( n2435 & ~n2433 ) | ( n2435 & n2460 ) | ( ~n2433 & n2460 ) ;
  assign n2465 = n2368 &  n2457 ;
  assign n2485 = n2461 &  n2465 ;
  assign n2486 = n2484 | n2485 ;
  assign n2395 = ( n742 & ~n788 ) | ( n742 & n1951 ) | ( ~n788 & n1951 ) ;
  assign n2396 = ( n742 & n788 ) | ( n742 & n1951 ) | ( n788 & n1951 ) ;
  assign n2397 = ( n2395 & ~n2396 ) | ( n2395 & 1'b0 ) | ( ~n2396 & 1'b0 ) ;
  assign n2402 = ( n2398 & n2400 ) | ( n2398 & n2401 ) | ( n2400 & n2401 ) ;
  assign n2404 = ( n2394 & n2397 ) | ( n2394 & n2402 ) | ( n2397 & n2402 ) ;
  assign n2403 = ( n2397 & ~n2394 ) | ( n2397 & n2402 ) | ( ~n2394 & n2402 ) ;
  assign n2405 = ( n2394 & ~n2404 ) | ( n2394 & n2403 ) | ( ~n2404 & n2403 ) ;
  assign n2373 = ( n162 & ~n827 ) | ( n162 & n310 ) | ( ~n827 & n310 ) ;
  assign n2374 = ( n827 & ~n309 ) | ( n827 & n2373 ) | ( ~n309 & n2373 ) ;
  assign n2375 = n309 | n2374 ;
  assign n2376 = n501 | n2375 ;
  assign n231 = n229 | n230 ;
  assign n2377 = ~n124 & n378 ;
  assign n2378 = ( n672 & ~n1734 ) | ( n672 & n2377 ) | ( ~n1734 & n2377 ) ;
  assign n2379 = ( n231 & ~n672 ) | ( n231 & n2378 ) | ( ~n672 & n2378 ) ;
  assign n2380 = ~n231 & n2379 ;
  assign n2381 = ( n2376 & ~n611 ) | ( n2376 & n2380 ) | ( ~n611 & n2380 ) ;
  assign n2382 = ~n2376 & n2381 ;
  assign n2370 = ( n276 & ~n142 ) | ( n276 & n2128 ) | ( ~n142 & n2128 ) ;
  assign n2371 = n142 | n2370 ;
  assign n2372 = n612 | n2371 ;
  assign n2383 = ( n496 & ~n2382 ) | ( n496 & n2372 ) | ( ~n2382 & n2372 ) ;
  assign n2384 = ( n496 & ~n2383 ) | ( n496 & 1'b0 ) | ( ~n2383 & 1'b0 ) ;
  assign n2385 = ( n452 & ~n911 ) | ( n452 & n2384 ) | ( ~n911 & n2384 ) ;
  assign n2386 = ( n182 & ~n452 ) | ( n182 & n2385 ) | ( ~n452 & n2385 ) ;
  assign n2387 = ~n182 & n2386 ;
  assign n2388 = ~n110 & n2387 ;
  assign n2436 = ( n2388 & n2405 ) | ( n2388 & n2435 ) | ( n2405 & n2435 ) ;
  assign n2463 = ( n2388 & ~n2405 ) | ( n2388 & n2435 ) | ( ~n2405 & n2435 ) ;
  assign n2464 = ( n2405 & ~n2436 ) | ( n2405 & n2463 ) | ( ~n2436 & n2463 ) ;
  assign n2487 = ~n2369 & n2464 ;
  assign n2488 = ( n2369 & ~n2486 ) | ( n2369 & n2487 ) | ( ~n2486 & n2487 ) ;
  assign n2470 = ( n2360 & ~n2368 ) | ( n2360 & 1'b0 ) | ( ~n2368 & 1'b0 ) ;
  assign n2471 = ( n2210 & ~n2187 ) | ( n2210 & n2341 ) | ( ~n2187 & n2341 ) ;
  assign n2472 = ( n2341 & ~n2461 ) | ( n2341 & n2471 ) | ( ~n2461 & n2471 ) ;
  assign n2473 = ( n2464 & ~n2461 ) | ( n2464 & n2472 ) | ( ~n2461 & n2472 ) ;
  assign n2489 = ( n2461 & ~n2472 ) | ( n2461 & n2464 ) | ( ~n2472 & n2464 ) ;
  assign n2490 = ( n2473 & ~n2464 ) | ( n2473 & n2489 ) | ( ~n2464 & n2489 ) ;
  assign n2491 = n2470 &  n2490 ;
  assign n2492 = ( n2488 & ~n2491 ) | ( n2488 & 1'b0 ) | ( ~n2491 & 1'b0 ) ;
  assign n2493 = ( x5 & ~n1074 ) | ( x5 & n2492 ) | ( ~n1074 & n2492 ) ;
  assign n2494 = ( x5 & ~n2492 ) | ( x5 & n1074 ) | ( ~n2492 & n1074 ) ;
  assign n2495 = ( n2493 & ~x5 ) | ( n2493 & n2494 ) | ( ~x5 & n2494 ) ;
  assign n2496 = ( n2231 & ~n2304 ) | ( n2231 & n2233 ) | ( ~n2304 & n2233 ) ;
  assign n2497 = ( n2233 & ~n2231 ) | ( n2233 & n2304 ) | ( ~n2231 & n2304 ) ;
  assign n2498 = ( n2496 & ~n2233 ) | ( n2496 & n2497 ) | ( ~n2233 & n2497 ) ;
  assign n2504 = ( n2341 & ~n2471 ) | ( n2341 & n2461 ) | ( ~n2471 & n2461 ) ;
  assign n2505 = ( n2472 & ~n2341 ) | ( n2472 & n2504 ) | ( ~n2341 & n2504 ) ;
  assign n2499 = n2369 &  n2461 ;
  assign n2500 = n2187 &  n2459 ;
  assign n2501 = ~n2341 & n2465 ;
  assign n2502 = n2500 | n2501 ;
  assign n2503 = ( n2461 & ~n2499 ) | ( n2461 & n2502 ) | ( ~n2499 & n2502 ) ;
  assign n2506 = ( n2470 & ~n2505 ) | ( n2470 & n2503 ) | ( ~n2505 & n2503 ) ;
  assign n2507 = ( n2470 & ~n2506 ) | ( n2470 & 1'b0 ) | ( ~n2506 & 1'b0 ) ;
  assign n2508 = ( n1077 & n2503 ) | ( n1077 & n2507 ) | ( n2503 & n2507 ) ;
  assign n2509 = ( n1077 & ~n2507 ) | ( n1077 & n2503 ) | ( ~n2507 & n2503 ) ;
  assign n2510 = ( n2507 & ~n2508 ) | ( n2507 & n2509 ) | ( ~n2508 & n2509 ) ;
  assign n2511 = ( n2235 & ~n2303 ) | ( n2235 & n2245 ) | ( ~n2303 & n2245 ) ;
  assign n2512 = ( n2245 & ~n2235 ) | ( n2245 & n2303 ) | ( ~n2235 & n2303 ) ;
  assign n2513 = ( n2511 & ~n2245 ) | ( n2511 & n2512 ) | ( ~n2245 & n2512 ) ;
  assign n2514 = ~n2203 & n2459 ;
  assign n2515 = n2187 &  n2465 ;
  assign n2516 = n2514 | n2515 ;
  assign n2517 = ~n2341 & n2369 ;
  assign n2518 = ( n2341 & ~n2516 ) | ( n2341 & n2517 ) | ( ~n2516 & n2517 ) ;
  assign n2519 = ( n2470 & ~n2344 ) | ( n2470 & n2518 ) | ( ~n2344 & n2518 ) ;
  assign n2520 = n2344 &  n2519 ;
  assign n2521 = ( n1077 & ~n2518 ) | ( n1077 & n2520 ) | ( ~n2518 & n2520 ) ;
  assign n2522 = ( n2518 & ~n1077 ) | ( n2518 & n2520 ) | ( ~n1077 & n2520 ) ;
  assign n2523 = ( n2521 & ~n2520 ) | ( n2521 & n2522 ) | ( ~n2520 & n2522 ) ;
  assign n2530 = n2187 &  n2369 ;
  assign n2527 = ~n1896 & n2459 ;
  assign n2528 = ~n2203 & n2465 ;
  assign n2529 = n2527 | n2528 ;
  assign n2531 = ( n2187 & ~n2530 ) | ( n2187 & n2529 ) | ( ~n2530 & n2529 ) ;
  assign n2532 = ( n2212 & ~n2470 ) | ( n2212 & n2531 ) | ( ~n2470 & n2531 ) ;
  assign n2533 = ( n2212 & ~n2532 ) | ( n2212 & 1'b0 ) | ( ~n2532 & 1'b0 ) ;
  assign n2534 = ( n1077 & n2531 ) | ( n1077 & n2533 ) | ( n2531 & n2533 ) ;
  assign n2535 = ( n1077 & ~n2533 ) | ( n1077 & n2531 ) | ( ~n2533 & n2531 ) ;
  assign n2536 = ( n2533 & ~n2534 ) | ( n2533 & n2535 ) | ( ~n2534 & n2535 ) ;
  assign n2524 = ( n2255 & n2257 ) | ( n2255 & n2302 ) | ( n2257 & n2302 ) ;
  assign n2525 = ( n2255 & ~n2302 ) | ( n2255 & n2257 ) | ( ~n2302 & n2257 ) ;
  assign n2526 = ( n2302 & ~n2524 ) | ( n2302 & n2525 ) | ( ~n2524 & n2525 ) ;
  assign n2537 = ~n1910 & n2459 ;
  assign n2538 = ~n1896 & n2465 ;
  assign n2539 = n2537 | n2538 ;
  assign n2540 = ~n2203 & n2369 ;
  assign n2541 = ( n2203 & ~n2539 ) | ( n2203 & n2540 ) | ( ~n2539 & n2540 ) ;
  assign n2542 = ~n2226 & n2470 ;
  assign n2543 = ( n2541 & ~n2542 ) | ( n2541 & 1'b0 ) | ( ~n2542 & 1'b0 ) ;
  assign n2544 = ( x5 & ~n1074 ) | ( x5 & n2543 ) | ( ~n1074 & n2543 ) ;
  assign n2545 = ( x5 & ~n2543 ) | ( x5 & n1074 ) | ( ~n2543 & n1074 ) ;
  assign n2546 = ( n2544 & ~x5 ) | ( n2544 & n2545 ) | ( ~x5 & n2545 ) ;
  assign n2547 = ( n2271 & ~n2261 ) | ( n2271 & n2301 ) | ( ~n2261 & n2301 ) ;
  assign n2548 = ( n2302 & ~n2271 ) | ( n2302 & n2547 ) | ( ~n2271 & n2547 ) ;
  assign n2550 = ( n2010 & n2290 ) | ( n2010 & n2300 ) | ( n2290 & n2300 ) ;
  assign n2549 = ( n2010 & ~n2290 ) | ( n2010 & n2300 ) | ( ~n2290 & n2300 ) ;
  assign n2551 = ( n2290 & ~n2550 ) | ( n2290 & n2549 ) | ( ~n2550 & n2549 ) ;
  assign n2552 = ~n1901 & n2459 ;
  assign n2553 = ~n1910 & n2465 ;
  assign n2554 = n2552 | n2553 ;
  assign n2555 = ~n1896 & n2369 ;
  assign n2556 = ( n1896 & ~n2554 ) | ( n1896 & n2555 ) | ( ~n2554 & n2555 ) ;
  assign n2557 = ( n1938 & n2470 ) | ( n1938 & n2556 ) | ( n2470 & n2556 ) ;
  assign n2558 = ~n1938 & n2557 ;
  assign n2559 = ( n1077 & ~n2556 ) | ( n1077 & n2558 ) | ( ~n2556 & n2558 ) ;
  assign n2560 = ( n2556 & ~n1077 ) | ( n2556 & n2558 ) | ( ~n1077 & n2558 ) ;
  assign n2561 = ( n2559 & ~n2558 ) | ( n2559 & n2560 ) | ( ~n2558 & n2560 ) ;
  assign n2562 = ~n1922 & n2459 ;
  assign n2563 = ~n1901 & n2465 ;
  assign n2564 = n2562 | n2563 ;
  assign n2565 = ~n1910 & n2369 ;
  assign n2566 = ( n1910 & ~n2564 ) | ( n1910 & n2565 ) | ( ~n2564 & n2565 ) ;
  assign n2567 = ~n2048 & n2470 ;
  assign n2568 = ( n2566 & ~n2567 ) | ( n2566 & 1'b0 ) | ( ~n2567 & 1'b0 ) ;
  assign n2569 = ( x5 & ~n1074 ) | ( x5 & n2568 ) | ( ~n1074 & n2568 ) ;
  assign n2570 = ( x5 & ~n2568 ) | ( x5 & n1074 ) | ( ~n2568 & n1074 ) ;
  assign n2571 = ( n2569 & ~x5 ) | ( n2569 & n2570 ) | ( ~x5 & n2570 ) ;
  assign n2572 = ~n2279 & n2289 ;
  assign n2573 = n2290 | n2572 ;
  assign n2574 = ( n248 & ~n2277 ) | ( n248 & 1'b0 ) | ( ~n2277 & 1'b0 ) ;
  assign n2575 = n2276 &  n2574 ;
  assign n2576 = n2276 | n2574 ;
  assign n2577 = ~n2575 & n2576 ;
  assign n2583 = n2004 | n2470 ;
  assign n2578 = ~n1924 & n2459 ;
  assign n2579 = ~n1922 & n2465 ;
  assign n2580 = n2578 | n2579 ;
  assign n2581 = ~n1901 & n2369 ;
  assign n2582 = ( n1901 & ~n2580 ) | ( n1901 & n2581 ) | ( ~n2580 & n2581 ) ;
  assign n2584 = ( n2004 & ~n2583 ) | ( n2004 & n2582 ) | ( ~n2583 & n2582 ) ;
  assign n2586 = ( x5 & n1074 ) | ( x5 & n2584 ) | ( n1074 & n2584 ) ;
  assign n2585 = ( x5 & ~n2584 ) | ( x5 & n1074 ) | ( ~n2584 & n1074 ) ;
  assign n2587 = ( n2584 & ~n2586 ) | ( n2584 & n2585 ) | ( ~n2586 & n2585 ) ;
  assign n2589 = ~n1928 & n2465 ;
  assign n2590 = ( n1930 & ~n2369 ) | ( n1930 & 1'b0 ) | ( ~n2369 & 1'b0 ) ;
  assign n2591 = n2589 | n2590 ;
  assign n2592 = n1957 | n2470 ;
  assign n2593 = ( n2591 & ~n1957 ) | ( n2591 & n2592 ) | ( ~n1957 & n2592 ) ;
  assign n2588 = n1928 | n2368 ;
  assign n2594 = ( n1077 & ~n2593 ) | ( n1077 & n2588 ) | ( ~n2593 & n2588 ) ;
  assign n2595 = ~n1077 & n2594 ;
  assign n2596 = ~n1928 & n2459 ;
  assign n2597 = n1930 &  n2465 ;
  assign n2598 = n2596 | n2597 ;
  assign n2599 = ~n1924 & n2369 ;
  assign n2600 = ( n1924 & ~n2598 ) | ( n1924 & n2599 ) | ( ~n2598 & n2599 ) ;
  assign n2601 = ( n1964 & n2470 ) | ( n1964 & n2600 ) | ( n2470 & n2600 ) ;
  assign n2602 = ~n1964 & n2601 ;
  assign n2603 = ( n1077 & ~n2600 ) | ( n1077 & n2602 ) | ( ~n2600 & n2602 ) ;
  assign n2604 = ( n2600 & ~n1077 ) | ( n2600 & n2602 ) | ( ~n1077 & n2602 ) ;
  assign n2605 = ( n2603 & ~n2602 ) | ( n2603 & n2604 ) | ( ~n2602 & n2604 ) ;
  assign n2606 = n2595 &  n2605 ;
  assign n2607 = ~n1924 & n2465 ;
  assign n2608 = n1930 &  n2459 ;
  assign n2609 = n2607 | n2608 ;
  assign n2610 = ~n1922 & n2369 ;
  assign n2611 = ( n1922 & ~n2609 ) | ( n1922 & n2610 ) | ( ~n2609 & n2610 ) ;
  assign n2612 = n1985 &  n2470 ;
  assign n2613 = ( n2611 & ~n2612 ) | ( n2611 & 1'b0 ) | ( ~n2612 & 1'b0 ) ;
  assign n2614 = ( x5 & ~n1074 ) | ( x5 & n2613 ) | ( ~n1074 & n2613 ) ;
  assign n2615 = ( x5 & ~n2613 ) | ( x5 & n1074 ) | ( ~n2613 & n1074 ) ;
  assign n2616 = ( n2614 & ~x5 ) | ( n2614 & n2615 ) | ( ~x5 & n2615 ) ;
  assign n2617 = ( n2277 & ~n2606 ) | ( n2277 & n2616 ) | ( ~n2606 & n2616 ) ;
  assign n2618 = ( n2577 & n2587 ) | ( n2577 & n2617 ) | ( n2587 & n2617 ) ;
  assign n2619 = ( n2571 & n2573 ) | ( n2571 & n2618 ) | ( n2573 & n2618 ) ;
  assign n2620 = ( n2551 & ~n2561 ) | ( n2551 & n2619 ) | ( ~n2561 & n2619 ) ;
  assign n2621 = ( n2546 & ~n2548 ) | ( n2546 & n2620 ) | ( ~n2548 & n2620 ) ;
  assign n2622 = ( n2536 & ~n2526 ) | ( n2536 & n2621 ) | ( ~n2526 & n2621 ) ;
  assign n2623 = ( n2513 & ~n2523 ) | ( n2513 & n2622 ) | ( ~n2523 & n2622 ) ;
  assign n2624 = ( n2498 & n2510 ) | ( n2498 & n2623 ) | ( n2510 & n2623 ) ;
  assign n2625 = ( n2483 & n2495 ) | ( n2483 & n2624 ) | ( n2495 & n2624 ) ;
  assign n2462 = n2459 &  n2461 ;
  assign n2466 = ~n2464 & n2465 ;
  assign n2467 = n2462 | n2466 ;
  assign n2437 = ( n104 & ~n614 ) | ( n104 & n816 ) | ( ~n614 & n816 ) ;
  assign n2438 = ( n200 & ~n149 ) | ( n200 & n2437 ) | ( ~n149 & n2437 ) ;
  assign n2439 = n149 | n2438 ;
  assign n2440 = n278 | n2439 ;
  assign n2441 = n693 | n890 ;
  assign n2442 = ( n1201 & n1699 ) | ( n1201 & n2441 ) | ( n1699 & n2441 ) ;
  assign n2443 = ( n1201 & ~n2442 ) | ( n1201 & 1'b0 ) | ( ~n2442 & 1'b0 ) ;
  assign n2444 = ( n654 & ~n2440 ) | ( n654 & n2443 ) | ( ~n2440 & n2443 ) ;
  assign n2445 = ~n654 & n2444 ;
  assign n2446 = ( n123 & ~n467 ) | ( n123 & n2445 ) | ( ~n467 & n2445 ) ;
  assign n2447 = ~n123 & n2446 ;
  assign n2448 = ( n437 & ~n499 ) | ( n437 & n2447 ) | ( ~n499 & n2447 ) ;
  assign n2449 = ~n437 & n2448 ;
  assign n2450 = ( n197 & ~n555 ) | ( n197 & n2449 ) | ( ~n555 & n2449 ) ;
  assign n2451 = ~n197 & n2450 ;
  assign n2452 = n2436 &  n2451 ;
  assign n2453 = n2436 | n2451 ;
  assign n2454 = ~n2452 & n2453 ;
  assign n2468 = ~n2369 & n2454 ;
  assign n2469 = ( n2369 & ~n2467 ) | ( n2369 & n2468 ) | ( ~n2467 & n2468 ) ;
  assign n2474 = ( n2464 & ~n2454 ) | ( n2464 & n2473 ) | ( ~n2454 & n2473 ) ;
  assign n2475 = ( n2454 & ~n2473 ) | ( n2454 & n2464 ) | ( ~n2473 & n2464 ) ;
  assign n2476 = ( n2474 & ~n2464 ) | ( n2474 & n2475 ) | ( ~n2464 & n2475 ) ;
  assign n2477 = ( n2469 & n2470 ) | ( n2469 & n2476 ) | ( n2470 & n2476 ) ;
  assign n2478 = ~n2476 & n2477 ;
  assign n2479 = ( n1077 & ~n2469 ) | ( n1077 & n2478 ) | ( ~n2469 & n2478 ) ;
  assign n2480 = ( n2469 & ~n1077 ) | ( n2469 & n2478 ) | ( ~n1077 & n2478 ) ;
  assign n2481 = ( n2479 & ~n2478 ) | ( n2479 & n2480 ) | ( ~n2478 & n2480 ) ;
  assign n2626 = ( n2357 & ~n2625 ) | ( n2357 & n2481 ) | ( ~n2625 & n2481 ) ;
  assign n2627 = ( n2357 & ~n2481 ) | ( n2357 & n2625 ) | ( ~n2481 & n2625 ) ;
  assign n2628 = ( n2626 & ~n2357 ) | ( n2626 & n2627 ) | ( ~n2357 & n2627 ) ;
  assign n2629 = ( x0 & x1 ) | ( x0 & x2 ) | ( x1 & x2 ) ;
  assign n2630 = ( x1 & ~x0 ) | ( x1 & x2 ) | ( ~x0 & x2 ) ;
  assign n2631 = ( n2629 & ~n2630 ) | ( n2629 & 1'b0 ) | ( ~n2630 & 1'b0 ) ;
  assign n2632 = ( n495 & ~n831 ) | ( n495 & 1'b0 ) | ( ~n831 & 1'b0 ) ;
  assign n2633 = ~n699 & n2632 ;
  assign n2634 = ( n1693 & ~n2633 ) | ( n1693 & n2118 ) | ( ~n2633 & n2118 ) ;
  assign n2635 = ( n776 & ~n1693 ) | ( n776 & n2634 ) | ( ~n1693 & n2634 ) ;
  assign n2636 = ( n776 & ~n2635 ) | ( n776 & 1'b0 ) | ( ~n2635 & 1'b0 ) ;
  assign n2637 = ( n303 & ~n1798 ) | ( n303 & n2636 ) | ( ~n1798 & n2636 ) ;
  assign n2638 = ~n303 & n2637 ;
  assign n2639 = ( n353 & ~n354 ) | ( n353 & n2638 ) | ( ~n354 & n2638 ) ;
  assign n2640 = ~n353 & n2639 ;
  assign n2641 = ( n186 & ~n230 ) | ( n186 & n2640 ) | ( ~n230 & n2640 ) ;
  assign n2642 = ~n186 & n2641 ;
  assign n2643 = ~n211 & n2642 ;
  assign n183 = ( n181 & ~n180 ) | ( n181 & n182 ) | ( ~n180 & n182 ) ;
  assign n184 = n180 | n183 ;
  assign n2658 = n369 | n1736 ;
  assign n2659 = ( n410 & ~n130 ) | ( n410 & n2658 ) | ( ~n130 & n2658 ) ;
  assign n2660 = n130 | n2659 ;
  assign n171 = ( n94 & ~n102 ) | ( n94 & 1'b0 ) | ( ~n102 & 1'b0 ) ;
  assign n170 = n167 | n169 ;
  assign n172 = ( n94 & ~n171 ) | ( n94 & n170 ) | ( ~n171 & n170 ) ;
  assign n173 = ( n165 & ~n164 ) | ( n165 & n172 ) | ( ~n164 & n172 ) ;
  assign n174 = n164 | n173 ;
  assign n2644 = n422 | n828 ;
  assign n2645 = n612 | n2644 ;
  assign n2646 = ( n2126 & ~n174 ) | ( n2126 & n2645 ) | ( ~n174 & n2645 ) ;
  assign n2647 = n174 | n2646 ;
  assign n2648 = ( n381 & ~n311 ) | ( n381 & n2647 ) | ( ~n311 & n2647 ) ;
  assign n2649 = n311 | n2648 ;
  assign n2650 = ( n318 & n645 ) | ( n318 & n2649 ) | ( n645 & n2649 ) ;
  assign n2651 = ( n645 & ~n2650 ) | ( n645 & 1'b0 ) | ( ~n2650 & 1'b0 ) ;
  assign n2652 = ( n501 & ~n292 ) | ( n501 & n2651 ) | ( ~n292 & n2651 ) ;
  assign n2653 = ~n501 & n2652 ;
  assign n2654 = ( n85 & ~n723 ) | ( n85 & n2653 ) | ( ~n723 & n2653 ) ;
  assign n2655 = ~n85 & n2654 ;
  assign n2656 = ( n69 & ~n487 ) | ( n69 & n2655 ) | ( ~n487 & n2655 ) ;
  assign n2657 = ~n69 & n2656 ;
  assign n2661 = ( n184 & ~n2660 ) | ( n184 & n2657 ) | ( ~n2660 & n2657 ) ;
  assign n2662 = ~n184 & n2661 ;
  assign n2663 = ( n124 & ~n478 ) | ( n124 & n2662 ) | ( ~n478 & n2662 ) ;
  assign n2664 = ~n124 & n2663 ;
  assign n2665 = ( n503 & ~n200 ) | ( n503 & n2664 ) | ( ~n200 & n2664 ) ;
  assign n2666 = ~n503 & n2665 ;
  assign n2667 = ( n160 & ~n277 ) | ( n160 & n2666 ) | ( ~n277 & n2666 ) ;
  assign n2668 = ~n160 & n2667 ;
  assign n2669 = ( n595 & ~n643 ) | ( n595 & n2668 ) | ( ~n643 & n2668 ) ;
  assign n2670 = ~n595 & n2669 ;
  assign n2671 = n2452 &  n2670 ;
  assign n2672 = n2643 &  n2671 ;
  assign n2673 = n2643 | n2671 ;
  assign n2674 = ~n2672 & n2673 ;
  assign n2675 = n110 | n419 ;
  assign n2676 = n672 | n768 ;
  assign n2677 = ( n982 & ~n747 ) | ( n982 & n2676 ) | ( ~n747 & n2676 ) ;
  assign n2678 = n747 | n2677 ;
  assign n2679 = ( n781 & ~n444 ) | ( n781 & n2678 ) | ( ~n444 & n2678 ) ;
  assign n2680 = n444 | n2679 ;
  assign n2681 = ( n729 & ~n699 ) | ( n729 & n2680 ) | ( ~n699 & n2680 ) ;
  assign n2682 = n699 | n2681 ;
  assign n2683 = ( n671 & ~n2675 ) | ( n671 & n2682 ) | ( ~n2675 & n2682 ) ;
  assign n2684 = ( n2675 & ~n114 ) | ( n2675 & n2683 ) | ( ~n114 & n2683 ) ;
  assign n2685 = n114 | n2684 ;
  assign n2687 = n2672 &  n2685 ;
  assign n2686 = ~n2672 & n2685 ;
  assign n2688 = ( n2672 & ~n2687 ) | ( n2672 & n2686 ) | ( ~n2687 & n2686 ) ;
  assign n2689 = ~n2452 & n2670 ;
  assign n2690 = ( n2452 & ~n2670 ) | ( n2452 & 1'b0 ) | ( ~n2670 & 1'b0 ) ;
  assign n2691 = n2689 | n2690 ;
  assign n2692 = ( n2454 & n2464 ) | ( n2454 & n2473 ) | ( n2464 & n2473 ) ;
  assign n2693 = ( n2454 & n2691 ) | ( n2454 & n2692 ) | ( n2691 & n2692 ) ;
  assign n2694 = ( n2674 & n2691 ) | ( n2674 & n2693 ) | ( n2691 & n2693 ) ;
  assign n2695 = ( n2674 & ~n2688 ) | ( n2674 & n2694 ) | ( ~n2688 & n2694 ) ;
  assign n2696 = ( n2674 & ~n2694 ) | ( n2674 & n2688 ) | ( ~n2694 & n2688 ) ;
  assign n2697 = ( n2695 & ~n2674 ) | ( n2695 & n2696 ) | ( ~n2674 & n2696 ) ;
  assign n2708 = ~n2697 & n2631 ;
  assign n2698 = ( x0 & ~x1 ) | ( x0 & x2 ) | ( ~x1 & x2 ) ;
  assign n2699 = ( x0 & ~x2 ) | ( x0 & x1 ) | ( ~x2 & x1 ) ;
  assign n2700 = n2698 &  n2699 ;
  assign n2706 = ~n2700 & n2688 ;
  assign n2701 = ~x0 & n2698 ;
  assign n2702 = ~n2691 & n2701 ;
  assign n2703 = ~x0 & x1 ;
  assign n2704 = ~n2674 & n2703 ;
  assign n2705 = n2702 | n2704 ;
  assign n2707 = ( n2688 & ~n2706 ) | ( n2688 & n2705 ) | ( ~n2706 & n2705 ) ;
  assign n2709 = ( n2631 & ~n2708 ) | ( n2631 & n2707 ) | ( ~n2708 & n2707 ) ;
  assign n2710 = ( n2365 & ~n2709 ) | ( n2365 & 1'b0 ) | ( ~n2709 & 1'b0 ) ;
  assign n2711 = ~n2365 & n2709 ;
  assign n2712 = n2710 | n2711 ;
  assign n2713 = ( n2483 & ~n2624 ) | ( n2483 & n2495 ) | ( ~n2624 & n2495 ) ;
  assign n2714 = ( n2495 & ~n2483 ) | ( n2495 & n2624 ) | ( ~n2483 & n2624 ) ;
  assign n2715 = ( n2713 & ~n2495 ) | ( n2713 & n2714 ) | ( ~n2495 & n2714 ) ;
  assign n2716 = ~n2454 & n2701 ;
  assign n2717 = ~n2691 & n2703 ;
  assign n2718 = n2716 | n2717 ;
  assign n2719 = n2674 | n2700 ;
  assign n2720 = ( n2718 & ~n2674 ) | ( n2718 & n2719 ) | ( ~n2674 & n2719 ) ;
  assign n2721 = ( n2691 & ~n2674 ) | ( n2691 & n2693 ) | ( ~n2674 & n2693 ) ;
  assign n2722 = ( n2674 & ~n2694 ) | ( n2674 & n2721 ) | ( ~n2694 & n2721 ) ;
  assign n2723 = ( n2631 & n2720 ) | ( n2631 & n2722 ) | ( n2720 & n2722 ) ;
  assign n2724 = ( n2631 & ~n2723 ) | ( n2631 & 1'b0 ) | ( ~n2723 & 1'b0 ) ;
  assign n2725 = ( n2365 & n2720 ) | ( n2365 & n2724 ) | ( n2720 & n2724 ) ;
  assign n2726 = ( n2365 & ~n2724 ) | ( n2365 & n2720 ) | ( ~n2724 & n2720 ) ;
  assign n2727 = ( n2724 & ~n2725 ) | ( n2724 & n2726 ) | ( ~n2725 & n2726 ) ;
  assign n2728 = ~n2464 & n2701 ;
  assign n2729 = ~n2454 & n2703 ;
  assign n2730 = n2728 | n2729 ;
  assign n2731 = n2691 | n2700 ;
  assign n2732 = ( n2730 & ~n2691 ) | ( n2730 & n2731 ) | ( ~n2691 & n2731 ) ;
  assign n2733 = ( n2454 & ~n2691 ) | ( n2454 & n2692 ) | ( ~n2691 & n2692 ) ;
  assign n2734 = ( n2691 & ~n2693 ) | ( n2691 & n2733 ) | ( ~n2693 & n2733 ) ;
  assign n2735 = ( n2631 & n2732 ) | ( n2631 & n2734 ) | ( n2732 & n2734 ) ;
  assign n2736 = ( n2631 & ~n2735 ) | ( n2631 & 1'b0 ) | ( ~n2735 & 1'b0 ) ;
  assign n2737 = ( n2365 & n2732 ) | ( n2365 & n2736 ) | ( n2732 & n2736 ) ;
  assign n2738 = ( n2365 & ~n2736 ) | ( n2365 & n2732 ) | ( ~n2736 & n2732 ) ;
  assign n2739 = ( n2736 & ~n2737 ) | ( n2736 & n2738 ) | ( ~n2737 & n2738 ) ;
  assign n2740 = ( n2498 & ~n2510 ) | ( n2498 & n2623 ) | ( ~n2510 & n2623 ) ;
  assign n2741 = ( n2510 & ~n2624 ) | ( n2510 & n2740 ) | ( ~n2624 & n2740 ) ;
  assign n2742 = ~n2365 & n2631 ;
  assign n2743 = n2505 &  n2742 ;
  assign n2744 = n2344 &  n2742 ;
  assign n2745 = ( n2571 & ~n2618 ) | ( n2571 & n2573 ) | ( ~n2618 & n2573 ) ;
  assign n2746 = ( n2618 & ~n2619 ) | ( n2618 & n2745 ) | ( ~n2619 & n2745 ) ;
  assign n2747 = ~n1938 & n2742 ;
  assign n2748 = ~n2004 & n2742 ;
  assign n2749 = ( x0 & ~n1928 ) | ( x0 & 1'b0 ) | ( ~n1928 & 1'b0 ) ;
  assign n2750 = ~n1928 & n2701 ;
  assign n2751 = n1930 &  n2703 ;
  assign n2752 = n2750 | n2751 ;
  assign n2753 = n1924 | n2700 ;
  assign n2754 = ( n2752 & ~n1924 ) | ( n2752 & n2753 ) | ( ~n1924 & n2753 ) ;
  assign n2766 = n2754 | n2365 ;
  assign n2755 = ( n1956 & ~n1924 ) | ( n1956 & n2631 ) | ( ~n1924 & n2631 ) ;
  assign n2756 = ( n1956 & ~n1924 ) | ( n1956 & n2365 ) | ( ~n1924 & n2365 ) ;
  assign n2757 = ( n2755 & ~n2756 ) | ( n2755 & 1'b0 ) | ( ~n2756 & 1'b0 ) ;
  assign n2760 = ~n2700 & n1930 ;
  assign n2758 = ~n1928 & n2703 ;
  assign n2759 = n2365 | n2758 ;
  assign n2761 = ( n1930 & ~n2760 ) | ( n1930 & n2759 ) | ( ~n2760 & n2759 ) ;
  assign n2762 = ~n1928 & n1930 ;
  assign n2763 = ( n1930 & ~n1928 ) | ( n1930 & n2742 ) | ( ~n1928 & n2742 ) ;
  assign n2764 = ( n2761 & ~n2762 ) | ( n2761 & n2763 ) | ( ~n2762 & n2763 ) ;
  assign n2765 = n2757 | n2764 ;
  assign n2767 = ( n2766 & ~n2365 ) | ( n2766 & n2765 ) | ( ~n2365 & n2765 ) ;
  assign n2768 = n2749 | n2767 ;
  assign n2769 = n2588 | n2768 ;
  assign n2770 = ~n1924 & n2703 ;
  assign n2771 = n1930 &  n2701 ;
  assign n2772 = n2770 | n2771 ;
  assign n2773 = n1922 | n2700 ;
  assign n2774 = ( n2772 & ~n1922 ) | ( n2772 & n2773 ) | ( ~n1922 & n2773 ) ;
  assign n2775 = n1985 &  n2631 ;
  assign n2776 = n2774 | n2775 ;
  assign n2777 = ( n2365 & ~n2776 ) | ( n2365 & 1'b0 ) | ( ~n2776 & 1'b0 ) ;
  assign n2778 = n2588 &  n2768 ;
  assign n2779 = ( n2776 & ~n2365 ) | ( n2776 & n2778 ) | ( ~n2365 & n2778 ) ;
  assign n2780 = ( n2769 & n2777 ) | ( n2769 & n2779 ) | ( n2777 & n2779 ) ;
  assign n2781 = n1077 | n2588 ;
  assign n2782 = ( n2593 & ~n2781 ) | ( n2593 & 1'b0 ) | ( ~n2781 & 1'b0 ) ;
  assign n2783 = ~n2593 & n2781 ;
  assign n2784 = n2782 | n2783 ;
  assign n2785 = n2780 &  n2784 ;
  assign n2786 = n2748 | n2785 ;
  assign n2790 = n2700 | n1901 ;
  assign n2787 = ~n1924 & n2701 ;
  assign n2788 = ~n1922 & n2703 ;
  assign n2789 = n2787 | n2788 ;
  assign n2791 = ( n2790 & ~n1901 ) | ( n2790 & n2789 ) | ( ~n1901 & n2789 ) ;
  assign n2792 = ~n2004 & n2631 ;
  assign n2793 = n2791 | n2792 ;
  assign n2794 = n2365 &  n2793 ;
  assign n2795 = n2365 | n2791 ;
  assign n2796 = ( n2786 & ~n2794 ) | ( n2786 & n2795 ) | ( ~n2794 & n2795 ) ;
  assign n2797 = n2780 | n2784 ;
  assign n2798 = n2796 &  n2797 ;
  assign n2809 = n2595 | n2605 ;
  assign n2810 = ~n2606 & n2809 ;
  assign n2799 = ~n1922 & n2701 ;
  assign n2800 = ~n1901 & n2703 ;
  assign n2801 = n2799 | n2800 ;
  assign n2802 = n1910 | n2700 ;
  assign n2803 = ( n2801 & ~n1910 ) | ( n2801 & n2802 ) | ( ~n1910 & n2802 ) ;
  assign n2804 = ( n2048 & n2631 ) | ( n2048 & n2803 ) | ( n2631 & n2803 ) ;
  assign n2805 = ( n2631 & ~n2804 ) | ( n2631 & 1'b0 ) | ( ~n2804 & 1'b0 ) ;
  assign n2806 = ( n2365 & n2803 ) | ( n2365 & n2805 ) | ( n2803 & n2805 ) ;
  assign n2807 = ( n2365 & ~n2805 ) | ( n2365 & n2803 ) | ( ~n2805 & n2803 ) ;
  assign n2808 = ( n2805 & ~n2806 ) | ( n2805 & n2807 ) | ( ~n2806 & n2807 ) ;
  assign n2811 = ( n2798 & ~n2810 ) | ( n2798 & n2808 ) | ( ~n2810 & n2808 ) ;
  assign n2812 = ( n2606 & ~n2277 ) | ( n2606 & n2616 ) | ( ~n2277 & n2616 ) ;
  assign n2813 = ( n2617 & ~n2616 ) | ( n2617 & n2812 ) | ( ~n2616 & n2812 ) ;
  assign n2814 = ( n2811 & ~n2813 ) | ( n2811 & 1'b0 ) | ( ~n2813 & 1'b0 ) ;
  assign n2815 = n2747 | n2814 ;
  assign n2819 = n2700 | n1896 ;
  assign n2816 = ~n1901 & n2701 ;
  assign n2817 = ~n1910 & n2703 ;
  assign n2818 = n2816 | n2817 ;
  assign n2820 = ( n2819 & ~n1896 ) | ( n2819 & n2818 ) | ( ~n1896 & n2818 ) ;
  assign n2821 = ~n1938 & n2631 ;
  assign n2822 = n2820 | n2821 ;
  assign n2823 = n2365 &  n2822 ;
  assign n2824 = n2365 | n2820 ;
  assign n2825 = ( n2815 & ~n2823 ) | ( n2815 & n2824 ) | ( ~n2823 & n2824 ) ;
  assign n2826 = ~n2811 & n2813 ;
  assign n2827 = ( n2825 & ~n2826 ) | ( n2825 & 1'b0 ) | ( ~n2826 & 1'b0 ) ;
  assign n2828 = ( n1077 & n2577 ) | ( n1077 & n2584 ) | ( n2577 & n2584 ) ;
  assign n2829 = ( n1077 & ~n2577 ) | ( n1077 & n2584 ) | ( ~n2577 & n2584 ) ;
  assign n2830 = ( n2577 & ~n2828 ) | ( n2577 & n2829 ) | ( ~n2828 & n2829 ) ;
  assign n2831 = ( n2617 & ~n2830 ) | ( n2617 & 1'b0 ) | ( ~n2830 & 1'b0 ) ;
  assign n2832 = ~n2617 & n2830 ;
  assign n2833 = n2831 | n2832 ;
  assign n2837 = n2700 | n2203 ;
  assign n2834 = ~n1910 & n2701 ;
  assign n2835 = ~n1896 & n2703 ;
  assign n2836 = n2834 | n2835 ;
  assign n2838 = ( n2837 & ~n2203 ) | ( n2837 & n2836 ) | ( ~n2203 & n2836 ) ;
  assign n2839 = ~n2226 & n2631 ;
  assign n2840 = n2838 | n2839 ;
  assign n2841 = ( n2365 & ~n2840 ) | ( n2365 & 1'b0 ) | ( ~n2840 & 1'b0 ) ;
  assign n2842 = ~n2365 & n2840 ;
  assign n2843 = n2841 | n2842 ;
  assign n2844 = ( n2827 & ~n2833 ) | ( n2827 & n2843 ) | ( ~n2833 & n2843 ) ;
  assign n2855 = ( n2746 & ~n2844 ) | ( n2746 & 1'b0 ) | ( ~n2844 & 1'b0 ) ;
  assign n2851 = ~n2631 & n2212 ;
  assign n2848 = ( n2187 & ~n2700 ) | ( n2187 & 1'b0 ) | ( ~n2700 & 1'b0 ) ;
  assign n2845 = ~n1896 & n2701 ;
  assign n2846 = ~n2203 & n2703 ;
  assign n2847 = n2845 | n2846 ;
  assign n2849 = ( n2187 & ~n2848 ) | ( n2187 & n2847 ) | ( ~n2848 & n2847 ) ;
  assign n2850 = ( n2365 & ~n2849 ) | ( n2365 & 1'b0 ) | ( ~n2849 & 1'b0 ) ;
  assign n2852 = ( n2851 & ~n2212 ) | ( n2851 & n2850 ) | ( ~n2212 & n2850 ) ;
  assign n2853 = n2212 &  n2742 ;
  assign n2854 = n2852 | n2853 ;
  assign n2856 = ( n2746 & ~n2855 ) | ( n2746 & n2854 ) | ( ~n2855 & n2854 ) ;
  assign n2859 = ~n2844 & n2746 ;
  assign n2857 = ~n2365 & n2849 ;
  assign n2858 = ~n2854 & n2857 ;
  assign n2860 = ( n2859 & ~n2746 ) | ( n2859 & n2858 ) | ( ~n2746 & n2858 ) ;
  assign n2861 = n2746 | n2844 ;
  assign n2862 = ( n2561 & ~n2551 ) | ( n2561 & n2619 ) | ( ~n2551 & n2619 ) ;
  assign n2863 = ( n2551 & ~n2619 ) | ( n2551 & n2561 ) | ( ~n2619 & n2561 ) ;
  assign n2864 = ( n2862 & ~n2561 ) | ( n2862 & n2863 ) | ( ~n2561 & n2863 ) ;
  assign n2865 = ( n2861 & ~n2864 ) | ( n2861 & 1'b0 ) | ( ~n2864 & 1'b0 ) ;
  assign n2866 = ( n2856 & n2860 ) | ( n2856 & n2865 ) | ( n2860 & n2865 ) ;
  assign n2867 = n2744 | n2866 ;
  assign n2871 = n2700 | n2341 ;
  assign n2868 = ~n2203 & n2701 ;
  assign n2869 = n2187 &  n2703 ;
  assign n2870 = n2868 | n2869 ;
  assign n2872 = ( n2871 & ~n2341 ) | ( n2871 & n2870 ) | ( ~n2341 & n2870 ) ;
  assign n2873 = n2344 &  n2631 ;
  assign n2874 = n2872 | n2873 ;
  assign n2875 = n2365 &  n2874 ;
  assign n2876 = n2365 | n2872 ;
  assign n2877 = ( n2867 & ~n2875 ) | ( n2867 & n2876 ) | ( ~n2875 & n2876 ) ;
  assign n2878 = ( n2857 & ~n2856 ) | ( n2857 & n2861 ) | ( ~n2856 & n2861 ) ;
  assign n2879 = ~n2857 & n2878 ;
  assign n2880 = ( n2864 & ~n2861 ) | ( n2864 & n2879 ) | ( ~n2861 & n2879 ) ;
  assign n2881 = ( n2877 & ~n2880 ) | ( n2877 & 1'b0 ) | ( ~n2880 & 1'b0 ) ;
  assign n2882 = ( n2546 & n2548 ) | ( n2546 & n2620 ) | ( n2548 & n2620 ) ;
  assign n2883 = ( n2548 & ~n2882 ) | ( n2548 & n2621 ) | ( ~n2882 & n2621 ) ;
  assign n2884 = ( n2881 & ~n2883 ) | ( n2881 & 1'b0 ) | ( ~n2883 & 1'b0 ) ;
  assign n2885 = n2743 | n2884 ;
  assign n2889 = ( n2461 & ~n2700 ) | ( n2461 & 1'b0 ) | ( ~n2700 & 1'b0 ) ;
  assign n2886 = n2187 &  n2701 ;
  assign n2887 = ~n2341 & n2703 ;
  assign n2888 = n2886 | n2887 ;
  assign n2890 = ( n2461 & ~n2889 ) | ( n2461 & n2888 ) | ( ~n2889 & n2888 ) ;
  assign n2891 = n2505 &  n2631 ;
  assign n2892 = n2890 | n2891 ;
  assign n2893 = n2365 &  n2892 ;
  assign n2894 = n2365 | n2890 ;
  assign n2895 = ( n2885 & ~n2893 ) | ( n2885 & n2894 ) | ( ~n2893 & n2894 ) ;
  assign n2896 = ~n2881 & n2883 ;
  assign n2897 = ( n2895 & ~n2896 ) | ( n2895 & 1'b0 ) | ( ~n2896 & 1'b0 ) ;
  assign n2899 = ( n2526 & n2536 ) | ( n2526 & n2621 ) | ( n2536 & n2621 ) ;
  assign n2898 = ( n2526 & ~n2536 ) | ( n2526 & n2621 ) | ( ~n2536 & n2621 ) ;
  assign n2900 = ( n2536 & ~n2899 ) | ( n2536 & n2898 ) | ( ~n2899 & n2898 ) ;
  assign n2904 = n2700 | n2464 ;
  assign n2901 = ~n2341 & n2701 ;
  assign n2902 = n2461 &  n2703 ;
  assign n2903 = n2901 | n2902 ;
  assign n2905 = ( n2904 & ~n2464 ) | ( n2904 & n2903 ) | ( ~n2464 & n2903 ) ;
  assign n2906 = n2490 &  n2631 ;
  assign n2907 = n2905 | n2906 ;
  assign n2908 = ( n2365 & ~n2907 ) | ( n2365 & 1'b0 ) | ( ~n2907 & 1'b0 ) ;
  assign n2909 = ~n2365 & n2907 ;
  assign n2910 = n2908 | n2909 ;
  assign n2911 = ( n2897 & ~n2900 ) | ( n2897 & n2910 ) | ( ~n2900 & n2910 ) ;
  assign n2912 = ( n2523 & ~n2513 ) | ( n2523 & n2622 ) | ( ~n2513 & n2622 ) ;
  assign n2913 = ( n2513 & ~n2622 ) | ( n2513 & n2523 ) | ( ~n2622 & n2523 ) ;
  assign n2914 = ( n2912 & ~n2523 ) | ( n2912 & n2913 ) | ( ~n2523 & n2913 ) ;
  assign n2918 = n2700 | n2454 ;
  assign n2915 = n2461 &  n2701 ;
  assign n2916 = ~n2464 & n2703 ;
  assign n2917 = n2915 | n2916 ;
  assign n2919 = ( n2918 & ~n2454 ) | ( n2918 & n2917 ) | ( ~n2454 & n2917 ) ;
  assign n2920 = ~n2476 & n2631 ;
  assign n2921 = n2919 | n2920 ;
  assign n2922 = ( n2365 & ~n2921 ) | ( n2365 & 1'b0 ) | ( ~n2921 & 1'b0 ) ;
  assign n2923 = ~n2365 & n2921 ;
  assign n2924 = n2922 | n2923 ;
  assign n2925 = ( n2911 & ~n2914 ) | ( n2911 & n2924 ) | ( ~n2914 & n2924 ) ;
  assign n2926 = ( n2739 & n2741 ) | ( n2739 & n2925 ) | ( n2741 & n2925 ) ;
  assign n2927 = ( n2715 & n2727 ) | ( n2715 & n2926 ) | ( n2727 & n2926 ) ;
  assign n2928 = ( n2628 & n2712 ) | ( n2628 & n2927 ) | ( n2712 & n2927 ) ;
  assign n2936 = ( n100 & ~n161 ) | ( n100 & 1'b0 ) | ( ~n161 & 1'b0 ) ;
  assign n2929 = n391 | n729 ;
  assign n2930 = n122 | n2929 ;
  assign n2931 = ( n736 & ~n699 ) | ( n736 & n2930 ) | ( ~n699 & n2930 ) ;
  assign n2932 = n699 | n2931 ;
  assign n2933 = ( n761 & ~n754 ) | ( n761 & n2932 ) | ( ~n754 & n2932 ) ;
  assign n2934 = n754 | n2933 ;
  assign n2935 = n198 | n2934 ;
  assign n2937 = ( n100 & ~n2936 ) | ( n100 & n2935 ) | ( ~n2936 & n2935 ) ;
  assign n2938 = ( n2672 & ~n2685 ) | ( n2672 & 1'b0 ) | ( ~n2685 & 1'b0 ) ;
  assign n2939 = ( n2937 & ~n2938 ) | ( n2937 & 1'b0 ) | ( ~n2938 & 1'b0 ) ;
  assign n2940 = n2937 | n2938 ;
  assign n2941 = ( n2939 & ~n2937 ) | ( n2939 & n2940 ) | ( ~n2937 & n2940 ) ;
  assign n2942 = ( n2688 & ~n2695 ) | ( n2688 & n2941 ) | ( ~n2695 & n2941 ) ;
  assign n2943 = ( n2695 & ~n2688 ) | ( n2695 & n2941 ) | ( ~n2688 & n2941 ) ;
  assign n2944 = ( n2942 & ~n2941 ) | ( n2942 & n2943 ) | ( ~n2941 & n2943 ) ;
  assign n2950 = n2631 &  n2944 ;
  assign n2948 = ~n2941 & n2700 ;
  assign n2945 = ~n2674 & n2701 ;
  assign n2946 = n2688 &  n2703 ;
  assign n2947 = n2945 | n2946 ;
  assign n2949 = ( n2700 & ~n2948 ) | ( n2700 & n2947 ) | ( ~n2948 & n2947 ) ;
  assign n2951 = ( n2631 & ~n2950 ) | ( n2631 & n2949 ) | ( ~n2950 & n2949 ) ;
  assign n2952 = ( n2365 & ~n2951 ) | ( n2365 & 1'b0 ) | ( ~n2951 & 1'b0 ) ;
  assign n2953 = ~n2365 & n2951 ;
  assign n2954 = n2952 | n2953 ;
  assign n2956 = ( n2459 & ~n2464 ) | ( n2459 & 1'b0 ) | ( ~n2464 & 1'b0 ) ;
  assign n2957 = ~n2454 & n2465 ;
  assign n2958 = n2956 | n2957 ;
  assign n2955 = ( n2369 & ~n2691 ) | ( n2369 & 1'b0 ) | ( ~n2691 & 1'b0 ) ;
  assign n2959 = ( n2691 & ~n2958 ) | ( n2691 & n2955 ) | ( ~n2958 & n2955 ) ;
  assign n2960 = ( n2470 & ~n2734 ) | ( n2470 & 1'b0 ) | ( ~n2734 & 1'b0 ) ;
  assign n2961 = ( n2959 & ~n2960 ) | ( n2959 & 1'b0 ) | ( ~n2960 & 1'b0 ) ;
  assign n2962 = ( x5 & ~n1074 ) | ( x5 & n2961 ) | ( ~n1074 & n2961 ) ;
  assign n2963 = ( x5 & ~n2961 ) | ( x5 & n1074 ) | ( ~n2961 & n1074 ) ;
  assign n2964 = ( n2962 & ~x5 ) | ( n2962 & n2963 ) | ( ~x5 & n2963 ) ;
  assign n2996 = n2461 | n2194 ;
  assign n2993 = n2187 &  n2200 ;
  assign n2994 = ( n2204 & ~n2341 ) | ( n2204 & 1'b0 ) | ( ~n2341 & 1'b0 ) ;
  assign n2995 = n2993 | n2994 ;
  assign n2997 = ( n2996 & ~n2194 ) | ( n2996 & n2995 ) | ( ~n2194 & n2995 ) ;
  assign n2998 = ( n2213 & n2505 ) | ( n2213 & n2997 ) | ( n2505 & n2997 ) ;
  assign n2999 = ( n2505 & ~n2998 ) | ( n2505 & 1'b0 ) | ( ~n2998 & 1'b0 ) ;
  assign n3000 = ( n2997 & ~n248 ) | ( n2997 & n2999 ) | ( ~n248 & n2999 ) ;
  assign n3001 = ( n248 & ~n2997 ) | ( n248 & n2999 ) | ( ~n2997 & n2999 ) ;
  assign n3002 = ( n3000 & ~n2999 ) | ( n3000 & n3001 ) | ( ~n2999 & n3001 ) ;
  assign n2965 = ( n1906 & ~n1910 ) | ( n1906 & 1'b0 ) | ( ~n1910 & 1'b0 ) ;
  assign n2966 = ~n1896 & n1911 ;
  assign n2967 = n2965 | n2966 ;
  assign n2968 = ~n260 & n2203 ;
  assign n2969 = ( n260 & ~n2967 ) | ( n260 & n2968 ) | ( ~n2967 & n2968 ) ;
  assign n2970 = n1916 | n2226 ;
  assign n2971 = n2969 &  n2970 ;
  assign n2972 = ( x11 & ~n252 ) | ( x11 & n2971 ) | ( ~n252 & n2971 ) ;
  assign n2973 = ( x11 & ~n2971 ) | ( x11 & n252 ) | ( ~n2971 & n252 ) ;
  assign n2974 = ( n2972 & ~x11 ) | ( n2972 & n2973 ) | ( ~x11 & n2973 ) ;
  assign n2975 = ~n883 & n1940 ;
  assign n2976 = n2060 | n2975 ;
  assign n2977 = ( n1993 & ~n2059 ) | ( n1993 & n2976 ) | ( ~n2059 & n2976 ) ;
  assign n2978 = ( n1976 & n1977 ) | ( n1976 & n1990 ) | ( n1977 & n1990 ) ;
  assign n2979 = ( n540 & ~n1930 ) | ( n540 & 1'b0 ) | ( ~n1930 & 1'b0 ) ;
  assign n2983 = n1952 | n1901 ;
  assign n2980 = ~n1924 & n1967 ;
  assign n2981 = ~n1922 & n1947 ;
  assign n2982 = n2980 | n2981 ;
  assign n2984 = ( n2983 & ~n1901 ) | ( n2983 & n2982 ) | ( ~n1901 & n2982 ) ;
  assign n2985 = n1958 | n2004 ;
  assign n2986 = ~n2984 & n2985 ;
  assign n2988 = ( n2978 & n2979 ) | ( n2978 & n2986 ) | ( n2979 & n2986 ) ;
  assign n2987 = ( n2979 & ~n2978 ) | ( n2979 & n2986 ) | ( ~n2978 & n2986 ) ;
  assign n2989 = ( n2978 & ~n2988 ) | ( n2978 & n2987 ) | ( ~n2988 & n2987 ) ;
  assign n2991 = ( n2974 & n2977 ) | ( n2974 & n2989 ) | ( n2977 & n2989 ) ;
  assign n2990 = ( n2977 & ~n2974 ) | ( n2977 & n2989 ) | ( ~n2974 & n2989 ) ;
  assign n2992 = ( n2974 & ~n2991 ) | ( n2974 & n2990 ) | ( ~n2991 & n2990 ) ;
  assign n3003 = ( n2355 & ~n3002 ) | ( n2355 & n2992 ) | ( ~n3002 & n2992 ) ;
  assign n3004 = ( n2992 & ~n2355 ) | ( n2992 & n3002 ) | ( ~n2355 & n3002 ) ;
  assign n3005 = ( n3003 & ~n2992 ) | ( n3003 & n3004 ) | ( ~n2992 & n3004 ) ;
  assign n3006 = ( n2964 & ~n2626 ) | ( n2964 & n3005 ) | ( ~n2626 & n3005 ) ;
  assign n3007 = ( n2626 & ~n3005 ) | ( n2626 & n2964 ) | ( ~n3005 & n2964 ) ;
  assign n3008 = ( n3006 & ~n2964 ) | ( n3006 & n3007 ) | ( ~n2964 & n3007 ) ;
  assign n3009 = ( n2928 & ~n2954 ) | ( n2928 & n3008 ) | ( ~n2954 & n3008 ) ;
  assign n3010 = ( n2928 & ~n3008 ) | ( n2928 & n2954 ) | ( ~n3008 & n2954 ) ;
  assign n3011 = ( n3009 & ~n2928 ) | ( n3009 & n3010 ) | ( ~n2928 & n3010 ) ;
  assign n175 = ( n163 & ~n159 ) | ( n163 & n174 ) | ( ~n159 & n174 ) ;
  assign n176 = n159 | n175 ;
  assign n177 = ( n141 & ~n140 ) | ( n141 & n176 ) | ( ~n140 & n176 ) ;
  assign n178 = n140 | n177 ;
  assign n193 = ( n101 & ~n161 ) | ( n101 & n107 ) | ( ~n161 & n107 ) ;
  assign n194 = n161 | n193 ;
  assign n203 = n148 &  n68 ;
  assign n202 = n200 | n201 ;
  assign n204 = ( n68 & ~n203 ) | ( n68 & n202 ) | ( ~n203 & n202 ) ;
  assign n205 = ( n199 & ~n198 ) | ( n199 & n204 ) | ( ~n198 & n204 ) ;
  assign n206 = n198 | n205 ;
  assign n207 = n197 | n206 ;
  assign n213 = n211 | n212 ;
  assign n214 = ( n210 & ~n207 ) | ( n210 & n213 ) | ( ~n207 & n213 ) ;
  assign n215 = n207 | n214 ;
  assign n216 = ( n196 & ~n195 ) | ( n196 & n215 ) | ( ~n195 & n215 ) ;
  assign n217 = n195 | n216 ;
  assign n218 = ( n194 & ~n101 ) | ( n194 & n217 ) | ( ~n101 & n217 ) ;
  assign n219 = ( n192 & ~n191 ) | ( n192 & n218 ) | ( ~n191 & n218 ) ;
  assign n220 = n191 | n219 ;
  assign n221 = ( n190 & ~n189 ) | ( n190 & n220 ) | ( ~n189 & n220 ) ;
  assign n222 = n189 | n221 ;
  assign n187 = ( n101 & ~n148 ) | ( n101 & n146 ) | ( ~n148 & n146 ) ;
  assign n188 = ( n101 & ~n187 ) | ( n101 & 1'b0 ) | ( ~n187 & 1'b0 ) ;
  assign n223 = ( n146 & ~n222 ) | ( n146 & n188 ) | ( ~n222 & n188 ) ;
  assign n224 = ( n185 & ~n186 ) | ( n185 & n223 ) | ( ~n186 & n223 ) ;
  assign n225 = ~n185 & n224 ;
  assign n232 = ( n225 & n228 ) | ( n225 & n231 ) | ( n228 & n231 ) ;
  assign n233 = ( n225 & ~n232 ) | ( n225 & 1'b0 ) | ( ~n232 & 1'b0 ) ;
  assign n234 = ( n178 & ~n184 ) | ( n178 & n233 ) | ( ~n184 & n233 ) ;
  assign n235 = ~n178 & n234 ;
  assign n236 = ( n105 & ~n139 ) | ( n105 & n235 ) | ( ~n139 & n235 ) ;
  assign n237 = ~n105 & n236 ;
  assign n238 = ( n97 & ~n103 ) | ( n97 & n237 ) | ( ~n103 & n237 ) ;
  assign n239 = ~n97 & n238 ;
  assign n240 = ( n85 & ~n91 ) | ( n85 & n239 ) | ( ~n91 & n239 ) ;
  assign n241 = ~n85 & n240 ;
  assign n242 = ( n69 & ~n78 ) | ( n69 & n241 ) | ( ~n78 & n241 ) ;
  assign n243 = ~n69 & n242 ;
  assign n3012 = n85 | n363 ;
  assign n3013 = ( n807 & ~n106 ) | ( n807 & n3012 ) | ( ~n106 & n3012 ) ;
  assign n3014 = n128 | n3013 ;
  assign n3015 = ( n826 & ~n113 ) | ( n826 & n3014 ) | ( ~n113 & n3014 ) ;
  assign n3016 = n113 | n3015 ;
  assign n3017 = ( n160 & ~n124 ) | ( n160 & n3016 ) | ( ~n124 & n3016 ) ;
  assign n3018 = n124 | n3017 ;
  assign n3019 = ( n412 & ~n109 ) | ( n412 & n3018 ) | ( ~n109 & n3018 ) ;
  assign n3020 = n109 | n3019 ;
  assign n3021 = ( n290 & ~n116 ) | ( n290 & n3020 ) | ( ~n116 & n3020 ) ;
  assign n3022 = n116 | n3021 ;
  assign n3023 = n69 | n3022 ;
  assign n3024 = n615 | n1725 ;
  assign n3025 = ( n941 & ~n191 ) | ( n941 & n3024 ) | ( ~n191 & n3024 ) ;
  assign n3026 = n191 | n3025 ;
  assign n3027 = ( n364 & ~n227 ) | ( n364 & n3026 ) | ( ~n227 & n3026 ) ;
  assign n3028 = n227 | n3027 ;
  assign n3029 = ( n554 & ~n316 ) | ( n554 & n3028 ) | ( ~n316 & n3028 ) ;
  assign n3030 = n316 | n3029 ;
  assign n3031 = ( n282 & ~n189 ) | ( n282 & n3030 ) | ( ~n189 & n3030 ) ;
  assign n3032 = n189 | n3031 ;
  assign n3033 = ( n809 & ~n323 ) | ( n809 & n3032 ) | ( ~n323 & n3032 ) ;
  assign n3034 = n323 | n3033 ;
  assign n3035 = n398 | n3034 ;
  assign n3036 = ( n1834 & ~n3023 ) | ( n1834 & n3035 ) | ( ~n3023 & n3035 ) ;
  assign n3037 = ( n3023 & ~n326 ) | ( n3023 & n3036 ) | ( ~n326 & n3036 ) ;
  assign n3038 = n326 | n3037 ;
  assign n3039 = ( n226 & ~n411 ) | ( n226 & n3038 ) | ( ~n411 & n3038 ) ;
  assign n3040 = n411 | n3039 ;
  assign n3041 = ( n277 & ~n276 ) | ( n277 & n3040 ) | ( ~n276 & n3040 ) ;
  assign n3042 = n276 | n3041 ;
  assign n3043 = ( n353 & ~n120 ) | ( n353 & n3042 ) | ( ~n120 & n3042 ) ;
  assign n3044 = n120 | n3043 ;
  assign n3045 = ( n487 & ~n379 ) | ( n487 & n3044 ) | ( ~n379 & n3044 ) ;
  assign n3046 = ( n379 & ~n501 ) | ( n379 & n3045 ) | ( ~n501 & n3045 ) ;
  assign n3047 = n501 | n3046 ;
  assign n3048 = ( n2628 & ~n2927 ) | ( n2628 & n2712 ) | ( ~n2927 & n2712 ) ;
  assign n3049 = ( n2927 & ~n2928 ) | ( n2927 & n3048 ) | ( ~n2928 & n3048 ) ;
  assign n3072 = n2715 &  n2727 ;
  assign n3073 = ~n2715 & n2727 ;
  assign n3074 = ( n2715 & ~n3072 ) | ( n2715 & n3073 ) | ( ~n3072 & n3073 ) ;
  assign n3050 = n835 | n2376 ;
  assign n3051 = ( n129 & ~n411 ) | ( n129 & n3050 ) | ( ~n411 & n3050 ) ;
  assign n3052 = n411 | n3051 ;
  assign n3053 = n747 | n1803 ;
  assign n3054 = ( n1665 & ~n118 ) | ( n1665 & n3053 ) | ( ~n118 & n3053 ) ;
  assign n3055 = n118 | n3054 ;
  assign n3056 = ( n362 & ~n266 ) | ( n362 & n3055 ) | ( ~n266 & n3055 ) ;
  assign n3057 = n266 | n3056 ;
  assign n3058 = n643 | n3057 ;
  assign n3059 = n680 | n1804 ;
  assign n3060 = ( n1815 & ~n611 ) | ( n1815 & n3059 ) | ( ~n611 & n3059 ) ;
  assign n3061 = n611 | n3060 ;
  assign n3062 = ( n3058 & ~n3052 ) | ( n3058 & n3061 ) | ( ~n3052 & n3061 ) ;
  assign n3063 = ( n3052 & ~n1723 ) | ( n3052 & n3062 ) | ( ~n1723 & n3062 ) ;
  assign n3064 = n1723 | n3063 ;
  assign n3065 = ( n381 & ~n124 ) | ( n381 & n3064 ) | ( ~n124 & n3064 ) ;
  assign n3066 = n124 | n3065 ;
  assign n3067 = ( n446 & ~n380 ) | ( n446 & n3066 ) | ( ~n380 & n3066 ) ;
  assign n3068 = n380 | n3067 ;
  assign n3069 = ( n192 & ~n149 ) | ( n192 & n3068 ) | ( ~n149 & n3068 ) ;
  assign n3070 = n149 | n3069 ;
  assign n3071 = n302 | n3070 ;
  assign n3075 = ( n2926 & ~n3074 ) | ( n2926 & n3071 ) | ( ~n3074 & n3071 ) ;
  assign n3076 = ( n3071 & ~n2926 ) | ( n3071 & n3074 ) | ( ~n2926 & n3074 ) ;
  assign n3077 = n3075 &  n3076 ;
  assign n3078 = ( n3047 & ~n3049 ) | ( n3047 & n3077 ) | ( ~n3049 & n3077 ) ;
  assign n3079 = ( n3011 & ~n243 ) | ( n3011 & n3078 ) | ( ~n243 & n3078 ) ;
  assign n3080 = n213 | n888 ;
  assign n3081 = ( n1192 & ~n826 ) | ( n1192 & n3080 ) | ( ~n826 & n3080 ) ;
  assign n3082 = n826 | n3081 ;
  assign n3083 = ( n642 & ~n3082 ) | ( n642 & n1674 ) | ( ~n3082 & n1674 ) ;
  assign n3084 = ~n642 & n3083 ;
  assign n3085 = ( n184 & ~n624 ) | ( n184 & n3084 ) | ( ~n624 & n3084 ) ;
  assign n3086 = ~n184 & n3085 ;
  assign n3087 = ( n122 & ~n227 ) | ( n122 & n3086 ) | ( ~n227 & n3086 ) ;
  assign n3088 = ~n122 & n3087 ;
  assign n3089 = n378 &  n3088 ;
  assign n3169 = ~n2454 & n2459 ;
  assign n3170 = ( n2465 & ~n2691 ) | ( n2465 & 1'b0 ) | ( ~n2691 & 1'b0 ) ;
  assign n3171 = n3169 | n3170 ;
  assign n3168 = ( n2369 & ~n2674 ) | ( n2369 & 1'b0 ) | ( ~n2674 & 1'b0 ) ;
  assign n3172 = ( n2674 & ~n3171 ) | ( n2674 & n3168 ) | ( ~n3171 & n3168 ) ;
  assign n3173 = ( n2470 & n2722 ) | ( n2470 & n3172 ) | ( n2722 & n3172 ) ;
  assign n3174 = ~n2722 & n3173 ;
  assign n3175 = ( n1077 & ~n3172 ) | ( n1077 & n3174 ) | ( ~n3172 & n3174 ) ;
  assign n3176 = ( n3172 & ~n1077 ) | ( n3172 & n3174 ) | ( ~n1077 & n3174 ) ;
  assign n3177 = ( n3175 & ~n3174 ) | ( n3175 & n3176 ) | ( ~n3174 & n3176 ) ;
  assign n3128 = n540 &  n2986 ;
  assign n3129 = ( n2978 & ~n2988 ) | ( n2978 & n3128 ) | ( ~n2988 & n3128 ) ;
  assign n3130 = ~n1922 & n1967 ;
  assign n3131 = ~n1901 & n1947 ;
  assign n3132 = n3130 | n3131 ;
  assign n3133 = n1910 | n1952 ;
  assign n3134 = ( n3132 & ~n1910 ) | ( n3132 & n3133 ) | ( ~n1910 & n3133 ) ;
  assign n3135 = n1958 | n2048 ;
  assign n3136 = ~n3134 & n3135 ;
  assign n3137 = n540 &  n1924 ;
  assign n3138 = ( n3129 & n3136 ) | ( n3129 & n3137 ) | ( n3136 & n3137 ) ;
  assign n3139 = ( n3136 & ~n3129 ) | ( n3136 & n3137 ) | ( ~n3129 & n3137 ) ;
  assign n3140 = ( n3129 & ~n3138 ) | ( n3129 & n3139 ) | ( ~n3138 & n3139 ) ;
  assign n3147 = n2212 | n1916 ;
  assign n3145 = n2187 | n260 ;
  assign n3142 = ~n1896 & n1906 ;
  assign n3143 = ( n1911 & ~n2203 ) | ( n1911 & 1'b0 ) | ( ~n2203 & 1'b0 ) ;
  assign n3144 = n3142 | n3143 ;
  assign n3146 = ( n3145 & ~n260 ) | ( n3145 & n3144 ) | ( ~n260 & n3144 ) ;
  assign n3148 = ( n3147 & ~n1916 ) | ( n3147 & n3146 ) | ( ~n1916 & n3146 ) ;
  assign n3149 = ( x11 & n252 ) | ( x11 & n3148 ) | ( n252 & n3148 ) ;
  assign n3150 = ( x11 & ~n3148 ) | ( x11 & n252 ) | ( ~n3148 & n252 ) ;
  assign n3151 = ( n3148 & ~n3149 ) | ( n3148 & n3150 ) | ( ~n3149 & n3150 ) ;
  assign n3141 = ( n2974 & ~n2977 ) | ( n2974 & n2989 ) | ( ~n2977 & n2989 ) ;
  assign n3152 = ( n3140 & ~n3151 ) | ( n3140 & n3141 ) | ( ~n3151 & n3141 ) ;
  assign n3153 = ( n3140 & ~n3141 ) | ( n3140 & n3151 ) | ( ~n3141 & n3151 ) ;
  assign n3154 = ( n3152 & ~n3140 ) | ( n3152 & n3153 ) | ( ~n3140 & n3153 ) ;
  assign n3155 = ( n2200 & ~n2341 ) | ( n2200 & 1'b0 ) | ( ~n2341 & 1'b0 ) ;
  assign n3156 = n2204 &  n2461 ;
  assign n3157 = n3155 | n3156 ;
  assign n3158 = ~n2194 & n2464 ;
  assign n3159 = ( n2194 & ~n3157 ) | ( n2194 & n3158 ) | ( ~n3157 & n3158 ) ;
  assign n3160 = ~n2213 & n2490 ;
  assign n3161 = ( n3159 & ~n3160 ) | ( n3159 & 1'b0 ) | ( ~n3160 & 1'b0 ) ;
  assign n3162 = ~n248 & n3161 ;
  assign n3163 = ( n248 & ~n3161 ) | ( n248 & 1'b0 ) | ( ~n3161 & 1'b0 ) ;
  assign n3164 = n3162 | n3163 ;
  assign n3165 = ( n3004 & n3154 ) | ( n3004 & n3164 ) | ( n3154 & n3164 ) ;
  assign n3166 = ( n3004 & ~n3154 ) | ( n3004 & n3164 ) | ( ~n3154 & n3164 ) ;
  assign n3167 = ( n3154 & ~n3165 ) | ( n3154 & n3166 ) | ( ~n3165 & n3166 ) ;
  assign n3178 = ( n3006 & ~n3177 ) | ( n3006 & n3167 ) | ( ~n3177 & n3167 ) ;
  assign n3179 = ( n3167 & ~n3006 ) | ( n3167 & n3177 ) | ( ~n3006 & n3177 ) ;
  assign n3180 = ( n3178 & ~n3167 ) | ( n3178 & n3179 ) | ( ~n3167 & n3179 ) ;
  assign n3090 = ~n2937 & n2938 ;
  assign n3091 = n213 | n584 ;
  assign n3092 = ( n291 & ~n97 ) | ( n291 & n3091 ) | ( ~n97 & n3091 ) ;
  assign n3093 = n97 | n3092 ;
  assign n3094 = ( n412 & ~n181 ) | ( n412 & n3093 ) | ( ~n181 & n3093 ) ;
  assign n3095 = n181 | n3094 ;
  assign n3096 = ( n281 & ~n316 ) | ( n281 & n3095 ) | ( ~n316 & n3095 ) ;
  assign n3097 = n316 | n3096 ;
  assign n3098 = n319 | n547 ;
  assign n3099 = n2372 | n3098 ;
  assign n3100 = ( n1798 & ~n3097 ) | ( n1798 & n3099 ) | ( ~n3097 & n3099 ) ;
  assign n3101 = ( n973 & n3097 ) | ( n973 & n3100 ) | ( n3097 & n3100 ) ;
  assign n3102 = ( n973 & ~n3101 ) | ( n973 & 1'b0 ) | ( ~n3101 & 1'b0 ) ;
  assign n3103 = ( n196 & ~n446 ) | ( n196 & n3102 ) | ( ~n446 & n3102 ) ;
  assign n3104 = ~n196 & n3103 ;
  assign n3105 = ( n152 & ~n192 ) | ( n152 & n3104 ) | ( ~n192 & n3104 ) ;
  assign n3106 = ~n152 & n3105 ;
  assign n3107 = ( n185 & ~n555 ) | ( n185 & n3106 ) | ( ~n555 & n3106 ) ;
  assign n3108 = ~n185 & n3107 ;
  assign n3109 = ( n108 & ~n197 ) | ( n108 & n3108 ) | ( ~n197 & n3108 ) ;
  assign n3110 = ~n108 & n3109 ;
  assign n3111 = n3090 | n3110 ;
  assign n3112 = ( n3090 & ~n3110 ) | ( n3090 & 1'b0 ) | ( ~n3110 & 1'b0 ) ;
  assign n3113 = ( n3111 & ~n3090 ) | ( n3111 & n3112 ) | ( ~n3090 & n3112 ) ;
  assign n3117 = n3113 &  n2700 ;
  assign n3114 = n2688 &  n2701 ;
  assign n3115 = n2703 &  n2941 ;
  assign n3116 = n3114 | n3115 ;
  assign n3118 = ( n2700 & ~n3117 ) | ( n2700 & n3116 ) | ( ~n3117 & n3116 ) ;
  assign n3119 = ( n2939 & ~n3110 ) | ( n2939 & 1'b0 ) | ( ~n3110 & 1'b0 ) ;
  assign n3120 = ~n2939 & n3110 ;
  assign n3121 = n3119 | n3120 ;
  assign n3122 = ( n2942 & ~n3121 ) | ( n2942 & 1'b0 ) | ( ~n3121 & 1'b0 ) ;
  assign n3123 = ( n2631 & ~n3121 ) | ( n2631 & n2942 ) | ( ~n3121 & n2942 ) ;
  assign n3124 = ( n3118 & ~n3122 ) | ( n3118 & n3123 ) | ( ~n3122 & n3123 ) ;
  assign n3125 = n2365 &  n3124 ;
  assign n3126 = n2365 | n3124 ;
  assign n3127 = ~n3125 & n3126 ;
  assign n3181 = ( n3010 & n3127 ) | ( n3010 & n3180 ) | ( n3127 & n3180 ) ;
  assign n3182 = ( n3010 & ~n3180 ) | ( n3010 & n3127 ) | ( ~n3180 & n3127 ) ;
  assign n3183 = ( n3180 & ~n3181 ) | ( n3180 & n3182 ) | ( ~n3181 & n3182 ) ;
  assign n3184 = ( n3079 & ~n3089 ) | ( n3079 & n3183 ) | ( ~n3089 & n3183 ) ;
  assign n3185 = ( n3079 & ~n3183 ) | ( n3079 & n3089 ) | ( ~n3183 & n3089 ) ;
  assign n3186 = ( n3184 & ~n3079 ) | ( n3184 & n3185 ) | ( ~n3079 & n3185 ) ;
  assign n3188 = ( n243 & n3011 ) | ( n243 & n3078 ) | ( n3011 & n3078 ) ;
  assign n3187 = ( n243 & ~n3011 ) | ( n243 & n3078 ) | ( ~n3011 & n3078 ) ;
  assign n3189 = ( n3011 & ~n3188 ) | ( n3011 & n3187 ) | ( ~n3188 & n3187 ) ;
  assign n3190 = ~n3186 & n3189 ;
  assign n3191 = ( n3186 & ~n3189 ) | ( n3186 & 1'b0 ) | ( ~n3189 & 1'b0 ) ;
  assign n3192 = n3190 | n3191 ;
  assign n3193 = ( x22 & ~x23 ) | ( x22 & 1'b0 ) | ( ~x23 & 1'b0 ) ;
  assign n3194 = ~x22 & x23 ;
  assign n3195 = ~n3193 &  ~n3194 ;
  assign n3196 = ( n3186 & n3189 ) | ( n3186 & n3195 ) | ( n3189 & n3195 ) ;
  assign n3197 = n114 | n419 ;
  assign n3198 = ( n595 & ~n230 ) | ( n595 & n3197 ) | ( ~n230 & n3197 ) ;
  assign n3199 = n230 | n3198 ;
  assign n3200 = n637 | n1700 ;
  assign n3201 = n2159 | n3200 ;
  assign n3202 = ( n399 & ~n3199 ) | ( n399 & n3201 ) | ( ~n3199 & n3201 ) ;
  assign n3203 = ( n3199 & ~n222 ) | ( n3199 & n3202 ) | ( ~n222 & n3202 ) ;
  assign n3204 = n222 | n3203 ;
  assign n3205 = ( n2645 & ~n184 ) | ( n2645 & n3204 ) | ( ~n184 & n3204 ) ;
  assign n3206 = n184 | n3205 ;
  assign n3207 = ( n309 & ~n129 ) | ( n309 & n3206 ) | ( ~n129 & n3206 ) ;
  assign n3208 = n129 | n3207 ;
  assign n3209 = ( n276 & ~n165 ) | ( n276 & n3208 ) | ( ~n165 & n3208 ) ;
  assign n3210 = n165 | n3209 ;
  assign n3211 = n91 | n3210 ;
  assign n3212 = n316 | n3211 ;
  assign n3251 = n1952 | n1896 ;
  assign n3248 = ~n1901 & n1967 ;
  assign n3249 = ~n1910 & n1947 ;
  assign n3250 = n3248 | n3249 ;
  assign n3252 = ( n3251 & ~n1896 ) | ( n3251 & n3250 ) | ( ~n1896 & n3250 ) ;
  assign n3253 = n1938 | n1958 ;
  assign n3254 = ~n3252 & n3253 ;
  assign n3255 = n540 &  n3136 ;
  assign n3256 = ( n3129 & ~n3138 ) | ( n3129 & n3255 ) | ( ~n3138 & n3255 ) ;
  assign n3257 = n540 &  n1922 ;
  assign n3258 = ( n3254 & n3256 ) | ( n3254 & n3257 ) | ( n3256 & n3257 ) ;
  assign n3259 = ( n3256 & ~n3254 ) | ( n3256 & n3257 ) | ( ~n3254 & n3257 ) ;
  assign n3260 = ( n3254 & ~n3258 ) | ( n3254 & n3259 ) | ( ~n3258 & n3259 ) ;
  assign n3266 = n2344 | n1916 ;
  assign n3261 = ( n1906 & ~n2203 ) | ( n1906 & 1'b0 ) | ( ~n2203 & 1'b0 ) ;
  assign n3262 = n1911 &  n2187 ;
  assign n3263 = n3261 | n3262 ;
  assign n3264 = ~n260 & n2341 ;
  assign n3265 = ( n260 & ~n3263 ) | ( n260 & n3264 ) | ( ~n3263 & n3264 ) ;
  assign n3267 = ( n1916 & ~n3266 ) | ( n1916 & n3265 ) | ( ~n3266 & n3265 ) ;
  assign n3269 = ( x11 & n252 ) | ( x11 & n3267 ) | ( n252 & n3267 ) ;
  assign n3268 = ( x11 & ~n3267 ) | ( x11 & n252 ) | ( ~n3267 & n252 ) ;
  assign n3270 = ( n3267 & ~n3269 ) | ( n3267 & n3268 ) | ( ~n3269 & n3268 ) ;
  assign n3272 = ( n3152 & n3260 ) | ( n3152 & n3270 ) | ( n3260 & n3270 ) ;
  assign n3271 = ( n3152 & ~n3260 ) | ( n3152 & n3270 ) | ( ~n3260 & n3270 ) ;
  assign n3273 = ( n3260 & ~n3272 ) | ( n3260 & n3271 ) | ( ~n3272 & n3271 ) ;
  assign n3274 = n2200 &  n2461 ;
  assign n3275 = ( n2204 & ~n2464 ) | ( n2204 & 1'b0 ) | ( ~n2464 & 1'b0 ) ;
  assign n3276 = n3274 | n3275 ;
  assign n3277 = ~n2194 & n2454 ;
  assign n3278 = ( n2194 & ~n3276 ) | ( n2194 & n3277 ) | ( ~n3276 & n3277 ) ;
  assign n3279 = n2213 | n2476 ;
  assign n3280 = n3278 &  n3279 ;
  assign n3281 = ~n248 & n3280 ;
  assign n3282 = ( n248 & ~n3280 ) | ( n248 & 1'b0 ) | ( ~n3280 & 1'b0 ) ;
  assign n3283 = n3281 | n3282 ;
  assign n3284 = ( n3004 & ~n3164 ) | ( n3004 & n3154 ) | ( ~n3164 & n3154 ) ;
  assign n3286 = ( n3273 & n3283 ) | ( n3273 & n3284 ) | ( n3283 & n3284 ) ;
  assign n3285 = ( n3283 & ~n3273 ) | ( n3283 & n3284 ) | ( ~n3273 & n3284 ) ;
  assign n3287 = ( n3273 & ~n3286 ) | ( n3273 & n3285 ) | ( ~n3286 & n3285 ) ;
  assign n3291 = n2688 | n2369 ;
  assign n3288 = ( n2459 & ~n2691 ) | ( n2459 & 1'b0 ) | ( ~n2691 & 1'b0 ) ;
  assign n3289 = ( n2465 & ~n2674 ) | ( n2465 & 1'b0 ) | ( ~n2674 & 1'b0 ) ;
  assign n3290 = n3288 | n3289 ;
  assign n3292 = ( n3291 & ~n2369 ) | ( n3291 & n3290 ) | ( ~n2369 & n3290 ) ;
  assign n3293 = ( n2697 & ~n2470 ) | ( n2697 & n3292 ) | ( ~n2470 & n3292 ) ;
  assign n3294 = ( n2697 & ~n3293 ) | ( n2697 & 1'b0 ) | ( ~n3293 & 1'b0 ) ;
  assign n3295 = ( n1077 & n3292 ) | ( n1077 & n3294 ) | ( n3292 & n3294 ) ;
  assign n3296 = ( n1077 & ~n3294 ) | ( n1077 & n3292 ) | ( ~n3294 & n3292 ) ;
  assign n3297 = ( n3294 & ~n3295 ) | ( n3294 & n3296 ) | ( ~n3295 & n3296 ) ;
  assign n3299 = ( n3178 & n3287 ) | ( n3178 & n3297 ) | ( n3287 & n3297 ) ;
  assign n3298 = ( n3178 & ~n3287 ) | ( n3178 & n3297 ) | ( ~n3287 & n3297 ) ;
  assign n3300 = ( n3287 & ~n3299 ) | ( n3287 & n3298 ) | ( ~n3299 & n3298 ) ;
  assign n3213 = n3090 &  n3110 ;
  assign n3221 = n445 | n556 ;
  assign n3222 = ( n837 & ~n3221 ) | ( n837 & n1209 ) | ( ~n3221 & n1209 ) ;
  assign n3223 = ~n837 & n3222 ;
  assign n3214 = n210 | n1815 ;
  assign n3215 = ( n399 & ~n677 ) | ( n399 & n3214 ) | ( ~n677 & n3214 ) ;
  assign n3216 = n677 | n3215 ;
  assign n3217 = ( n143 & ~n91 ) | ( n143 & n3216 ) | ( ~n91 & n3216 ) ;
  assign n3218 = n91 | n3217 ;
  assign n3219 = ( n142 & ~n140 ) | ( n142 & n3218 ) | ( ~n140 & n3218 ) ;
  assign n3220 = n140 | n3219 ;
  assign n3224 = ( n1814 & ~n3223 ) | ( n1814 & n3220 ) | ( ~n3223 & n3220 ) ;
  assign n3225 = ( n1814 & ~n3224 ) | ( n1814 & 1'b0 ) | ( ~n3224 & 1'b0 ) ;
  assign n3226 = ( n364 & ~n303 ) | ( n364 & n3225 ) | ( ~n303 & n3225 ) ;
  assign n3227 = ~n364 & n3226 ;
  assign n3228 = ( n261 & ~n379 ) | ( n261 & n3227 ) | ( ~n379 & n3227 ) ;
  assign n3229 = ~n261 & n3228 ;
  assign n3230 = ~n612 & n3229 ;
  assign n3231 = n3213 &  n3230 ;
  assign n3232 = n3213 | n3230 ;
  assign n3233 = ~n3231 & n3232 ;
  assign n3237 = n3233 &  n2700 ;
  assign n3234 = n2701 &  n2941 ;
  assign n3235 = ( n2703 & ~n3113 ) | ( n2703 & 1'b0 ) | ( ~n3113 & 1'b0 ) ;
  assign n3236 = n3234 | n3235 ;
  assign n3238 = ( n2700 & ~n3237 ) | ( n2700 & n3236 ) | ( ~n3237 & n3236 ) ;
  assign n3239 = ( n2941 & ~n3113 ) | ( n2941 & n2942 ) | ( ~n3113 & n2942 ) ;
  assign n3240 = ( n3233 & ~n3113 ) | ( n3233 & n3239 ) | ( ~n3113 & n3239 ) ;
  assign n3241 = ( n3113 & ~n3239 ) | ( n3113 & n3233 ) | ( ~n3239 & n3233 ) ;
  assign n3242 = ( n3240 & ~n3233 ) | ( n3240 & n3241 ) | ( ~n3233 & n3241 ) ;
  assign n3243 = n2631 &  n3242 ;
  assign n3244 = n3238 | n3243 ;
  assign n3245 = n2365 &  n3244 ;
  assign n3246 = n2365 | n3244 ;
  assign n3247 = ~n3245 & n3246 ;
  assign n3301 = ( n3182 & n3247 ) | ( n3182 & n3300 ) | ( n3247 & n3300 ) ;
  assign n3302 = ( n3182 & ~n3300 ) | ( n3182 & n3247 ) | ( ~n3300 & n3247 ) ;
  assign n3303 = ( n3300 & ~n3301 ) | ( n3300 & n3302 ) | ( ~n3301 & n3302 ) ;
  assign n3304 = ( n3184 & n3212 ) | ( n3184 & n3303 ) | ( n3212 & n3303 ) ;
  assign n3305 = ( n3212 & ~n3184 ) | ( n3212 & n3303 ) | ( ~n3184 & n3303 ) ;
  assign n3306 = ( n3184 & ~n3304 ) | ( n3184 & n3305 ) | ( ~n3304 & n3305 ) ;
  assign n3307 = ~n3196 & n3306 ;
  assign n3308 = ( n3196 & ~n3306 ) | ( n3196 & 1'b0 ) | ( ~n3306 & 1'b0 ) ;
  assign n3309 = n3307 | n3308 ;
  assign n3310 = n3186 | n3189 ;
  assign n3312 = ( n3190 & n3306 ) | ( n3190 & n3310 ) | ( n3306 & n3310 ) ;
  assign n3313 = n3189 | n3306 ;
  assign n3314 = ~n3312 & n3313 ;
  assign n3315 = n3195 | n3314 ;
  assign n3311 = ( n3306 & ~n3310 ) | ( n3306 & 1'b0 ) | ( ~n3310 & 1'b0 ) ;
  assign n3345 = ( n3273 & ~n3284 ) | ( n3273 & n3283 ) | ( ~n3284 & n3283 ) ;
  assign n3380 = n3272 &  n3345 ;
  assign n3379 = ~n3272 & n3345 ;
  assign n3381 = ( n3272 & ~n3380 ) | ( n3272 & n3379 ) | ( ~n3380 & n3379 ) ;
  assign n3347 = ( n2200 & ~n2464 ) | ( n2200 & 1'b0 ) | ( ~n2464 & 1'b0 ) ;
  assign n3348 = ( n2204 & ~n2454 ) | ( n2204 & 1'b0 ) | ( ~n2454 & 1'b0 ) ;
  assign n3349 = n3347 | n3348 ;
  assign n3346 = ( n2194 & ~n2691 ) | ( n2194 & 1'b0 ) | ( ~n2691 & 1'b0 ) ;
  assign n3350 = ( n2691 & ~n3349 ) | ( n2691 & n3346 ) | ( ~n3349 & n3346 ) ;
  assign n3351 = n2213 | n2734 ;
  assign n3352 = n3350 &  n3351 ;
  assign n3353 = ~n248 & n3352 ;
  assign n3354 = ( n248 & ~n3352 ) | ( n248 & 1'b0 ) | ( ~n3352 & 1'b0 ) ;
  assign n3355 = n3353 | n3354 ;
  assign n3356 = n540 &  n3254 ;
  assign n3357 = ( n3256 & ~n3258 ) | ( n3256 & n3356 ) | ( ~n3258 & n3356 ) ;
  assign n3358 = n540 &  n1901 ;
  assign n3362 = n2203 &  n1952 ;
  assign n3359 = ~n1910 & n1967 ;
  assign n3360 = ~n1896 & n1947 ;
  assign n3361 = n3359 | n3360 ;
  assign n3363 = ( n1952 & ~n3362 ) | ( n1952 & n3361 ) | ( ~n3362 & n3361 ) ;
  assign n3364 = n1958 | n2226 ;
  assign n3365 = ~n3363 & n3364 ;
  assign n3367 = ( n3357 & n3358 ) | ( n3357 & n3365 ) | ( n3358 & n3365 ) ;
  assign n3366 = ( n3358 & ~n3357 ) | ( n3358 & n3365 ) | ( ~n3357 & n3365 ) ;
  assign n3368 = ( n3357 & ~n3367 ) | ( n3357 & n3366 ) | ( ~n3367 & n3366 ) ;
  assign n3374 = n2505 | n1916 ;
  assign n3372 = n2461 | n260 ;
  assign n3369 = n1906 &  n2187 ;
  assign n3370 = ( n1911 & ~n2341 ) | ( n1911 & 1'b0 ) | ( ~n2341 & 1'b0 ) ;
  assign n3371 = n3369 | n3370 ;
  assign n3373 = ( n3372 & ~n260 ) | ( n3372 & n3371 ) | ( ~n260 & n3371 ) ;
  assign n3375 = ( n3374 & ~n1916 ) | ( n3374 & n3373 ) | ( ~n1916 & n3373 ) ;
  assign n3376 = ( n3368 & ~n883 ) | ( n3368 & n3375 ) | ( ~n883 & n3375 ) ;
  assign n3377 = ( n883 & ~n3375 ) | ( n883 & n3368 ) | ( ~n3375 & n3368 ) ;
  assign n3378 = ( n3376 & ~n3368 ) | ( n3376 & n3377 ) | ( ~n3368 & n3377 ) ;
  assign n3382 = ( n3355 & n3378 ) | ( n3355 & n3381 ) | ( n3378 & n3381 ) ;
  assign n3383 = ( n3355 & ~n3381 ) | ( n3355 & n3378 ) | ( ~n3381 & n3378 ) ;
  assign n3384 = ( n3381 & ~n3382 ) | ( n3381 & n3383 ) | ( ~n3382 & n3383 ) ;
  assign n3388 = n2941 | n2369 ;
  assign n3385 = ( n2459 & ~n2674 ) | ( n2459 & 1'b0 ) | ( ~n2674 & 1'b0 ) ;
  assign n3386 = n2465 &  n2688 ;
  assign n3387 = n3385 | n3386 ;
  assign n3389 = ( n3388 & ~n2369 ) | ( n3388 & n3387 ) | ( ~n2369 & n3387 ) ;
  assign n3390 = ( n2470 & ~n3389 ) | ( n2470 & n2944 ) | ( ~n3389 & n2944 ) ;
  assign n3391 = ~n2944 & n3390 ;
  assign n3392 = ( n1077 & n3389 ) | ( n1077 & n3391 ) | ( n3389 & n3391 ) ;
  assign n3393 = ( n1077 & ~n3391 ) | ( n1077 & n3389 ) | ( ~n3391 & n3389 ) ;
  assign n3394 = ( n3391 & ~n3392 ) | ( n3391 & n3393 ) | ( ~n3392 & n3393 ) ;
  assign n3395 = ( n3298 & n3384 ) | ( n3298 & n3394 ) | ( n3384 & n3394 ) ;
  assign n3396 = ( n3298 & ~n3384 ) | ( n3298 & n3394 ) | ( ~n3384 & n3394 ) ;
  assign n3397 = ( n3384 & ~n3395 ) | ( n3384 & n3396 ) | ( ~n3395 & n3396 ) ;
  assign n3335 = n3239 &  n3113 ;
  assign n3336 = ( n3113 & ~n3335 ) | ( n3113 & n3233 ) | ( ~n3335 & n3233 ) ;
  assign n3337 = n3239 | n3113 ;
  assign n3338 = ( n3113 & ~n3337 ) | ( n3113 & n3233 ) | ( ~n3337 & n3233 ) ;
  assign n3339 = ( n3336 & ~n3338 ) | ( n3336 & 1'b0 ) | ( ~n3338 & 1'b0 ) ;
  assign n3340 = ( n2631 & ~n3339 ) | ( n2631 & 1'b0 ) | ( ~n3339 & 1'b0 ) ;
  assign n3332 = ( n2701 & ~n3113 ) | ( n2701 & 1'b0 ) | ( ~n3113 & 1'b0 ) ;
  assign n3333 = ( n2703 & ~n3233 ) | ( n2703 & 1'b0 ) | ( ~n3233 & 1'b0 ) ;
  assign n3334 = n3332 | n3333 ;
  assign n3341 = ( n2631 & ~n3340 ) | ( n2631 & n3334 ) | ( ~n3340 & n3334 ) ;
  assign n3342 = n2365 &  n3341 ;
  assign n3343 = n2365 | n3341 ;
  assign n3344 = ~n3342 & n3343 ;
  assign n3399 = ( n3302 & n3344 ) | ( n3302 & n3397 ) | ( n3344 & n3397 ) ;
  assign n3398 = ( n3302 & ~n3397 ) | ( n3302 & n3344 ) | ( ~n3397 & n3344 ) ;
  assign n3400 = ( n3397 & ~n3399 ) | ( n3397 & n3398 ) | ( ~n3399 & n3398 ) ;
  assign n3316 = ~n352 & n2377 ;
  assign n3317 = ( n105 & ~n201 ) | ( n105 & n3316 ) | ( ~n201 & n3316 ) ;
  assign n3318 = ~n105 & n3317 ;
  assign n3319 = ( n108 & ~n116 ) | ( n108 & n3318 ) | ( ~n116 & n3318 ) ;
  assign n3320 = ~n108 & n3319 ;
  assign n3321 = n609 | n755 ;
  assign n3322 = ( n3058 & n3320 ) | ( n3058 & n3321 ) | ( n3320 & n3321 ) ;
  assign n3323 = ( n825 & ~n3322 ) | ( n825 & n3320 ) | ( ~n3322 & n3320 ) ;
  assign n3324 = ~n825 & n3323 ;
  assign n3325 = ( n412 & ~n647 ) | ( n412 & n3324 ) | ( ~n647 & n3324 ) ;
  assign n3326 = ~n412 & n3325 ;
  assign n3327 = ( n398 & ~n354 ) | ( n398 & n3326 ) | ( ~n354 & n3326 ) ;
  assign n3328 = ~n398 & n3327 ;
  assign n3329 = ( n120 & ~n363 ) | ( n120 & n3328 ) | ( ~n363 & n3328 ) ;
  assign n3330 = ~n120 & n3329 ;
  assign n3331 = ~n612 & n3330 ;
  assign n3401 = ( n3304 & n3331 ) | ( n3304 & n3400 ) | ( n3331 & n3400 ) ;
  assign n3402 = ( n3304 & ~n3400 ) | ( n3304 & n3331 ) | ( ~n3400 & n3331 ) ;
  assign n3403 = ( n3400 & ~n3401 ) | ( n3400 & n3402 ) | ( ~n3401 & n3402 ) ;
  assign n3404 = ( n3315 & ~n3311 ) | ( n3315 & n3403 ) | ( ~n3311 & n3403 ) ;
  assign n3405 = ( n3311 & ~n3315 ) | ( n3311 & n3403 ) | ( ~n3315 & n3403 ) ;
  assign n3406 = ( n3404 & ~n3403 ) | ( n3404 & n3405 ) | ( ~n3403 & n3405 ) ;
  assign n3407 = n3311 &  n3403 ;
  assign n3408 = n3311 | n3403 ;
  assign n3409 = ( n3314 & ~n3408 ) | ( n3314 & n3407 ) | ( ~n3408 & n3407 ) ;
  assign n3410 = n3195 | n3409 ;
  assign n3412 = n1700 | n3014 ;
  assign n3413 = ( n500 & ~n747 ) | ( n500 & n3412 ) | ( ~n747 & n3412 ) ;
  assign n3414 = n747 | n3413 ;
  assign n3415 = ( n1201 & n2165 ) | ( n1201 & n3414 ) | ( n2165 & n3414 ) ;
  assign n3416 = ( n1201 & ~n3415 ) | ( n1201 & 1'b0 ) | ( ~n3415 & 1'b0 ) ;
  assign n3417 = ( n388 & n549 ) | ( n388 & n3416 ) | ( n549 & n3416 ) ;
  assign n3418 = ~n549 & n3417 ;
  assign n3419 = ( n309 & ~n446 ) | ( n309 & n3418 ) | ( ~n446 & n3418 ) ;
  assign n3420 = ~n309 & n3419 ;
  assign n3421 = ( n78 & ~n318 ) | ( n78 & n3420 ) | ( ~n318 & n3420 ) ;
  assign n3422 = ~n78 & n3421 ;
  assign n3423 = ~n230 & n3422 ;
  assign n3424 = ~n212 & n3423 ;
  assign n3411 = ( n3331 & ~n3304 ) | ( n3331 & n3400 ) | ( ~n3304 & n3400 ) ;
  assign n3425 = ( n2701 & ~n3233 ) | ( n2701 & 1'b0 ) | ( ~n3233 & 1'b0 ) ;
  assign n3426 = ( n2631 & ~n3336 ) | ( n2631 & 1'b0 ) | ( ~n3336 & 1'b0 ) ;
  assign n3427 = n3425 | n3426 ;
  assign n3428 = n2365 | n3427 ;
  assign n3429 = n2365 &  n3427 ;
  assign n3430 = ( n3428 & ~n3429 ) | ( n3428 & 1'b0 ) | ( ~n3429 & 1'b0 ) ;
  assign n3478 = n2459 &  n2688 ;
  assign n3479 = n2465 &  n2941 ;
  assign n3480 = n3478 | n3479 ;
  assign n3481 = ~n2369 & n3113 ;
  assign n3482 = ( n2369 & ~n3480 ) | ( n2369 & n3481 ) | ( ~n3480 & n3481 ) ;
  assign n3483 = ~n2942 & n3121 ;
  assign n3484 = n3122 | n3483 ;
  assign n3485 = ( n2470 & n3482 ) | ( n2470 & n3484 ) | ( n3482 & n3484 ) ;
  assign n3486 = ~n3484 & n3485 ;
  assign n3487 = ( n1077 & ~n3482 ) | ( n1077 & n3486 ) | ( ~n3482 & n3486 ) ;
  assign n3488 = ( n3482 & ~n1077 ) | ( n3482 & n3486 ) | ( ~n1077 & n3486 ) ;
  assign n3489 = ( n3487 & ~n3486 ) | ( n3487 & n3488 ) | ( ~n3486 & n3488 ) ;
  assign n3434 = ~n2187 & n1952 ;
  assign n3431 = ~n1896 & n1967 ;
  assign n3432 = ( n1947 & ~n2203 ) | ( n1947 & 1'b0 ) | ( ~n2203 & 1'b0 ) ;
  assign n3433 = n3431 | n3432 ;
  assign n3435 = ( n1952 & ~n3434 ) | ( n1952 & n3433 ) | ( ~n3434 & n3433 ) ;
  assign n3436 = ~n1958 & n2212 ;
  assign n3437 = n3435 | n3436 ;
  assign n3438 = n540 &  n3365 ;
  assign n3439 = ( n3357 & ~n3367 ) | ( n3357 & n3438 ) | ( ~n3367 & n3438 ) ;
  assign n3440 = n540 &  n1910 ;
  assign n3442 = ( n3437 & n3439 ) | ( n3437 & n3440 ) | ( n3439 & n3440 ) ;
  assign n3441 = ( n3439 & ~n3437 ) | ( n3439 & n3440 ) | ( ~n3437 & n3440 ) ;
  assign n3443 = ( n3437 & ~n3442 ) | ( n3437 & n3441 ) | ( ~n3442 & n3441 ) ;
  assign n3448 = ( n1906 & ~n2341 ) | ( n1906 & 1'b0 ) | ( ~n2341 & 1'b0 ) ;
  assign n3449 = n1911 &  n2461 ;
  assign n3450 = n3448 | n3449 ;
  assign n3451 = ~n260 & n2464 ;
  assign n3452 = ( n260 & ~n3450 ) | ( n260 & n3451 ) | ( ~n3450 & n3451 ) ;
  assign n3453 = ( n1916 & ~n3452 ) | ( n1916 & n2490 ) | ( ~n3452 & n2490 ) ;
  assign n3454 = ( n2490 & ~n3453 ) | ( n2490 & 1'b0 ) | ( ~n3453 & 1'b0 ) ;
  assign n3455 = ( n883 & ~n3452 ) | ( n883 & n3454 ) | ( ~n3452 & n3454 ) ;
  assign n3456 = ( n3452 & ~n883 ) | ( n3452 & n3454 ) | ( ~n883 & n3454 ) ;
  assign n3457 = ( n3455 & ~n3454 ) | ( n3455 & n3456 ) | ( ~n3454 & n3456 ) ;
  assign n3444 = ( x11 & n252 ) | ( x11 & n3375 ) | ( n252 & n3375 ) ;
  assign n3445 = ( x11 & ~n3375 ) | ( x11 & n252 ) | ( ~n3375 & n252 ) ;
  assign n3446 = ( n3375 & ~n3444 ) | ( n3375 & n3445 ) | ( ~n3444 & n3445 ) ;
  assign n3447 = ( n3272 & ~n3446 ) | ( n3272 & n3368 ) | ( ~n3446 & n3368 ) ;
  assign n3458 = ( n3443 & ~n3457 ) | ( n3443 & n3447 ) | ( ~n3457 & n3447 ) ;
  assign n3459 = ( n3443 & ~n3447 ) | ( n3443 & n3457 ) | ( ~n3447 & n3457 ) ;
  assign n3460 = ( n3458 & ~n3443 ) | ( n3458 & n3459 ) | ( ~n3443 & n3459 ) ;
  assign n3471 = n3272 | n3378 ;
  assign n3472 = n3272 &  n3378 ;
  assign n3473 = ( n3471 & ~n3472 ) | ( n3471 & 1'b0 ) | ( ~n3472 & 1'b0 ) ;
  assign n3474 = ( n3345 & n3355 ) | ( n3345 & n3473 ) | ( n3355 & n3473 ) ;
  assign n3462 = ( n2200 & ~n2454 ) | ( n2200 & 1'b0 ) | ( ~n2454 & 1'b0 ) ;
  assign n3463 = ( n2204 & ~n2691 ) | ( n2204 & 1'b0 ) | ( ~n2691 & 1'b0 ) ;
  assign n3464 = n3462 | n3463 ;
  assign n3461 = ( n2194 & ~n2674 ) | ( n2194 & 1'b0 ) | ( ~n2674 & 1'b0 ) ;
  assign n3465 = ( n2674 & ~n3464 ) | ( n2674 & n3461 ) | ( ~n3464 & n3461 ) ;
  assign n3466 = n2213 | n2722 ;
  assign n3467 = n3465 &  n3466 ;
  assign n3468 = ~n248 & n3467 ;
  assign n3469 = ( n248 & ~n3467 ) | ( n248 & 1'b0 ) | ( ~n3467 & 1'b0 ) ;
  assign n3470 = n3468 | n3469 ;
  assign n3475 = ( n3460 & ~n3474 ) | ( n3460 & n3470 ) | ( ~n3474 & n3470 ) ;
  assign n3476 = ( n3460 & ~n3470 ) | ( n3460 & n3474 ) | ( ~n3470 & n3474 ) ;
  assign n3477 = ( n3475 & ~n3460 ) | ( n3475 & n3476 ) | ( ~n3460 & n3476 ) ;
  assign n3490 = ( n3430 & ~n3489 ) | ( n3430 & n3477 ) | ( ~n3489 & n3477 ) ;
  assign n3491 = ( n3477 & ~n3430 ) | ( n3477 & n3489 ) | ( ~n3430 & n3489 ) ;
  assign n3492 = ( n3490 & ~n3477 ) | ( n3490 & n3491 ) | ( ~n3477 & n3491 ) ;
  assign n3493 = ( n3395 & n3399 ) | ( n3395 & n3492 ) | ( n3399 & n3492 ) ;
  assign n3494 = ( n3395 & ~n3399 ) | ( n3395 & n3492 ) | ( ~n3399 & n3492 ) ;
  assign n3495 = ( n3399 & ~n3493 ) | ( n3399 & n3494 ) | ( ~n3493 & n3494 ) ;
  assign n3496 = ( n3424 & ~n3411 ) | ( n3424 & n3495 ) | ( ~n3411 & n3495 ) ;
  assign n3497 = ( n3411 & ~n3424 ) | ( n3411 & n3495 ) | ( ~n3424 & n3495 ) ;
  assign n3498 = ( n3496 & ~n3495 ) | ( n3496 & n3497 ) | ( ~n3495 & n3497 ) ;
  assign n3499 = ( n3407 & ~n3410 ) | ( n3407 & n3498 ) | ( ~n3410 & n3498 ) ;
  assign n3500 = ( n3407 & ~n3498 ) | ( n3407 & n3410 ) | ( ~n3498 & n3410 ) ;
  assign n3501 = ( n3499 & ~n3407 ) | ( n3499 & n3500 ) | ( ~n3407 & n3500 ) ;
  assign n3502 = n3407 &  n3498 ;
  assign n3503 = n3407 | n3498 ;
  assign n3504 = ( n3409 & ~n3503 ) | ( n3409 & n3502 ) | ( ~n3503 & n3502 ) ;
  assign n3505 = n3195 | n3504 ;
  assign n3507 = ~n502 & n2377 ;
  assign n3508 = ( n830 & ~n1844 ) | ( n830 & n3507 ) | ( ~n1844 & n3507 ) ;
  assign n3509 = ~n830 & n3508 ;
  assign n3510 = ( n377 & ~n288 ) | ( n377 & n3509 ) | ( ~n288 & n3509 ) ;
  assign n3511 = ~n377 & n3510 ;
  assign n3512 = ( n646 & ~n3511 ) | ( n646 & n1798 ) | ( ~n3511 & n1798 ) ;
  assign n3513 = ( n646 & ~n3512 ) | ( n646 & 1'b0 ) | ( ~n3512 & 1'b0 ) ;
  assign n3514 = ( n153 & ~n167 ) | ( n153 & n3513 ) | ( ~n167 & n3513 ) ;
  assign n3515 = ~n153 & n3514 ;
  assign n3516 = ~n468 & n3515 ;
  assign n3506 = ( n3411 & ~n3495 ) | ( n3411 & n3424 ) | ( ~n3495 & n3424 ) ;
  assign n3517 = ( n3395 & ~n3492 ) | ( n3395 & n3399 ) | ( ~n3492 & n3399 ) ;
  assign n3518 = ( n540 & ~n3437 ) | ( n540 & 1'b0 ) | ( ~n3437 & 1'b0 ) ;
  assign n3519 = ( n3439 & ~n3441 ) | ( n3439 & n3518 ) | ( ~n3441 & n3518 ) ;
  assign n3520 = n540 &  n1896 ;
  assign n3524 = n2341 &  n1952 ;
  assign n3521 = ( n1967 & ~n2203 ) | ( n1967 & 1'b0 ) | ( ~n2203 & 1'b0 ) ;
  assign n3522 = n1947 &  n2187 ;
  assign n3523 = n3521 | n3522 ;
  assign n3525 = ( n1952 & ~n3524 ) | ( n1952 & n3523 ) | ( ~n3524 & n3523 ) ;
  assign n3526 = ~n1958 & n2344 ;
  assign n3527 = n3525 | n3526 ;
  assign n3528 = ( n2365 & ~n3520 ) | ( n2365 & n3527 ) | ( ~n3520 & n3527 ) ;
  assign n3529 = ( n3520 & ~n2365 ) | ( n3520 & n3527 ) | ( ~n2365 & n3527 ) ;
  assign n3530 = ( n3528 & ~n3527 ) | ( n3528 & n3529 ) | ( ~n3527 & n3529 ) ;
  assign n3531 = n1906 &  n2461 ;
  assign n3532 = ( n1911 & ~n2464 ) | ( n1911 & 1'b0 ) | ( ~n2464 & 1'b0 ) ;
  assign n3533 = n3531 | n3532 ;
  assign n3534 = ~n260 & n2454 ;
  assign n3535 = ( n260 & ~n3533 ) | ( n260 & n3534 ) | ( ~n3533 & n3534 ) ;
  assign n3536 = n1916 | n2476 ;
  assign n3537 = n3535 &  n3536 ;
  assign n3538 = ( x11 & ~n252 ) | ( x11 & n3537 ) | ( ~n252 & n3537 ) ;
  assign n3539 = ( x11 & ~n3537 ) | ( x11 & n252 ) | ( ~n3537 & n252 ) ;
  assign n3540 = ( n3538 & ~x11 ) | ( n3538 & n3539 ) | ( ~x11 & n3539 ) ;
  assign n3541 = ( n3519 & n3530 ) | ( n3519 & n3540 ) | ( n3530 & n3540 ) ;
  assign n3542 = ( n3530 & ~n3519 ) | ( n3530 & n3540 ) | ( ~n3519 & n3540 ) ;
  assign n3543 = ( n3519 & ~n3541 ) | ( n3519 & n3542 ) | ( ~n3541 & n3542 ) ;
  assign n3547 = n2688 | n2194 ;
  assign n3544 = ( n2200 & ~n2691 ) | ( n2200 & 1'b0 ) | ( ~n2691 & 1'b0 ) ;
  assign n3545 = ( n2204 & ~n2674 ) | ( n2204 & 1'b0 ) | ( ~n2674 & 1'b0 ) ;
  assign n3546 = n3544 | n3545 ;
  assign n3548 = ( n3547 & ~n2194 ) | ( n3547 & n3546 ) | ( ~n2194 & n3546 ) ;
  assign n3549 = ~n2213 & n2697 ;
  assign n3550 = n3548 | n3549 ;
  assign n3551 = n248 | n3550 ;
  assign n3552 = n248 &  n3550 ;
  assign n3553 = ( n3551 & ~n3552 ) | ( n3551 & 1'b0 ) | ( ~n3552 & 1'b0 ) ;
  assign n3554 = ( n3543 & ~n3459 ) | ( n3543 & n3553 ) | ( ~n3459 & n3553 ) ;
  assign n3555 = ( n3459 & ~n3553 ) | ( n3459 & n3543 ) | ( ~n3553 & n3543 ) ;
  assign n3556 = ( n3554 & ~n3543 ) | ( n3554 & n3555 ) | ( ~n3543 & n3555 ) ;
  assign n3557 = ( n3460 & n3470 ) | ( n3460 & n3474 ) | ( n3470 & n3474 ) ;
  assign n3559 = n2459 &  n2941 ;
  assign n3560 = ( n2465 & ~n3113 ) | ( n2465 & 1'b0 ) | ( ~n3113 & 1'b0 ) ;
  assign n3561 = n3559 | n3560 ;
  assign n3558 = ( n2369 & ~n3233 ) | ( n2369 & 1'b0 ) | ( ~n3233 & 1'b0 ) ;
  assign n3562 = ( n3233 & ~n3561 ) | ( n3233 & n3558 ) | ( ~n3561 & n3558 ) ;
  assign n3563 = n2470 &  n3242 ;
  assign n3564 = ( n3562 & ~n3563 ) | ( n3562 & 1'b0 ) | ( ~n3563 & 1'b0 ) ;
  assign n3565 = ( x5 & ~n1074 ) | ( x5 & n3564 ) | ( ~n1074 & n3564 ) ;
  assign n3566 = ( x5 & ~n3564 ) | ( x5 & n1074 ) | ( ~n3564 & n1074 ) ;
  assign n3567 = ( n3565 & ~x5 ) | ( n3565 & n3566 ) | ( ~x5 & n3566 ) ;
  assign n3569 = ( n3556 & n3557 ) | ( n3556 & n3567 ) | ( n3557 & n3567 ) ;
  assign n3568 = ( n3557 & ~n3556 ) | ( n3557 & n3567 ) | ( ~n3556 & n3567 ) ;
  assign n3570 = ( n3556 & ~n3569 ) | ( n3556 & n3568 ) | ( ~n3569 & n3568 ) ;
  assign n3571 = ( n3490 & n3517 ) | ( n3490 & n3570 ) | ( n3517 & n3570 ) ;
  assign n3572 = ( n3490 & ~n3517 ) | ( n3490 & n3570 ) | ( ~n3517 & n3570 ) ;
  assign n3573 = ( n3517 & ~n3571 ) | ( n3517 & n3572 ) | ( ~n3571 & n3572 ) ;
  assign n3574 = ( n3516 & ~n3506 ) | ( n3516 & n3573 ) | ( ~n3506 & n3573 ) ;
  assign n3575 = ( n3506 & ~n3516 ) | ( n3506 & n3573 ) | ( ~n3516 & n3573 ) ;
  assign n3576 = ( n3574 & ~n3573 ) | ( n3574 & n3575 ) | ( ~n3573 & n3575 ) ;
  assign n3577 = ( n3502 & ~n3505 ) | ( n3502 & n3576 ) | ( ~n3505 & n3576 ) ;
  assign n3578 = ( n3502 & ~n3576 ) | ( n3502 & n3505 ) | ( ~n3576 & n3505 ) ;
  assign n3579 = ( n3577 & ~n3502 ) | ( n3577 & n3578 ) | ( ~n3502 & n3578 ) ;
  assign n3580 = n3502 &  n3576 ;
  assign n3581 = n3502 | n3576 ;
  assign n3582 = ( n3504 & ~n3581 ) | ( n3504 & n3580 ) | ( ~n3581 & n3580 ) ;
  assign n3583 = n3195 | n3582 ;
  assign n3584 = ( n3506 & ~n3573 ) | ( n3506 & n3516 ) | ( ~n3573 & n3516 ) ;
  assign n3585 = n290 | n446 ;
  assign n3586 = n402 | n3585 ;
  assign n3587 = n163 | n829 ;
  assign n3588 = ( n3586 & ~n1680 ) | ( n3586 & n3587 ) | ( ~n1680 & n3587 ) ;
  assign n3589 = n1680 | n3588 ;
  assign n3590 = ( n3220 & ~n444 ) | ( n3220 & n3589 ) | ( ~n444 & n3589 ) ;
  assign n3591 = n444 | n3590 ;
  assign n3592 = ( n2657 & n3199 ) | ( n2657 & n3591 ) | ( n3199 & n3591 ) ;
  assign n3593 = ( n2657 & ~n3592 ) | ( n2657 & 1'b0 ) | ( ~n3592 & 1'b0 ) ;
  assign n3594 = ( n153 & ~n1666 ) | ( n153 & n3593 ) | ( ~n1666 & n3593 ) ;
  assign n3595 = ~n153 & n3594 ;
  assign n3596 = ( n467 & ~n323 ) | ( n467 & n3595 ) | ( ~n323 & n3595 ) ;
  assign n3597 = ~n467 & n3596 ;
  assign n3598 = ~n211 & n3597 ;
  assign n3600 = ( n3459 & n3543 ) | ( n3459 & n3553 ) | ( n3543 & n3553 ) ;
  assign n3604 = n2941 | n2194 ;
  assign n3601 = ( n2200 & ~n2674 ) | ( n2200 & 1'b0 ) | ( ~n2674 & 1'b0 ) ;
  assign n3602 = n2204 &  n2688 ;
  assign n3603 = n3601 | n3602 ;
  assign n3605 = ( n3604 & ~n2194 ) | ( n3604 & n3603 ) | ( ~n2194 & n3603 ) ;
  assign n3606 = n2213 | n2944 ;
  assign n3607 = ~n3605 & n3606 ;
  assign n3608 = ~n248 & n3607 ;
  assign n3609 = ( n248 & ~n3607 ) | ( n248 & 1'b0 ) | ( ~n3607 & 1'b0 ) ;
  assign n3610 = n3608 | n3609 ;
  assign n3614 = ~n2461 & n1952 ;
  assign n3611 = n1967 &  n2187 ;
  assign n3612 = ( n1947 & ~n2341 ) | ( n1947 & 1'b0 ) | ( ~n2341 & 1'b0 ) ;
  assign n3613 = n3611 | n3612 ;
  assign n3615 = ( n1952 & ~n3614 ) | ( n1952 & n3613 ) | ( ~n3614 & n3613 ) ;
  assign n3616 = ( n1958 & n2505 ) | ( n1958 & n3615 ) | ( n2505 & n3615 ) ;
  assign n3617 = ( n2505 & ~n3616 ) | ( n2505 & 1'b0 ) | ( ~n3616 & 1'b0 ) ;
  assign n3618 = ( n3615 & ~n540 ) | ( n3615 & n3617 ) | ( ~n540 & n3617 ) ;
  assign n3619 = ( n540 & ~n3615 ) | ( n540 & n3617 ) | ( ~n3615 & n3617 ) ;
  assign n3620 = ( n3618 & ~n3617 ) | ( n3618 & n3619 ) | ( ~n3617 & n3619 ) ;
  assign n3622 = ( n540 & ~n3527 ) | ( n540 & 1'b0 ) | ( ~n3527 & 1'b0 ) ;
  assign n3623 = ( n3528 & ~n2365 ) | ( n3528 & n3622 ) | ( ~n2365 & n3622 ) ;
  assign n3621 = ( n540 & ~n2203 ) | ( n540 & 1'b0 ) | ( ~n2203 & 1'b0 ) ;
  assign n3625 = ( n2365 & n3621 ) | ( n2365 & n3623 ) | ( n3621 & n3623 ) ;
  assign n3624 = ( n2365 & ~n3623 ) | ( n2365 & n3621 ) | ( ~n3623 & n3621 ) ;
  assign n3626 = ( n3623 & ~n3625 ) | ( n3623 & n3624 ) | ( ~n3625 & n3624 ) ;
  assign n3628 = ( n1906 & ~n2464 ) | ( n1906 & 1'b0 ) | ( ~n2464 & 1'b0 ) ;
  assign n3629 = ( n1911 & ~n2454 ) | ( n1911 & 1'b0 ) | ( ~n2454 & 1'b0 ) ;
  assign n3630 = n3628 | n3629 ;
  assign n3627 = ( n260 & ~n2691 ) | ( n260 & 1'b0 ) | ( ~n2691 & 1'b0 ) ;
  assign n3631 = ( n2691 & ~n3630 ) | ( n2691 & n3627 ) | ( ~n3630 & n3627 ) ;
  assign n3632 = n1916 | n2734 ;
  assign n3633 = n3631 &  n3632 ;
  assign n3634 = ( x11 & ~n252 ) | ( x11 & n3633 ) | ( ~n252 & n3633 ) ;
  assign n3635 = ( x11 & ~n3633 ) | ( x11 & n252 ) | ( ~n3633 & n252 ) ;
  assign n3636 = ( n3634 & ~x11 ) | ( n3634 & n3635 ) | ( ~x11 & n3635 ) ;
  assign n3638 = ( n3620 & n3626 ) | ( n3620 & n3636 ) | ( n3626 & n3636 ) ;
  assign n3637 = ( n3626 & ~n3620 ) | ( n3626 & n3636 ) | ( ~n3620 & n3636 ) ;
  assign n3639 = ( n3620 & ~n3638 ) | ( n3620 & n3637 ) | ( ~n3638 & n3637 ) ;
  assign n3640 = ( n3542 & ~n3610 ) | ( n3542 & n3639 ) | ( ~n3610 & n3639 ) ;
  assign n3641 = ( n3542 & ~n3639 ) | ( n3542 & n3610 ) | ( ~n3639 & n3610 ) ;
  assign n3642 = ( n3640 & ~n3542 ) | ( n3640 & n3641 ) | ( ~n3542 & n3641 ) ;
  assign n3646 = ~n3339 & n2470 ;
  assign n3643 = ( n2459 & ~n3113 ) | ( n2459 & 1'b0 ) | ( ~n3113 & 1'b0 ) ;
  assign n3644 = ( n2465 & ~n3233 ) | ( n2465 & 1'b0 ) | ( ~n3233 & 1'b0 ) ;
  assign n3645 = n3643 | n3644 ;
  assign n3647 = ( n2470 & ~n3646 ) | ( n2470 & n3645 ) | ( ~n3646 & n3645 ) ;
  assign n3648 = ~n1077 & n3647 ;
  assign n3649 = ( n1077 & ~n3647 ) | ( n1077 & 1'b0 ) | ( ~n3647 & 1'b0 ) ;
  assign n3650 = n3648 | n3649 ;
  assign n3651 = ( n3600 & n3642 ) | ( n3600 & n3650 ) | ( n3642 & n3650 ) ;
  assign n3652 = ( n3642 & ~n3600 ) | ( n3642 & n3650 ) | ( ~n3600 & n3650 ) ;
  assign n3653 = ( n3600 & ~n3651 ) | ( n3600 & n3652 ) | ( ~n3651 & n3652 ) ;
  assign n3599 = ( n3490 & ~n3570 ) | ( n3490 & n3517 ) | ( ~n3570 & n3517 ) ;
  assign n3654 = ( n3568 & ~n3653 ) | ( n3568 & n3599 ) | ( ~n3653 & n3599 ) ;
  assign n3655 = ( n3599 & ~n3568 ) | ( n3599 & n3653 ) | ( ~n3568 & n3653 ) ;
  assign n3656 = ( n3654 & ~n3599 ) | ( n3654 & n3655 ) | ( ~n3599 & n3655 ) ;
  assign n3657 = ( n3584 & ~n3598 ) | ( n3584 & n3656 ) | ( ~n3598 & n3656 ) ;
  assign n3658 = ( n3598 & ~n3584 ) | ( n3598 & n3656 ) | ( ~n3584 & n3656 ) ;
  assign n3659 = ( n3657 & ~n3656 ) | ( n3657 & n3658 ) | ( ~n3656 & n3658 ) ;
  assign n3661 = ( n3580 & n3583 ) | ( n3580 & n3659 ) | ( n3583 & n3659 ) ;
  assign n3660 = ( n3583 & ~n3580 ) | ( n3583 & n3659 ) | ( ~n3580 & n3659 ) ;
  assign n3662 = ( n3580 & ~n3661 ) | ( n3580 & n3660 ) | ( ~n3661 & n3660 ) ;
  assign n3663 = ( n3580 & ~n3659 ) | ( n3580 & 1'b0 ) | ( ~n3659 & 1'b0 ) ;
  assign n3664 = ~n3580 & n3659 ;
  assign n3665 = ( n3582 & n3663 ) | ( n3582 & n3664 ) | ( n3663 & n3664 ) ;
  assign n3666 = n3195 | n3665 ;
  assign n3668 = n445 | n924 ;
  assign n3669 = ( n1801 & ~n581 ) | ( n1801 & n3668 ) | ( ~n581 & n3668 ) ;
  assign n3670 = n581 | n3669 ;
  assign n3671 = ( n1700 & ~n130 ) | ( n1700 & n3670 ) | ( ~n130 & n3670 ) ;
  assign n3672 = n130 | n3671 ;
  assign n3673 = ( n303 & ~n1666 ) | ( n303 & n3672 ) | ( ~n1666 & n3672 ) ;
  assign n3674 = n1666 | n3673 ;
  assign n3675 = n289 | n3674 ;
  assign n3676 = ( n283 & ~n1838 ) | ( n283 & n2675 ) | ( ~n1838 & n2675 ) ;
  assign n3677 = ( n225 & n1838 ) | ( n225 & n3676 ) | ( n1838 & n3676 ) ;
  assign n3678 = ( n225 & ~n3677 ) | ( n225 & 1'b0 ) | ( ~n3677 & 1'b0 ) ;
  assign n3679 = ( n310 & ~n3675 ) | ( n310 & n3678 ) | ( ~n3675 & n3678 ) ;
  assign n3680 = ~n310 & n3679 ;
  assign n3681 = ( n124 & ~n147 ) | ( n124 & n3680 ) | ( ~n147 & n3680 ) ;
  assign n3682 = ~n124 & n3681 ;
  assign n3683 = ( n143 & ~n292 ) | ( n143 & n3682 ) | ( ~n292 & n3682 ) ;
  assign n3684 = ~n143 & n3683 ;
  assign n3685 = ~n122 & n3684 ;
  assign n3667 = ( n3584 & n3598 ) | ( n3584 & n3656 ) | ( n3598 & n3656 ) ;
  assign n3686 = ( n3568 & n3599 ) | ( n3568 & n3653 ) | ( n3599 & n3653 ) ;
  assign n3687 = ( n3600 & ~n3650 ) | ( n3600 & n3642 ) | ( ~n3650 & n3642 ) ;
  assign n3694 = n2200 &  n2688 ;
  assign n3695 = n2204 &  n2941 ;
  assign n3696 = n3694 | n3695 ;
  assign n3697 = ~n2194 & n3113 ;
  assign n3698 = ( n2194 & ~n3696 ) | ( n2194 & n3697 ) | ( ~n3696 & n3697 ) ;
  assign n3699 = n2213 | n3484 ;
  assign n3700 = n3698 &  n3699 ;
  assign n3701 = ~n248 & n3700 ;
  assign n3702 = ( n248 & ~n3700 ) | ( n248 & 1'b0 ) | ( ~n3700 & 1'b0 ) ;
  assign n3703 = n3701 | n3702 ;
  assign n3707 = n2464 &  n1952 ;
  assign n3704 = ( n1967 & ~n2341 ) | ( n1967 & 1'b0 ) | ( ~n2341 & 1'b0 ) ;
  assign n3705 = n1947 &  n2461 ;
  assign n3706 = n3704 | n3705 ;
  assign n3708 = ( n1952 & ~n3707 ) | ( n1952 & n3706 ) | ( ~n3707 & n3706 ) ;
  assign n3709 = ( n1958 & n2490 ) | ( n1958 & n3708 ) | ( n2490 & n3708 ) ;
  assign n3710 = ( n2490 & ~n3709 ) | ( n2490 & 1'b0 ) | ( ~n3709 & 1'b0 ) ;
  assign n3711 = ( n3708 & ~n540 ) | ( n3708 & n3710 ) | ( ~n540 & n3710 ) ;
  assign n3712 = ( n540 & ~n3708 ) | ( n540 & n3710 ) | ( ~n3708 & n3710 ) ;
  assign n3713 = ( n3711 & ~n3710 ) | ( n3711 & n3712 ) | ( ~n3710 & n3712 ) ;
  assign n3714 = n540 &  n2187 ;
  assign n3715 = ( n3621 & ~n2365 ) | ( n3621 & n3623 ) | ( ~n2365 & n3623 ) ;
  assign n3716 = ( n2365 & ~n3714 ) | ( n2365 & n3715 ) | ( ~n3714 & n3715 ) ;
  assign n3717 = ( n3714 & ~n2365 ) | ( n3714 & n3715 ) | ( ~n2365 & n3715 ) ;
  assign n3718 = ( n3716 & ~n3715 ) | ( n3716 & n3717 ) | ( ~n3715 & n3717 ) ;
  assign n3720 = ( n1906 & ~n2454 ) | ( n1906 & 1'b0 ) | ( ~n2454 & 1'b0 ) ;
  assign n3721 = ( n1911 & ~n2691 ) | ( n1911 & 1'b0 ) | ( ~n2691 & 1'b0 ) ;
  assign n3722 = n3720 | n3721 ;
  assign n3719 = ( n260 & ~n2674 ) | ( n260 & 1'b0 ) | ( ~n2674 & 1'b0 ) ;
  assign n3723 = ( n2674 & ~n3722 ) | ( n2674 & n3719 ) | ( ~n3722 & n3719 ) ;
  assign n3724 = n1916 | n2722 ;
  assign n3725 = n3723 &  n3724 ;
  assign n3726 = ( x11 & ~n252 ) | ( x11 & n3725 ) | ( ~n252 & n3725 ) ;
  assign n3727 = ( x11 & ~n3725 ) | ( x11 & n252 ) | ( ~n3725 & n252 ) ;
  assign n3728 = ( n3726 & ~x11 ) | ( n3726 & n3727 ) | ( ~x11 & n3727 ) ;
  assign n3730 = ( n3713 & n3718 ) | ( n3713 & n3728 ) | ( n3718 & n3728 ) ;
  assign n3729 = ( n3718 & ~n3713 ) | ( n3718 & n3728 ) | ( ~n3713 & n3728 ) ;
  assign n3731 = ( n3713 & ~n3730 ) | ( n3713 & n3729 ) | ( ~n3730 & n3729 ) ;
  assign n3732 = ( n3637 & ~n3703 ) | ( n3637 & n3731 ) | ( ~n3703 & n3731 ) ;
  assign n3733 = ( n3637 & ~n3731 ) | ( n3637 & n3703 ) | ( ~n3731 & n3703 ) ;
  assign n3734 = ( n3732 & ~n3637 ) | ( n3732 & n3733 ) | ( ~n3637 & n3733 ) ;
  assign n3688 = ( n2459 & ~n3233 ) | ( n2459 & 1'b0 ) | ( ~n3233 & 1'b0 ) ;
  assign n3689 = ( n2470 & ~n3336 ) | ( n2470 & 1'b0 ) | ( ~n3336 & 1'b0 ) ;
  assign n3690 = n3688 | n3689 ;
  assign n3691 = ( x5 & ~n3690 ) | ( x5 & n1074 ) | ( ~n3690 & n1074 ) ;
  assign n3692 = ( x5 & ~n1074 ) | ( x5 & n3690 ) | ( ~n1074 & n3690 ) ;
  assign n3693 = ( n3691 & ~x5 ) | ( n3691 & n3692 ) | ( ~x5 & n3692 ) ;
  assign n3735 = ( n3641 & ~n3734 ) | ( n3641 & n3693 ) | ( ~n3734 & n3693 ) ;
  assign n3736 = ( n3693 & ~n3641 ) | ( n3693 & n3734 ) | ( ~n3641 & n3734 ) ;
  assign n3737 = ( n3735 & ~n3693 ) | ( n3735 & n3736 ) | ( ~n3693 & n3736 ) ;
  assign n3739 = ( n3686 & n3687 ) | ( n3686 & n3737 ) | ( n3687 & n3737 ) ;
  assign n3738 = ( n3687 & ~n3686 ) | ( n3687 & n3737 ) | ( ~n3686 & n3737 ) ;
  assign n3740 = ( n3686 & ~n3739 ) | ( n3686 & n3738 ) | ( ~n3739 & n3738 ) ;
  assign n3741 = ( n3685 & ~n3667 ) | ( n3685 & n3740 ) | ( ~n3667 & n3740 ) ;
  assign n3742 = ( n3667 & ~n3685 ) | ( n3667 & n3740 ) | ( ~n3685 & n3740 ) ;
  assign n3743 = ( n3741 & ~n3740 ) | ( n3741 & n3742 ) | ( ~n3740 & n3742 ) ;
  assign n3744 = ( n3663 & ~n3666 ) | ( n3663 & n3743 ) | ( ~n3666 & n3743 ) ;
  assign n3745 = ( n3663 & ~n3743 ) | ( n3663 & n3666 ) | ( ~n3743 & n3666 ) ;
  assign n3746 = ( n3744 & ~n3663 ) | ( n3744 & n3745 ) | ( ~n3663 & n3745 ) ;
  assign n3747 = n3663 &  n3743 ;
  assign n3748 = n3663 | n3743 ;
  assign n3749 = ( n3665 & ~n3748 ) | ( n3665 & n3747 ) | ( ~n3748 & n3747 ) ;
  assign n3750 = n3195 | n3749 ;
  assign n3751 = ( n3667 & ~n3740 ) | ( n3667 & n3685 ) | ( ~n3740 & n3685 ) ;
  assign n3752 = n475 | n2168 ;
  assign n3753 = ( n3586 & ~n831 ) | ( n3586 & n3752 ) | ( ~n831 & n3752 ) ;
  assign n3754 = n831 | n3753 ;
  assign n3755 = ( n3675 & ~n105 ) | ( n3675 & n3754 ) | ( ~n105 & n3754 ) ;
  assign n3756 = n105 | n3755 ;
  assign n3757 = ( n167 & ~n411 ) | ( n167 & n3756 ) | ( ~n411 & n3756 ) ;
  assign n3758 = n411 | n3757 ;
  assign n3759 = ( n889 & ~n192 ) | ( n889 & n3758 ) | ( ~n192 & n3758 ) ;
  assign n3760 = n192 | n3759 ;
  assign n3761 = n142 | n3760 ;
  assign n3762 = n316 | n3761 ;
  assign n3764 = n2200 &  n2941 ;
  assign n3765 = ( n2204 & ~n3113 ) | ( n2204 & 1'b0 ) | ( ~n3113 & 1'b0 ) ;
  assign n3766 = n3764 | n3765 ;
  assign n3763 = ( n2194 & ~n3233 ) | ( n2194 & 1'b0 ) | ( ~n3233 & 1'b0 ) ;
  assign n3767 = ( n3233 & ~n3766 ) | ( n3233 & n3763 ) | ( ~n3766 & n3763 ) ;
  assign n3768 = ( n2213 & ~n3767 ) | ( n2213 & n3242 ) | ( ~n3767 & n3242 ) ;
  assign n3769 = ( n3242 & ~n3768 ) | ( n3242 & 1'b0 ) | ( ~n3768 & 1'b0 ) ;
  assign n3771 = ( n248 & n3767 ) | ( n248 & n3769 ) | ( n3767 & n3769 ) ;
  assign n3770 = ( n248 & ~n3769 ) | ( n248 & n3767 ) | ( ~n3769 & n3767 ) ;
  assign n3772 = ( n3769 & ~n3771 ) | ( n3769 & n3770 ) | ( ~n3771 & n3770 ) ;
  assign n3776 = n2454 &  n1952 ;
  assign n3773 = n1967 &  n2461 ;
  assign n3774 = ( n1947 & ~n2464 ) | ( n1947 & 1'b0 ) | ( ~n2464 & 1'b0 ) ;
  assign n3775 = n3773 | n3774 ;
  assign n3777 = ( n1952 & ~n3776 ) | ( n1952 & n3775 ) | ( ~n3776 & n3775 ) ;
  assign n3778 = n1958 | n2476 ;
  assign n3779 = ~n3777 & n3778 ;
  assign n3780 = ( n540 & ~n2341 ) | ( n540 & 1'b0 ) | ( ~n2341 & 1'b0 ) ;
  assign n3781 = ( n2365 & ~n1077 ) | ( n2365 & n3780 ) | ( ~n1077 & n3780 ) ;
  assign n3782 = ( n1077 & ~n3780 ) | ( n1077 & n2365 ) | ( ~n3780 & n2365 ) ;
  assign n3783 = ( n3781 & ~n2365 ) | ( n3781 & n3782 ) | ( ~n2365 & n3782 ) ;
  assign n3784 = ( n540 & n3779 ) | ( n540 & n3783 ) | ( n3779 & n3783 ) ;
  assign n3785 = ( n540 & ~n3779 ) | ( n540 & n3783 ) | ( ~n3779 & n3783 ) ;
  assign n3786 = ( n3779 & ~n3784 ) | ( n3779 & n3785 ) | ( ~n3784 & n3785 ) ;
  assign n3787 = ( n3717 & ~n3786 ) | ( n3717 & 1'b0 ) | ( ~n3786 & 1'b0 ) ;
  assign n3788 = n3717 | n3786 ;
  assign n3789 = ( n3787 & ~n3717 ) | ( n3787 & n3788 ) | ( ~n3717 & n3788 ) ;
  assign n3795 = n2697 | n1916 ;
  assign n3793 = n2688 | n260 ;
  assign n3790 = ( n1906 & ~n2691 ) | ( n1906 & 1'b0 ) | ( ~n2691 & 1'b0 ) ;
  assign n3791 = ( n1911 & ~n2674 ) | ( n1911 & 1'b0 ) | ( ~n2674 & 1'b0 ) ;
  assign n3792 = n3790 | n3791 ;
  assign n3794 = ( n3793 & ~n260 ) | ( n3793 & n3792 ) | ( ~n260 & n3792 ) ;
  assign n3796 = ( n3795 & ~n1916 ) | ( n3795 & n3794 ) | ( ~n1916 & n3794 ) ;
  assign n3797 = ( n883 & ~n3796 ) | ( n883 & 1'b0 ) | ( ~n3796 & 1'b0 ) ;
  assign n3798 = ~n883 & n3796 ;
  assign n3799 = n3797 | n3798 ;
  assign n3801 = ( n3729 & n3789 ) | ( n3729 & n3799 ) | ( n3789 & n3799 ) ;
  assign n3800 = ( n3729 & ~n3789 ) | ( n3729 & n3799 ) | ( ~n3789 & n3799 ) ;
  assign n3802 = ( n3789 & ~n3801 ) | ( n3789 & n3800 ) | ( ~n3801 & n3800 ) ;
  assign n3804 = ( n3733 & n3772 ) | ( n3733 & n3802 ) | ( n3772 & n3802 ) ;
  assign n3803 = ( n3733 & ~n3772 ) | ( n3733 & n3802 ) | ( ~n3772 & n3802 ) ;
  assign n3805 = ( n3772 & ~n3804 ) | ( n3772 & n3803 ) | ( ~n3804 & n3803 ) ;
  assign n3806 = ( n3686 & ~n3687 ) | ( n3686 & n3737 ) | ( ~n3687 & n3737 ) ;
  assign n3807 = ( n3805 & ~n3736 ) | ( n3805 & n3806 ) | ( ~n3736 & n3806 ) ;
  assign n3808 = ( n3736 & ~n3805 ) | ( n3736 & n3806 ) | ( ~n3805 & n3806 ) ;
  assign n3809 = ( n3807 & ~n3806 ) | ( n3807 & n3808 ) | ( ~n3806 & n3808 ) ;
  assign n3811 = ( n3751 & n3762 ) | ( n3751 & n3809 ) | ( n3762 & n3809 ) ;
  assign n3810 = ( n3762 & ~n3751 ) | ( n3762 & n3809 ) | ( ~n3751 & n3809 ) ;
  assign n3812 = ( n3751 & ~n3811 ) | ( n3751 & n3810 ) | ( ~n3811 & n3810 ) ;
  assign n3814 = ( n3747 & n3750 ) | ( n3747 & n3812 ) | ( n3750 & n3812 ) ;
  assign n3813 = ( n3750 & ~n3747 ) | ( n3750 & n3812 ) | ( ~n3747 & n3812 ) ;
  assign n3815 = ( n3747 & ~n3814 ) | ( n3747 & n3813 ) | ( ~n3814 & n3813 ) ;
  assign n3816 = ( n3747 & ~n3812 ) | ( n3747 & 1'b0 ) | ( ~n3812 & 1'b0 ) ;
  assign n3817 = ~n3747 & n3812 ;
  assign n3818 = ( n3749 & n3816 ) | ( n3749 & n3817 ) | ( n3816 & n3817 ) ;
  assign n3819 = n3195 | n3818 ;
  assign n3878 = n248 &  n3801 ;
  assign n3877 = ( n248 & ~n3801 ) | ( n248 & 1'b0 ) | ( ~n3801 & 1'b0 ) ;
  assign n3879 = ( n3801 & ~n3878 ) | ( n3801 & n3877 ) | ( ~n3878 & n3877 ) ;
  assign n3840 = ( n1077 & n2365 ) | ( n1077 & n3780 ) | ( n2365 & n3780 ) ;
  assign n3841 = n540 &  n2461 ;
  assign n3842 = n1952 | n2691 ;
  assign n3843 = ( n1967 & ~n2464 ) | ( n1967 & 1'b0 ) | ( ~n2464 & 1'b0 ) ;
  assign n3844 = ( n1947 & ~n2454 ) | ( n1947 & 1'b0 ) | ( ~n2454 & 1'b0 ) ;
  assign n3845 = n3843 | n3844 ;
  assign n3846 = ( n3842 & ~n2691 ) | ( n3842 & n3845 ) | ( ~n2691 & n3845 ) ;
  assign n3847 = ( n1958 & ~n2734 ) | ( n1958 & n3846 ) | ( ~n2734 & n3846 ) ;
  assign n3848 = n2734 | n3847 ;
  assign n3849 = ( n540 & ~n3846 ) | ( n540 & n3848 ) | ( ~n3846 & n3848 ) ;
  assign n3850 = ( n3846 & ~n540 ) | ( n3846 & n3848 ) | ( ~n540 & n3848 ) ;
  assign n3851 = ( n3849 & ~n3848 ) | ( n3849 & n3850 ) | ( ~n3848 & n3850 ) ;
  assign n3852 = ( n3840 & n3841 ) | ( n3840 & n3851 ) | ( n3841 & n3851 ) ;
  assign n3853 = ( n3841 & ~n3840 ) | ( n3841 & n3851 ) | ( ~n3840 & n3851 ) ;
  assign n3854 = ( n3840 & ~n3852 ) | ( n3840 & n3853 ) | ( ~n3852 & n3853 ) ;
  assign n3862 = n2941 | n260 ;
  assign n3859 = ( n1906 & ~n2674 ) | ( n1906 & 1'b0 ) | ( ~n2674 & 1'b0 ) ;
  assign n3860 = n1911 &  n2688 ;
  assign n3861 = n3859 | n3860 ;
  assign n3863 = ( n3862 & ~n260 ) | ( n3862 & n3861 ) | ( ~n260 & n3861 ) ;
  assign n3864 = n1916 | n2944 ;
  assign n3865 = ~n3863 & n3864 ;
  assign n3866 = ( x11 & ~n252 ) | ( x11 & n3865 ) | ( ~n252 & n3865 ) ;
  assign n3867 = ( x11 & ~n3865 ) | ( x11 & n252 ) | ( ~n3865 & n252 ) ;
  assign n3868 = ( n3866 & ~x11 ) | ( n3866 & n3867 ) | ( ~x11 & n3867 ) ;
  assign n3855 = ( x14 & n537 ) | ( x14 & n3779 ) | ( n537 & n3779 ) ;
  assign n3856 = ( x14 & ~n3779 ) | ( x14 & n537 ) | ( ~n3779 & n537 ) ;
  assign n3857 = ( n3779 & ~n3855 ) | ( n3779 & n3856 ) | ( ~n3855 & n3856 ) ;
  assign n3858 = ( n3717 & ~n3857 ) | ( n3717 & n3783 ) | ( ~n3857 & n3783 ) ;
  assign n3869 = ( n3854 & ~n3868 ) | ( n3854 & n3858 ) | ( ~n3868 & n3858 ) ;
  assign n3870 = ( n3854 & ~n3858 ) | ( n3854 & n3868 ) | ( ~n3858 & n3868 ) ;
  assign n3871 = ( n3869 & ~n3854 ) | ( n3869 & n3870 ) | ( ~n3854 & n3870 ) ;
  assign n3875 = n3339 | n2213 ;
  assign n3872 = ( n2200 & ~n3113 ) | ( n2200 & 1'b0 ) | ( ~n3113 & 1'b0 ) ;
  assign n3873 = ( n2204 & ~n3233 ) | ( n2204 & 1'b0 ) | ( ~n3233 & 1'b0 ) ;
  assign n3874 = n3872 | n3873 ;
  assign n3876 = ( n3875 & ~n2213 ) | ( n3875 & n3874 ) | ( ~n2213 & n3874 ) ;
  assign n3881 = ( n3871 & n3876 ) | ( n3871 & n3879 ) | ( n3876 & n3879 ) ;
  assign n3880 = ( n3871 & ~n3879 ) | ( n3871 & n3876 ) | ( ~n3879 & n3876 ) ;
  assign n3882 = ( n3879 & ~n3881 ) | ( n3879 & n3880 ) | ( ~n3881 & n3880 ) ;
  assign n3883 = ( n3804 & n3807 ) | ( n3804 & n3882 ) | ( n3807 & n3882 ) ;
  assign n3884 = ( n3804 & ~n3807 ) | ( n3804 & n3882 ) | ( ~n3807 & n3882 ) ;
  assign n3885 = ( n3807 & ~n3883 ) | ( n3807 & n3884 ) | ( ~n3883 & n3884 ) ;
  assign n3829 = n295 | n1702 ;
  assign n3830 = ( n3035 & ~n306 ) | ( n3035 & n3829 ) | ( ~n306 & n3829 ) ;
  assign n3831 = n306 | n3830 ;
  assign n3820 = ~n268 & n1866 ;
  assign n3821 = ( n195 & ~n380 ) | ( n195 & n3820 ) | ( ~n380 & n3820 ) ;
  assign n3822 = ( n139 & ~n195 ) | ( n139 & n3821 ) | ( ~n195 & n3821 ) ;
  assign n3823 = ~n139 & n3822 ;
  assign n3824 = ( n141 & ~n199 ) | ( n141 & n3823 ) | ( ~n199 & n3823 ) ;
  assign n3825 = ~n141 & n3824 ;
  assign n3826 = ( n78 & ~n277 ) | ( n78 & n3825 ) | ( ~n277 & n3825 ) ;
  assign n3827 = ~n78 & n3826 ;
  assign n3828 = ~n185 & n3827 ;
  assign n3832 = ( n352 & ~n3831 ) | ( n352 & n3828 ) | ( ~n3831 & n3828 ) ;
  assign n3833 = ~n352 & n3832 ;
  assign n3834 = ( n181 & ~n229 ) | ( n181 & n3833 ) | ( ~n229 & n3833 ) ;
  assign n3835 = ~n181 & n3834 ;
  assign n3836 = ( n198 & ~n595 ) | ( n198 & n3835 ) | ( ~n595 & n3835 ) ;
  assign n3837 = ~n198 & n3836 ;
  assign n3838 = ~n612 & n3837 ;
  assign n3839 = ~n281 & n3838 ;
  assign n3886 = ( n3810 & n3839 ) | ( n3810 & n3885 ) | ( n3839 & n3885 ) ;
  assign n3887 = ( n3810 & ~n3885 ) | ( n3810 & n3839 ) | ( ~n3885 & n3839 ) ;
  assign n3888 = ( n3885 & ~n3886 ) | ( n3885 & n3887 ) | ( ~n3886 & n3887 ) ;
  assign n3890 = ( n3816 & n3819 ) | ( n3816 & n3888 ) | ( n3819 & n3888 ) ;
  assign n3889 = ( n3819 & ~n3816 ) | ( n3819 & n3888 ) | ( ~n3816 & n3888 ) ;
  assign n3891 = ( n3816 & ~n3890 ) | ( n3816 & n3889 ) | ( ~n3890 & n3889 ) ;
  assign n3892 = ( n3816 & ~n3888 ) | ( n3816 & 1'b0 ) | ( ~n3888 & 1'b0 ) ;
  assign n3893 = ~n3816 & n3888 ;
  assign n3894 = ( n3818 & n3892 ) | ( n3818 & n3893 ) | ( n3892 & n3893 ) ;
  assign n3895 = n3195 | n3894 ;
  assign n3914 = n1952 | n2674 ;
  assign n3915 = ( n1967 & ~n2454 ) | ( n1967 & 1'b0 ) | ( ~n2454 & 1'b0 ) ;
  assign n3916 = ( n1947 & ~n2691 ) | ( n1947 & 1'b0 ) | ( ~n2691 & 1'b0 ) ;
  assign n3917 = n3915 | n3916 ;
  assign n3918 = ( n3914 & ~n2674 ) | ( n3914 & n3917 ) | ( ~n2674 & n3917 ) ;
  assign n3919 = n1958 | n2722 ;
  assign n3920 = ~n3918 & n3919 ;
  assign n3921 = ( n540 & ~n2461 ) | ( n540 & 1'b0 ) | ( ~n2461 & 1'b0 ) ;
  assign n3922 = ( n540 & ~n2464 ) | ( n540 & 1'b0 ) | ( ~n2464 & 1'b0 ) ;
  assign n3923 = ( n3920 & ~n3921 ) | ( n3920 & n3922 ) | ( ~n3921 & n3922 ) ;
  assign n3924 = ( n3921 & ~n3920 ) | ( n3921 & n3922 ) | ( ~n3920 & n3922 ) ;
  assign n3925 = ( n3923 & ~n3922 ) | ( n3923 & n3924 ) | ( ~n3922 & n3924 ) ;
  assign n3926 = n1906 &  n2688 ;
  assign n3927 = n1911 &  n2941 ;
  assign n3928 = n3926 | n3927 ;
  assign n3929 = ~n260 & n3113 ;
  assign n3930 = ( n260 & ~n3928 ) | ( n260 & n3929 ) | ( ~n3928 & n3929 ) ;
  assign n3931 = n1916 | n3484 ;
  assign n3932 = n3930 &  n3931 ;
  assign n3933 = ( x11 & ~n252 ) | ( x11 & n3932 ) | ( ~n252 & n3932 ) ;
  assign n3934 = ( x11 & ~n3932 ) | ( x11 & n252 ) | ( ~n3932 & n252 ) ;
  assign n3935 = ( n3933 & ~x11 ) | ( n3933 & n3934 ) | ( ~x11 & n3934 ) ;
  assign n3936 = ( n3853 & n3925 ) | ( n3853 & n3935 ) | ( n3925 & n3935 ) ;
  assign n3937 = ( n3853 & ~n3925 ) | ( n3853 & n3935 ) | ( ~n3925 & n3935 ) ;
  assign n3938 = ( n3925 & ~n3936 ) | ( n3925 & n3937 ) | ( ~n3936 & n3937 ) ;
  assign n3939 = ( n2200 & ~n3233 ) | ( n2200 & 1'b0 ) | ( ~n3233 & 1'b0 ) ;
  assign n3940 = n2213 | n3336 ;
  assign n3941 = ~n3939 & n3940 ;
  assign n3942 = n248 &  n3941 ;
  assign n3943 = n248 | n3941 ;
  assign n3944 = ~n3942 & n3943 ;
  assign n3946 = ( n3869 & n3938 ) | ( n3869 & n3944 ) | ( n3938 & n3944 ) ;
  assign n3945 = ( n3938 & ~n3869 ) | ( n3938 & n3944 ) | ( ~n3869 & n3944 ) ;
  assign n3947 = ( n3869 & ~n3946 ) | ( n3869 & n3945 ) | ( ~n3946 & n3945 ) ;
  assign n3909 = ~n248 & n3876 ;
  assign n3910 = ( n248 & ~n3876 ) | ( n248 & 1'b0 ) | ( ~n3876 & 1'b0 ) ;
  assign n3911 = n3909 | n3910 ;
  assign n3912 = ( n3801 & ~n3911 ) | ( n3801 & n3871 ) | ( ~n3911 & n3871 ) ;
  assign n3913 = ( n3804 & ~n3882 ) | ( n3804 & n3807 ) | ( ~n3882 & n3807 ) ;
  assign n3949 = ( n3912 & n3913 ) | ( n3912 & n3947 ) | ( n3913 & n3947 ) ;
  assign n3948 = ( n3912 & ~n3947 ) | ( n3912 & n3913 ) | ( ~n3947 & n3913 ) ;
  assign n3950 = ( n3947 & ~n3949 ) | ( n3947 & n3948 ) | ( ~n3949 & n3948 ) ;
  assign n3896 = ( n3810 & ~n3839 ) | ( n3810 & n3885 ) | ( ~n3839 & n3885 ) ;
  assign n3897 = n397 | n831 ;
  assign n3898 = ( n2645 & ~n178 ) | ( n2645 & n3897 ) | ( ~n178 & n3897 ) ;
  assign n3899 = n178 | n3898 ;
  assign n3900 = ( n1814 & n2675 ) | ( n1814 & n3899 ) | ( n2675 & n3899 ) ;
  assign n3901 = ( n1814 & ~n3900 ) | ( n1814 & 1'b0 ) | ( ~n3900 & 1'b0 ) ;
  assign n3902 = ( n276 & ~n310 ) | ( n276 & n3901 ) | ( ~n310 & n3901 ) ;
  assign n3903 = ~n276 & n3902 ;
  assign n3904 = ( n109 & ~n199 ) | ( n109 & n3903 ) | ( ~n199 & n3903 ) ;
  assign n3905 = ~n109 & n3904 ;
  assign n3906 = ( n208 & ~n266 ) | ( n208 & n3905 ) | ( ~n266 & n3905 ) ;
  assign n3907 = ~n208 & n3906 ;
  assign n3908 = ~n190 & n3907 ;
  assign n3952 = ( n3896 & n3908 ) | ( n3896 & n3950 ) | ( n3908 & n3950 ) ;
  assign n3951 = ( n3896 & ~n3950 ) | ( n3896 & n3908 ) | ( ~n3950 & n3908 ) ;
  assign n3953 = ( n3950 & ~n3952 ) | ( n3950 & n3951 ) | ( ~n3952 & n3951 ) ;
  assign n3954 = ( n3892 & ~n3895 ) | ( n3892 & n3953 ) | ( ~n3895 & n3953 ) ;
  assign n3955 = ( n3892 & ~n3953 ) | ( n3892 & n3895 ) | ( ~n3953 & n3895 ) ;
  assign n3956 = ( n3954 & ~n3892 ) | ( n3954 & n3955 ) | ( ~n3892 & n3955 ) ;
  assign n3957 = n3892 &  n3953 ;
  assign n3958 = n3892 | n3953 ;
  assign n3959 = ( n3894 & ~n3958 ) | ( n3894 & n3957 ) | ( ~n3958 & n3957 ) ;
  assign n3960 = n3195 | n3959 ;
  assign n3973 = ( n3869 & ~n3944 ) | ( n3869 & n3938 ) | ( ~n3944 & n3938 ) ;
  assign n3974 = ( n540 & ~n2454 ) | ( n540 & 1'b0 ) | ( ~n2454 & 1'b0 ) ;
  assign n3975 = ( n248 & n3841 ) | ( n248 & n3974 ) | ( n3841 & n3974 ) ;
  assign n3976 = ( n248 & ~n3974 ) | ( n248 & n3841 ) | ( ~n3974 & n3841 ) ;
  assign n3977 = ( n3974 & ~n3975 ) | ( n3974 & n3976 ) | ( ~n3975 & n3976 ) ;
  assign n3978 = ( n2461 & ~n3920 ) | ( n2461 & n2464 ) | ( ~n3920 & n2464 ) ;
  assign n3979 = ( n540 & ~n3978 ) | ( n540 & 1'b0 ) | ( ~n3978 & 1'b0 ) ;
  assign n3980 = ~n540 & n3920 ;
  assign n3981 = ( n540 & ~n3979 ) | ( n540 & n3980 ) | ( ~n3979 & n3980 ) ;
  assign n3985 = ~n2688 & n1952 ;
  assign n3982 = ( n1967 & ~n2691 ) | ( n1967 & 1'b0 ) | ( ~n2691 & 1'b0 ) ;
  assign n3983 = ( n1947 & ~n2674 ) | ( n1947 & 1'b0 ) | ( ~n2674 & 1'b0 ) ;
  assign n3984 = n3982 | n3983 ;
  assign n3986 = ( n1952 & ~n3985 ) | ( n1952 & n3984 ) | ( ~n3985 & n3984 ) ;
  assign n3987 = ~n1958 & n2697 ;
  assign n3988 = n3986 | n3987 ;
  assign n3989 = n540 | n3988 ;
  assign n3990 = n540 &  n3988 ;
  assign n3991 = ( n3989 & ~n3990 ) | ( n3989 & 1'b0 ) | ( ~n3990 & 1'b0 ) ;
  assign n3993 = ( n3977 & n3981 ) | ( n3977 & n3991 ) | ( n3981 & n3991 ) ;
  assign n3992 = ( n3981 & ~n3977 ) | ( n3981 & n3991 ) | ( ~n3977 & n3991 ) ;
  assign n3994 = ( n3977 & ~n3993 ) | ( n3977 & n3992 ) | ( ~n3993 & n3992 ) ;
  assign n3996 = n1906 &  n2941 ;
  assign n3997 = ( n1911 & ~n3113 ) | ( n1911 & 1'b0 ) | ( ~n3113 & 1'b0 ) ;
  assign n3998 = n3996 | n3997 ;
  assign n3995 = ( n260 & ~n3233 ) | ( n260 & 1'b0 ) | ( ~n3233 & 1'b0 ) ;
  assign n3999 = ( n3233 & ~n3998 ) | ( n3233 & n3995 ) | ( ~n3998 & n3995 ) ;
  assign n4000 = ( n1916 & ~n3999 ) | ( n1916 & n3242 ) | ( ~n3999 & n3242 ) ;
  assign n4001 = ( n3242 & ~n4000 ) | ( n3242 & 1'b0 ) | ( ~n4000 & 1'b0 ) ;
  assign n4002 = ( n883 & ~n3999 ) | ( n883 & n4001 ) | ( ~n3999 & n4001 ) ;
  assign n4003 = ( n3999 & ~n883 ) | ( n3999 & n4001 ) | ( ~n883 & n4001 ) ;
  assign n4004 = ( n4002 & ~n4001 ) | ( n4002 & n4003 ) | ( ~n4001 & n4003 ) ;
  assign n4005 = ( n3937 & n3994 ) | ( n3937 & n4004 ) | ( n3994 & n4004 ) ;
  assign n4006 = ( n3994 & ~n3937 ) | ( n3994 & n4004 ) | ( ~n3937 & n4004 ) ;
  assign n4007 = ( n3937 & ~n4005 ) | ( n3937 & n4006 ) | ( ~n4005 & n4006 ) ;
  assign n4009 = ( n3949 & n3973 ) | ( n3949 & n4007 ) | ( n3973 & n4007 ) ;
  assign n4008 = ( n3973 & ~n3949 ) | ( n3973 & n4007 ) | ( ~n3949 & n4007 ) ;
  assign n4010 = ( n3949 & ~n4009 ) | ( n3949 & n4008 ) | ( ~n4009 & n4008 ) ;
  assign n3961 = ( n3908 & ~n3896 ) | ( n3908 & n3950 ) | ( ~n3896 & n3950 ) ;
  assign n3962 = n231 | n656 ;
  assign n3963 = ( n615 & ~n360 ) | ( n615 & n3962 ) | ( ~n360 & n3962 ) ;
  assign n3964 = n360 | n3963 ;
  assign n3965 = ( n3023 & ~n184 ) | ( n3023 & n3964 ) | ( ~n184 & n3964 ) ;
  assign n3966 = n184 | n3965 ;
  assign n3967 = ( n2675 & ~n902 ) | ( n2675 & n3966 ) | ( ~n902 & n3966 ) ;
  assign n3968 = n902 | n3967 ;
  assign n3969 = ( n304 & ~n443 ) | ( n304 & n3968 ) | ( ~n443 & n3968 ) ;
  assign n3970 = n443 | n3969 ;
  assign n3971 = n488 | n3970 ;
  assign n3972 = n275 | n3971 ;
  assign n4012 = ( n3961 & n3972 ) | ( n3961 & n4010 ) | ( n3972 & n4010 ) ;
  assign n4011 = ( n3961 & ~n4010 ) | ( n3961 & n3972 ) | ( ~n4010 & n3972 ) ;
  assign n4013 = ( n4010 & ~n4012 ) | ( n4010 & n4011 ) | ( ~n4012 & n4011 ) ;
  assign n4015 = ( n3957 & n3960 ) | ( n3957 & n4013 ) | ( n3960 & n4013 ) ;
  assign n4014 = ( n3960 & ~n3957 ) | ( n3960 & n4013 ) | ( ~n3957 & n4013 ) ;
  assign n4016 = ( n3957 & ~n4015 ) | ( n3957 & n4014 ) | ( ~n4015 & n4014 ) ;
  assign n4017 = ( n3957 & ~n4013 ) | ( n3957 & 1'b0 ) | ( ~n4013 & 1'b0 ) ;
  assign n4018 = ~n3957 & n4013 ;
  assign n4019 = ( n3959 & n4017 ) | ( n3959 & n4018 ) | ( n4017 & n4018 ) ;
  assign n4020 = n3195 | n4019 ;
  assign n4028 = ( n3949 & ~n3973 ) | ( n3949 & n4007 ) | ( ~n3973 & n4007 ) ;
  assign n4029 = ( n3977 & ~n3991 ) | ( n3977 & n3981 ) | ( ~n3991 & n3981 ) ;
  assign n4030 = ( n540 & ~n2691 ) | ( n540 & 1'b0 ) | ( ~n2691 & 1'b0 ) ;
  assign n4035 = ~n2941 & n1952 ;
  assign n4032 = ( n1967 & ~n2674 ) | ( n1967 & 1'b0 ) | ( ~n2674 & 1'b0 ) ;
  assign n4033 = n1947 &  n2688 ;
  assign n4034 = n4032 | n4033 ;
  assign n4036 = ( n1952 & ~n4035 ) | ( n1952 & n4034 ) | ( ~n4035 & n4034 ) ;
  assign n4037 = ( n1958 & ~n2944 ) | ( n1958 & n4036 ) | ( ~n2944 & n4036 ) ;
  assign n4038 = n2944 | n4037 ;
  assign n4039 = ( n540 & ~n4036 ) | ( n540 & n4038 ) | ( ~n4036 & n4038 ) ;
  assign n4040 = ( n4036 & ~n540 ) | ( n4036 & n4038 ) | ( ~n540 & n4038 ) ;
  assign n4041 = ( n4039 & ~n4038 ) | ( n4039 & n4040 ) | ( ~n4038 & n4040 ) ;
  assign n4031 = ( n3841 & ~n248 ) | ( n3841 & n3974 ) | ( ~n248 & n3974 ) ;
  assign n4042 = ( n4030 & ~n4041 ) | ( n4030 & n4031 ) | ( ~n4041 & n4031 ) ;
  assign n4043 = ( n4030 & ~n4031 ) | ( n4030 & n4041 ) | ( ~n4031 & n4041 ) ;
  assign n4044 = ( n4042 & ~n4030 ) | ( n4042 & n4043 ) | ( ~n4030 & n4043 ) ;
  assign n4048 = n3339 | n1916 ;
  assign n4045 = ( n1906 & ~n3113 ) | ( n1906 & 1'b0 ) | ( ~n3113 & 1'b0 ) ;
  assign n4046 = ( n1911 & ~n3233 ) | ( n1911 & 1'b0 ) | ( ~n3233 & 1'b0 ) ;
  assign n4047 = n4045 | n4046 ;
  assign n4049 = ( n4048 & ~n1916 ) | ( n4048 & n4047 ) | ( ~n1916 & n4047 ) ;
  assign n4050 = ~n883 & n4049 ;
  assign n4051 = ( n883 & ~n4049 ) | ( n883 & 1'b0 ) | ( ~n4049 & 1'b0 ) ;
  assign n4052 = n4050 | n4051 ;
  assign n4054 = ( n4029 & n4044 ) | ( n4029 & n4052 ) | ( n4044 & n4052 ) ;
  assign n4053 = ( n4044 & ~n4029 ) | ( n4044 & n4052 ) | ( ~n4029 & n4052 ) ;
  assign n4055 = ( n4029 & ~n4054 ) | ( n4029 & n4053 ) | ( ~n4054 & n4053 ) ;
  assign n4056 = ( n4028 & ~n4006 ) | ( n4028 & n4055 ) | ( ~n4006 & n4055 ) ;
  assign n4057 = ( n4006 & ~n4055 ) | ( n4006 & n4028 ) | ( ~n4055 & n4028 ) ;
  assign n4058 = ( n4056 & ~n4028 ) | ( n4056 & n4057 ) | ( ~n4028 & n4057 ) ;
  assign n4021 = ( n3972 & ~n3961 ) | ( n3972 & n4010 ) | ( ~n3961 & n4010 ) ;
  assign n4022 = n280 | n454 ;
  assign n4023 = ( n3097 & ~n726 ) | ( n3097 & n4022 ) | ( ~n726 & n4022 ) ;
  assign n4024 = n726 | n4023 ;
  assign n4025 = ( n671 & ~n827 ) | ( n671 & n4024 ) | ( ~n827 & n4024 ) ;
  assign n4026 = ( n636 & n827 ) | ( n636 & n4025 ) | ( n827 & n4025 ) ;
  assign n4027 = ( n636 & ~n4026 ) | ( n636 & 1'b0 ) | ( ~n4026 & 1'b0 ) ;
  assign n4060 = ( n4021 & n4027 ) | ( n4021 & n4058 ) | ( n4027 & n4058 ) ;
  assign n4059 = ( n4021 & ~n4058 ) | ( n4021 & n4027 ) | ( ~n4058 & n4027 ) ;
  assign n4061 = ( n4058 & ~n4060 ) | ( n4058 & n4059 ) | ( ~n4060 & n4059 ) ;
  assign n4062 = ( n4017 & ~n4020 ) | ( n4017 & n4061 ) | ( ~n4020 & n4061 ) ;
  assign n4063 = ( n4017 & ~n4061 ) | ( n4017 & n4020 ) | ( ~n4061 & n4020 ) ;
  assign n4064 = ( n4062 & ~n4017 ) | ( n4062 & n4063 ) | ( ~n4017 & n4063 ) ;
  assign n4065 = n4017 &  n4061 ;
  assign n4066 = n4017 | n4061 ;
  assign n4067 = ( n4019 & ~n4066 ) | ( n4019 & n4065 ) | ( ~n4066 & n4065 ) ;
  assign n4068 = n3195 | n4067 ;
  assign n4069 = ( n4027 & ~n4021 ) | ( n4027 & n4058 ) | ( ~n4021 & n4058 ) ;
  assign n4070 = n152 | n160 ;
  assign n4071 = ( n208 & ~n181 ) | ( n208 & n4070 ) | ( ~n181 & n4070 ) ;
  assign n4072 = n181 | n4071 ;
  assign n4073 = n501 | n4072 ;
  assign n4074 = ( n1737 & ~n500 ) | ( n1737 & n4073 ) | ( ~n500 & n4073 ) ;
  assign n4075 = n500 | n4074 ;
  assign n4076 = ( n2124 & ~n3320 ) | ( n2124 & n4075 ) | ( ~n3320 & n4075 ) ;
  assign n4077 = ( n2124 & ~n4076 ) | ( n2124 & 1'b0 ) | ( ~n4076 & 1'b0 ) ;
  assign n4078 = ( n1732 & ~n113 ) | ( n1732 & n4077 ) | ( ~n113 & n4077 ) ;
  assign n4079 = ( n110 & ~n1732 ) | ( n110 & n4078 ) | ( ~n1732 & n4078 ) ;
  assign n4080 = ~n110 & n4079 ;
  assign n4081 = ~n185 & n4080 ;
  assign n4092 = n3113 &  n1952 ;
  assign n4089 = n1967 &  n2688 ;
  assign n4090 = n1947 &  n2941 ;
  assign n4091 = n4089 | n4090 ;
  assign n4093 = ( n1952 & ~n4092 ) | ( n1952 & n4091 ) | ( ~n4092 & n4091 ) ;
  assign n4094 = n1958 | n3484 ;
  assign n4095 = ~n4093 & n4094 ;
  assign n4096 = ~n540 & n4095 ;
  assign n4097 = ( n540 & ~n4095 ) | ( n540 & 1'b0 ) | ( ~n4095 & 1'b0 ) ;
  assign n4098 = n4096 | n4097 ;
  assign n4083 = ( n1906 & ~n3233 ) | ( n1906 & 1'b0 ) | ( ~n3233 & 1'b0 ) ;
  assign n4084 = n1916 | n3336 ;
  assign n4085 = ~n4083 & n4084 ;
  assign n4086 = ( x11 & n252 ) | ( x11 & n4085 ) | ( n252 & n4085 ) ;
  assign n4087 = ( n252 & ~x11 ) | ( n252 & n4085 ) | ( ~x11 & n4085 ) ;
  assign n4088 = ( x11 & ~n4086 ) | ( x11 & n4087 ) | ( ~n4086 & n4087 ) ;
  assign n4099 = ( n540 & ~n2674 ) | ( n540 & 1'b0 ) | ( ~n2674 & 1'b0 ) ;
  assign n4100 = ( n4030 & n4043 ) | ( n4030 & n4099 ) | ( n4043 & n4099 ) ;
  assign n4101 = ( n4030 & ~n4043 ) | ( n4030 & n4099 ) | ( ~n4043 & n4099 ) ;
  assign n4102 = ( n4043 & ~n4100 ) | ( n4043 & n4101 ) | ( ~n4100 & n4101 ) ;
  assign n4104 = ( n4088 & n4098 ) | ( n4088 & n4102 ) | ( n4098 & n4102 ) ;
  assign n4103 = ( n4088 & ~n4098 ) | ( n4088 & n4102 ) | ( ~n4098 & n4102 ) ;
  assign n4105 = ( n4098 & ~n4104 ) | ( n4098 & n4103 ) | ( ~n4104 & n4103 ) ;
  assign n4082 = ( n4029 & ~n4044 ) | ( n4029 & n4052 ) | ( ~n4044 & n4052 ) ;
  assign n4106 = ( n4006 & ~n4028 ) | ( n4006 & n4055 ) | ( ~n4028 & n4055 ) ;
  assign n4107 = ( n4105 & ~n4082 ) | ( n4105 & n4106 ) | ( ~n4082 & n4106 ) ;
  assign n4108 = ( n4082 & ~n4105 ) | ( n4082 & n4106 ) | ( ~n4105 & n4106 ) ;
  assign n4109 = ( n4107 & ~n4106 ) | ( n4107 & n4108 ) | ( ~n4106 & n4108 ) ;
  assign n4110 = ( n4069 & ~n4081 ) | ( n4069 & n4109 ) | ( ~n4081 & n4109 ) ;
  assign n4111 = ( n4081 & ~n4069 ) | ( n4081 & n4109 ) | ( ~n4069 & n4109 ) ;
  assign n4112 = ( n4110 & ~n4109 ) | ( n4110 & n4111 ) | ( ~n4109 & n4111 ) ;
  assign n4114 = ( n4065 & n4068 ) | ( n4065 & n4112 ) | ( n4068 & n4112 ) ;
  assign n4113 = ( n4068 & ~n4065 ) | ( n4068 & n4112 ) | ( ~n4065 & n4112 ) ;
  assign n4115 = ( n4065 & ~n4114 ) | ( n4065 & n4113 ) | ( ~n4114 & n4113 ) ;
  assign n4116 = ( n4065 & ~n4112 ) | ( n4065 & 1'b0 ) | ( ~n4112 & 1'b0 ) ;
  assign n4117 = ~n4065 & n4112 ;
  assign n4118 = ( n4067 & n4116 ) | ( n4067 & n4117 ) | ( n4116 & n4117 ) ;
  assign n4119 = n3195 | n4118 ;
  assign n4138 = ( n4088 & ~n4102 ) | ( n4088 & n4098 ) | ( ~n4102 & n4098 ) ;
  assign n4139 = n1952 | n3233 ;
  assign n4140 = n1967 &  n2941 ;
  assign n4141 = ( n1947 & ~n3113 ) | ( n1947 & 1'b0 ) | ( ~n3113 & 1'b0 ) ;
  assign n4142 = n4140 | n4141 ;
  assign n4143 = ( n4139 & ~n3233 ) | ( n4139 & n4142 ) | ( ~n3233 & n4142 ) ;
  assign n4144 = ~n1958 & n3242 ;
  assign n4145 = n4143 | n4144 ;
  assign n4146 = n540 | n4145 ;
  assign n4147 = n540 &  n4145 ;
  assign n4148 = ( n4146 & ~n4147 ) | ( n4146 & 1'b0 ) | ( ~n4147 & 1'b0 ) ;
  assign n4150 = n540 &  n2688 ;
  assign n4151 = ( n4099 & ~n883 ) | ( n4099 & n4150 ) | ( ~n883 & n4150 ) ;
  assign n4152 = ( n883 & ~n4150 ) | ( n883 & n4099 ) | ( ~n4150 & n4099 ) ;
  assign n4153 = ( n4151 & ~n4099 ) | ( n4151 & n4152 ) | ( ~n4099 & n4152 ) ;
  assign n4149 = ( n4043 & ~n4030 ) | ( n4043 & n4099 ) | ( ~n4030 & n4099 ) ;
  assign n4154 = ( n4148 & ~n4153 ) | ( n4148 & n4149 ) | ( ~n4153 & n4149 ) ;
  assign n4155 = ( n4148 & ~n4149 ) | ( n4148 & n4153 ) | ( ~n4149 & n4153 ) ;
  assign n4156 = ( n4154 & ~n4148 ) | ( n4154 & n4155 ) | ( ~n4148 & n4155 ) ;
  assign n4158 = ( n4107 & n4138 ) | ( n4107 & n4156 ) | ( n4138 & n4156 ) ;
  assign n4157 = ( n4138 & ~n4107 ) | ( n4138 & n4156 ) | ( ~n4107 & n4156 ) ;
  assign n4159 = ( n4107 & ~n4158 ) | ( n4107 & n4157 ) | ( ~n4158 & n4157 ) ;
  assign n4120 = n167 | n324 ;
  assign n4121 = ( n293 & ~n227 ) | ( n293 & n4120 ) | ( ~n227 & n4120 ) ;
  assign n4122 = n227 | n4121 ;
  assign n4123 = n91 | n4122 ;
  assign n4124 = ( n3199 & ~n130 ) | ( n3199 & n4123 ) | ( ~n130 & n4123 ) ;
  assign n4125 = n130 | n4124 ;
  assign n4126 = ( n2417 & ~n911 ) | ( n2417 & n4125 ) | ( ~n911 & n4125 ) ;
  assign n4127 = n911 | n4126 ;
  assign n4128 = ( n3058 & ~n326 ) | ( n3058 & n4127 ) | ( ~n326 & n4127 ) ;
  assign n4129 = n326 | n4128 ;
  assign n4130 = ( n610 & ~n169 ) | ( n610 & n4129 ) | ( ~n169 & n4129 ) ;
  assign n4131 = n169 | n4130 ;
  assign n4132 = ( n229 & ~n143 ) | ( n229 & n4131 ) | ( ~n143 & n4131 ) ;
  assign n4133 = n143 | n4132 ;
  assign n4134 = ( n379 & ~n116 ) | ( n379 & n4133 ) | ( ~n116 & n4133 ) ;
  assign n4135 = n116 | n4134 ;
  assign n4136 = n361 | n4135 ;
  assign n4137 = ( n4069 & n4081 ) | ( n4069 & n4109 ) | ( n4081 & n4109 ) ;
  assign n4160 = ( n4136 & n4137 ) | ( n4136 & n4159 ) | ( n4137 & n4159 ) ;
  assign n4161 = ( n4136 & ~n4159 ) | ( n4136 & n4137 ) | ( ~n4159 & n4137 ) ;
  assign n4162 = ( n4159 & ~n4160 ) | ( n4159 & n4161 ) | ( ~n4160 & n4161 ) ;
  assign n4163 = ( n4116 & ~n4119 ) | ( n4116 & n4162 ) | ( ~n4119 & n4162 ) ;
  assign n4164 = ( n4116 & ~n4162 ) | ( n4116 & n4119 ) | ( ~n4162 & n4119 ) ;
  assign n4165 = ( n4163 & ~n4116 ) | ( n4163 & n4164 ) | ( ~n4116 & n4164 ) ;
  assign n4166 = ( n4116 & ~n4162 ) | ( n4116 & 1'b0 ) | ( ~n4162 & 1'b0 ) ;
  assign n4167 = ~n4116 & n4162 ;
  assign n4168 = ( n4118 & n4166 ) | ( n4118 & n4167 ) | ( n4166 & n4167 ) ;
  assign n4169 = n3195 | n4168 ;
  assign n4185 = ( n883 & n4099 ) | ( n883 & n4150 ) | ( n4099 & n4150 ) ;
  assign n4191 = ( n540 & ~n2941 ) | ( n540 & 1'b0 ) | ( ~n2941 & 1'b0 ) ;
  assign n4189 = n3339 | n1958 ;
  assign n4186 = ( n1967 & ~n3113 ) | ( n1967 & 1'b0 ) | ( ~n3113 & 1'b0 ) ;
  assign n4187 = ( n1947 & ~n3233 ) | ( n1947 & 1'b0 ) | ( ~n3233 & 1'b0 ) ;
  assign n4188 = n4186 | n4187 ;
  assign n4190 = ( n4189 & ~n1958 ) | ( n4189 & n4188 ) | ( ~n1958 & n4188 ) ;
  assign n4192 = ( n4185 & ~n4191 ) | ( n4185 & n4190 ) | ( ~n4191 & n4190 ) ;
  assign n4193 = ( n4185 & ~n4190 ) | ( n4185 & n4191 ) | ( ~n4190 & n4191 ) ;
  assign n4194 = ( n4192 & ~n4185 ) | ( n4192 & n4193 ) | ( ~n4185 & n4193 ) ;
  assign n4196 = ( n4155 & n4157 ) | ( n4155 & n4194 ) | ( n4157 & n4194 ) ;
  assign n4195 = ( n4155 & ~n4157 ) | ( n4155 & n4194 ) | ( ~n4157 & n4194 ) ;
  assign n4197 = ( n4157 & ~n4196 ) | ( n4157 & n4195 ) | ( ~n4196 & n4195 ) ;
  assign n4170 = ( n4136 & ~n4137 ) | ( n4136 & n4159 ) | ( ~n4137 & n4159 ) ;
  assign n4171 = n1737 | n1815 ;
  assign n4172 = ( n301 & ~n691 ) | ( n301 & n4171 ) | ( ~n691 & n4171 ) ;
  assign n4173 = n691 | n4172 ;
  assign n4174 = ( n1190 & ~n4173 ) | ( n1190 & n1875 ) | ( ~n4173 & n1875 ) ;
  assign n4175 = ~n1190 & n4174 ;
  assign n4176 = ( n329 & ~n2675 ) | ( n329 & n4175 ) | ( ~n2675 & n4175 ) ;
  assign n4177 = ~n329 & n4176 ;
  assign n4178 = ( n392 & ~n478 ) | ( n392 & n4177 ) | ( ~n478 & n4177 ) ;
  assign n4179 = ~n392 & n4178 ;
  assign n4180 = ( n103 & ~n610 ) | ( n103 & n4179 ) | ( ~n610 & n4179 ) ;
  assign n4181 = ~n103 & n4180 ;
  assign n4182 = ( n827 & ~n318 ) | ( n827 & n4181 ) | ( ~n318 & n4181 ) ;
  assign n4183 = ~n827 & n4182 ;
  assign n4184 = ~n363 & n4183 ;
  assign n4198 = ( n4170 & n4184 ) | ( n4170 & n4197 ) | ( n4184 & n4197 ) ;
  assign n4199 = ( n4170 & ~n4197 ) | ( n4170 & n4184 ) | ( ~n4197 & n4184 ) ;
  assign n4200 = ( n4197 & ~n4198 ) | ( n4197 & n4199 ) | ( ~n4198 & n4199 ) ;
  assign n4202 = ( n4166 & n4169 ) | ( n4166 & n4200 ) | ( n4169 & n4200 ) ;
  assign n4201 = ( n4169 & ~n4166 ) | ( n4169 & n4200 ) | ( ~n4166 & n4200 ) ;
  assign n4203 = ( n4166 & ~n4202 ) | ( n4166 & n4201 ) | ( ~n4202 & n4201 ) ;
  assign n4204 = ( n4166 & ~n4200 ) | ( n4166 & 1'b0 ) | ( ~n4200 & 1'b0 ) ;
  assign n4205 = ~n4166 & n4200 ;
  assign n4206 = ( n4168 & n4204 ) | ( n4168 & n4205 ) | ( n4204 & n4205 ) ;
  assign n4207 = n3195 | n4206 ;
  assign n4223 = ( n1967 & ~n3233 ) | ( n1967 & 1'b0 ) | ( ~n3233 & 1'b0 ) ;
  assign n4224 = n1958 | n3336 ;
  assign n4225 = ~n4223 & n4224 ;
  assign n4226 = ( n540 & ~n3121 ) | ( n540 & 1'b0 ) | ( ~n3121 & 1'b0 ) ;
  assign n4227 = ( n540 & n4225 ) | ( n540 & n4226 ) | ( n4225 & n4226 ) ;
  assign n4228 = ( n540 & ~n4225 ) | ( n540 & n4226 ) | ( ~n4225 & n4226 ) ;
  assign n4229 = ( n4225 & ~n4227 ) | ( n4225 & n4228 ) | ( ~n4227 & n4228 ) ;
  assign n4233 = ( n4157 & ~n4155 ) | ( n4157 & n4194 ) | ( ~n4155 & n4194 ) ;
  assign n4231 = n540 &  n4190 ;
  assign n4230 = ( n4190 & ~n4185 ) | ( n4190 & n4191 ) | ( ~n4185 & n4191 ) ;
  assign n4232 = ( n4185 & ~n4231 ) | ( n4185 & n4230 ) | ( ~n4231 & n4230 ) ;
  assign n4234 = ( n4229 & ~n4233 ) | ( n4229 & n4232 ) | ( ~n4233 & n4232 ) ;
  assign n4235 = ( n4229 & ~n4232 ) | ( n4229 & n4233 ) | ( ~n4232 & n4233 ) ;
  assign n4236 = ( n4234 & ~n4229 ) | ( n4234 & n4235 ) | ( ~n4229 & n4235 ) ;
  assign n4208 = ~n310 & n952 ;
  assign n4209 = ( n226 & ~n315 ) | ( n226 & n4208 ) | ( ~n315 & n4208 ) ;
  assign n4210 = ~n226 & n4209 ;
  assign n4211 = ( n611 & ~n283 ) | ( n611 & n4210 ) | ( ~n283 & n4210 ) ;
  assign n4212 = ~n611 & n4211 ;
  assign n4213 = ( n1744 & ~n4073 ) | ( n1744 & n4212 ) | ( ~n4073 & n4212 ) ;
  assign n4214 = ~n1744 & n4213 ;
  assign n4215 = ( n103 & n918 ) | ( n103 & n4214 ) | ( n918 & n4214 ) ;
  assign n4216 = ~n103 & n4215 ;
  assign n4217 = ( n191 & ~n311 ) | ( n191 & n4216 ) | ( ~n311 & n4216 ) ;
  assign n4218 = ~n191 & n4217 ;
  assign n4219 = ( n266 & ~n363 ) | ( n266 & n4218 ) | ( ~n363 & n4218 ) ;
  assign n4220 = ~n266 & n4219 ;
  assign n4221 = ~n355 & n4220 ;
  assign n4222 = ( n4170 & ~n4184 ) | ( n4170 & n4197 ) | ( ~n4184 & n4197 ) ;
  assign n4237 = ( n4221 & n4222 ) | ( n4221 & n4236 ) | ( n4222 & n4236 ) ;
  assign n4238 = ( n4221 & ~n4236 ) | ( n4221 & n4222 ) | ( ~n4236 & n4222 ) ;
  assign n4239 = ( n4236 & ~n4237 ) | ( n4236 & n4238 ) | ( ~n4237 & n4238 ) ;
  assign n4241 = ( n4204 & n4207 ) | ( n4204 & n4239 ) | ( n4207 & n4239 ) ;
  assign n4240 = ( n4207 & ~n4204 ) | ( n4207 & n4239 ) | ( ~n4204 & n4239 ) ;
  assign n4242 = ( n4204 & ~n4241 ) | ( n4204 & n4240 ) | ( ~n4241 & n4240 ) ;
  assign n4243 = n4204 &  n4239 ;
  assign n4244 = n4204 | n4239 ;
  assign n4245 = ( n4206 & ~n4244 ) | ( n4206 & n4243 ) | ( ~n4244 & n4243 ) ;
  assign n4246 = n3195 | n4245 ;
  assign n4247 = ( n4221 & ~n4222 ) | ( n4221 & n4236 ) | ( ~n4222 & n4236 ) ;
  assign n4248 = ~n479 & n1676 ;
  assign n4249 = ( n2140 & ~n4123 ) | ( n2140 & n4248 ) | ( ~n4123 & n4248 ) ;
  assign n4250 = ~n2140 & n4249 ;
  assign n4251 = ( n207 & ~n359 ) | ( n207 & n4250 ) | ( ~n359 & n4250 ) ;
  assign n4252 = ~n207 & n4251 ;
  assign n4253 = ( n182 & ~n3052 ) | ( n182 & n4252 ) | ( ~n3052 & n4252 ) ;
  assign n4254 = ~n182 & n4253 ;
  assign n4255 = ~n292 & n4254 ;
  assign n4256 = ~n643 & n4255 ;
  assign n4257 = ( n2941 & ~n3213 ) | ( n2941 & n3230 ) | ( ~n3213 & n3230 ) ;
  assign n4258 = ( n2941 & ~n3230 ) | ( n2941 & n3213 ) | ( ~n3230 & n3213 ) ;
  assign n4259 = ( n4257 & ~n2941 ) | ( n4257 & n4258 ) | ( ~n2941 & n4258 ) ;
  assign n4260 = n540 &  n4259 ;
  assign n4262 = ~n540 & n4225 ;
  assign n4261 = ( n2941 & ~n4225 ) | ( n2941 & n3113 ) | ( ~n4225 & n3113 ) ;
  assign n4263 = n540 &  n4261 ;
  assign n4264 = n4262 | n4263 ;
  assign n4265 = ( n4234 & ~n4260 ) | ( n4234 & n4264 ) | ( ~n4260 & n4264 ) ;
  assign n4266 = ( n4234 & ~n4264 ) | ( n4234 & n4260 ) | ( ~n4264 & n4260 ) ;
  assign n4267 = ( n4265 & ~n4234 ) | ( n4265 & n4266 ) | ( ~n4234 & n4266 ) ;
  assign n4268 = ( n4247 & ~n4256 ) | ( n4247 & n4267 ) | ( ~n4256 & n4267 ) ;
  assign n4269 = ( n4256 & ~n4247 ) | ( n4256 & n4267 ) | ( ~n4247 & n4267 ) ;
  assign n4270 = ( n4268 & ~n4267 ) | ( n4268 & n4269 ) | ( ~n4267 & n4269 ) ;
  assign n4272 = ( n4243 & n4246 ) | ( n4243 & n4270 ) | ( n4246 & n4270 ) ;
  assign n4271 = ( n4246 & ~n4243 ) | ( n4246 & n4270 ) | ( ~n4243 & n4270 ) ;
  assign n4273 = ( n4243 & ~n4272 ) | ( n4243 & n4271 ) | ( ~n4272 & n4271 ) ;
  assign n4274 = n4243 &  n4270 ;
  assign n4275 = n4243 | n4270 ;
  assign n4276 = ( n4245 & ~n4275 ) | ( n4245 & n4274 ) | ( ~n4275 & n4274 ) ;
  assign n4277 = n3195 | n4276 ;
  assign n4278 = ( n4247 & ~n4267 ) | ( n4247 & n4256 ) | ( ~n4267 & n4256 ) ;
  assign n4279 = ( n231 & n421 ) | ( n231 & n438 ) | ( n421 & n438 ) ;
  assign n4280 = ( n132 & ~n4279 ) | ( n132 & n421 ) | ( ~n4279 & n421 ) ;
  assign n4281 = ~n132 & n4280 ;
  assign n4282 = ( n570 & n2657 ) | ( n570 & n4281 ) | ( n2657 & n4281 ) ;
  assign n4283 = ~n570 & n4282 ;
  assign n4284 = ( n113 & ~n326 ) | ( n113 & n4283 ) | ( ~n326 & n4283 ) ;
  assign n4285 = ~n113 & n4284 ;
  assign n4286 = ( n181 & ~n353 ) | ( n181 & n4285 ) | ( ~n353 & n4285 ) ;
  assign n4287 = ~n181 & n4286 ;
  assign n4288 = ( n189 & ~n278 ) | ( n189 & n4287 ) | ( ~n278 & n4287 ) ;
  assign n4289 = ~n189 & n4288 ;
  assign n4290 = n4278 | n4289 ;
  assign n4291 = n4278 &  n4289 ;
  assign n4292 = ( n4290 & ~n4291 ) | ( n4290 & 1'b0 ) | ( ~n4291 & 1'b0 ) ;
  assign n4293 = ( n4274 & ~n4277 ) | ( n4274 & n4292 ) | ( ~n4277 & n4292 ) ;
  assign n4294 = ( n4274 & ~n4292 ) | ( n4274 & n4277 ) | ( ~n4292 & n4277 ) ;
  assign n4295 = ( n4293 & ~n4274 ) | ( n4293 & n4294 ) | ( ~n4274 & n4294 ) ;
  assign n4296 = n4274 &  n4292 ;
  assign n4297 = ( n609 & n965 ) | ( n609 & n2409 ) | ( n965 & n2409 ) ;
  assign n4298 = ( n583 & ~n4297 ) | ( n583 & n965 ) | ( ~n4297 & n965 ) ;
  assign n4299 = ~n583 & n4298 ;
  assign n4300 = ( n334 & ~n922 ) | ( n334 & n4299 ) | ( ~n922 & n4299 ) ;
  assign n4301 = ~n334 & n4300 ;
  assign n4302 = ( n478 & ~n3032 ) | ( n478 & n4301 ) | ( ~n3032 & n4301 ) ;
  assign n4303 = ~n478 & n4302 ;
  assign n4304 = ( n181 & ~n200 ) | ( n181 & n4303 ) | ( ~n200 & n4303 ) ;
  assign n4305 = ~n181 & n4304 ;
  assign n4306 = ( n212 & ~n289 ) | ( n212 & n4305 ) | ( ~n289 & n4305 ) ;
  assign n4307 = ~n212 & n4306 ;
  assign n4309 = n4290 &  n4307 ;
  assign n4308 = n4290 | n4307 ;
  assign n4310 = ( n4296 & ~n4309 ) | ( n4296 & n4308 ) | ( ~n4309 & n4308 ) ;
  assign n4311 = ( n4296 & ~n4309 ) | ( n4296 & 1'b0 ) | ( ~n4309 & 1'b0 ) ;
  assign n4312 = ( n4310 & ~n4311 ) | ( n4310 & 1'b0 ) | ( ~n4311 & 1'b0 ) ;
  assign n4313 = n4274 | n4292 ;
  assign n4314 = ( n4276 & ~n4313 ) | ( n4276 & n4296 ) | ( ~n4313 & n4296 ) ;
  assign n4315 = n3195 | n4314 ;
  assign n4316 = n4312 | n4315 ;
  assign n4317 = n4312 &  n4315 ;
  assign n4318 = ( n4316 & ~n4317 ) | ( n4316 & 1'b0 ) | ( ~n4317 & 1'b0 ) ;
  assign n4319 = ~n4312 & n4314 ;
  assign n4320 = n3195 | n4319 ;
  assign n4321 = ~n3586 & n4210 ;
  assign n4322 = ( n600 & ~n2440 ) | ( n600 & n4321 ) | ( ~n2440 & n4321 ) ;
  assign n4323 = ~n600 & n4322 ;
  assign n4324 = ( n118 & ~n486 ) | ( n118 & n4323 ) | ( ~n486 & n4323 ) ;
  assign n4325 = ~n118 & n4324 ;
  assign n4326 = ( n126 & ~n182 ) | ( n126 & n4325 ) | ( ~n182 & n4325 ) ;
  assign n4327 = ~n126 & n4326 ;
  assign n4328 = ( n114 & ~n277 ) | ( n114 & n4327 ) | ( ~n277 & n4327 ) ;
  assign n4329 = ~n114 & n4328 ;
  assign n4330 = ( n180 & ~n398 ) | ( n180 & n4329 ) | ( ~n398 & n4329 ) ;
  assign n4331 = ~n180 & n4330 ;
  assign n4332 = n4308 &  n4331 ;
  assign n4333 = n4308 | n4331 ;
  assign n4334 = ~n4332 & n4333 ;
  assign n4335 = ( n4311 & ~n4320 ) | ( n4311 & n4334 ) | ( ~n4320 & n4334 ) ;
  assign n4336 = ( n4311 & ~n4334 ) | ( n4311 & n4320 ) | ( ~n4334 & n4320 ) ;
  assign n4337 = ( n4335 & ~n4311 ) | ( n4335 & n4336 ) | ( ~n4311 & n4336 ) ;
  assign n4338 = n4311 &  n4334 ;
  assign n4339 = n163 | n673 ;
  assign n4340 = ( n345 & ~n729 ) | ( n345 & n4339 ) | ( ~n729 & n4339 ) ;
  assign n4341 = n729 | n4340 ;
  assign n4342 = ( n1666 & ~n4341 ) | ( n1666 & n3828 ) | ( ~n4341 & n3828 ) ;
  assign n4343 = ~n1666 & n4342 ;
  assign n4344 = ( n167 & ~n200 ) | ( n167 & n4343 ) | ( ~n200 & n4343 ) ;
  assign n4345 = ~n167 & n4344 ;
  assign n4346 = ( n192 & ~n443 ) | ( n192 & n4345 ) | ( ~n443 & n4345 ) ;
  assign n4347 = ~n192 & n4346 ;
  assign n4348 = ( n186 & n645 ) | ( n186 & n4347 ) | ( n645 & n4347 ) ;
  assign n4349 = ~n186 & n4348 ;
  assign n4350 = ~n555 & n4349 ;
  assign n4352 = n4333 &  n4350 ;
  assign n4351 = n4333 | n4350 ;
  assign n4353 = ( n4338 & ~n4352 ) | ( n4338 & n4351 ) | ( ~n4352 & n4351 ) ;
  assign n4354 = ( n4338 & ~n4352 ) | ( n4338 & 1'b0 ) | ( ~n4352 & 1'b0 ) ;
  assign n4355 = ( n4353 & ~n4354 ) | ( n4353 & 1'b0 ) | ( ~n4354 & 1'b0 ) ;
  assign n4356 = ~n4308 & n4331 ;
  assign n4357 = ( n4309 & ~n4308 ) | ( n4309 & n4331 ) | ( ~n4308 & n4331 ) ;
  assign n4358 = ( n4296 & ~n4357 ) | ( n4296 & n4308 ) | ( ~n4357 & n4308 ) ;
  assign n4359 = ( n4356 & ~n4311 ) | ( n4356 & n4358 ) | ( ~n4311 & n4358 ) ;
  assign n4360 = ( n4314 & ~n4311 ) | ( n4314 & n4334 ) | ( ~n4311 & n4334 ) ;
  assign n4361 = ~n4359 & n4360 ;
  assign n4362 = n3195 | n4361 ;
  assign n4363 = n4355 | n4362 ;
  assign n4364 = n4355 &  n4362 ;
  assign n4365 = ( n4363 & ~n4364 ) | ( n4363 & 1'b0 ) | ( ~n4364 & 1'b0 ) ;
  assign n4366 = ~n4355 & n4361 ;
  assign n4367 = n3195 | n4366 ;
  assign n4368 = n703 | n2930 ;
  assign n4369 = ( n293 & n788 ) | ( n293 & n4368 ) | ( n788 & n4368 ) ;
  assign n4370 = ( n610 & ~n4369 ) | ( n610 & n788 ) | ( ~n4369 & n788 ) ;
  assign n4371 = ~n610 & n4370 ;
  assign n4372 = n4351 &  n4371 ;
  assign n4373 = n4351 | n4371 ;
  assign n4374 = ~n4372 & n4373 ;
  assign n4375 = ( n4354 & ~n4367 ) | ( n4354 & n4374 ) | ( ~n4367 & n4374 ) ;
  assign n4376 = ( n4354 & ~n4374 ) | ( n4354 & n4367 ) | ( ~n4374 & n4367 ) ;
  assign n4377 = ( n4375 & ~n4354 ) | ( n4375 & n4376 ) | ( ~n4354 & n4376 ) ;
  assign n4378 = ~n739 & n788 ;
  assign n4389 = n4373 &  n4378 ;
  assign n4380 = ~n4351 & n4371 ;
  assign n4381 = ( n4352 & ~n4351 ) | ( n4352 & n4371 ) | ( ~n4351 & n4371 ) ;
  assign n4382 = ( n4338 & ~n4381 ) | ( n4338 & n4351 ) | ( ~n4381 & n4351 ) ;
  assign n4383 = ( n4380 & ~n4354 ) | ( n4380 & n4382 ) | ( ~n4354 & n4382 ) ;
  assign n4384 = ( n4361 & ~n4354 ) | ( n4361 & n4374 ) | ( ~n4354 & n4374 ) ;
  assign n4385 = ~n4383 & n4384 ;
  assign n4386 = n3195 | n4385 ;
  assign n4379 = n4354 &  n4374 ;
  assign n4387 = ~n4373 & n4378 ;
  assign n4388 = ( n4373 & ~n4379 ) | ( n4373 & n4387 ) | ( ~n4379 & n4387 ) ;
  assign n4391 = ( n4386 & n4388 ) | ( n4386 & n4389 ) | ( n4388 & n4389 ) ;
  assign n4390 = ( n4386 & ~n4389 ) | ( n4386 & n4388 ) | ( ~n4389 & n4388 ) ;
  assign n4392 = ( n4389 & ~n4391 ) | ( n4389 & n4390 ) | ( ~n4391 & n4390 ) ;
  assign n4393 = ( n4373 & ~n4379 ) | ( n4373 & n4378 ) | ( ~n4379 & n4378 ) ;
  assign n4397 = ( n4351 & ~n4354 ) | ( n4351 & n4371 ) | ( ~n4354 & n4371 ) ;
  assign n4398 = n4378 &  n4397 ;
  assign n4399 = ( n4385 & ~n4393 ) | ( n4385 & n4398 ) | ( ~n4393 & n4398 ) ;
  assign n4400 = n3195 | n4399 ;
  assign n4394 = ( x21 & ~x20 ) | ( x21 & n43 ) | ( ~x20 & n43 ) ;
  assign n4395 = x20 | n4394 ;
  assign n4396 = x22 | n4395 ;
  assign n4401 = ( n4393 & ~n4400 ) | ( n4393 & n4396 ) | ( ~n4400 & n4396 ) ;
  assign n4402 = ( n4396 & ~n4393 ) | ( n4396 & n4400 ) | ( ~n4393 & n4400 ) ;
  assign n4403 = n4401 &  n4402 ;
  assign n4404 = n4393 &  n4399 ;
  assign n4405 = ~n4396 & n4404 ;
  assign n4406 = ( n3195 & ~n4405 ) | ( n3195 & n4404 ) | ( ~n4405 & n4404 ) ;
  assign y0 = n3192 ;
  assign y1 = ~n3309 ;
  assign y2 = ~n3406 ;
  assign y3 = ~n3501 ;
  assign y4 = ~n3579 ;
  assign y5 = n3662 ;
  assign y6 = ~n3746 ;
  assign y7 = n3815 ;
  assign y8 = n3891 ;
  assign y9 = ~n3956 ;
  assign y10 = n4016 ;
  assign y11 = ~n4064 ;
  assign y12 = n4115 ;
  assign y13 = n4165 ;
  assign y14 = n4203 ;
  assign y15 = ~n4242 ;
  assign y16 = ~n4273 ;
  assign y17 = ~n4295 ;
  assign y18 = ~n4318 ;
  assign y19 = ~n4337 ;
  assign y20 = ~n4365 ;
  assign y21 = ~n4377 ;
  assign y22 = ~n4392 ;
  assign y23 = ~n4403 ;
  assign y24 = ~n4406 ;
endmodule
