module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 ;
  assign n257 = ( x0 & ~x128 ) | ( x0 & 1'b0 ) | ( ~x128 & 1'b0 ) ;
  assign n258 = ~x0 & x128 ;
  assign n259 = n257 | n258 ;
  assign n260 = x0 &  x128 ;
  assign n261 = ( x129 & ~x1 ) | ( x129 & n260 ) | ( ~x1 & n260 ) ;
  assign n262 = ( x1 & ~n260 ) | ( x1 & x129 ) | ( ~n260 & x129 ) ;
  assign n263 = ( n261 & ~x129 ) | ( n261 & n262 ) | ( ~x129 & n262 ) ;
  assign n264 = ( x1 & x129 ) | ( x1 & n260 ) | ( x129 & n260 ) ;
  assign n266 = ( x2 & x130 ) | ( x2 & n264 ) | ( x130 & n264 ) ;
  assign n265 = ( x2 & ~x130 ) | ( x2 & n264 ) | ( ~x130 & n264 ) ;
  assign n267 = ( x130 & ~n266 ) | ( x130 & n265 ) | ( ~n266 & n265 ) ;
  assign n269 = ( x3 & x131 ) | ( x3 & n266 ) | ( x131 & n266 ) ;
  assign n268 = ( x3 & ~x131 ) | ( x3 & n266 ) | ( ~x131 & n266 ) ;
  assign n270 = ( x131 & ~n269 ) | ( x131 & n268 ) | ( ~n269 & n268 ) ;
  assign n272 = ( x4 & x132 ) | ( x4 & n269 ) | ( x132 & n269 ) ;
  assign n271 = ( x4 & ~x132 ) | ( x4 & n269 ) | ( ~x132 & n269 ) ;
  assign n273 = ( x132 & ~n272 ) | ( x132 & n271 ) | ( ~n272 & n271 ) ;
  assign n275 = ( x5 & x133 ) | ( x5 & n272 ) | ( x133 & n272 ) ;
  assign n274 = ( x5 & ~x133 ) | ( x5 & n272 ) | ( ~x133 & n272 ) ;
  assign n276 = ( x133 & ~n275 ) | ( x133 & n274 ) | ( ~n275 & n274 ) ;
  assign n278 = ( x6 & x134 ) | ( x6 & n275 ) | ( x134 & n275 ) ;
  assign n277 = ( x6 & ~x134 ) | ( x6 & n275 ) | ( ~x134 & n275 ) ;
  assign n279 = ( x134 & ~n278 ) | ( x134 & n277 ) | ( ~n278 & n277 ) ;
  assign n281 = ( x7 & x135 ) | ( x7 & n278 ) | ( x135 & n278 ) ;
  assign n280 = ( x7 & ~x135 ) | ( x7 & n278 ) | ( ~x135 & n278 ) ;
  assign n282 = ( x135 & ~n281 ) | ( x135 & n280 ) | ( ~n281 & n280 ) ;
  assign n284 = ( x8 & x136 ) | ( x8 & n281 ) | ( x136 & n281 ) ;
  assign n283 = ( x8 & ~x136 ) | ( x8 & n281 ) | ( ~x136 & n281 ) ;
  assign n285 = ( x136 & ~n284 ) | ( x136 & n283 ) | ( ~n284 & n283 ) ;
  assign n287 = ( x9 & x137 ) | ( x9 & n284 ) | ( x137 & n284 ) ;
  assign n286 = ( x9 & ~x137 ) | ( x9 & n284 ) | ( ~x137 & n284 ) ;
  assign n288 = ( x137 & ~n287 ) | ( x137 & n286 ) | ( ~n287 & n286 ) ;
  assign n290 = ( x10 & x138 ) | ( x10 & n287 ) | ( x138 & n287 ) ;
  assign n289 = ( x10 & ~x138 ) | ( x10 & n287 ) | ( ~x138 & n287 ) ;
  assign n291 = ( x138 & ~n290 ) | ( x138 & n289 ) | ( ~n290 & n289 ) ;
  assign n293 = ( x11 & x139 ) | ( x11 & n290 ) | ( x139 & n290 ) ;
  assign n292 = ( x11 & ~x139 ) | ( x11 & n290 ) | ( ~x139 & n290 ) ;
  assign n294 = ( x139 & ~n293 ) | ( x139 & n292 ) | ( ~n293 & n292 ) ;
  assign n296 = ( x12 & x140 ) | ( x12 & n293 ) | ( x140 & n293 ) ;
  assign n295 = ( x12 & ~x140 ) | ( x12 & n293 ) | ( ~x140 & n293 ) ;
  assign n297 = ( x140 & ~n296 ) | ( x140 & n295 ) | ( ~n296 & n295 ) ;
  assign n299 = ( x13 & x141 ) | ( x13 & n296 ) | ( x141 & n296 ) ;
  assign n298 = ( x13 & ~x141 ) | ( x13 & n296 ) | ( ~x141 & n296 ) ;
  assign n300 = ( x141 & ~n299 ) | ( x141 & n298 ) | ( ~n299 & n298 ) ;
  assign n302 = ( x14 & x142 ) | ( x14 & n299 ) | ( x142 & n299 ) ;
  assign n301 = ( x14 & ~x142 ) | ( x14 & n299 ) | ( ~x142 & n299 ) ;
  assign n303 = ( x142 & ~n302 ) | ( x142 & n301 ) | ( ~n302 & n301 ) ;
  assign n305 = ( x15 & x143 ) | ( x15 & n302 ) | ( x143 & n302 ) ;
  assign n304 = ( x15 & ~x143 ) | ( x15 & n302 ) | ( ~x143 & n302 ) ;
  assign n306 = ( x143 & ~n305 ) | ( x143 & n304 ) | ( ~n305 & n304 ) ;
  assign n308 = ( x16 & x144 ) | ( x16 & n305 ) | ( x144 & n305 ) ;
  assign n307 = ( x16 & ~x144 ) | ( x16 & n305 ) | ( ~x144 & n305 ) ;
  assign n309 = ( x144 & ~n308 ) | ( x144 & n307 ) | ( ~n308 & n307 ) ;
  assign n311 = ( x17 & x145 ) | ( x17 & n308 ) | ( x145 & n308 ) ;
  assign n310 = ( x17 & ~x145 ) | ( x17 & n308 ) | ( ~x145 & n308 ) ;
  assign n312 = ( x145 & ~n311 ) | ( x145 & n310 ) | ( ~n311 & n310 ) ;
  assign n314 = ( x18 & x146 ) | ( x18 & n311 ) | ( x146 & n311 ) ;
  assign n313 = ( x18 & ~x146 ) | ( x18 & n311 ) | ( ~x146 & n311 ) ;
  assign n315 = ( x146 & ~n314 ) | ( x146 & n313 ) | ( ~n314 & n313 ) ;
  assign n317 = ( x19 & x147 ) | ( x19 & n314 ) | ( x147 & n314 ) ;
  assign n316 = ( x19 & ~x147 ) | ( x19 & n314 ) | ( ~x147 & n314 ) ;
  assign n318 = ( x147 & ~n317 ) | ( x147 & n316 ) | ( ~n317 & n316 ) ;
  assign n320 = ( x20 & x148 ) | ( x20 & n317 ) | ( x148 & n317 ) ;
  assign n319 = ( x20 & ~x148 ) | ( x20 & n317 ) | ( ~x148 & n317 ) ;
  assign n321 = ( x148 & ~n320 ) | ( x148 & n319 ) | ( ~n320 & n319 ) ;
  assign n323 = ( x21 & x149 ) | ( x21 & n320 ) | ( x149 & n320 ) ;
  assign n322 = ( x21 & ~x149 ) | ( x21 & n320 ) | ( ~x149 & n320 ) ;
  assign n324 = ( x149 & ~n323 ) | ( x149 & n322 ) | ( ~n323 & n322 ) ;
  assign n326 = ( x22 & x150 ) | ( x22 & n323 ) | ( x150 & n323 ) ;
  assign n325 = ( x22 & ~x150 ) | ( x22 & n323 ) | ( ~x150 & n323 ) ;
  assign n327 = ( x150 & ~n326 ) | ( x150 & n325 ) | ( ~n326 & n325 ) ;
  assign n329 = ( x23 & x151 ) | ( x23 & n326 ) | ( x151 & n326 ) ;
  assign n328 = ( x23 & ~x151 ) | ( x23 & n326 ) | ( ~x151 & n326 ) ;
  assign n330 = ( x151 & ~n329 ) | ( x151 & n328 ) | ( ~n329 & n328 ) ;
  assign n332 = ( x24 & x152 ) | ( x24 & n329 ) | ( x152 & n329 ) ;
  assign n331 = ( x24 & ~x152 ) | ( x24 & n329 ) | ( ~x152 & n329 ) ;
  assign n333 = ( x152 & ~n332 ) | ( x152 & n331 ) | ( ~n332 & n331 ) ;
  assign n335 = ( x25 & x153 ) | ( x25 & n332 ) | ( x153 & n332 ) ;
  assign n334 = ( x25 & ~x153 ) | ( x25 & n332 ) | ( ~x153 & n332 ) ;
  assign n336 = ( x153 & ~n335 ) | ( x153 & n334 ) | ( ~n335 & n334 ) ;
  assign n338 = ( x26 & x154 ) | ( x26 & n335 ) | ( x154 & n335 ) ;
  assign n337 = ( x26 & ~x154 ) | ( x26 & n335 ) | ( ~x154 & n335 ) ;
  assign n339 = ( x154 & ~n338 ) | ( x154 & n337 ) | ( ~n338 & n337 ) ;
  assign n341 = ( x27 & x155 ) | ( x27 & n338 ) | ( x155 & n338 ) ;
  assign n340 = ( x27 & ~x155 ) | ( x27 & n338 ) | ( ~x155 & n338 ) ;
  assign n342 = ( x155 & ~n341 ) | ( x155 & n340 ) | ( ~n341 & n340 ) ;
  assign n344 = ( x28 & x156 ) | ( x28 & n341 ) | ( x156 & n341 ) ;
  assign n343 = ( x28 & ~x156 ) | ( x28 & n341 ) | ( ~x156 & n341 ) ;
  assign n345 = ( x156 & ~n344 ) | ( x156 & n343 ) | ( ~n344 & n343 ) ;
  assign n347 = ( x29 & x157 ) | ( x29 & n344 ) | ( x157 & n344 ) ;
  assign n346 = ( x29 & ~x157 ) | ( x29 & n344 ) | ( ~x157 & n344 ) ;
  assign n348 = ( x157 & ~n347 ) | ( x157 & n346 ) | ( ~n347 & n346 ) ;
  assign n350 = ( x30 & x158 ) | ( x30 & n347 ) | ( x158 & n347 ) ;
  assign n349 = ( x30 & ~x158 ) | ( x30 & n347 ) | ( ~x158 & n347 ) ;
  assign n351 = ( x158 & ~n350 ) | ( x158 & n349 ) | ( ~n350 & n349 ) ;
  assign n353 = ( x31 & x159 ) | ( x31 & n350 ) | ( x159 & n350 ) ;
  assign n352 = ( x31 & ~x159 ) | ( x31 & n350 ) | ( ~x159 & n350 ) ;
  assign n354 = ( x159 & ~n353 ) | ( x159 & n352 ) | ( ~n353 & n352 ) ;
  assign n356 = ( x32 & x160 ) | ( x32 & n353 ) | ( x160 & n353 ) ;
  assign n355 = ( x32 & ~x160 ) | ( x32 & n353 ) | ( ~x160 & n353 ) ;
  assign n357 = ( x160 & ~n356 ) | ( x160 & n355 ) | ( ~n356 & n355 ) ;
  assign n359 = ( x33 & x161 ) | ( x33 & n356 ) | ( x161 & n356 ) ;
  assign n358 = ( x33 & ~x161 ) | ( x33 & n356 ) | ( ~x161 & n356 ) ;
  assign n360 = ( x161 & ~n359 ) | ( x161 & n358 ) | ( ~n359 & n358 ) ;
  assign n362 = ( x34 & x162 ) | ( x34 & n359 ) | ( x162 & n359 ) ;
  assign n361 = ( x34 & ~x162 ) | ( x34 & n359 ) | ( ~x162 & n359 ) ;
  assign n363 = ( x162 & ~n362 ) | ( x162 & n361 ) | ( ~n362 & n361 ) ;
  assign n365 = ( x35 & x163 ) | ( x35 & n362 ) | ( x163 & n362 ) ;
  assign n364 = ( x35 & ~x163 ) | ( x35 & n362 ) | ( ~x163 & n362 ) ;
  assign n366 = ( x163 & ~n365 ) | ( x163 & n364 ) | ( ~n365 & n364 ) ;
  assign n368 = ( x36 & x164 ) | ( x36 & n365 ) | ( x164 & n365 ) ;
  assign n367 = ( x36 & ~x164 ) | ( x36 & n365 ) | ( ~x164 & n365 ) ;
  assign n369 = ( x164 & ~n368 ) | ( x164 & n367 ) | ( ~n368 & n367 ) ;
  assign n371 = ( x37 & x165 ) | ( x37 & n368 ) | ( x165 & n368 ) ;
  assign n370 = ( x37 & ~x165 ) | ( x37 & n368 ) | ( ~x165 & n368 ) ;
  assign n372 = ( x165 & ~n371 ) | ( x165 & n370 ) | ( ~n371 & n370 ) ;
  assign n374 = ( x38 & x166 ) | ( x38 & n371 ) | ( x166 & n371 ) ;
  assign n373 = ( x38 & ~x166 ) | ( x38 & n371 ) | ( ~x166 & n371 ) ;
  assign n375 = ( x166 & ~n374 ) | ( x166 & n373 ) | ( ~n374 & n373 ) ;
  assign n377 = ( x39 & x167 ) | ( x39 & n374 ) | ( x167 & n374 ) ;
  assign n376 = ( x39 & ~x167 ) | ( x39 & n374 ) | ( ~x167 & n374 ) ;
  assign n378 = ( x167 & ~n377 ) | ( x167 & n376 ) | ( ~n377 & n376 ) ;
  assign n380 = ( x40 & x168 ) | ( x40 & n377 ) | ( x168 & n377 ) ;
  assign n379 = ( x40 & ~x168 ) | ( x40 & n377 ) | ( ~x168 & n377 ) ;
  assign n381 = ( x168 & ~n380 ) | ( x168 & n379 ) | ( ~n380 & n379 ) ;
  assign n383 = ( x41 & x169 ) | ( x41 & n380 ) | ( x169 & n380 ) ;
  assign n382 = ( x41 & ~x169 ) | ( x41 & n380 ) | ( ~x169 & n380 ) ;
  assign n384 = ( x169 & ~n383 ) | ( x169 & n382 ) | ( ~n383 & n382 ) ;
  assign n386 = ( x42 & x170 ) | ( x42 & n383 ) | ( x170 & n383 ) ;
  assign n385 = ( x42 & ~x170 ) | ( x42 & n383 ) | ( ~x170 & n383 ) ;
  assign n387 = ( x170 & ~n386 ) | ( x170 & n385 ) | ( ~n386 & n385 ) ;
  assign n389 = ( x43 & x171 ) | ( x43 & n386 ) | ( x171 & n386 ) ;
  assign n388 = ( x43 & ~x171 ) | ( x43 & n386 ) | ( ~x171 & n386 ) ;
  assign n390 = ( x171 & ~n389 ) | ( x171 & n388 ) | ( ~n389 & n388 ) ;
  assign n392 = ( x44 & x172 ) | ( x44 & n389 ) | ( x172 & n389 ) ;
  assign n391 = ( x44 & ~x172 ) | ( x44 & n389 ) | ( ~x172 & n389 ) ;
  assign n393 = ( x172 & ~n392 ) | ( x172 & n391 ) | ( ~n392 & n391 ) ;
  assign n395 = ( x45 & x173 ) | ( x45 & n392 ) | ( x173 & n392 ) ;
  assign n394 = ( x45 & ~x173 ) | ( x45 & n392 ) | ( ~x173 & n392 ) ;
  assign n396 = ( x173 & ~n395 ) | ( x173 & n394 ) | ( ~n395 & n394 ) ;
  assign n398 = ( x46 & x174 ) | ( x46 & n395 ) | ( x174 & n395 ) ;
  assign n397 = ( x46 & ~x174 ) | ( x46 & n395 ) | ( ~x174 & n395 ) ;
  assign n399 = ( x174 & ~n398 ) | ( x174 & n397 ) | ( ~n398 & n397 ) ;
  assign n401 = ( x47 & x175 ) | ( x47 & n398 ) | ( x175 & n398 ) ;
  assign n400 = ( x47 & ~x175 ) | ( x47 & n398 ) | ( ~x175 & n398 ) ;
  assign n402 = ( x175 & ~n401 ) | ( x175 & n400 ) | ( ~n401 & n400 ) ;
  assign n404 = ( x48 & x176 ) | ( x48 & n401 ) | ( x176 & n401 ) ;
  assign n403 = ( x48 & ~x176 ) | ( x48 & n401 ) | ( ~x176 & n401 ) ;
  assign n405 = ( x176 & ~n404 ) | ( x176 & n403 ) | ( ~n404 & n403 ) ;
  assign n407 = ( x49 & x177 ) | ( x49 & n404 ) | ( x177 & n404 ) ;
  assign n406 = ( x49 & ~x177 ) | ( x49 & n404 ) | ( ~x177 & n404 ) ;
  assign n408 = ( x177 & ~n407 ) | ( x177 & n406 ) | ( ~n407 & n406 ) ;
  assign n410 = ( x50 & x178 ) | ( x50 & n407 ) | ( x178 & n407 ) ;
  assign n409 = ( x50 & ~x178 ) | ( x50 & n407 ) | ( ~x178 & n407 ) ;
  assign n411 = ( x178 & ~n410 ) | ( x178 & n409 ) | ( ~n410 & n409 ) ;
  assign n413 = ( x51 & x179 ) | ( x51 & n410 ) | ( x179 & n410 ) ;
  assign n412 = ( x51 & ~x179 ) | ( x51 & n410 ) | ( ~x179 & n410 ) ;
  assign n414 = ( x179 & ~n413 ) | ( x179 & n412 ) | ( ~n413 & n412 ) ;
  assign n416 = ( x52 & x180 ) | ( x52 & n413 ) | ( x180 & n413 ) ;
  assign n415 = ( x52 & ~x180 ) | ( x52 & n413 ) | ( ~x180 & n413 ) ;
  assign n417 = ( x180 & ~n416 ) | ( x180 & n415 ) | ( ~n416 & n415 ) ;
  assign n419 = ( x53 & x181 ) | ( x53 & n416 ) | ( x181 & n416 ) ;
  assign n418 = ( x53 & ~x181 ) | ( x53 & n416 ) | ( ~x181 & n416 ) ;
  assign n420 = ( x181 & ~n419 ) | ( x181 & n418 ) | ( ~n419 & n418 ) ;
  assign n422 = ( x54 & x182 ) | ( x54 & n419 ) | ( x182 & n419 ) ;
  assign n421 = ( x54 & ~x182 ) | ( x54 & n419 ) | ( ~x182 & n419 ) ;
  assign n423 = ( x182 & ~n422 ) | ( x182 & n421 ) | ( ~n422 & n421 ) ;
  assign n425 = ( x55 & x183 ) | ( x55 & n422 ) | ( x183 & n422 ) ;
  assign n424 = ( x55 & ~x183 ) | ( x55 & n422 ) | ( ~x183 & n422 ) ;
  assign n426 = ( x183 & ~n425 ) | ( x183 & n424 ) | ( ~n425 & n424 ) ;
  assign n428 = ( x56 & x184 ) | ( x56 & n425 ) | ( x184 & n425 ) ;
  assign n427 = ( x56 & ~x184 ) | ( x56 & n425 ) | ( ~x184 & n425 ) ;
  assign n429 = ( x184 & ~n428 ) | ( x184 & n427 ) | ( ~n428 & n427 ) ;
  assign n431 = ( x57 & x185 ) | ( x57 & n428 ) | ( x185 & n428 ) ;
  assign n430 = ( x57 & ~x185 ) | ( x57 & n428 ) | ( ~x185 & n428 ) ;
  assign n432 = ( x185 & ~n431 ) | ( x185 & n430 ) | ( ~n431 & n430 ) ;
  assign n434 = ( x58 & x186 ) | ( x58 & n431 ) | ( x186 & n431 ) ;
  assign n433 = ( x58 & ~x186 ) | ( x58 & n431 ) | ( ~x186 & n431 ) ;
  assign n435 = ( x186 & ~n434 ) | ( x186 & n433 ) | ( ~n434 & n433 ) ;
  assign n437 = ( x59 & x187 ) | ( x59 & n434 ) | ( x187 & n434 ) ;
  assign n436 = ( x59 & ~x187 ) | ( x59 & n434 ) | ( ~x187 & n434 ) ;
  assign n438 = ( x187 & ~n437 ) | ( x187 & n436 ) | ( ~n437 & n436 ) ;
  assign n440 = ( x60 & x188 ) | ( x60 & n437 ) | ( x188 & n437 ) ;
  assign n439 = ( x60 & ~x188 ) | ( x60 & n437 ) | ( ~x188 & n437 ) ;
  assign n441 = ( x188 & ~n440 ) | ( x188 & n439 ) | ( ~n440 & n439 ) ;
  assign n443 = ( x61 & x189 ) | ( x61 & n440 ) | ( x189 & n440 ) ;
  assign n442 = ( x61 & ~x189 ) | ( x61 & n440 ) | ( ~x189 & n440 ) ;
  assign n444 = ( x189 & ~n443 ) | ( x189 & n442 ) | ( ~n443 & n442 ) ;
  assign n446 = ( x62 & x190 ) | ( x62 & n443 ) | ( x190 & n443 ) ;
  assign n445 = ( x62 & ~x190 ) | ( x62 & n443 ) | ( ~x190 & n443 ) ;
  assign n447 = ( x190 & ~n446 ) | ( x190 & n445 ) | ( ~n446 & n445 ) ;
  assign n449 = ( x63 & x191 ) | ( x63 & n446 ) | ( x191 & n446 ) ;
  assign n448 = ( x63 & ~x191 ) | ( x63 & n446 ) | ( ~x191 & n446 ) ;
  assign n450 = ( x191 & ~n449 ) | ( x191 & n448 ) | ( ~n449 & n448 ) ;
  assign n452 = ( x64 & x192 ) | ( x64 & n449 ) | ( x192 & n449 ) ;
  assign n451 = ( x64 & ~x192 ) | ( x64 & n449 ) | ( ~x192 & n449 ) ;
  assign n453 = ( x192 & ~n452 ) | ( x192 & n451 ) | ( ~n452 & n451 ) ;
  assign n455 = ( x65 & x193 ) | ( x65 & n452 ) | ( x193 & n452 ) ;
  assign n454 = ( x65 & ~x193 ) | ( x65 & n452 ) | ( ~x193 & n452 ) ;
  assign n456 = ( x193 & ~n455 ) | ( x193 & n454 ) | ( ~n455 & n454 ) ;
  assign n458 = ( x66 & x194 ) | ( x66 & n455 ) | ( x194 & n455 ) ;
  assign n457 = ( x66 & ~x194 ) | ( x66 & n455 ) | ( ~x194 & n455 ) ;
  assign n459 = ( x194 & ~n458 ) | ( x194 & n457 ) | ( ~n458 & n457 ) ;
  assign n461 = ( x67 & x195 ) | ( x67 & n458 ) | ( x195 & n458 ) ;
  assign n460 = ( x67 & ~x195 ) | ( x67 & n458 ) | ( ~x195 & n458 ) ;
  assign n462 = ( x195 & ~n461 ) | ( x195 & n460 ) | ( ~n461 & n460 ) ;
  assign n464 = ( x68 & x196 ) | ( x68 & n461 ) | ( x196 & n461 ) ;
  assign n463 = ( x68 & ~x196 ) | ( x68 & n461 ) | ( ~x196 & n461 ) ;
  assign n465 = ( x196 & ~n464 ) | ( x196 & n463 ) | ( ~n464 & n463 ) ;
  assign n467 = ( x69 & x197 ) | ( x69 & n464 ) | ( x197 & n464 ) ;
  assign n466 = ( x69 & ~x197 ) | ( x69 & n464 ) | ( ~x197 & n464 ) ;
  assign n468 = ( x197 & ~n467 ) | ( x197 & n466 ) | ( ~n467 & n466 ) ;
  assign n470 = ( x70 & x198 ) | ( x70 & n467 ) | ( x198 & n467 ) ;
  assign n469 = ( x70 & ~x198 ) | ( x70 & n467 ) | ( ~x198 & n467 ) ;
  assign n471 = ( x198 & ~n470 ) | ( x198 & n469 ) | ( ~n470 & n469 ) ;
  assign n473 = ( x71 & x199 ) | ( x71 & n470 ) | ( x199 & n470 ) ;
  assign n472 = ( x71 & ~x199 ) | ( x71 & n470 ) | ( ~x199 & n470 ) ;
  assign n474 = ( x199 & ~n473 ) | ( x199 & n472 ) | ( ~n473 & n472 ) ;
  assign n476 = ( x72 & x200 ) | ( x72 & n473 ) | ( x200 & n473 ) ;
  assign n475 = ( x72 & ~x200 ) | ( x72 & n473 ) | ( ~x200 & n473 ) ;
  assign n477 = ( x200 & ~n476 ) | ( x200 & n475 ) | ( ~n476 & n475 ) ;
  assign n479 = ( x73 & x201 ) | ( x73 & n476 ) | ( x201 & n476 ) ;
  assign n478 = ( x73 & ~x201 ) | ( x73 & n476 ) | ( ~x201 & n476 ) ;
  assign n480 = ( x201 & ~n479 ) | ( x201 & n478 ) | ( ~n479 & n478 ) ;
  assign n482 = ( x74 & x202 ) | ( x74 & n479 ) | ( x202 & n479 ) ;
  assign n481 = ( x74 & ~x202 ) | ( x74 & n479 ) | ( ~x202 & n479 ) ;
  assign n483 = ( x202 & ~n482 ) | ( x202 & n481 ) | ( ~n482 & n481 ) ;
  assign n485 = ( x75 & x203 ) | ( x75 & n482 ) | ( x203 & n482 ) ;
  assign n484 = ( x75 & ~x203 ) | ( x75 & n482 ) | ( ~x203 & n482 ) ;
  assign n486 = ( x203 & ~n485 ) | ( x203 & n484 ) | ( ~n485 & n484 ) ;
  assign n488 = ( x76 & x204 ) | ( x76 & n485 ) | ( x204 & n485 ) ;
  assign n487 = ( x76 & ~x204 ) | ( x76 & n485 ) | ( ~x204 & n485 ) ;
  assign n489 = ( x204 & ~n488 ) | ( x204 & n487 ) | ( ~n488 & n487 ) ;
  assign n491 = ( x77 & x205 ) | ( x77 & n488 ) | ( x205 & n488 ) ;
  assign n490 = ( x77 & ~x205 ) | ( x77 & n488 ) | ( ~x205 & n488 ) ;
  assign n492 = ( x205 & ~n491 ) | ( x205 & n490 ) | ( ~n491 & n490 ) ;
  assign n494 = ( x78 & x206 ) | ( x78 & n491 ) | ( x206 & n491 ) ;
  assign n493 = ( x78 & ~x206 ) | ( x78 & n491 ) | ( ~x206 & n491 ) ;
  assign n495 = ( x206 & ~n494 ) | ( x206 & n493 ) | ( ~n494 & n493 ) ;
  assign n497 = ( x79 & x207 ) | ( x79 & n494 ) | ( x207 & n494 ) ;
  assign n496 = ( x79 & ~x207 ) | ( x79 & n494 ) | ( ~x207 & n494 ) ;
  assign n498 = ( x207 & ~n497 ) | ( x207 & n496 ) | ( ~n497 & n496 ) ;
  assign n500 = ( x80 & x208 ) | ( x80 & n497 ) | ( x208 & n497 ) ;
  assign n499 = ( x80 & ~x208 ) | ( x80 & n497 ) | ( ~x208 & n497 ) ;
  assign n501 = ( x208 & ~n500 ) | ( x208 & n499 ) | ( ~n500 & n499 ) ;
  assign n503 = ( x81 & x209 ) | ( x81 & n500 ) | ( x209 & n500 ) ;
  assign n502 = ( x81 & ~x209 ) | ( x81 & n500 ) | ( ~x209 & n500 ) ;
  assign n504 = ( x209 & ~n503 ) | ( x209 & n502 ) | ( ~n503 & n502 ) ;
  assign n506 = ( x82 & x210 ) | ( x82 & n503 ) | ( x210 & n503 ) ;
  assign n505 = ( x82 & ~x210 ) | ( x82 & n503 ) | ( ~x210 & n503 ) ;
  assign n507 = ( x210 & ~n506 ) | ( x210 & n505 ) | ( ~n506 & n505 ) ;
  assign n509 = ( x83 & x211 ) | ( x83 & n506 ) | ( x211 & n506 ) ;
  assign n508 = ( x83 & ~x211 ) | ( x83 & n506 ) | ( ~x211 & n506 ) ;
  assign n510 = ( x211 & ~n509 ) | ( x211 & n508 ) | ( ~n509 & n508 ) ;
  assign n512 = ( x84 & x212 ) | ( x84 & n509 ) | ( x212 & n509 ) ;
  assign n511 = ( x84 & ~x212 ) | ( x84 & n509 ) | ( ~x212 & n509 ) ;
  assign n513 = ( x212 & ~n512 ) | ( x212 & n511 ) | ( ~n512 & n511 ) ;
  assign n515 = ( x85 & x213 ) | ( x85 & n512 ) | ( x213 & n512 ) ;
  assign n514 = ( x85 & ~x213 ) | ( x85 & n512 ) | ( ~x213 & n512 ) ;
  assign n516 = ( x213 & ~n515 ) | ( x213 & n514 ) | ( ~n515 & n514 ) ;
  assign n518 = ( x86 & x214 ) | ( x86 & n515 ) | ( x214 & n515 ) ;
  assign n517 = ( x86 & ~x214 ) | ( x86 & n515 ) | ( ~x214 & n515 ) ;
  assign n519 = ( x214 & ~n518 ) | ( x214 & n517 ) | ( ~n518 & n517 ) ;
  assign n521 = ( x87 & x215 ) | ( x87 & n518 ) | ( x215 & n518 ) ;
  assign n520 = ( x87 & ~x215 ) | ( x87 & n518 ) | ( ~x215 & n518 ) ;
  assign n522 = ( x215 & ~n521 ) | ( x215 & n520 ) | ( ~n521 & n520 ) ;
  assign n524 = ( x88 & x216 ) | ( x88 & n521 ) | ( x216 & n521 ) ;
  assign n523 = ( x88 & ~x216 ) | ( x88 & n521 ) | ( ~x216 & n521 ) ;
  assign n525 = ( x216 & ~n524 ) | ( x216 & n523 ) | ( ~n524 & n523 ) ;
  assign n527 = ( x89 & x217 ) | ( x89 & n524 ) | ( x217 & n524 ) ;
  assign n526 = ( x89 & ~x217 ) | ( x89 & n524 ) | ( ~x217 & n524 ) ;
  assign n528 = ( x217 & ~n527 ) | ( x217 & n526 ) | ( ~n527 & n526 ) ;
  assign n530 = ( x90 & x218 ) | ( x90 & n527 ) | ( x218 & n527 ) ;
  assign n529 = ( x90 & ~x218 ) | ( x90 & n527 ) | ( ~x218 & n527 ) ;
  assign n531 = ( x218 & ~n530 ) | ( x218 & n529 ) | ( ~n530 & n529 ) ;
  assign n533 = ( x91 & x219 ) | ( x91 & n530 ) | ( x219 & n530 ) ;
  assign n532 = ( x91 & ~x219 ) | ( x91 & n530 ) | ( ~x219 & n530 ) ;
  assign n534 = ( x219 & ~n533 ) | ( x219 & n532 ) | ( ~n533 & n532 ) ;
  assign n536 = ( x92 & x220 ) | ( x92 & n533 ) | ( x220 & n533 ) ;
  assign n535 = ( x92 & ~x220 ) | ( x92 & n533 ) | ( ~x220 & n533 ) ;
  assign n537 = ( x220 & ~n536 ) | ( x220 & n535 ) | ( ~n536 & n535 ) ;
  assign n539 = ( x93 & x221 ) | ( x93 & n536 ) | ( x221 & n536 ) ;
  assign n538 = ( x93 & ~x221 ) | ( x93 & n536 ) | ( ~x221 & n536 ) ;
  assign n540 = ( x221 & ~n539 ) | ( x221 & n538 ) | ( ~n539 & n538 ) ;
  assign n542 = ( x94 & x222 ) | ( x94 & n539 ) | ( x222 & n539 ) ;
  assign n541 = ( x94 & ~x222 ) | ( x94 & n539 ) | ( ~x222 & n539 ) ;
  assign n543 = ( x222 & ~n542 ) | ( x222 & n541 ) | ( ~n542 & n541 ) ;
  assign n545 = ( x95 & x223 ) | ( x95 & n542 ) | ( x223 & n542 ) ;
  assign n544 = ( x95 & ~x223 ) | ( x95 & n542 ) | ( ~x223 & n542 ) ;
  assign n546 = ( x223 & ~n545 ) | ( x223 & n544 ) | ( ~n545 & n544 ) ;
  assign n548 = ( x96 & x224 ) | ( x96 & n545 ) | ( x224 & n545 ) ;
  assign n547 = ( x96 & ~x224 ) | ( x96 & n545 ) | ( ~x224 & n545 ) ;
  assign n549 = ( x224 & ~n548 ) | ( x224 & n547 ) | ( ~n548 & n547 ) ;
  assign n551 = ( x97 & x225 ) | ( x97 & n548 ) | ( x225 & n548 ) ;
  assign n550 = ( x97 & ~x225 ) | ( x97 & n548 ) | ( ~x225 & n548 ) ;
  assign n552 = ( x225 & ~n551 ) | ( x225 & n550 ) | ( ~n551 & n550 ) ;
  assign n554 = ( x98 & x226 ) | ( x98 & n551 ) | ( x226 & n551 ) ;
  assign n553 = ( x98 & ~x226 ) | ( x98 & n551 ) | ( ~x226 & n551 ) ;
  assign n555 = ( x226 & ~n554 ) | ( x226 & n553 ) | ( ~n554 & n553 ) ;
  assign n557 = ( x99 & x227 ) | ( x99 & n554 ) | ( x227 & n554 ) ;
  assign n556 = ( x99 & ~x227 ) | ( x99 & n554 ) | ( ~x227 & n554 ) ;
  assign n558 = ( x227 & ~n557 ) | ( x227 & n556 ) | ( ~n557 & n556 ) ;
  assign n560 = ( x100 & x228 ) | ( x100 & n557 ) | ( x228 & n557 ) ;
  assign n559 = ( x100 & ~x228 ) | ( x100 & n557 ) | ( ~x228 & n557 ) ;
  assign n561 = ( x228 & ~n560 ) | ( x228 & n559 ) | ( ~n560 & n559 ) ;
  assign n563 = ( x101 & x229 ) | ( x101 & n560 ) | ( x229 & n560 ) ;
  assign n562 = ( x101 & ~x229 ) | ( x101 & n560 ) | ( ~x229 & n560 ) ;
  assign n564 = ( x229 & ~n563 ) | ( x229 & n562 ) | ( ~n563 & n562 ) ;
  assign n566 = ( x102 & x230 ) | ( x102 & n563 ) | ( x230 & n563 ) ;
  assign n565 = ( x102 & ~x230 ) | ( x102 & n563 ) | ( ~x230 & n563 ) ;
  assign n567 = ( x230 & ~n566 ) | ( x230 & n565 ) | ( ~n566 & n565 ) ;
  assign n569 = ( x103 & x231 ) | ( x103 & n566 ) | ( x231 & n566 ) ;
  assign n568 = ( x103 & ~x231 ) | ( x103 & n566 ) | ( ~x231 & n566 ) ;
  assign n570 = ( x231 & ~n569 ) | ( x231 & n568 ) | ( ~n569 & n568 ) ;
  assign n572 = ( x104 & x232 ) | ( x104 & n569 ) | ( x232 & n569 ) ;
  assign n571 = ( x104 & ~x232 ) | ( x104 & n569 ) | ( ~x232 & n569 ) ;
  assign n573 = ( x232 & ~n572 ) | ( x232 & n571 ) | ( ~n572 & n571 ) ;
  assign n575 = ( x105 & x233 ) | ( x105 & n572 ) | ( x233 & n572 ) ;
  assign n574 = ( x105 & ~x233 ) | ( x105 & n572 ) | ( ~x233 & n572 ) ;
  assign n576 = ( x233 & ~n575 ) | ( x233 & n574 ) | ( ~n575 & n574 ) ;
  assign n578 = ( x106 & x234 ) | ( x106 & n575 ) | ( x234 & n575 ) ;
  assign n577 = ( x106 & ~x234 ) | ( x106 & n575 ) | ( ~x234 & n575 ) ;
  assign n579 = ( x234 & ~n578 ) | ( x234 & n577 ) | ( ~n578 & n577 ) ;
  assign n581 = ( x107 & x235 ) | ( x107 & n578 ) | ( x235 & n578 ) ;
  assign n580 = ( x107 & ~x235 ) | ( x107 & n578 ) | ( ~x235 & n578 ) ;
  assign n582 = ( x235 & ~n581 ) | ( x235 & n580 ) | ( ~n581 & n580 ) ;
  assign n584 = ( x108 & x236 ) | ( x108 & n581 ) | ( x236 & n581 ) ;
  assign n583 = ( x108 & ~x236 ) | ( x108 & n581 ) | ( ~x236 & n581 ) ;
  assign n585 = ( x236 & ~n584 ) | ( x236 & n583 ) | ( ~n584 & n583 ) ;
  assign n587 = ( x109 & x237 ) | ( x109 & n584 ) | ( x237 & n584 ) ;
  assign n586 = ( x109 & ~x237 ) | ( x109 & n584 ) | ( ~x237 & n584 ) ;
  assign n588 = ( x237 & ~n587 ) | ( x237 & n586 ) | ( ~n587 & n586 ) ;
  assign n590 = ( x110 & x238 ) | ( x110 & n587 ) | ( x238 & n587 ) ;
  assign n589 = ( x110 & ~x238 ) | ( x110 & n587 ) | ( ~x238 & n587 ) ;
  assign n591 = ( x238 & ~n590 ) | ( x238 & n589 ) | ( ~n590 & n589 ) ;
  assign n593 = ( x111 & x239 ) | ( x111 & n590 ) | ( x239 & n590 ) ;
  assign n592 = ( x111 & ~x239 ) | ( x111 & n590 ) | ( ~x239 & n590 ) ;
  assign n594 = ( x239 & ~n593 ) | ( x239 & n592 ) | ( ~n593 & n592 ) ;
  assign n596 = ( x112 & x240 ) | ( x112 & n593 ) | ( x240 & n593 ) ;
  assign n595 = ( x112 & ~x240 ) | ( x112 & n593 ) | ( ~x240 & n593 ) ;
  assign n597 = ( x240 & ~n596 ) | ( x240 & n595 ) | ( ~n596 & n595 ) ;
  assign n599 = ( x113 & x241 ) | ( x113 & n596 ) | ( x241 & n596 ) ;
  assign n598 = ( x113 & ~x241 ) | ( x113 & n596 ) | ( ~x241 & n596 ) ;
  assign n600 = ( x241 & ~n599 ) | ( x241 & n598 ) | ( ~n599 & n598 ) ;
  assign n602 = ( x114 & x242 ) | ( x114 & n599 ) | ( x242 & n599 ) ;
  assign n601 = ( x114 & ~x242 ) | ( x114 & n599 ) | ( ~x242 & n599 ) ;
  assign n603 = ( x242 & ~n602 ) | ( x242 & n601 ) | ( ~n602 & n601 ) ;
  assign n605 = ( x115 & x243 ) | ( x115 & n602 ) | ( x243 & n602 ) ;
  assign n604 = ( x115 & ~x243 ) | ( x115 & n602 ) | ( ~x243 & n602 ) ;
  assign n606 = ( x243 & ~n605 ) | ( x243 & n604 ) | ( ~n605 & n604 ) ;
  assign n608 = ( x116 & x244 ) | ( x116 & n605 ) | ( x244 & n605 ) ;
  assign n607 = ( x116 & ~x244 ) | ( x116 & n605 ) | ( ~x244 & n605 ) ;
  assign n609 = ( x244 & ~n608 ) | ( x244 & n607 ) | ( ~n608 & n607 ) ;
  assign n611 = ( x117 & x245 ) | ( x117 & n608 ) | ( x245 & n608 ) ;
  assign n610 = ( x117 & ~x245 ) | ( x117 & n608 ) | ( ~x245 & n608 ) ;
  assign n612 = ( x245 & ~n611 ) | ( x245 & n610 ) | ( ~n611 & n610 ) ;
  assign n614 = ( x118 & x246 ) | ( x118 & n611 ) | ( x246 & n611 ) ;
  assign n613 = ( x118 & ~x246 ) | ( x118 & n611 ) | ( ~x246 & n611 ) ;
  assign n615 = ( x246 & ~n614 ) | ( x246 & n613 ) | ( ~n614 & n613 ) ;
  assign n617 = ( x119 & x247 ) | ( x119 & n614 ) | ( x247 & n614 ) ;
  assign n616 = ( x119 & ~x247 ) | ( x119 & n614 ) | ( ~x247 & n614 ) ;
  assign n618 = ( x247 & ~n617 ) | ( x247 & n616 ) | ( ~n617 & n616 ) ;
  assign n620 = ( x120 & x248 ) | ( x120 & n617 ) | ( x248 & n617 ) ;
  assign n619 = ( x120 & ~x248 ) | ( x120 & n617 ) | ( ~x248 & n617 ) ;
  assign n621 = ( x248 & ~n620 ) | ( x248 & n619 ) | ( ~n620 & n619 ) ;
  assign n623 = ( x121 & x249 ) | ( x121 & n620 ) | ( x249 & n620 ) ;
  assign n622 = ( x121 & ~x249 ) | ( x121 & n620 ) | ( ~x249 & n620 ) ;
  assign n624 = ( x249 & ~n623 ) | ( x249 & n622 ) | ( ~n623 & n622 ) ;
  assign n626 = ( x122 & x250 ) | ( x122 & n623 ) | ( x250 & n623 ) ;
  assign n625 = ( x122 & ~x250 ) | ( x122 & n623 ) | ( ~x250 & n623 ) ;
  assign n627 = ( x250 & ~n626 ) | ( x250 & n625 ) | ( ~n626 & n625 ) ;
  assign n629 = ( x123 & x251 ) | ( x123 & n626 ) | ( x251 & n626 ) ;
  assign n628 = ( x123 & ~x251 ) | ( x123 & n626 ) | ( ~x251 & n626 ) ;
  assign n630 = ( x251 & ~n629 ) | ( x251 & n628 ) | ( ~n629 & n628 ) ;
  assign n632 = ( x124 & x252 ) | ( x124 & n629 ) | ( x252 & n629 ) ;
  assign n631 = ( x124 & ~x252 ) | ( x124 & n629 ) | ( ~x252 & n629 ) ;
  assign n633 = ( x252 & ~n632 ) | ( x252 & n631 ) | ( ~n632 & n631 ) ;
  assign n635 = ( x125 & x253 ) | ( x125 & n632 ) | ( x253 & n632 ) ;
  assign n634 = ( x125 & ~x253 ) | ( x125 & n632 ) | ( ~x253 & n632 ) ;
  assign n636 = ( x253 & ~n635 ) | ( x253 & n634 ) | ( ~n635 & n634 ) ;
  assign n638 = ( x126 & x254 ) | ( x126 & n635 ) | ( x254 & n635 ) ;
  assign n637 = ( x126 & ~x254 ) | ( x126 & n635 ) | ( ~x254 & n635 ) ;
  assign n639 = ( x254 & ~n638 ) | ( x254 & n637 ) | ( ~n638 & n637 ) ;
  assign n640 = x127 | x255 ;
  assign n641 = x127 &  x255 ;
  assign n642 = ( n640 & ~n641 ) | ( n640 & 1'b0 ) | ( ~n641 & 1'b0 ) ;
  assign n643 = n638 &  n642 ;
  assign n644 = n638 | n642 ;
  assign n645 = ~n643 & n644 ;
  assign n646 = ( x127 & x255 ) | ( x127 & n638 ) | ( x255 & n638 ) ;
  assign y0 = n259 ;
  assign y1 = n263 ;
  assign y2 = n267 ;
  assign y3 = n270 ;
  assign y4 = n273 ;
  assign y5 = n276 ;
  assign y6 = n279 ;
  assign y7 = n282 ;
  assign y8 = n285 ;
  assign y9 = n288 ;
  assign y10 = n291 ;
  assign y11 = n294 ;
  assign y12 = n297 ;
  assign y13 = n300 ;
  assign y14 = n303 ;
  assign y15 = n306 ;
  assign y16 = n309 ;
  assign y17 = n312 ;
  assign y18 = n315 ;
  assign y19 = n318 ;
  assign y20 = n321 ;
  assign y21 = n324 ;
  assign y22 = n327 ;
  assign y23 = n330 ;
  assign y24 = n333 ;
  assign y25 = n336 ;
  assign y26 = n339 ;
  assign y27 = n342 ;
  assign y28 = n345 ;
  assign y29 = n348 ;
  assign y30 = n351 ;
  assign y31 = n354 ;
  assign y32 = n357 ;
  assign y33 = n360 ;
  assign y34 = n363 ;
  assign y35 = n366 ;
  assign y36 = n369 ;
  assign y37 = n372 ;
  assign y38 = n375 ;
  assign y39 = n378 ;
  assign y40 = n381 ;
  assign y41 = n384 ;
  assign y42 = n387 ;
  assign y43 = n390 ;
  assign y44 = n393 ;
  assign y45 = n396 ;
  assign y46 = n399 ;
  assign y47 = n402 ;
  assign y48 = n405 ;
  assign y49 = n408 ;
  assign y50 = n411 ;
  assign y51 = n414 ;
  assign y52 = n417 ;
  assign y53 = n420 ;
  assign y54 = n423 ;
  assign y55 = n426 ;
  assign y56 = n429 ;
  assign y57 = n432 ;
  assign y58 = n435 ;
  assign y59 = n438 ;
  assign y60 = n441 ;
  assign y61 = n444 ;
  assign y62 = n447 ;
  assign y63 = n450 ;
  assign y64 = n453 ;
  assign y65 = n456 ;
  assign y66 = n459 ;
  assign y67 = n462 ;
  assign y68 = n465 ;
  assign y69 = n468 ;
  assign y70 = n471 ;
  assign y71 = n474 ;
  assign y72 = n477 ;
  assign y73 = n480 ;
  assign y74 = n483 ;
  assign y75 = n486 ;
  assign y76 = n489 ;
  assign y77 = n492 ;
  assign y78 = n495 ;
  assign y79 = n498 ;
  assign y80 = n501 ;
  assign y81 = n504 ;
  assign y82 = n507 ;
  assign y83 = n510 ;
  assign y84 = n513 ;
  assign y85 = n516 ;
  assign y86 = n519 ;
  assign y87 = n522 ;
  assign y88 = n525 ;
  assign y89 = n528 ;
  assign y90 = n531 ;
  assign y91 = n534 ;
  assign y92 = n537 ;
  assign y93 = n540 ;
  assign y94 = n543 ;
  assign y95 = n546 ;
  assign y96 = n549 ;
  assign y97 = n552 ;
  assign y98 = n555 ;
  assign y99 = n558 ;
  assign y100 = n561 ;
  assign y101 = n564 ;
  assign y102 = n567 ;
  assign y103 = n570 ;
  assign y104 = n573 ;
  assign y105 = n576 ;
  assign y106 = n579 ;
  assign y107 = n582 ;
  assign y108 = n585 ;
  assign y109 = n588 ;
  assign y110 = n591 ;
  assign y111 = n594 ;
  assign y112 = n597 ;
  assign y113 = n600 ;
  assign y114 = n603 ;
  assign y115 = n606 ;
  assign y116 = n609 ;
  assign y117 = n612 ;
  assign y118 = n615 ;
  assign y119 = n618 ;
  assign y120 = n621 ;
  assign y121 = n624 ;
  assign y122 = n627 ;
  assign y123 = n630 ;
  assign y124 = n633 ;
  assign y125 = n636 ;
  assign y126 = n639 ;
  assign y127 = n645 ;
  assign y128 = n646 ;
endmodule
